module gpio (clk_i,
    rst_ni,
    alert_rx_i,
    alert_tx_o,
    cio_gpio_en_o,
    cio_gpio_i,
    cio_gpio_o,
    intr_gpio_o,
    tl_i,
    tl_o);
 input clk_i;
 input rst_ni;
 input [3:0] alert_rx_i;
 output [1:0] alert_tx_o;
 output [31:0] cio_gpio_en_o;
 input [31:0] cio_gpio_i;
 output [31:0] cio_gpio_o;
 output [31:0] intr_gpio_o;
 input [108:0] tl_i;
 output [65:0] tl_o;

 wire N113;
 wire N114;
 wire N115;
 wire N116;
 wire N117;
 wire N118;
 wire N119;
 wire N120;
 wire N121;
 wire N122;
 wire N123;
 wire N124;
 wire N125;
 wire N126;
 wire N127;
 wire N128;
 wire N129;
 wire N130;
 wire N131;
 wire N132;
 wire N133;
 wire N134;
 wire N135;
 wire N136;
 wire N137;
 wire N138;
 wire N139;
 wire N140;
 wire N141;
 wire N142;
 wire N143;
 wire N144;
 wire N145;
 wire N146;
 wire N38;
 wire N39;
 wire N40;
 wire N41;
 wire N42;
 wire N43;
 wire N44;
 wire N45;
 wire N46;
 wire N47;
 wire N48;
 wire N49;
 wire N50;
 wire N51;
 wire N52;
 wire N53;
 wire N54;
 wire N55;
 wire N56;
 wire N57;
 wire N58;
 wire N59;
 wire N60;
 wire N61;
 wire N62;
 wire N63;
 wire N64;
 wire N65;
 wire N66;
 wire N67;
 wire N68;
 wire N69;
 wire N70;
 wire N71;
 wire eq_x_101_n25;
 wire eq_x_106_n25;
 wire eq_x_111_n25;
 wire eq_x_116_n25;
 wire eq_x_121_n25;
 wire eq_x_126_n25;
 wire eq_x_131_n25;
 wire eq_x_136_n25;
 wire eq_x_141_n25;
 wire eq_x_146_n25;
 wire eq_x_151_n25;
 wire eq_x_156_n25;
 wire eq_x_161_n25;
 wire eq_x_166_n25;
 wire eq_x_171_n25;
 wire eq_x_176_n25;
 wire eq_x_181_n25;
 wire eq_x_26_n25;
 wire eq_x_31_n25;
 wire eq_x_36_n25;
 wire eq_x_41_n25;
 wire eq_x_46_n25;
 wire eq_x_51_n25;
 wire eq_x_56_n25;
 wire eq_x_61_n25;
 wire eq_x_66_n25;
 wire eq_x_71_n25;
 wire eq_x_76_n25;
 wire eq_x_81_n25;
 wire eq_x_86_n25;
 wire eq_x_91_n25;
 wire eq_x_96_n25;
 wire gen_alert_tx_0__u_prim_alert_sender_ack_level;
 wire gen_alert_tx_0__u_prim_alert_sender_alert_nd;
 wire gen_alert_tx_0__u_prim_alert_sender_alert_pd;
 wire gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger;
 wire gen_alert_tx_0__u_prim_alert_sender_alert_test_set_d;
 wire gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q;
 wire gen_alert_tx_0__u_prim_alert_sender_n1;
 wire gen_alert_tx_0__u_prim_alert_sender_ping_set_d;
 wire gen_alert_tx_0__u_prim_alert_sender_ping_set_q;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_intq_0_;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_intq_0_;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_intq_0_;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_intq_0_;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_n3;
 wire gen_filter_0__u_filter_filter_q;
 wire gen_filter_0__u_filter_filter_synced;
 wire gen_filter_0__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_0__u_filter_stored_value_q;
 wire gen_filter_10__u_filter_filter_q;
 wire gen_filter_10__u_filter_filter_synced;
 wire gen_filter_10__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_10__u_filter_stored_value_q;
 wire gen_filter_11__u_filter_filter_q;
 wire gen_filter_11__u_filter_filter_synced;
 wire gen_filter_11__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_11__u_filter_stored_value_q;
 wire gen_filter_12__u_filter_filter_q;
 wire gen_filter_12__u_filter_filter_synced;
 wire gen_filter_12__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_12__u_filter_stored_value_q;
 wire gen_filter_13__u_filter_filter_q;
 wire gen_filter_13__u_filter_filter_synced;
 wire gen_filter_13__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_13__u_filter_stored_value_q;
 wire gen_filter_14__u_filter_filter_q;
 wire gen_filter_14__u_filter_filter_synced;
 wire gen_filter_14__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_14__u_filter_stored_value_q;
 wire gen_filter_15__u_filter_filter_q;
 wire gen_filter_15__u_filter_filter_synced;
 wire gen_filter_15__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_15__u_filter_stored_value_q;
 wire gen_filter_16__u_filter_filter_q;
 wire gen_filter_16__u_filter_filter_synced;
 wire gen_filter_16__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_16__u_filter_stored_value_q;
 wire gen_filter_17__u_filter_filter_q;
 wire gen_filter_17__u_filter_filter_synced;
 wire gen_filter_17__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_17__u_filter_stored_value_q;
 wire gen_filter_18__u_filter_filter_q;
 wire gen_filter_18__u_filter_filter_synced;
 wire gen_filter_18__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_18__u_filter_stored_value_q;
 wire gen_filter_19__u_filter_filter_q;
 wire gen_filter_19__u_filter_filter_synced;
 wire gen_filter_19__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_19__u_filter_stored_value_q;
 wire gen_filter_1__u_filter_filter_q;
 wire gen_filter_1__u_filter_filter_synced;
 wire gen_filter_1__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_1__u_filter_stored_value_q;
 wire gen_filter_20__u_filter_filter_q;
 wire gen_filter_20__u_filter_filter_synced;
 wire gen_filter_20__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_20__u_filter_stored_value_q;
 wire gen_filter_21__u_filter_filter_q;
 wire gen_filter_21__u_filter_filter_synced;
 wire gen_filter_21__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_21__u_filter_stored_value_q;
 wire gen_filter_22__u_filter_filter_q;
 wire gen_filter_22__u_filter_filter_synced;
 wire gen_filter_22__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_22__u_filter_stored_value_q;
 wire gen_filter_23__u_filter_filter_q;
 wire gen_filter_23__u_filter_filter_synced;
 wire gen_filter_23__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_23__u_filter_stored_value_q;
 wire gen_filter_24__u_filter_filter_q;
 wire gen_filter_24__u_filter_filter_synced;
 wire gen_filter_24__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_24__u_filter_stored_value_q;
 wire gen_filter_25__u_filter_filter_q;
 wire gen_filter_25__u_filter_filter_synced;
 wire gen_filter_25__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_25__u_filter_stored_value_q;
 wire gen_filter_26__u_filter_filter_q;
 wire gen_filter_26__u_filter_filter_synced;
 wire gen_filter_26__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_26__u_filter_stored_value_q;
 wire gen_filter_27__u_filter_filter_q;
 wire gen_filter_27__u_filter_filter_synced;
 wire gen_filter_27__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_27__u_filter_stored_value_q;
 wire gen_filter_28__u_filter_filter_q;
 wire gen_filter_28__u_filter_filter_synced;
 wire gen_filter_28__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_28__u_filter_stored_value_q;
 wire gen_filter_29__u_filter_filter_q;
 wire gen_filter_29__u_filter_filter_synced;
 wire gen_filter_29__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_29__u_filter_stored_value_q;
 wire gen_filter_2__u_filter_filter_q;
 wire gen_filter_2__u_filter_filter_synced;
 wire gen_filter_2__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_2__u_filter_stored_value_q;
 wire gen_filter_30__u_filter_filter_q;
 wire gen_filter_30__u_filter_filter_synced;
 wire gen_filter_30__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_30__u_filter_stored_value_q;
 wire gen_filter_31__u_filter_filter_q;
 wire gen_filter_31__u_filter_filter_synced;
 wire gen_filter_31__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_31__u_filter_stored_value_q;
 wire gen_filter_3__u_filter_filter_q;
 wire gen_filter_3__u_filter_filter_synced;
 wire gen_filter_3__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_3__u_filter_stored_value_q;
 wire gen_filter_4__u_filter_filter_q;
 wire gen_filter_4__u_filter_filter_synced;
 wire gen_filter_4__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_4__u_filter_stored_value_q;
 wire gen_filter_5__u_filter_filter_q;
 wire gen_filter_5__u_filter_filter_synced;
 wire gen_filter_5__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_5__u_filter_stored_value_q;
 wire gen_filter_6__u_filter_filter_q;
 wire gen_filter_6__u_filter_filter_synced;
 wire gen_filter_6__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_6__u_filter_stored_value_q;
 wire gen_filter_7__u_filter_filter_q;
 wire gen_filter_7__u_filter_filter_synced;
 wire gen_filter_7__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_7__u_filter_stored_value_q;
 wire gen_filter_8__u_filter_filter_q;
 wire gen_filter_8__u_filter_filter_synced;
 wire gen_filter_8__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_8__u_filter_stored_value_q;
 wire gen_filter_9__u_filter_filter_q;
 wire gen_filter_9__u_filter_filter_synced;
 wire gen_filter_9__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_9__u_filter_stored_value_q;
 wire intr_hw_N1;
 wire intr_hw_N10;
 wire intr_hw_N11;
 wire intr_hw_N12;
 wire intr_hw_N13;
 wire intr_hw_N14;
 wire intr_hw_N15;
 wire intr_hw_N16;
 wire intr_hw_N17;
 wire intr_hw_N18;
 wire intr_hw_N19;
 wire intr_hw_N2;
 wire intr_hw_N20;
 wire intr_hw_N21;
 wire intr_hw_N22;
 wire intr_hw_N23;
 wire intr_hw_N24;
 wire intr_hw_N25;
 wire intr_hw_N26;
 wire intr_hw_N27;
 wire intr_hw_N28;
 wire intr_hw_N29;
 wire intr_hw_N3;
 wire intr_hw_N30;
 wire intr_hw_N31;
 wire intr_hw_N32;
 wire intr_hw_N4;
 wire intr_hw_N5;
 wire intr_hw_N6;
 wire intr_hw_N7;
 wire intr_hw_N8;
 wire intr_hw_N9;
 wire n1429;
 wire n1432;
 wire n1439;
 wire n2695;
 wire n2696;
 wire n2697;
 wire n2698;
 wire n2699;
 wire n2700;
 wire n2701;
 wire n2702;
 wire n2703;
 wire n2704;
 wire n2705;
 wire n2706;
 wire n2707;
 wire n2708;
 wire n2709;
 wire n2710;
 wire n2711;
 wire n2712;
 wire n2713;
 wire n2714;
 wire n2715;
 wire n2716;
 wire n2717;
 wire n2718;
 wire n2719;
 wire n2720;
 wire n2721;
 wire n2722;
 wire n2723;
 wire n2724;
 wire n2725;
 wire n2726;
 wire n2727;
 wire n2728;
 wire n2729;
 wire n2730;
 wire n2731;
 wire n2732;
 wire n2733;
 wire n2734;
 wire n2735;
 wire n2736;
 wire n2737;
 wire n2738;
 wire n2739;
 wire n2740;
 wire n2741;
 wire n2742;
 wire n2743;
 wire n2744;
 wire n2745;
 wire n2746;
 wire n2747;
 wire n2748;
 wire n2749;
 wire n2750;
 wire n2751;
 wire n2752;
 wire n2753;
 wire n2754;
 wire n2755;
 wire n2756;
 wire n2757;
 wire n2758;
 wire n2759;
 wire n2760;
 wire n2761;
 wire n2762;
 wire n2763;
 wire n2764;
 wire n2765;
 wire n2766;
 wire n2767;
 wire n2768;
 wire n2769;
 wire n2770;
 wire n2771;
 wire n2772;
 wire n2773;
 wire n2774;
 wire n2775;
 wire n2776;
 wire n2777;
 wire n2778;
 wire n2779;
 wire n2780;
 wire n2781;
 wire n2782;
 wire n2783;
 wire n2784;
 wire n2785;
 wire n2786;
 wire n2787;
 wire n2788;
 wire n2789;
 wire n2790;
 wire n2791;
 wire n2792;
 wire n2793;
 wire n2794;
 wire n2795;
 wire n2796;
 wire n2797;
 wire n2798;
 wire n2799;
 wire n2800;
 wire n2801;
 wire n2802;
 wire n2803;
 wire n2804;
 wire n2805;
 wire n2806;
 wire n2807;
 wire n2808;
 wire n2809;
 wire n2810;
 wire n2811;
 wire n2812;
 wire n2813;
 wire n2814;
 wire n2815;
 wire n2816;
 wire n2817;
 wire n2818;
 wire n2819;
 wire n2820;
 wire n2821;
 wire n2822;
 wire n2823;
 wire n2824;
 wire n2825;
 wire n2826;
 wire n2827;
 wire n2828;
 wire n2829;
 wire n2830;
 wire n2831;
 wire n2832;
 wire n2833;
 wire n2834;
 wire n2835;
 wire n2836;
 wire n2837;
 wire n2838;
 wire n2839;
 wire n2840;
 wire n2841;
 wire n2842;
 wire n2843;
 wire n2844;
 wire n2845;
 wire n2846;
 wire n2847;
 wire n2848;
 wire n2849;
 wire n2850;
 wire n2851;
 wire n2852;
 wire n2853;
 wire n2854;
 wire n2855;
 wire n2856;
 wire n2857;
 wire n2858;
 wire n2859;
 wire n2860;
 wire n2861;
 wire n2862;
 wire n2863;
 wire n2864;
 wire n2865;
 wire n2866;
 wire n2867;
 wire n2868;
 wire n2869;
 wire n2870;
 wire n2871;
 wire n2872;
 wire n2873;
 wire n2874;
 wire n2875;
 wire n2876;
 wire n2877;
 wire n2878;
 wire n2879;
 wire n2880;
 wire n2881;
 wire n2882;
 wire n2883;
 wire n2884;
 wire n2885;
 wire n2886;
 wire n2887;
 wire n2888;
 wire n2889;
 wire n2890;
 wire n2891;
 wire n2892;
 wire n2893;
 wire n2894;
 wire n2895;
 wire n2896;
 wire n2897;
 wire n2898;
 wire n2899;
 wire n2900;
 wire n2901;
 wire n2902;
 wire n2903;
 wire n2904;
 wire n2905;
 wire n2906;
 wire n2907;
 wire n2908;
 wire n2909;
 wire n2910;
 wire n2911;
 wire n2912;
 wire n2913;
 wire n2914;
 wire n2915;
 wire n2916;
 wire n2917;
 wire n2918;
 wire n2919;
 wire n2920;
 wire n2921;
 wire n2922;
 wire n2923;
 wire n2924;
 wire n2925;
 wire n2926;
 wire n2927;
 wire n2928;
 wire n2929;
 wire n2930;
 wire n2931;
 wire n2932;
 wire n2933;
 wire n2934;
 wire n2935;
 wire n2936;
 wire n2937;
 wire n2938;
 wire n2939;
 wire n2940;
 wire n2941;
 wire n2942;
 wire n2943;
 wire n2944;
 wire n2945;
 wire n2946;
 wire n2947;
 wire n2948;
 wire n2949;
 wire n2950;
 wire n2951;
 wire n2952;
 wire n2953;
 wire n2954;
 wire n2955;
 wire n2956;
 wire n2957;
 wire n2958;
 wire n2959;
 wire n2960;
 wire n2961;
 wire n2962;
 wire n2963;
 wire n2964;
 wire n2965;
 wire n2966;
 wire n2967;
 wire n2968;
 wire n2969;
 wire n2970;
 wire n2971;
 wire n2972;
 wire n2973;
 wire n2974;
 wire n2975;
 wire n2976;
 wire n2977;
 wire n2978;
 wire n2979;
 wire n2980;
 wire n2981;
 wire n2982;
 wire n2983;
 wire n2984;
 wire n2985;
 wire n2986;
 wire n2987;
 wire n2988;
 wire n2989;
 wire n2990;
 wire n2991;
 wire n2992;
 wire n2993;
 wire n2994;
 wire n2995;
 wire n2996;
 wire n2997;
 wire n2998;
 wire n2999;
 wire n3000;
 wire n3001;
 wire n3002;
 wire n3003;
 wire n3004;
 wire n3005;
 wire n3006;
 wire n3007;
 wire n3008;
 wire n3009;
 wire n3010;
 wire n3011;
 wire n3012;
 wire n3013;
 wire n3014;
 wire n3015;
 wire n3016;
 wire n3017;
 wire n3018;
 wire n3019;
 wire n3020;
 wire n3021;
 wire n3022;
 wire n3023;
 wire n3024;
 wire n3025;
 wire n3026;
 wire n3027;
 wire n3028;
 wire n3029;
 wire n3030;
 wire n3031;
 wire n3032;
 wire n3033;
 wire n3034;
 wire n3035;
 wire n3036;
 wire n3037;
 wire n3038;
 wire n3039;
 wire n3040;
 wire n3041;
 wire n3042;
 wire n3043;
 wire n3044;
 wire n3045;
 wire n3046;
 wire n3047;
 wire n3048;
 wire n3049;
 wire n3050;
 wire n3051;
 wire n3052;
 wire n3053;
 wire n3054;
 wire n3055;
 wire n3056;
 wire n3057;
 wire n3058;
 wire n3059;
 wire n3060;
 wire n3061;
 wire n3062;
 wire n3063;
 wire n3064;
 wire n3065;
 wire n3066;
 wire n3067;
 wire n3068;
 wire n3069;
 wire n3070;
 wire n3071;
 wire n3072;
 wire n3073;
 wire n3074;
 wire n3075;
 wire n3076;
 wire n3077;
 wire n3078;
 wire n3079;
 wire n3080;
 wire n3081;
 wire n3082;
 wire n3083;
 wire n3084;
 wire n3085;
 wire n3086;
 wire n3087;
 wire n3088;
 wire n3089;
 wire n3090;
 wire n3091;
 wire n3092;
 wire n3093;
 wire n3094;
 wire n3095;
 wire n3096;
 wire n3097;
 wire n3098;
 wire n3099;
 wire n3100;
 wire n3101;
 wire n3102;
 wire n3103;
 wire n3104;
 wire n3105;
 wire n3106;
 wire n3107;
 wire n3108;
 wire n3109;
 wire n3110;
 wire n3111;
 wire n3112;
 wire n3113;
 wire n3114;
 wire n3115;
 wire n3116;
 wire n3117;
 wire n3118;
 wire n3119;
 wire n3120;
 wire n3121;
 wire n3122;
 wire n3123;
 wire n3124;
 wire n3125;
 wire n3126;
 wire n3127;
 wire n3128;
 wire n3129;
 wire n3130;
 wire n3131;
 wire n3132;
 wire n3133;
 wire n3134;
 wire n3135;
 wire n3136;
 wire n3137;
 wire n3138;
 wire n3139;
 wire n3140;
 wire n3141;
 wire n3142;
 wire n3143;
 wire n3144;
 wire n3145;
 wire n3146;
 wire n3147;
 wire n3148;
 wire n3149;
 wire n3150;
 wire n3151;
 wire n3152;
 wire n3153;
 wire n3154;
 wire n3155;
 wire n3156;
 wire n3157;
 wire n3158;
 wire n3159;
 wire n3160;
 wire n3161;
 wire n3162;
 wire n3163;
 wire n3164;
 wire n3165;
 wire n3166;
 wire n3167;
 wire n3168;
 wire n3169;
 wire n3170;
 wire n3171;
 wire n3172;
 wire n3173;
 wire n3174;
 wire n3175;
 wire n3176;
 wire n3177;
 wire n3178;
 wire n3179;
 wire n3180;
 wire n3181;
 wire n3182;
 wire n3183;
 wire n3184;
 wire n3185;
 wire n3186;
 wire n3187;
 wire n3188;
 wire n3189;
 wire n3190;
 wire n3191;
 wire n3192;
 wire n3193;
 wire n3194;
 wire n3195;
 wire n3196;
 wire n3197;
 wire n3198;
 wire n3199;
 wire n3200;
 wire n3201;
 wire n3202;
 wire n3203;
 wire n3204;
 wire n3205;
 wire n3206;
 wire n3207;
 wire n3208;
 wire n3209;
 wire n3210;
 wire n3211;
 wire n3212;
 wire n3213;
 wire n3214;
 wire n3215;
 wire n3216;
 wire n3217;
 wire n3218;
 wire n3219;
 wire n3220;
 wire n3221;
 wire n3222;
 wire n3223;
 wire n3224;
 wire n3225;
 wire n3226;
 wire n3227;
 wire n3228;
 wire n3229;
 wire n3230;
 wire n3231;
 wire n3232;
 wire n3233;
 wire n3234;
 wire n3235;
 wire n3236;
 wire n3237;
 wire n3238;
 wire n3239;
 wire n3240;
 wire n3241;
 wire n3242;
 wire n3243;
 wire n3244;
 wire n3245;
 wire n3246;
 wire n3247;
 wire n3248;
 wire n3249;
 wire n3250;
 wire n3251;
 wire n3252;
 wire n3253;
 wire n3254;
 wire n3255;
 wire n3256;
 wire n3257;
 wire n3258;
 wire n3259;
 wire n3260;
 wire n3261;
 wire n3262;
 wire n3263;
 wire n3264;
 wire n3265;
 wire n3266;
 wire n3267;
 wire n3268;
 wire n3269;
 wire n3270;
 wire n3271;
 wire n3272;
 wire n3273;
 wire n3274;
 wire n3275;
 wire n3276;
 wire n3277;
 wire n3278;
 wire n3279;
 wire n3280;
 wire n3281;
 wire n3282;
 wire n3283;
 wire n3284;
 wire n3285;
 wire n3286;
 wire n3287;
 wire n3288;
 wire n3289;
 wire n3290;
 wire n3291;
 wire n3292;
 wire n3293;
 wire n3294;
 wire n3295;
 wire n3296;
 wire n3297;
 wire n3298;
 wire n3299;
 wire n3300;
 wire n3301;
 wire n3302;
 wire n3303;
 wire n3304;
 wire n3305;
 wire n3306;
 wire n3307;
 wire n3308;
 wire n3309;
 wire n3311;
 wire n3312;
 wire n3313;
 wire n3314;
 wire n3315;
 wire n3316;
 wire n3317;
 wire n3318;
 wire n3319;
 wire n3320;
 wire n3321;
 wire n3322;
 wire n3323;
 wire n3324;
 wire n3325;
 wire n3326;
 wire n3343;
 wire n3344;
 wire n3347;
 wire n3348;
 wire n3349;
 wire n3350;
 wire n3351;
 wire n3352;
 wire n3353;
 wire n3354;
 wire n3355;
 wire n3356;
 wire n3357;
 wire n3358;
 wire n3359;
 wire n3360;
 wire n3361;
 wire n3362;
 wire n3363;
 wire n3364;
 wire n3365;
 wire n3367;
 wire n3368;
 wire n3369;
 wire n3371;
 wire n3372;
 wire n3373;
 wire n3374;
 wire n3375;
 wire n3376;
 wire n3377;
 wire n3378;
 wire n3379;
 wire n3380;
 wire n3381;
 wire n3382;
 wire n3383;
 wire n3384;
 wire n3385;
 wire n3386;
 wire n3387;
 wire n3388;
 wire n3389;
 wire n3390;
 wire n3391;
 wire n3392;
 wire n3393;
 wire n3394;
 wire n3395;
 wire n3396;
 wire n3397;
 wire n3398;
 wire n3399;
 wire n3400;
 wire n3401;
 wire n3402;
 wire n3403;
 wire n3404;
 wire n3405;
 wire n3406;
 wire n3407;
 wire n3408;
 wire n3409;
 wire n3410;
 wire n3411;
 wire n3412;
 wire n3413;
 wire n3415;
 wire n3416;
 wire n3417;
 wire n3418;
 wire n3419;
 wire n3421;
 wire n3422;
 wire n3423;
 wire n3424;
 wire n3425;
 wire n3426;
 wire n3427;
 wire n3428;
 wire n3429;
 wire n3430;
 wire n3432;
 wire n3433;
 wire n3434;
 wire n3435;
 wire n3437;
 wire n3438;
 wire n3439;
 wire n3440;
 wire n3441;
 wire n3442;
 wire n3443;
 wire n3444;
 wire n3448;
 wire n3456;
 wire n3457;
 wire n3458;
 wire n3459;
 wire n3460;
 wire n3461;
 wire n3462;
 wire n3463;
 wire n3464;
 wire n3465;
 wire n3466;
 wire n3467;
 wire n3468;
 wire n3469;
 wire n3470;
 wire n3471;
 wire n3472;
 wire n3473;
 wire n3474;
 wire n3475;
 wire n3476;
 wire n3477;
 wire n3478;
 wire n3479;
 wire n3480;
 wire n3481;
 wire n3482;
 wire n3483;
 wire n3484;
 wire n3485;
 wire n3486;
 wire n3487;
 wire n3488;
 wire n3490;
 wire n3491;
 wire n3492;
 wire n3494;
 wire n3495;
 wire n3496;
 wire n3497;
 wire n3498;
 wire n3499;
 wire n3500;
 wire n3501;
 wire n3502;
 wire n3503;
 wire n3504;
 wire n3505;
 wire n3506;
 wire n3507;
 wire n3508;
 wire n3509;
 wire n3510;
 wire n3511;
 wire n3512;
 wire n3513;
 wire n3515;
 wire n3516;
 wire n3517;
 wire n3518;
 wire n3519;
 wire n3520;
 wire n3521;
 wire n3522;
 wire n3523;
 wire n3524;
 wire n3525;
 wire n3526;
 wire n3527;
 wire n3528;
 wire n3529;
 wire n3530;
 wire n3531;
 wire n3532;
 wire n3533;
 wire n3534;
 wire n3535;
 wire n3536;
 wire n3537;
 wire n3538;
 wire n3539;
 wire n3540;
 wire n3541;
 wire n3542;
 wire n3543;
 wire n3544;
 wire n3545;
 wire n3546;
 wire n3547;
 wire n3548;
 wire n3549;
 wire n3550;
 wire n3551;
 wire n3552;
 wire n3553;
 wire n3554;
 wire n3555;
 wire n3556;
 wire n3557;
 wire n3558;
 wire n3559;
 wire n3560;
 wire n3561;
 wire n3562;
 wire n3563;
 wire n3564;
 wire n3565;
 wire n3566;
 wire n3567;
 wire n3568;
 wire n3569;
 wire n3570;
 wire n3571;
 wire n3572;
 wire n3573;
 wire n3574;
 wire n3576;
 wire n3577;
 wire n3578;
 wire n3579;
 wire n3580;
 wire n3581;
 wire n3582;
 wire n3583;
 wire n3584;
 wire n3585;
 wire n3586;
 wire n3587;
 wire n3588;
 wire n3589;
 wire n3590;
 wire n3591;
 wire n3592;
 wire n3593;
 wire n3594;
 wire n3595;
 wire n3596;
 wire n3597;
 wire n3598;
 wire n3599;
 wire n3600;
 wire n3601;
 wire n3602;
 wire n3603;
 wire n3604;
 wire n3605;
 wire n3606;
 wire n3607;
 wire n3608;
 wire n3609;
 wire n3610;
 wire n3611;
 wire n3612;
 wire n3613;
 wire n3614;
 wire n3615;
 wire n3616;
 wire n3617;
 wire n3618;
 wire n3619;
 wire n3620;
 wire n3621;
 wire n3622;
 wire n3623;
 wire n3624;
 wire n3625;
 wire n3626;
 wire n3627;
 wire n3628;
 wire n3629;
 wire n3630;
 wire n3631;
 wire n3632;
 wire n3633;
 wire n3634;
 wire n3635;
 wire n3636;
 wire n3637;
 wire n3638;
 wire n3639;
 wire n3640;
 wire n3641;
 wire n3642;
 wire n3643;
 wire n3644;
 wire n3645;
 wire n3646;
 wire n3647;
 wire n3648;
 wire n3649;
 wire n3650;
 wire n3653;
 wire n3654;
 wire n3655;
 wire n3656;
 wire n3657;
 wire n3658;
 wire n3659;
 wire n3660;
 wire n3661;
 wire n3662;
 wire n3663;
 wire n3664;
 wire n3665;
 wire n3666;
 wire n3667;
 wire n3668;
 wire n3669;
 wire n3670;
 wire n3671;
 wire n3672;
 wire n3673;
 wire n3674;
 wire n3675;
 wire n3676;
 wire n3679;
 wire n3680;
 wire n3681;
 wire n3682;
 wire n3683;
 wire n3684;
 wire n3685;
 wire n3686;
 wire n3687;
 wire n3688;
 wire n3689;
 wire n3690;
 wire n3691;
 wire n3692;
 wire n3693;
 wire n3694;
 wire n3696;
 wire n3697;
 wire n3700;
 wire n3701;
 wire n3704;
 wire n3705;
 wire n3708;
 wire n3709;
 wire n3712;
 wire n3713;
 wire n3715;
 wire n3716;
 wire n3719;
 wire n3720;
 wire n3723;
 wire n3724;
 wire n3727;
 wire n3728;
 wire n3731;
 wire n3732;
 wire n3735;
 wire n3736;
 wire n3739;
 wire n3740;
 wire n3742;
 wire n3743;
 wire n3746;
 wire n3747;
 wire n3749;
 wire n3750;
 wire n3751;
 wire n3752;
 wire n3754;
 wire n3755;
 wire n3756;
 wire n3757;
 wire n3758;
 wire n3759;
 wire n3760;
 wire n3761;
 wire n3762;
 wire n3763;
 wire n3764;
 wire n3765;
 wire n3766;
 wire n3767;
 wire n3768;
 wire n3770;
 wire n3771;
 wire n3772;
 wire n3773;
 wire n3774;
 wire n3775;
 wire n3776;
 wire n3777;
 wire n3778;
 wire n3779;
 wire n3780;
 wire n3781;
 wire n3782;
 wire n3783;
 wire n3784;
 wire n3785;
 wire n3786;
 wire n3787;
 wire n3788;
 wire n3789;
 wire n3790;
 wire n3791;
 wire n3792;
 wire n3793;
 wire n3794;
 wire n3795;
 wire n3796;
 wire n3797;
 wire n3798;
 wire n3799;
 wire n3801;
 wire n3802;
 wire n3803;
 wire n3804;
 wire n3805;
 wire n3806;
 wire n3807;
 wire n3808;
 wire n3809;
 wire n3810;
 wire n3811;
 wire n3812;
 wire n3814;
 wire n3815;
 wire n3817;
 wire n3818;
 wire n3819;
 wire n3820;
 wire n3821;
 wire n3822;
 wire n3823;
 wire n3825;
 wire n3826;
 wire n3828;
 wire n3829;
 wire n3831;
 wire n3832;
 wire n3833;
 wire n3834;
 wire n3835;
 wire n3836;
 wire n3837;
 wire n3838;
 wire n3839;
 wire n3840;
 wire n3842;
 wire n3843;
 wire n3844;
 wire n3845;
 wire n3846;
 wire n3847;
 wire n3848;
 wire n3849;
 wire n3850;
 wire n3851;
 wire n3852;
 wire n3855;
 wire n3856;
 wire n3857;
 wire n3858;
 wire n3859;
 wire n3860;
 wire n3861;
 wire n3863;
 wire n3864;
 wire n3865;
 wire n3866;
 wire n3867;
 wire n3869;
 wire n3870;
 wire n3872;
 wire n3873;
 wire n3874;
 wire n3875;
 wire n3876;
 wire n3877;
 wire n3878;
 wire n3879;
 wire n3881;
 wire n3882;
 wire n3884;
 wire n3885;
 wire n3886;
 wire n3887;
 wire n3888;
 wire n3889;
 wire n3890;
 wire n3891;
 wire n3892;
 wire n3893;
 wire n3894;
 wire n3895;
 wire n3896;
 wire n3897;
 wire n3898;
 wire n3899;
 wire n3901;
 wire n3902;
 wire n3903;
 wire n3904;
 wire n3905;
 wire n3906;
 wire n3907;
 wire n3908;
 wire n3909;
 wire n3911;
 wire n3912;
 wire n3913;
 wire n3914;
 wire n3915;
 wire n3916;
 wire n3917;
 wire n3918;
 wire n3919;
 wire n3920;
 wire n3921;
 wire n3922;
 wire n3923;
 wire n3924;
 wire n3925;
 wire n3926;
 wire n3927;
 wire n3928;
 wire n3929;
 wire n3930;
 wire n3931;
 wire n3932;
 wire n3933;
 wire n3934;
 wire n3935;
 wire n3936;
 wire n3937;
 wire n3938;
 wire n3939;
 wire n3940;
 wire n3941;
 wire n3942;
 wire n3943;
 wire n3944;
 wire n3945;
 wire n3946;
 wire n3947;
 wire n3948;
 wire n3949;
 wire n3950;
 wire n3951;
 wire n3952;
 wire n3953;
 wire n3954;
 wire n3955;
 wire n3956;
 wire n3957;
 wire n3958;
 wire n3959;
 wire n3960;
 wire n3961;
 wire n3962;
 wire n3963;
 wire n3964;
 wire n3966;
 wire n3967;
 wire n3968;
 wire n3969;
 wire n3970;
 wire n3971;
 wire n3973;
 wire n3974;
 wire n3976;
 wire n3977;
 wire n3978;
 wire n3979;
 wire n3980;
 wire n3981;
 wire n3983;
 wire n3984;
 wire n3985;
 wire n3986;
 wire n3987;
 wire n3988;
 wire n3989;
 wire n3990;
 wire n3991;
 wire n3992;
 wire n3993;
 wire n3994;
 wire n3995;
 wire n3996;
 wire n3997;
 wire n3998;
 wire n3999;
 wire n4000;
 wire n4002;
 wire n4003;
 wire n4004;
 wire n4005;
 wire n4008;
 wire n4009;
 wire n4010;
 wire n4011;
 wire n4012;
 wire n4013;
 wire n4018;
 wire n4019;
 wire n4020;
 wire n4021;
 wire n4022;
 wire n4023;
 wire n4024;
 wire n4026;
 wire n4033;
 wire n4035;
 wire n4038;
 wire n4039;
 wire n4040;
 wire n4041;
 wire n4042;
 wire n4043;
 wire n4044;
 wire n4045;
 wire n4046;
 wire n4047;
 wire n4048;
 wire n4049;
 wire n4116;
 wire n4117;
 wire n4118;
 wire n4119;
 wire n4120;
 wire n4121;
 wire n4122;
 wire n4123;
 wire n4124;
 wire n4125;
 wire n4126;
 wire n4127;
 wire n4128;
 wire n4129;
 wire n4130;
 wire n4131;
 wire n4132;
 wire n4133;
 wire n4134;
 wire n4135;
 wire n4136;
 wire n4137;
 wire n4138;
 wire n4139;
 wire n4140;
 wire n4141;
 wire n4142;
 wire n4143;
 wire n4144;
 wire n4145;
 wire n4146;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire net66;
 wire net65;
 wire n4174;
 wire n4175;
 wire n4176;
 wire n4177;
 wire n4178;
 wire n4179;
 wire n4180;
 wire n4181;
 wire n4182;
 wire n4183;
 wire n4184;
 wire n4185;
 wire n4186;
 wire n4187;
 wire n4188;
 wire n4189;
 wire n4190;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire net20;
 wire net18;
 wire net17;
 wire net64;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire net12;
 wire net19;
 wire net2059;
 wire net2065;
 wire net2070;
 wire net2075;
 wire clknet_leaf_0_clk_i;
 wire reg2hw_ctrl_en_input_filter__q__0_;
 wire reg2hw_ctrl_en_input_filter__q__10_;
 wire reg2hw_ctrl_en_input_filter__q__11_;
 wire reg2hw_ctrl_en_input_filter__q__12_;
 wire reg2hw_ctrl_en_input_filter__q__13_;
 wire reg2hw_ctrl_en_input_filter__q__14_;
 wire reg2hw_ctrl_en_input_filter__q__15_;
 wire reg2hw_ctrl_en_input_filter__q__16_;
 wire reg2hw_ctrl_en_input_filter__q__17_;
 wire reg2hw_ctrl_en_input_filter__q__18_;
 wire reg2hw_ctrl_en_input_filter__q__19_;
 wire reg2hw_ctrl_en_input_filter__q__1_;
 wire reg2hw_ctrl_en_input_filter__q__20_;
 wire reg2hw_ctrl_en_input_filter__q__21_;
 wire reg2hw_ctrl_en_input_filter__q__22_;
 wire reg2hw_ctrl_en_input_filter__q__23_;
 wire reg2hw_ctrl_en_input_filter__q__24_;
 wire reg2hw_ctrl_en_input_filter__q__25_;
 wire reg2hw_ctrl_en_input_filter__q__26_;
 wire reg2hw_ctrl_en_input_filter__q__27_;
 wire reg2hw_ctrl_en_input_filter__q__28_;
 wire reg2hw_ctrl_en_input_filter__q__29_;
 wire reg2hw_ctrl_en_input_filter__q__2_;
 wire reg2hw_ctrl_en_input_filter__q__30_;
 wire reg2hw_ctrl_en_input_filter__q__31_;
 wire reg2hw_ctrl_en_input_filter__q__3_;
 wire reg2hw_ctrl_en_input_filter__q__4_;
 wire reg2hw_ctrl_en_input_filter__q__5_;
 wire reg2hw_ctrl_en_input_filter__q__6_;
 wire reg2hw_ctrl_en_input_filter__q__7_;
 wire reg2hw_ctrl_en_input_filter__q__8_;
 wire reg2hw_ctrl_en_input_filter__q__9_;
 wire reg2hw_intr_ctrl_en_falling__q__0_;
 wire reg2hw_intr_ctrl_en_falling__q__10_;
 wire reg2hw_intr_ctrl_en_falling__q__11_;
 wire reg2hw_intr_ctrl_en_falling__q__12_;
 wire reg2hw_intr_ctrl_en_falling__q__13_;
 wire reg2hw_intr_ctrl_en_falling__q__14_;
 wire reg2hw_intr_ctrl_en_falling__q__15_;
 wire reg2hw_intr_ctrl_en_falling__q__16_;
 wire reg2hw_intr_ctrl_en_falling__q__17_;
 wire reg2hw_intr_ctrl_en_falling__q__18_;
 wire reg2hw_intr_ctrl_en_falling__q__19_;
 wire reg2hw_intr_ctrl_en_falling__q__1_;
 wire reg2hw_intr_ctrl_en_falling__q__20_;
 wire reg2hw_intr_ctrl_en_falling__q__21_;
 wire reg2hw_intr_ctrl_en_falling__q__22_;
 wire reg2hw_intr_ctrl_en_falling__q__23_;
 wire reg2hw_intr_ctrl_en_falling__q__24_;
 wire reg2hw_intr_ctrl_en_falling__q__25_;
 wire reg2hw_intr_ctrl_en_falling__q__26_;
 wire reg2hw_intr_ctrl_en_falling__q__27_;
 wire reg2hw_intr_ctrl_en_falling__q__28_;
 wire reg2hw_intr_ctrl_en_falling__q__29_;
 wire reg2hw_intr_ctrl_en_falling__q__2_;
 wire reg2hw_intr_ctrl_en_falling__q__30_;
 wire reg2hw_intr_ctrl_en_falling__q__31_;
 wire reg2hw_intr_ctrl_en_falling__q__3_;
 wire reg2hw_intr_ctrl_en_falling__q__4_;
 wire reg2hw_intr_ctrl_en_falling__q__5_;
 wire reg2hw_intr_ctrl_en_falling__q__6_;
 wire reg2hw_intr_ctrl_en_falling__q__7_;
 wire reg2hw_intr_ctrl_en_falling__q__8_;
 wire reg2hw_intr_ctrl_en_falling__q__9_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__0_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__10_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__11_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__12_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__13_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__14_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__15_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__16_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__17_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__18_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__19_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__1_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__20_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__21_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__22_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__23_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__24_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__25_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__26_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__27_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__28_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__29_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__2_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__30_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__31_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__3_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__4_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__5_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__6_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__7_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__8_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__9_;
 wire reg2hw_intr_ctrl_en_lvllow__q__0_;
 wire reg2hw_intr_ctrl_en_lvllow__q__10_;
 wire reg2hw_intr_ctrl_en_lvllow__q__11_;
 wire reg2hw_intr_ctrl_en_lvllow__q__12_;
 wire reg2hw_intr_ctrl_en_lvllow__q__13_;
 wire reg2hw_intr_ctrl_en_lvllow__q__14_;
 wire reg2hw_intr_ctrl_en_lvllow__q__15_;
 wire reg2hw_intr_ctrl_en_lvllow__q__16_;
 wire reg2hw_intr_ctrl_en_lvllow__q__17_;
 wire reg2hw_intr_ctrl_en_lvllow__q__18_;
 wire reg2hw_intr_ctrl_en_lvllow__q__19_;
 wire reg2hw_intr_ctrl_en_lvllow__q__1_;
 wire reg2hw_intr_ctrl_en_lvllow__q__20_;
 wire reg2hw_intr_ctrl_en_lvllow__q__21_;
 wire reg2hw_intr_ctrl_en_lvllow__q__22_;
 wire reg2hw_intr_ctrl_en_lvllow__q__23_;
 wire reg2hw_intr_ctrl_en_lvllow__q__24_;
 wire reg2hw_intr_ctrl_en_lvllow__q__25_;
 wire reg2hw_intr_ctrl_en_lvllow__q__26_;
 wire reg2hw_intr_ctrl_en_lvllow__q__27_;
 wire reg2hw_intr_ctrl_en_lvllow__q__28_;
 wire reg2hw_intr_ctrl_en_lvllow__q__29_;
 wire reg2hw_intr_ctrl_en_lvllow__q__2_;
 wire reg2hw_intr_ctrl_en_lvllow__q__30_;
 wire reg2hw_intr_ctrl_en_lvllow__q__31_;
 wire reg2hw_intr_ctrl_en_lvllow__q__3_;
 wire reg2hw_intr_ctrl_en_lvllow__q__4_;
 wire reg2hw_intr_ctrl_en_lvllow__q__5_;
 wire reg2hw_intr_ctrl_en_lvllow__q__6_;
 wire reg2hw_intr_ctrl_en_lvllow__q__7_;
 wire reg2hw_intr_ctrl_en_lvllow__q__8_;
 wire reg2hw_intr_ctrl_en_lvllow__q__9_;
 wire reg2hw_intr_ctrl_en_rising__q__0_;
 wire reg2hw_intr_ctrl_en_rising__q__10_;
 wire reg2hw_intr_ctrl_en_rising__q__11_;
 wire reg2hw_intr_ctrl_en_rising__q__12_;
 wire reg2hw_intr_ctrl_en_rising__q__13_;
 wire reg2hw_intr_ctrl_en_rising__q__14_;
 wire reg2hw_intr_ctrl_en_rising__q__15_;
 wire reg2hw_intr_ctrl_en_rising__q__16_;
 wire reg2hw_intr_ctrl_en_rising__q__17_;
 wire reg2hw_intr_ctrl_en_rising__q__18_;
 wire reg2hw_intr_ctrl_en_rising__q__19_;
 wire reg2hw_intr_ctrl_en_rising__q__1_;
 wire reg2hw_intr_ctrl_en_rising__q__20_;
 wire reg2hw_intr_ctrl_en_rising__q__21_;
 wire reg2hw_intr_ctrl_en_rising__q__22_;
 wire reg2hw_intr_ctrl_en_rising__q__23_;
 wire reg2hw_intr_ctrl_en_rising__q__24_;
 wire reg2hw_intr_ctrl_en_rising__q__25_;
 wire reg2hw_intr_ctrl_en_rising__q__26_;
 wire reg2hw_intr_ctrl_en_rising__q__27_;
 wire reg2hw_intr_ctrl_en_rising__q__28_;
 wire reg2hw_intr_ctrl_en_rising__q__29_;
 wire reg2hw_intr_ctrl_en_rising__q__2_;
 wire reg2hw_intr_ctrl_en_rising__q__30_;
 wire reg2hw_intr_ctrl_en_rising__q__31_;
 wire reg2hw_intr_ctrl_en_rising__q__3_;
 wire reg2hw_intr_ctrl_en_rising__q__4_;
 wire reg2hw_intr_ctrl_en_rising__q__5_;
 wire reg2hw_intr_ctrl_en_rising__q__6_;
 wire reg2hw_intr_ctrl_en_rising__q__7_;
 wire reg2hw_intr_ctrl_en_rising__q__8_;
 wire reg2hw_intr_ctrl_en_rising__q__9_;
 wire reg2hw_intr_enable__q__0_;
 wire reg2hw_intr_enable__q__10_;
 wire reg2hw_intr_enable__q__11_;
 wire reg2hw_intr_enable__q__12_;
 wire reg2hw_intr_enable__q__13_;
 wire reg2hw_intr_enable__q__14_;
 wire reg2hw_intr_enable__q__15_;
 wire reg2hw_intr_enable__q__16_;
 wire reg2hw_intr_enable__q__17_;
 wire reg2hw_intr_enable__q__18_;
 wire reg2hw_intr_enable__q__19_;
 wire reg2hw_intr_enable__q__1_;
 wire reg2hw_intr_enable__q__20_;
 wire reg2hw_intr_enable__q__21_;
 wire reg2hw_intr_enable__q__22_;
 wire reg2hw_intr_enable__q__23_;
 wire reg2hw_intr_enable__q__24_;
 wire reg2hw_intr_enable__q__25_;
 wire reg2hw_intr_enable__q__26_;
 wire reg2hw_intr_enable__q__27_;
 wire reg2hw_intr_enable__q__28_;
 wire reg2hw_intr_enable__q__29_;
 wire reg2hw_intr_enable__q__2_;
 wire reg2hw_intr_enable__q__30_;
 wire reg2hw_intr_enable__q__31_;
 wire reg2hw_intr_enable__q__3_;
 wire reg2hw_intr_enable__q__4_;
 wire reg2hw_intr_enable__q__5_;
 wire reg2hw_intr_enable__q__6_;
 wire reg2hw_intr_enable__q__7_;
 wire reg2hw_intr_enable__q__8_;
 wire reg2hw_intr_enable__q__9_;
 wire reg2hw_intr_state__q__0_;
 wire reg2hw_intr_state__q__10_;
 wire reg2hw_intr_state__q__11_;
 wire reg2hw_intr_state__q__12_;
 wire reg2hw_intr_state__q__13_;
 wire reg2hw_intr_state__q__14_;
 wire reg2hw_intr_state__q__15_;
 wire reg2hw_intr_state__q__16_;
 wire reg2hw_intr_state__q__17_;
 wire reg2hw_intr_state__q__18_;
 wire reg2hw_intr_state__q__19_;
 wire reg2hw_intr_state__q__1_;
 wire reg2hw_intr_state__q__20_;
 wire reg2hw_intr_state__q__21_;
 wire reg2hw_intr_state__q__22_;
 wire reg2hw_intr_state__q__23_;
 wire reg2hw_intr_state__q__24_;
 wire reg2hw_intr_state__q__25_;
 wire reg2hw_intr_state__q__26_;
 wire reg2hw_intr_state__q__27_;
 wire reg2hw_intr_state__q__28_;
 wire reg2hw_intr_state__q__29_;
 wire reg2hw_intr_state__q__2_;
 wire reg2hw_intr_state__q__30_;
 wire reg2hw_intr_state__q__31_;
 wire reg2hw_intr_state__q__3_;
 wire reg2hw_intr_state__q__4_;
 wire reg2hw_intr_state__q__5_;
 wire reg2hw_intr_state__q__6_;
 wire reg2hw_intr_state__q__7_;
 wire reg2hw_intr_state__q__8_;
 wire reg2hw_intr_state__q__9_;
 wire u_reg_err_q;
 wire u_reg_reg_we_check_15_;
 wire u_reg_u_ctrl_en_input_filter_net2092;
 wire u_reg_u_ctrl_en_input_filter_net2098;
 wire u_reg_u_intr_ctrl_en_falling_net2092;
 wire u_reg_u_intr_ctrl_en_falling_net2098;
 wire u_reg_u_intr_ctrl_en_lvlhigh_net2092;
 wire u_reg_u_intr_ctrl_en_lvlhigh_net2098;
 wire u_reg_u_intr_ctrl_en_lvllow_net2092;
 wire u_reg_u_intr_ctrl_en_lvllow_net2098;
 wire u_reg_u_intr_ctrl_en_rising_net2092;
 wire u_reg_u_intr_ctrl_en_rising_net2098;
 wire u_reg_u_intr_enable_net2092;
 wire u_reg_u_intr_enable_net2098;
 wire u_reg_u_intr_state_n1;
 wire u_reg_u_intr_state_net2115;
 wire u_reg_u_intr_state_net2121;
 wire u_reg_u_reg_if_N14;
 wire u_reg_u_reg_if_N15;
 wire u_reg_u_reg_if_N16;
 wire u_reg_u_reg_if_N17;
 wire u_reg_u_reg_if_N18;
 wire u_reg_u_reg_if_N19;
 wire u_reg_u_reg_if_N20;
 wire u_reg_u_reg_if_N21;
 wire u_reg_u_reg_if_N22;
 wire u_reg_u_reg_if_N23;
 wire u_reg_u_reg_if_N24;
 wire u_reg_u_reg_if_N25;
 wire u_reg_u_reg_if_N26;
 wire u_reg_u_reg_if_N27;
 wire u_reg_u_reg_if_N28;
 wire u_reg_u_reg_if_N29;
 wire u_reg_u_reg_if_N30;
 wire u_reg_u_reg_if_N31;
 wire u_reg_u_reg_if_N32;
 wire u_reg_u_reg_if_N33;
 wire u_reg_u_reg_if_N34;
 wire u_reg_u_reg_if_N35;
 wire u_reg_u_reg_if_N36;
 wire u_reg_u_reg_if_N37;
 wire u_reg_u_reg_if_N38;
 wire u_reg_u_reg_if_N39;
 wire u_reg_u_reg_if_N40;
 wire u_reg_u_reg_if_N41;
 wire u_reg_u_reg_if_N42;
 wire u_reg_u_reg_if_N43;
 wire u_reg_u_reg_if_N44;
 wire u_reg_u_reg_if_N45;
 wire u_reg_u_reg_if_N46;
 wire u_reg_u_reg_if_N7;
 wire u_reg_u_reg_if_a_ack;
 wire u_reg_u_reg_if_net2138;
 wire u_reg_u_reg_if_net2144;
 wire u_reg_u_reg_if_net2149;
 wire u_reg_u_reg_if_rd_req;
 wire net1496;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_13_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_0_clk_i;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_1_1__leaf_clk_i;
 wire clknet_0_u_reg_u_reg_if_net2138;
 wire clknet_1_0__leaf_u_reg_u_reg_if_net2138;
 wire clknet_1_1__leaf_u_reg_u_reg_if_net2138;
 wire clknet_0_u_reg_u_reg_if_net2144;
 wire clknet_1_0__leaf_u_reg_u_reg_if_net2144;
 wire clknet_1_1__leaf_u_reg_u_reg_if_net2144;
 wire clknet_0_u_reg_u_reg_if_net2149;
 wire clknet_1_0__leaf_u_reg_u_reg_if_net2149;
 wire clknet_1_1__leaf_u_reg_u_reg_if_net2149;
 wire clknet_0_u_reg_u_intr_state_net2115;
 wire clknet_1_0__leaf_u_reg_u_intr_state_net2115;
 wire clknet_1_1__leaf_u_reg_u_intr_state_net2115;
 wire clknet_0_u_reg_u_intr_state_net2121;
 wire clknet_1_0__leaf_u_reg_u_intr_state_net2121;
 wire clknet_1_1__leaf_u_reg_u_intr_state_net2121;
 wire clknet_0_u_reg_u_intr_enable_net2092;
 wire clknet_1_0__leaf_u_reg_u_intr_enable_net2092;
 wire clknet_1_1__leaf_u_reg_u_intr_enable_net2092;
 wire clknet_0_u_reg_u_intr_enable_net2098;
 wire clknet_1_0__leaf_u_reg_u_intr_enable_net2098;
 wire clknet_1_1__leaf_u_reg_u_intr_enable_net2098;
 wire clknet_0_u_reg_u_intr_ctrl_en_rising_net2092;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2092;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2092;
 wire clknet_0_u_reg_u_intr_ctrl_en_rising_net2098;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2098;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2098;
 wire clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2092;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092;
 wire clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2098;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098;
 wire clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2092;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092;
 wire clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2098;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098;
 wire clknet_0_u_reg_u_intr_ctrl_en_falling_net2092;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2092;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2092;
 wire clknet_0_u_reg_u_intr_ctrl_en_falling_net2098;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2098;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2098;
 wire clknet_0_u_reg_u_ctrl_en_input_filter_net2092;
 wire clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2092;
 wire clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2092;
 wire clknet_0_u_reg_u_ctrl_en_input_filter_net2098;
 wire clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2098;
 wire clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2098;
 wire clknet_0_net2059;
 wire clknet_1_0__leaf_net2059;
 wire clknet_1_1__leaf_net2059;
 wire clknet_0_net2065;
 wire clknet_1_0__leaf_net2065;
 wire clknet_1_1__leaf_net2065;
 wire clknet_0_net2070;
 wire clknet_1_0__leaf_net2070;
 wire clknet_1_1__leaf_net2070;
 wire clknet_0_net2075;
 wire clknet_1_0__leaf_net2075;
 wire clknet_1_1__leaf_net2075;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire [31:0] data_in_q;
 wire [2:0] gen_alert_tx_0__u_prim_alert_sender_state_d;
 wire [2:0] gen_alert_tx_0__u_prim_alert_sender_state_q;
 wire [1:0] gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d;
 wire [1:0] gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q;
 wire [1:0] gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d;
 wire [1:0] gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q;
 wire [3:0] gen_filter_0__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_0__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_10__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_10__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_11__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_11__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_12__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_12__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_13__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_13__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_14__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_14__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_15__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_15__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_16__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_16__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_17__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_17__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_18__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_18__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_19__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_19__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_1__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_1__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_20__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_20__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_21__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_21__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_22__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_22__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_23__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_23__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_24__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_24__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_25__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_25__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_26__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_26__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_27__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_27__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_28__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_28__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_29__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_29__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_2__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_2__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_30__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_30__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_31__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_31__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_3__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_3__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_4__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_4__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_5__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_5__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_6__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_6__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_7__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_7__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_8__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_8__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_9__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_9__u_filter_diff_ctr_q;
 wire [31:0] u_reg_data_in_qs;
 wire [31:0] u_reg_u_ctrl_en_input_filter_wr_data;
 wire [31:0] u_reg_u_data_in_wr_data;
 wire [31:0] u_reg_u_intr_ctrl_en_falling_wr_data;
 wire [31:0] u_reg_u_intr_ctrl_en_lvlhigh_wr_data;
 wire [31:0] u_reg_u_intr_ctrl_en_lvllow_wr_data;
 wire [31:0] u_reg_u_intr_ctrl_en_rising_wr_data;
 wire [31:0] u_reg_u_intr_enable_wr_data;
 wire [31:0] u_reg_u_intr_state_wr_data;

 b15bfm201ah1n02x5 U3252 (.a(net1990),
    .o(net241));
 b15bfn000al1n02x5 U3253 (.a(net1919),
    .o(net243));
 b15inv040as1n36x5 U3254 (.a(net724),
    .o1(n4116));
 b15inv000as1n40x5 U3255 (.a(net723),
    .o1(n4117));
 b15inv000ah1n48x5 U3256 (.a(net722),
    .o1(n4118));
 b15and002al1n02x5 U3257 (.a(net516),
    .b(reg2hw_intr_enable__q__10_),
    .o(intr_hw_N22));
 b15and002ar1n08x5 U3258 (.a(reg2hw_intr_state__q__2_),
    .b(reg2hw_intr_enable__q__2_),
    .o(intr_hw_N30));
 b15and002ar1n02x5 U3259 (.a(net517),
    .b(reg2hw_intr_enable__q__1_),
    .o(intr_hw_N31));
 b15and002al1n16x5 U3260 (.a(reg2hw_intr_state__q__8_),
    .b(reg2hw_intr_enable__q__8_),
    .o(intr_hw_N24));
 b15and002ah1n04x5 U3261 (.a(net505),
    .b(reg2hw_intr_enable__q__6_),
    .o(intr_hw_N26));
 b15and002ar1n08x5 U3262 (.a(reg2hw_intr_state__q__14_),
    .b(reg2hw_intr_enable__q__14_),
    .o(intr_hw_N18));
 b15and002ar1n16x5 U3263 (.a(reg2hw_intr_state__q__9_),
    .b(reg2hw_intr_enable__q__9_),
    .o(intr_hw_N23));
 b15and002al1n08x5 U3264 (.a(reg2hw_intr_state__q__7_),
    .b(reg2hw_intr_enable__q__7_),
    .o(intr_hw_N25));
 b15and002an1n03x5 U3265 (.a(reg2hw_intr_state__q__18_),
    .b(reg2hw_intr_enable__q__18_),
    .o(intr_hw_N14));
 b15and002an1n08x5 U3266 (.a(net515),
    .b(reg2hw_intr_enable__q__11_),
    .o(intr_hw_N21));
 b15and002aq1n16x5 U3267 (.a(reg2hw_intr_state__q__3_),
    .b(reg2hw_intr_enable__q__3_),
    .o(intr_hw_N29));
 b15and002al1n04x5 U3268 (.a(reg2hw_intr_state__q__13_),
    .b(net523),
    .o(intr_hw_N19));
 b15and002as1n08x5 U3269 (.a(net508),
    .b(reg2hw_intr_enable__q__4_),
    .o(intr_hw_N28));
 b15and002al1n02x5 U3270 (.a(net507),
    .b(net518),
    .o(intr_hw_N27));
 b15and002aq1n02x5 U3271 (.a(reg2hw_intr_state__q__12_),
    .b(net524),
    .o(intr_hw_N20));
 b15and002aq1n12x5 U3272 (.a(net2474),
    .b(reg2hw_intr_state__q__30_),
    .o(intr_hw_N2));
 b15and002ar1n12x5 U3273 (.a(reg2hw_intr_enable__q__19_),
    .b(reg2hw_intr_state__q__19_),
    .o(intr_hw_N13));
 b15and002an1n02x5 U3274 (.a(reg2hw_intr_enable__q__29_),
    .b(net510),
    .o(intr_hw_N3));
 b15and002ar1n16x5 U3275 (.a(reg2hw_intr_enable__q__26_),
    .b(reg2hw_intr_state__q__26_),
    .o(intr_hw_N6));
 b15and002al1n08x5 U3276 (.a(net519),
    .b(reg2hw_intr_state__q__27_),
    .o(intr_hw_N5));
 b15and002al1n02x5 U3277 (.a(reg2hw_intr_enable__q__16_),
    .b(reg2hw_intr_state__q__16_),
    .o(intr_hw_N16));
 b15and002aq1n02x5 U3278 (.a(reg2hw_intr_enable__q__22_),
    .b(reg2hw_intr_state__q__22_),
    .o(intr_hw_N10));
 b15and002ar1n03x5 U3279 (.a(reg2hw_intr_enable__q__28_),
    .b(reg2hw_intr_state__q__28_),
    .o(intr_hw_N4));
 b15and002ar1n08x5 U3280 (.a(reg2hw_intr_enable__q__20_),
    .b(reg2hw_intr_state__q__20_),
    .o(intr_hw_N12));
 b15and002al1n08x5 U3281 (.a(net520),
    .b(reg2hw_intr_state__q__25_),
    .o(intr_hw_N7));
 b15and002al1n08x5 U3282 (.a(reg2hw_intr_enable__q__21_),
    .b(reg2hw_intr_state__q__21_),
    .o(intr_hw_N11));
 b15and002an1n04x5 U3283 (.a(reg2hw_intr_enable__q__17_),
    .b(reg2hw_intr_state__q__17_),
    .o(intr_hw_N15));
 b15and002aq1n12x5 U3284 (.a(reg2hw_intr_enable__q__31_),
    .b(reg2hw_intr_state__q__31_),
    .o(intr_hw_N1));
 b15and002ah1n04x5 U3285 (.a(net521),
    .b(reg2hw_intr_state__q__24_),
    .o(intr_hw_N8));
 b15and002al1n03x5 U3286 (.a(reg2hw_intr_enable__q__23_),
    .b(reg2hw_intr_state__q__23_),
    .o(intr_hw_N9));
 b15and002al1n02x5 U3287 (.a(reg2hw_intr_enable__q__15_),
    .b(net511),
    .o(intr_hw_N17));
 b15and002ah1n16x5 U3288 (.a(reg2hw_intr_enable__q__0_),
    .b(reg2hw_intr_state__q__0_),
    .o(intr_hw_N32));
 b15inv020aq1n64x5 U3289 (.a(net721),
    .o1(n4119));
 b15inv000as1n56x5 U3290 (.a(net720),
    .o1(n4120));
 b15inv020as1n64x5 U3291 (.a(net62),
    .o1(n4121));
 b15inv000as1n56x5 U3292 (.a(net63),
    .o1(n4122));
 b15inv020aq1n64x5 U3293 (.a(net719),
    .o1(n4123));
 b15inv000al1n80x5 U3294 (.a(net65),
    .o1(n4124));
 b15inv040as1n40x5 U3295 (.a(net66),
    .o1(n4125));
 b15inv040an1n60x5 U3296 (.a(net67),
    .o1(n4126));
 b15inv020as1n64x5 U3297 (.a(net68),
    .o1(n4127));
 b15inv000as1n28x5 U3298 (.a(net718),
    .o1(n4128));
 b15inv000as1n48x5 U3299 (.a(net717),
    .o1(n4129));
 b15inv020as1n64x5 U3300 (.a(net716),
    .o1(n4130));
 b15inv000as1n64x5 U3301 (.a(net715),
    .o1(n4131));
 b15inv020ah1n64x5 U3302 (.a(net75),
    .o1(n4132));
 b15inv040aq1n48x5 U3303 (.a(net714),
    .o1(n4133));
 b15inv000as1n80x5 U3304 (.a(net77),
    .o1(n4134));
 b15inv040as1n40x5 U3305 (.a(net713),
    .o1(n4135));
 b15inv000ah1n48x5 U3306 (.a(net79),
    .o1(n4136));
 b15inv000as1n48x5 U3307 (.a(net80),
    .o1(n4137));
 b15inv000ah1n64x5 U3308 (.a(net712),
    .o1(n4138));
 b15inv020as1n10x5 U3309 (.a(net82),
    .o1(n4139));
 b15inv000as1n56x5 U3310 (.a(net84),
    .o1(n4140));
 b15inv000as1n64x5 U3311 (.a(net85),
    .o1(n4141));
 b15inv000as1n64x5 U3312 (.a(net711),
    .o1(n4142));
 b15inv000as1n80x5 U3313 (.a(net87),
    .o1(n4143));
 b15inv040as1n40x5 U3314 (.a(net88),
    .o1(n4144));
 b15inv020an1n80x5 U3315 (.a(net89),
    .o1(n4145));
 b15inv040as1n28x5 U3316 (.a(net709),
    .o1(n4146));
 b15ztpn00an1n08x5 PHY_91 ();
 b15ztpn00an1n08x5 PHY_90 ();
 b15ztpn00an1n08x5 PHY_89 ();
 b15ztpn00an1n08x5 PHY_88 ();
 b15ztpn00an1n08x5 PHY_87 ();
 b15ztpn00an1n08x5 PHY_86 ();
 b15ztpn00an1n08x5 PHY_85 ();
 b15ztpn00an1n08x5 PHY_84 ();
 b15ztpn00an1n08x5 PHY_83 ();
 b15ztpn00an1n08x5 PHY_82 ();
 b15ztpn00an1n08x5 PHY_81 ();
 b15ztpn00an1n08x5 PHY_80 ();
 b15ztpn00an1n08x5 PHY_79 ();
 b15ztpn00an1n08x5 PHY_78 ();
 b15ztpn00an1n08x5 PHY_77 ();
 b15ztpn00an1n08x5 PHY_76 ();
 b15ztpn00an1n08x5 PHY_75 ();
 b15ztpn00an1n08x5 PHY_74 ();
 b15ztpn00an1n08x5 PHY_73 ();
 b15ztpn00an1n08x5 PHY_72 ();
 b15ztpn00an1n08x5 PHY_71 ();
 b15ztpn00an1n08x5 PHY_70 ();
 b15inv000ar1n03x5 U3339 (.a(net1496),
    .o1(tl_o[48]));
 b15ztpn00an1n08x5 PHY_69 ();
 b15ztpn00an1n08x5 PHY_68 ();
 b15ztpn00an1n08x5 PHY_67 ();
 b15ztpn00an1n08x5 PHY_66 ();
 b15inv000ar1n28x5 U3344 (.a(net433),
    .o1(n4174));
 b15inv000as1n80x5 U3345 (.a(net416),
    .o1(n4175));
 b15inv020ah1n64x5 U3346 (.a(net367),
    .o1(n4176));
 b15inv000ah1n10x5 U3347 (.a(net385),
    .o1(n4177));
 b15inv040as1n16x5 U3348 (.a(net357),
    .o1(n4178));
 b15inv020ar1n06x5 U3349 (.a(net359),
    .o1(n4179));
 b15inv000aq1n04x5 U3350 (.a(net334),
    .o1(n4180));
 b15inv000as1n48x5 U3351 (.a(n3749),
    .o1(n4181));
 b15inv040aq1n28x5 U3352 (.a(net336),
    .o1(n4182));
 b15inv020an1n16x5 U3353 (.a(net338),
    .o1(n4183));
 b15inv000as1n24x5 U3354 (.a(net346),
    .o1(n4184));
 b15inv040as1n20x5 U3355 (.a(net347),
    .o1(n4185));
 b15inv040as1n48x5 U3356 (.a(net328),
    .o1(n4186));
 b15inv020an1n28x5 U3357 (.a(u_reg_reg_we_check_15_),
    .o1(n4187));
 b15inv000as1n40x5 U3358 (.a(n3861),
    .o1(n4188));
 b15inv000al1n80x5 U3359 (.a(net304),
    .o1(n4189));
 b15inv000al1n20x5 U3360 (.a(net312),
    .o1(n4190));
 b15inv000ar1n03x5 U3362 (.a(net1497),
    .o1(tl_o[59]));
 b15inv000ar1n03x5 U3364 (.a(net1498),
    .o1(tl_o[60]));
 b15inv000ar1n03x5 U3366 (.a(net1499),
    .o1(tl_o[61]));
 b15ztpn00an1n08x5 PHY_65 ();
 b15nand03as1n06x5 U3369 (.a(gen_filter_19__u_filter_diff_ctr_q[1]),
    .b(gen_filter_19__u_filter_diff_ctr_q[3]),
    .c(net2306),
    .o1(n2788));
 b15xor002as1n06x5 U3370 (.a(net686),
    .b(net2276),
    .out0(n2785));
 b15aoi012aq1n02x5 U3371 (.a(n2785),
    .b(gen_filter_19__u_filter_diff_ctr_q[0]),
    .c(n2788),
    .o1(gen_filter_19__u_filter_diff_ctr_d[0]));
 b15inv000ar1n06x5 U3372 (.a(net1997),
    .o1(net237));
 b15xor002aq1n16x5 U3373 (.a(net683),
    .b(net2425),
    .out0(n2737));
 b15and002an1n02x5 U3374 (.a(net2381),
    .b(gen_filter_26__u_filter_diff_ctr_q[1]),
    .o(n2735));
 b15nand03as1n04x5 U3375 (.a(net2381),
    .b(gen_filter_26__u_filter_diff_ctr_q[1]),
    .c(gen_filter_26__u_filter_diff_ctr_q[2]),
    .o1(n2697));
 b15oai022ar1n02x5 U3376 (.a(n2735),
    .b(net2463),
    .c(gen_filter_26__u_filter_diff_ctr_q[3]),
    .d(n2697),
    .o1(n2695));
 b15norp02ar1n02x5 U3377 (.a(n2737),
    .b(n2695),
    .o1(gen_filter_26__u_filter_diff_ctr_d[2]));
 b15and002ar1n02x5 U3378 (.a(gen_filter_19__u_filter_diff_ctr_q[1]),
    .b(gen_filter_19__u_filter_diff_ctr_q[0]),
    .o(n2732));
 b15nandp3an1n04x5 U3379 (.a(gen_filter_19__u_filter_diff_ctr_q[1]),
    .b(net2294),
    .c(gen_filter_19__u_filter_diff_ctr_q[0]),
    .o1(n2786));
 b15oai022ar1n02x5 U3380 (.a(net2294),
    .b(n2732),
    .c(net2314),
    .d(n2786),
    .o1(n2696));
 b15norp02ar1n02x5 U3381 (.a(n2785),
    .b(n2696),
    .o1(gen_filter_19__u_filter_diff_ctr_d[2]));
 b15and003al1n04x5 U3382 (.a(gen_filter_9__u_filter_diff_ctr_q[0]),
    .b(gen_filter_9__u_filter_diff_ctr_q[1]),
    .c(net2358),
    .o(n2780));
 b15xor002ah1n08x5 U3383 (.a(gen_filter_9__u_filter_filter_synced),
    .b(net2332),
    .out0(n2808));
 b15oab012ar1n02x5 U3384 (.a(n2808),
    .b(net2279),
    .c(n2780),
    .out0(gen_filter_9__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3385 (.a(gen_filter_26__u_filter_diff_ctr_q[3]),
    .o1(n2698));
 b15aoi012ar1n02x5 U3386 (.a(n2737),
    .b(n2698),
    .c(n2697),
    .o1(gen_filter_26__u_filter_diff_ctr_d[3]));
 b15nand03ar1n16x5 U3387 (.a(gen_filter_26__u_filter_diff_ctr_q[3]),
    .b(gen_filter_26__u_filter_diff_ctr_q[1]),
    .c(gen_filter_26__u_filter_diff_ctr_q[2]),
    .o1(n2736));
 b15aoi012al1n04x5 U3388 (.a(n2737),
    .b(net2381),
    .c(n2736),
    .o1(gen_filter_26__u_filter_diff_ctr_d[0]));
 b15and003ah1n02x5 U3389 (.a(gen_filter_24__u_filter_diff_ctr_q[0]),
    .b(gen_filter_24__u_filter_diff_ctr_q[1]),
    .c(net2260),
    .o(n2741));
 b15xor002as1n06x5 U3390 (.a(gen_filter_24__u_filter_filter_synced),
    .b(net2241),
    .out0(n2810));
 b15oab012ar1n02x5 U3391 (.a(n2810),
    .b(net2281),
    .c(n2741),
    .out0(gen_filter_24__u_filter_diff_ctr_d[3]));
 b15and003aq1n03x5 U3392 (.a(gen_filter_0__u_filter_diff_ctr_q[2]),
    .b(net2402),
    .c(gen_filter_0__u_filter_diff_ctr_q[1]),
    .o(n2772));
 b15xor002as1n06x5 U3393 (.a(gen_filter_0__u_filter_filter_synced),
    .b(net2302),
    .out0(n2767));
 b15oab012al1n02x5 U3394 (.a(n2767),
    .b(gen_filter_0__u_filter_diff_ctr_q[3]),
    .c(n2772),
    .out0(gen_filter_0__u_filter_diff_ctr_d[3]));
 b15and003al1n04x5 U3395 (.a(gen_filter_6__u_filter_diff_ctr_q[0]),
    .b(net2566),
    .c(net2354),
    .o(n2740));
 b15xor002ah1n08x5 U3396 (.a(net679),
    .b(net2265),
    .out0(n2794));
 b15oab012an1n02x5 U3397 (.a(n2794),
    .b(gen_filter_6__u_filter_diff_ctr_q[3]),
    .c(n2740),
    .out0(gen_filter_6__u_filter_diff_ctr_d[3]));
 b15and003al1n04x5 U3398 (.a(gen_filter_28__u_filter_diff_ctr_q[0]),
    .b(gen_filter_28__u_filter_diff_ctr_q[1]),
    .c(net2420),
    .o(n2739));
 b15xor002al1n16x5 U3399 (.a(gen_filter_28__u_filter_filter_synced),
    .b(gen_filter_28__u_filter_filter_q),
    .out0(n2799));
 b15oab012al1n02x5 U3400 (.a(n2799),
    .b(net2461),
    .c(n2739),
    .out0(gen_filter_28__u_filter_diff_ctr_d[3]));
 b15and003aq1n04x5 U3401 (.a(gen_filter_21__u_filter_diff_ctr_q[0]),
    .b(gen_filter_21__u_filter_diff_ctr_q[1]),
    .c(gen_filter_21__u_filter_diff_ctr_q[2]),
    .o(n2738));
 b15xor002as1n16x5 U3402 (.a(gen_filter_21__u_filter_filter_synced),
    .b(gen_filter_21__u_filter_filter_q),
    .out0(n2804));
 b15oab012ar1n02x5 U3403 (.a(n2804),
    .b(gen_filter_21__u_filter_diff_ctr_q[3]),
    .c(n2738),
    .out0(gen_filter_21__u_filter_diff_ctr_d[3]));
 b15and003aq1n04x5 U3404 (.a(net2395),
    .b(gen_filter_13__u_filter_diff_ctr_q[0]),
    .c(gen_filter_13__u_filter_diff_ctr_q[1]),
    .o(n2762));
 b15xor002ah1n08x5 U3405 (.a(gen_filter_13__u_filter_filter_synced),
    .b(net2324),
    .out0(n2932));
 b15oab012al1n02x5 U3406 (.a(n2932),
    .b(gen_filter_13__u_filter_diff_ctr_q[3]),
    .c(n2762),
    .out0(gen_filter_13__u_filter_diff_ctr_d[3]));
 b15and003an1n04x5 U3407 (.a(net2318),
    .b(gen_filter_25__u_filter_diff_ctr_q[0]),
    .c(gen_filter_25__u_filter_diff_ctr_q[1]),
    .o(n2766));
 b15xor002an1n12x5 U3408 (.a(gen_filter_25__u_filter_filter_synced),
    .b(net2372),
    .out0(n2926));
 b15oab012ar1n02x5 U3409 (.a(n2926),
    .b(net2454),
    .c(n2766),
    .out0(gen_filter_25__u_filter_diff_ctr_d[3]));
 b15inv020ah1n12x5 U3410 (.a(gen_filter_20__u_filter_filter_synced),
    .o1(n3634));
 b15xor002as1n16x5 U3411 (.a(net2359),
    .b(n3634),
    .out0(n2781));
 b15inv040aq1n03x5 U3412 (.a(n2781),
    .o1(n2749));
 b15inv000al1n02x5 U3413 (.a(gen_filter_20__u_filter_diff_ctr_q[0]),
    .o1(n2699));
 b15aoi013al1n02x5 U3414 (.a(n2699),
    .b(gen_filter_20__u_filter_diff_ctr_q[3]),
    .c(gen_filter_20__u_filter_diff_ctr_q[1]),
    .d(gen_filter_20__u_filter_diff_ctr_q[2]),
    .o1(n2700));
 b15norp02ar1n02x5 U3415 (.a(n2749),
    .b(n2700),
    .o1(gen_filter_20__u_filter_diff_ctr_d[0]));
 b15inv000aq1n08x5 U3416 (.a(gen_filter_7__u_filter_filter_synced),
    .o1(n3568));
 b15xor002an1n16x5 U3417 (.a(gen_filter_7__u_filter_filter_q),
    .b(n3568),
    .out0(n2783));
 b15inv020ar1n06x5 U3418 (.a(n2783),
    .o1(n2754));
 b15inv000al1n02x5 U3419 (.a(gen_filter_7__u_filter_diff_ctr_q[0]),
    .o1(n2701));
 b15aoi013aq1n03x5 U3420 (.a(n2701),
    .b(net2478),
    .c(gen_filter_7__u_filter_diff_ctr_q[1]),
    .d(gen_filter_7__u_filter_diff_ctr_q[2]),
    .o1(n2702));
 b15nor002al1n02x5 U3421 (.a(n2754),
    .b(n2702),
    .o1(gen_filter_7__u_filter_diff_ctr_d[0]));
 b15and003aq1n04x5 U3422 (.a(net687),
    .b(gen_filter_14__u_filter_diff_ctr_q[0]),
    .c(gen_filter_14__u_filter_diff_ctr_q[1]),
    .o(n2964));
 b15inv000as1n12x5 U3423 (.a(gen_filter_14__u_filter_filter_synced),
    .o1(n3526));
 b15xor002as1n12x5 U3424 (.a(gen_filter_14__u_filter_filter_q),
    .b(n3526),
    .out0(n2963));
 b15inv000ah1n03x5 U3425 (.a(n2963),
    .o1(n2967));
 b15oab012an1n03x5 U3426 (.a(n2967),
    .b(net2442),
    .c(n2964),
    .out0(gen_filter_14__u_filter_diff_ctr_d[3]));
 b15and003ar1n03x5 U3427 (.a(gen_filter_8__u_filter_diff_ctr_q[2]),
    .b(gen_filter_8__u_filter_diff_ctr_q[0]),
    .c(gen_filter_8__u_filter_diff_ctr_q[1]),
    .o(n2958));
 b15inv020as1n10x5 U3428 (.a(net2216),
    .o1(n3492));
 b15qgbxo2an1n10x5 U3429 (.a(net2298),
    .b(n3492),
    .out0(n2957));
 b15inv040al1n02x5 U3430 (.a(n2957),
    .o1(n2961));
 b15oab012ar1n02x5 U3431 (.a(n2961),
    .b(net2326),
    .c(n2958),
    .out0(gen_filter_8__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3432 (.a(net2257),
    .o1(n2703));
 b15inv000aq1n06x5 U3433 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .o1(n2813));
 b15norp03aq1n08x5 U3434 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .c(n2813),
    .o1(n2980));
 b15inv040ah1n05x5 U3435 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .o1(n2814));
 b15nor003as1n06x5 U3436 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .c(n2814),
    .o1(n2979));
 b15oabi12aq1n02x5 U3437 (.a(n2979),
    .b(n2703),
    .c(n2980),
    .out0(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_n3));
 b15inv000al1n02x5 U3438 (.a(gen_filter_20__u_filter_diff_ctr_q[3]),
    .o1(n2745));
 b15nandp3as1n03x5 U3439 (.a(gen_filter_20__u_filter_diff_ctr_q[0]),
    .b(gen_filter_20__u_filter_diff_ctr_q[1]),
    .c(gen_filter_20__u_filter_diff_ctr_q[2]),
    .o1(n4049));
 b15aoi012an1n02x5 U3440 (.a(n2749),
    .b(n2745),
    .c(n4049),
    .o1(gen_filter_20__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3441 (.a(net2560),
    .o1(n2750));
 b15nandp3al1n04x5 U3442 (.a(gen_filter_7__u_filter_diff_ctr_q[0]),
    .b(gen_filter_7__u_filter_diff_ctr_q[1]),
    .c(gen_filter_7__u_filter_diff_ctr_q[2]),
    .o1(n4043));
 b15aoi012ar1n02x5 U3443 (.a(n2754),
    .b(n2750),
    .c(n4043),
    .o1(gen_filter_7__u_filter_diff_ctr_d[3]));
 b15inv020aq1n08x5 U3444 (.a(net2311),
    .o1(n2906));
 b15nandp3ar1n12x5 U3445 (.o1(n2904),
    .a(gen_filter_2__u_filter_diff_ctr_q[0]),
    .b(gen_filter_2__u_filter_diff_ctr_q[1]),
    .c(net2383));
 b15xor002aq1n16x5 U3446 (.a(gen_filter_2__u_filter_filter_synced),
    .b(net2329),
    .out0(n2903));
 b15aoi012ar1n02x5 U3447 (.a(n2903),
    .b(n2906),
    .c(n2904),
    .o1(gen_filter_2__u_filter_diff_ctr_d[3]));
 b15inv020as1n08x5 U3448 (.a(net2152),
    .o1(n2918));
 b15nandp3as1n08x5 U3449 (.a(gen_filter_15__u_filter_diff_ctr_q[0]),
    .b(net2202),
    .c(gen_filter_15__u_filter_diff_ctr_q[2]),
    .o1(n2916));
 b15xor002as1n08x5 U3450 (.a(gen_filter_15__u_filter_filter_synced),
    .b(net2180),
    .out0(n2915));
 b15aoi012an1n02x5 U3451 (.a(n2915),
    .b(n2918),
    .c(n2916),
    .o1(gen_filter_15__u_filter_diff_ctr_d[3]));
 b15inv040ah1n08x5 U3452 (.a(net2338),
    .o1(n2876));
 b15nand03as1n12x5 U3453 (.a(gen_filter_3__u_filter_diff_ctr_q[0]),
    .b(gen_filter_3__u_filter_diff_ctr_q[1]),
    .c(gen_filter_3__u_filter_diff_ctr_q[2]),
    .o1(n2874));
 b15xor002as1n16x5 U3454 (.a(net682),
    .b(gen_filter_3__u_filter_filter_q),
    .out0(n2873));
 b15aoi012ar1n02x5 U3455 (.a(n2873),
    .b(n2876),
    .c(n2874),
    .o1(gen_filter_3__u_filter_diff_ctr_d[3]));
 b15inv000al1n10x5 U3456 (.a(net2177),
    .o1(n2888));
 b15nandp3an1n12x5 U3457 (.o1(n2886),
    .a(gen_filter_23__u_filter_diff_ctr_q[0]),
    .b(gen_filter_23__u_filter_diff_ctr_q[1]),
    .c(gen_filter_23__u_filter_diff_ctr_q[2]));
 b15xor002aq1n12x5 U3458 (.a(gen_filter_23__u_filter_filter_synced),
    .b(net2161),
    .out0(n2885));
 b15aoi012an1n02x5 U3459 (.a(n2885),
    .b(n2888),
    .c(n2886),
    .o1(gen_filter_23__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3460 (.a(gen_filter_28__u_filter_diff_ctr_q[3]),
    .o1(n2705));
 b15aoi012ar1n02x5 U3461 (.a(net2420),
    .b(gen_filter_28__u_filter_diff_ctr_q[1]),
    .c(gen_filter_28__u_filter_diff_ctr_q[0]),
    .o1(n2704));
 b15aoi112an1n02x5 U3462 (.a(n2799),
    .b(n2704),
    .c(n2739),
    .d(n2705),
    .o1(gen_filter_28__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3463 (.a(gen_filter_21__u_filter_diff_ctr_q[3]),
    .o1(n2707));
 b15aoi012ar1n04x5 U3464 (.a(gen_filter_21__u_filter_diff_ctr_q[2]),
    .b(gen_filter_21__u_filter_diff_ctr_q[1]),
    .c(gen_filter_21__u_filter_diff_ctr_q[0]),
    .o1(n2706));
 b15aoi112al1n04x5 U3465 (.a(n2804),
    .b(n2706),
    .c(n2738),
    .d(n2707),
    .o1(gen_filter_21__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3466 (.a(gen_filter_6__u_filter_diff_ctr_q[3]),
    .o1(n2709));
 b15aoi012ar1n02x5 U3467 (.a(net2354),
    .b(gen_filter_6__u_filter_diff_ctr_q[1]),
    .c(gen_filter_6__u_filter_diff_ctr_q[0]),
    .o1(n2708));
 b15aoi112an1n02x5 U3468 (.a(n2794),
    .b(net2355),
    .c(n2740),
    .d(n2709),
    .o1(gen_filter_6__u_filter_diff_ctr_d[2]));
 b15inv040as1n06x5 U3469 (.a(net2333),
    .o1(n2894));
 b15nandp3ah1n08x5 U3470 (.a(gen_filter_16__u_filter_diff_ctr_q[0]),
    .b(net2346),
    .c(gen_filter_16__u_filter_diff_ctr_q[2]),
    .o1(n2892));
 b15xor002as1n08x5 U3471 (.a(gen_filter_16__u_filter_filter_synced),
    .b(net2321),
    .out0(n2891));
 b15aoi012al1n02x5 U3472 (.a(n2891),
    .b(n2894),
    .c(n2892),
    .o1(gen_filter_16__u_filter_diff_ctr_d[3]));
 b15inv020as1n08x5 U3473 (.a(net2155),
    .o1(n2882));
 b15nand03ar1n16x5 U3474 (.a(gen_filter_17__u_filter_diff_ctr_q[0]),
    .b(gen_filter_17__u_filter_diff_ctr_q[1]),
    .c(gen_filter_17__u_filter_diff_ctr_q[2]),
    .o1(n2880));
 b15xor002ah1n08x5 U3475 (.a(gen_filter_17__u_filter_filter_synced),
    .b(net2121),
    .out0(n2879));
 b15aoi012an1n02x5 U3476 (.a(n2879),
    .b(n2882),
    .c(n2880),
    .o1(gen_filter_17__u_filter_diff_ctr_d[3]));
 b15inv020aq1n10x5 U3477 (.a(net2374),
    .o1(n2924));
 b15nand03ah1n12x5 U3478 (.a(gen_filter_27__u_filter_diff_ctr_q[0]),
    .b(gen_filter_27__u_filter_diff_ctr_q[1]),
    .c(net2384),
    .o1(n2922));
 b15xor002an1n12x5 U3479 (.a(gen_filter_27__u_filter_filter_synced),
    .b(net2378),
    .out0(n2921));
 b15aoi012ar1n02x5 U3480 (.a(n2921),
    .b(n2924),
    .c(n2922),
    .o1(gen_filter_27__u_filter_diff_ctr_d[3]));
 b15inv000an1n08x5 U3481 (.a(net2288),
    .o1(n2912));
 b15nandp3as1n08x5 U3482 (.a(gen_filter_31__u_filter_diff_ctr_q[0]),
    .b(gen_filter_31__u_filter_diff_ctr_q[1]),
    .c(gen_filter_31__u_filter_diff_ctr_q[2]),
    .o1(n2910));
 b15xor002as1n08x5 U3483 (.a(gen_filter_31__u_filter_filter_synced),
    .b(net2286),
    .out0(n2909));
 b15aoi012ar1n02x5 U3484 (.a(n2909),
    .b(n2912),
    .c(n2910),
    .o1(gen_filter_31__u_filter_diff_ctr_d[3]));
 b15inv020aq1n12x5 U3485 (.a(net2410),
    .o1(n2900));
 b15nand03aq1n12x5 U3486 (.a(gen_filter_5__u_filter_diff_ctr_q[0]),
    .b(gen_filter_5__u_filter_diff_ctr_q[1]),
    .c(gen_filter_5__u_filter_diff_ctr_q[2]),
    .o1(n2898));
 b15xor002al1n16x5 U3487 (.a(net680),
    .b(net2433),
    .out0(n2897));
 b15aoi012aq1n02x5 U3488 (.a(n2897),
    .b(n2900),
    .c(n2898),
    .o1(gen_filter_5__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3489 (.a(gen_filter_24__u_filter_diff_ctr_q[3]),
    .o1(n2711));
 b15aoi012ar1n02x5 U3490 (.a(net2260),
    .b(gen_filter_24__u_filter_diff_ctr_q[1]),
    .c(gen_filter_24__u_filter_diff_ctr_q[0]),
    .o1(n2710));
 b15aoi112aq1n02x5 U3491 (.a(n2810),
    .b(n2710),
    .c(net2261),
    .d(n2711),
    .o1(gen_filter_24__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3492 (.a(n2880),
    .o1(n2713));
 b15aoi012ar1n02x5 U3493 (.a(gen_filter_17__u_filter_diff_ctr_q[2]),
    .b(gen_filter_17__u_filter_diff_ctr_q[1]),
    .c(gen_filter_17__u_filter_diff_ctr_q[0]),
    .o1(n2712));
 b15aoi112ar1n03x5 U3494 (.a(n2712),
    .b(net2122),
    .c(n2713),
    .d(n2882),
    .o1(gen_filter_17__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3495 (.a(n2910),
    .o1(n2715));
 b15aoi012ar1n02x5 U3496 (.a(gen_filter_31__u_filter_diff_ctr_q[2]),
    .b(gen_filter_31__u_filter_diff_ctr_q[1]),
    .c(gen_filter_31__u_filter_diff_ctr_q[0]),
    .o1(n2714));
 b15aoi112al1n02x5 U3497 (.a(n2714),
    .b(n2909),
    .c(n2715),
    .d(n2912),
    .o1(gen_filter_31__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3498 (.a(n2892),
    .o1(n2717));
 b15aoi012aq1n02x5 U3499 (.a(gen_filter_16__u_filter_diff_ctr_q[2]),
    .b(net2346),
    .c(gen_filter_16__u_filter_diff_ctr_q[0]),
    .o1(n2716));
 b15aoi112an1n02x5 U3500 (.a(n2716),
    .b(n2891),
    .c(n2717),
    .d(n2894),
    .o1(gen_filter_16__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3501 (.a(n2898),
    .o1(n2719));
 b15aoi012ar1n02x5 U3502 (.a(gen_filter_5__u_filter_diff_ctr_q[2]),
    .b(gen_filter_5__u_filter_diff_ctr_q[1]),
    .c(gen_filter_5__u_filter_diff_ctr_q[0]),
    .o1(n2718));
 b15aoi112as1n02x5 U3503 (.a(n2718),
    .b(n2897),
    .c(n2719),
    .d(n2900),
    .o1(gen_filter_5__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3504 (.a(n2886),
    .o1(n2721));
 b15aoi012ar1n02x5 U3505 (.a(gen_filter_23__u_filter_diff_ctr_q[2]),
    .b(gen_filter_23__u_filter_diff_ctr_q[1]),
    .c(gen_filter_23__u_filter_diff_ctr_q[0]),
    .o1(n2720));
 b15aoi112aq1n02x5 U3506 (.a(n2720),
    .b(net2162),
    .c(n2721),
    .d(n2888),
    .o1(gen_filter_23__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3507 (.a(n2874),
    .o1(n2723));
 b15aoi012al1n02x5 U3508 (.a(gen_filter_3__u_filter_diff_ctr_q[2]),
    .b(gen_filter_3__u_filter_diff_ctr_q[1]),
    .c(gen_filter_3__u_filter_diff_ctr_q[0]),
    .o1(n2722));
 b15aoi112ar1n02x5 U3509 (.a(n2722),
    .b(n2873),
    .c(n2723),
    .d(n2876),
    .o1(gen_filter_3__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3510 (.a(n2922),
    .o1(n2725));
 b15aoi012al1n02x5 U3511 (.a(net2382),
    .b(gen_filter_27__u_filter_diff_ctr_q[1]),
    .c(gen_filter_27__u_filter_diff_ctr_q[0]),
    .o1(n2724));
 b15aoi112ar1n04x5 U3512 (.a(n2724),
    .b(n2921),
    .c(n2725),
    .d(n2924),
    .o1(gen_filter_27__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3513 (.a(n2916),
    .o1(n2727));
 b15aoi012ar1n02x5 U3514 (.a(gen_filter_15__u_filter_diff_ctr_q[2]),
    .b(gen_filter_15__u_filter_diff_ctr_q[1]),
    .c(gen_filter_15__u_filter_diff_ctr_q[0]),
    .o1(n2726));
 b15aoi112al1n02x5 U3515 (.a(n2726),
    .b(net2181),
    .c(n2727),
    .d(n2918),
    .o1(gen_filter_15__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3516 (.a(n2904),
    .o1(n2729));
 b15aoi012ar1n02x5 U3517 (.a(net2368),
    .b(gen_filter_2__u_filter_diff_ctr_q[1]),
    .c(gen_filter_2__u_filter_diff_ctr_q[0]),
    .o1(n2728));
 b15aoi112ar1n02x5 U3518 (.a(n2728),
    .b(n2903),
    .c(n2729),
    .d(n2906),
    .o1(gen_filter_2__u_filter_diff_ctr_d[2]));
 b15nand02ar1n02x5 U3519 (.a(gen_filter_19__u_filter_diff_ctr_q[3]),
    .b(net2306),
    .o1(n2731));
 b15norp02ar1n02x5 U3520 (.a(gen_filter_19__u_filter_diff_ctr_q[1]),
    .b(gen_filter_19__u_filter_diff_ctr_q[0]),
    .o1(n2730));
 b15aoi112ar1n02x5 U3521 (.a(n2730),
    .b(n2785),
    .c(n2732),
    .d(n2731),
    .o1(gen_filter_19__u_filter_diff_ctr_d[1]));
 b15and003al1n04x5 U3522 (.a(net2308),
    .b(gen_filter_18__u_filter_diff_ctr_q[0]),
    .c(gen_filter_18__u_filter_diff_ctr_q[1]),
    .o(n2946));
 b15inv040aq1n08x5 U3523 (.a(gen_filter_18__u_filter_filter_synced),
    .o1(n3556));
 b15xor002as1n08x5 U3524 (.a(gen_filter_18__u_filter_filter_q),
    .b(n3556),
    .out0(n2948));
 b15inv040ah1n03x5 U3525 (.a(n2948),
    .o1(n2947));
 b15oab012ah1n03x5 U3526 (.a(n2947),
    .b(net2417),
    .c(n2946),
    .out0(gen_filter_18__u_filter_diff_ctr_d[3]));
 b15and003ah1n03x5 U3527 (.a(net2405),
    .b(gen_filter_11__u_filter_diff_ctr_q[0]),
    .c(gen_filter_11__u_filter_diff_ctr_q[1]),
    .o(n2938));
 b15inv000al1n20x5 U3528 (.a(gen_filter_11__u_filter_filter_synced),
    .o1(n3506));
 b15xor002ar1n16x5 U3529 (.a(gen_filter_11__u_filter_filter_q),
    .b(n3506),
    .out0(n2940));
 b15inv000aq1n06x5 U3530 (.a(n2940),
    .o1(n2939));
 b15oab012ah1n02x5 U3531 (.a(n2939),
    .b(net2348),
    .c(n2938),
    .out0(gen_filter_11__u_filter_diff_ctr_d[3]));
 b15nand02ar1n02x5 U3532 (.a(gen_filter_26__u_filter_diff_ctr_q[3]),
    .b(gen_filter_26__u_filter_diff_ctr_q[2]),
    .o1(n2734));
 b15norp02ar1n02x5 U3533 (.a(net2469),
    .b(gen_filter_26__u_filter_diff_ctr_q[1]),
    .o1(n2733));
 b15aoi112ar1n02x5 U3534 (.a(n2737),
    .b(n2733),
    .c(n2735),
    .d(n2734),
    .o1(gen_filter_26__u_filter_diff_ctr_d[1]));
 b15norp02ah1n12x5 U3535 (.a(n2737),
    .b(n2736),
    .o1(eq_x_51_n25));
 b15nandp2ah1n03x5 U3536 (.a(net2473),
    .b(n2738),
    .o1(n2806));
 b15aoi012an1n02x5 U3537 (.a(n2804),
    .b(net2390),
    .c(n2806),
    .o1(gen_filter_21__u_filter_diff_ctr_d[0]));
 b15nand02aq1n04x5 U3538 (.a(net2461),
    .b(n2739),
    .o1(n2801));
 b15aoi012ah1n02x5 U3539 (.a(n2799),
    .b(net2339),
    .c(n2801),
    .o1(gen_filter_28__u_filter_diff_ctr_d[0]));
 b15nandp2ah1n03x5 U3540 (.a(gen_filter_6__u_filter_diff_ctr_q[3]),
    .b(n2740),
    .o1(n2796));
 b15aoi012as1n02x5 U3541 (.a(n2794),
    .b(gen_filter_6__u_filter_diff_ctr_q[0]),
    .c(n2796),
    .o1(gen_filter_6__u_filter_diff_ctr_d[0]));
 b15nand02aq1n06x5 U3542 (.a(net2437),
    .b(n2772),
    .o1(n2816));
 b15aoi012ar1n02x5 U3543 (.a(n2767),
    .b(net2304),
    .c(n2816),
    .o1(gen_filter_0__u_filter_diff_ctr_d[0]));
 b15nandp2as1n05x5 U3544 (.a(gen_filter_13__u_filter_diff_ctr_q[3]),
    .b(n2762),
    .o1(n2936));
 b15aoi012an1n02x5 U3545 (.a(n2932),
    .b(net2364),
    .c(n2936),
    .o1(gen_filter_13__u_filter_diff_ctr_d[0]));
 b15nandp2an1n08x5 U3546 (.a(net2436),
    .b(n2766),
    .o1(n2930));
 b15aoi012ar1n06x5 U3547 (.a(n2926),
    .b(gen_filter_25__u_filter_diff_ctr_q[0]),
    .c(n2930),
    .o1(gen_filter_25__u_filter_diff_ctr_d[0]));
 b15inv000al1n02x5 U3548 (.a(net2450),
    .o1(n2831));
 b15nandp3ah1n02x5 U3549 (.a(gen_filter_30__u_filter_diff_ctr_q[0]),
    .b(gen_filter_30__u_filter_diff_ctr_q[1]),
    .c(net2414),
    .o1(n2773));
 b15inv040ah1n12x5 U3550 (.a(gen_filter_30__u_filter_filter_synced),
    .o1(n3483));
 b15xor002an1n12x5 U3551 (.a(gen_filter_30__u_filter_filter_q),
    .b(n3483),
    .out0(n2826));
 b15inv000as1n02x5 U3552 (.a(n2826),
    .o1(n2829));
 b15aoi012ar1n02x5 U3553 (.a(n2829),
    .b(n2831),
    .c(n2773),
    .o1(gen_filter_30__u_filter_diff_ctr_d[3]));
 b15inv000an1n02x5 U3554 (.a(gen_filter_12__u_filter_diff_ctr_q[3]),
    .o1(n2853));
 b15nand03an1n06x5 U3555 (.a(gen_filter_12__u_filter_diff_ctr_q[0]),
    .b(gen_filter_12__u_filter_diff_ctr_q[1]),
    .c(gen_filter_12__u_filter_diff_ctr_q[2]),
    .o1(n2774));
 b15inv020ah1n12x5 U3556 (.a(gen_filter_12__u_filter_filter_synced),
    .o1(n3628));
 b15xor002as1n06x5 U3557 (.a(net2360),
    .b(n3628),
    .out0(n2848));
 b15inv000as1n03x5 U3558 (.a(n2848),
    .o1(n2851));
 b15aoi012ar1n04x5 U3559 (.a(n2851),
    .b(n2853),
    .c(net2386),
    .o1(gen_filter_12__u_filter_diff_ctr_d[3]));
 b15inv040al1n02x5 U3560 (.a(net2282),
    .o1(n2838));
 b15nandp3ar1n04x5 U3561 (.a(gen_filter_22__u_filter_diff_ctr_q[0]),
    .b(gen_filter_22__u_filter_diff_ctr_q[1]),
    .c(gen_filter_22__u_filter_diff_ctr_q[2]),
    .o1(n2775));
 b15inv040al1n12x5 U3562 (.a(gen_filter_22__u_filter_filter_synced),
    .o1(n3654));
 b15xor002as1n16x5 U3563 (.a(gen_filter_22__u_filter_filter_q),
    .b(n3654),
    .out0(n2833));
 b15inv000as1n03x5 U3564 (.a(n2833),
    .o1(n2836));
 b15aoi012aq1n02x5 U3565 (.a(n2836),
    .b(n2838),
    .c(n2775),
    .o1(gen_filter_22__u_filter_diff_ctr_d[3]));
 b15inv040al1n02x5 U3566 (.a(gen_filter_4__u_filter_diff_ctr_q[3]),
    .o1(n2867));
 b15nand03an1n06x5 U3567 (.a(net2271),
    .b(gen_filter_4__u_filter_diff_ctr_q[1]),
    .c(gen_filter_4__u_filter_diff_ctr_q[2]),
    .o1(n2776));
 b15inv000as1n10x5 U3568 (.a(gen_filter_4__u_filter_filter_synced),
    .o1(n3598));
 b15xor002an1n12x5 U3569 (.a(net2392),
    .b(n3598),
    .out0(n2862));
 b15inv040ar1n03x5 U3570 (.a(n2862),
    .o1(n2865));
 b15aoi012al1n04x5 U3571 (.a(n2865),
    .b(n2867),
    .c(n2776),
    .o1(gen_filter_4__u_filter_diff_ctr_d[3]));
 b15inv040al1n02x5 U3572 (.a(net2470),
    .o1(n2860));
 b15nand03an1n06x5 U3573 (.a(gen_filter_1__u_filter_diff_ctr_q[0]),
    .b(gen_filter_1__u_filter_diff_ctr_q[1]),
    .c(net2369),
    .o1(n2777));
 b15inv000ar1n20x5 U3574 (.a(gen_filter_1__u_filter_filter_synced),
    .o1(n3592));
 b15xor002an1n12x5 U3575 (.a(gen_filter_1__u_filter_filter_q),
    .b(n3592),
    .out0(n2855));
 b15inv020al1n05x5 U3576 (.a(n2855),
    .o1(n2858));
 b15aoi012ar1n04x5 U3577 (.a(n2858),
    .b(n2860),
    .c(n2777),
    .o1(gen_filter_1__u_filter_diff_ctr_d[3]));
 b15and003as1n02x5 U3578 (.a(net2342),
    .b(net2336),
    .c(gen_filter_29__u_filter_diff_ctr_q[1]),
    .o(n2819));
 b15inv040ah1n06x5 U3579 (.a(gen_filter_29__u_filter_filter_synced),
    .o1(n3660));
 b15xor002an1n12x5 U3580 (.a(gen_filter_29__u_filter_filter_q),
    .b(n3660),
    .out0(n2818));
 b15inv040al1n03x5 U3581 (.a(n2818),
    .o1(n2822));
 b15oab012ar1n02x5 U3582 (.a(n2822),
    .b(net2452),
    .c(n2819),
    .out0(gen_filter_29__u_filter_diff_ctr_d[3]));
 b15and003aq1n04x5 U3583 (.a(gen_filter_10__u_filter_diff_ctr_q[2]),
    .b(gen_filter_10__u_filter_diff_ctr_q[0]),
    .c(gen_filter_10__u_filter_diff_ctr_q[1]),
    .o(n2841));
 b15inv020as1n10x5 U3584 (.a(net2424),
    .o1(n3520));
 b15xor002aq1n12x5 U3585 (.a(net2247),
    .b(n3520),
    .out0(n2840));
 b15inv020aq1n05x5 U3586 (.a(n2840),
    .o1(n2844));
 b15oab012al1n02x5 U3587 (.a(n2844),
    .b(net2231),
    .c(n2841),
    .out0(gen_filter_10__u_filter_diff_ctr_d[3]));
 b15nand02ar1n02x5 U3588 (.a(gen_filter_24__u_filter_diff_ctr_q[0]),
    .b(gen_filter_24__u_filter_diff_ctr_q[1]),
    .o1(n2743));
 b15nandp2an1n03x5 U3589 (.a(gen_filter_24__u_filter_diff_ctr_q[3]),
    .b(n2741),
    .o1(n2811));
 b15inv000al1n02x5 U3590 (.a(n2811),
    .o1(n2742));
 b15oaoi13ar1n02x5 U3591 (.a(n2742),
    .b(n2743),
    .c(gen_filter_24__u_filter_diff_ctr_q[0]),
    .d(gen_filter_24__u_filter_diff_ctr_q[1]),
    .o1(n2744));
 b15norp02al1n02x5 U3592 (.a(n2744),
    .b(n2810),
    .o1(gen_filter_24__u_filter_diff_ctr_d[1]));
 b15nand02ar1n02x5 U3593 (.a(gen_filter_20__u_filter_diff_ctr_q[0]),
    .b(gen_filter_20__u_filter_diff_ctr_q[1]),
    .o1(n2747));
 b15norp02an1n02x5 U3594 (.a(n2745),
    .b(n4049),
    .o1(n2746));
 b15oaoi13ar1n02x3 U3595 (.a(n2746),
    .b(n2747),
    .c(gen_filter_20__u_filter_diff_ctr_q[0]),
    .d(gen_filter_20__u_filter_diff_ctr_q[1]),
    .o1(n2748));
 b15norp02ar1n02x5 U3596 (.a(n2749),
    .b(n2748),
    .o1(gen_filter_20__u_filter_diff_ctr_d[1]));
 b15nand02ar1n02x5 U3597 (.a(gen_filter_7__u_filter_diff_ctr_q[0]),
    .b(gen_filter_7__u_filter_diff_ctr_q[1]),
    .o1(n2752));
 b15nor002ah1n02x5 U3598 (.a(n2750),
    .b(n4043),
    .o1(n2751));
 b15oaoi13ar1n02x3 U3599 (.a(n2751),
    .b(n2752),
    .c(gen_filter_7__u_filter_diff_ctr_q[0]),
    .d(gen_filter_7__u_filter_diff_ctr_q[1]),
    .o1(n2753));
 b15norp02ar1n02x5 U3600 (.a(n2754),
    .b(n2753),
    .o1(gen_filter_7__u_filter_diff_ctr_d[1]));
 b15nandp2ar1n03x5 U3601 (.a(net2567),
    .b(gen_filter_0__u_filter_diff_ctr_q[1]),
    .o1(n2768));
 b15inv000al1n02x5 U3602 (.a(n2816),
    .o1(n2755));
 b15oaoi13aq1n02x5 U3603 (.a(n2755),
    .b(n2768),
    .c(net2304),
    .d(net2345),
    .o1(n2756));
 b15norp02ar1n02x5 U3604 (.a(n2767),
    .b(n2756),
    .o1(gen_filter_0__u_filter_diff_ctr_d[1]));
 b15inv020as1n16x5 U3605 (.a(net44),
    .o1(n3347));
 b15norp02ah1n16x5 U3606 (.a(n3347),
    .b(net294),
    .o1(u_reg_u_reg_if_a_ack));
 b15inv020aq1n05x5 U3607 (.a(net1982),
    .o1(n2951));
 b15nor002ah1n04x5 U3608 (.a(net672),
    .b(n2951),
    .o1(n1432));
 b15inv000an1n32x5 U3609 (.a(net1919),
    .o1(n2953));
 b15nor002al1n06x5 U3610 (.a(net672),
    .b(n2953),
    .o1(n1429));
 b15nandp2ar1n03x5 U3611 (.a(gen_filter_9__u_filter_diff_ctr_q[0]),
    .b(gen_filter_9__u_filter_diff_ctr_q[1]),
    .o1(n2758));
 b15nandp2as1n03x5 U3612 (.a(net2279),
    .b(n2780),
    .o1(n2809));
 b15inv040ar1n02x5 U3613 (.a(n2809),
    .o1(n2757));
 b15oaoi13al1n08x5 U3614 (.a(n2757),
    .b(n2758),
    .c(gen_filter_9__u_filter_diff_ctr_q[0]),
    .d(gen_filter_9__u_filter_diff_ctr_q[1]),
    .o1(n4045));
 b15norp02ah1n02x5 U3615 (.a(n2808),
    .b(n4045),
    .o1(gen_filter_9__u_filter_diff_ctr_d[1]));
 b15inv000al1n02x5 U3616 (.a(gen_filter_13__u_filter_diff_ctr_q[2]),
    .o1(n2759));
 b15nandp2ar1n03x5 U3617 (.a(gen_filter_13__u_filter_diff_ctr_q[0]),
    .b(gen_filter_13__u_filter_diff_ctr_q[1]),
    .o1(n2931));
 b15aoi012ar1n04x5 U3618 (.a(n2932),
    .b(n2759),
    .c(n2931),
    .o1(n2760));
 b15inv000al1n02x5 U3619 (.a(n2760),
    .o1(n2761));
 b15nandp2ar1n05x5 U3620 (.a(n2760),
    .b(gen_filter_13__u_filter_diff_ctr_q[3]),
    .o1(n2935));
 b15oai012aq1n02x5 U3621 (.a(n2935),
    .b(net2396),
    .c(n2761),
    .o1(gen_filter_13__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3622 (.a(net2318),
    .o1(n2763));
 b15nand02al1n02x5 U3623 (.a(gen_filter_25__u_filter_diff_ctr_q[0]),
    .b(gen_filter_25__u_filter_diff_ctr_q[1]),
    .o1(n2925));
 b15aoi012aq1n02x5 U3624 (.a(n2926),
    .b(n2763),
    .c(n2925),
    .o1(n2764));
 b15inv000al1n02x5 U3625 (.a(n2764),
    .o1(n2765));
 b15nandp2as1n04x5 U3626 (.a(n2764),
    .b(gen_filter_25__u_filter_diff_ctr_q[3]),
    .o1(n2929));
 b15oai012as1n03x5 U3627 (.a(n2929),
    .b(net2319),
    .c(n2765),
    .o1(gen_filter_25__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3628 (.a(gen_filter_0__u_filter_diff_ctr_q[2]),
    .o1(n2769));
 b15aoi012an1n02x5 U3629 (.a(n2767),
    .b(n2769),
    .c(n2768),
    .o1(n2770));
 b15inv000al1n02x5 U3630 (.a(n2770),
    .o1(n2771));
 b15nandp2aq1n03x5 U3631 (.a(n2770),
    .b(net2437),
    .o1(n2815));
 b15oai012ar1n04x5 U3632 (.a(n2815),
    .b(net2403),
    .c(n2771),
    .o1(gen_filter_0__u_filter_diff_ctr_d[2]));
 b15nand02as1n06x5 U3633 (.a(gen_filter_18__u_filter_diff_ctr_q[3]),
    .b(n2948),
    .o1(n4046));
 b15aoi012aq1n04x5 U3634 (.a(net2308),
    .b(gen_filter_18__u_filter_diff_ctr_q[0]),
    .c(gen_filter_18__u_filter_diff_ctr_q[1]),
    .o1(n4047));
 b15oaoi13al1n02x5 U3635 (.a(n4047),
    .b(n4046),
    .c(n2947),
    .d(n2946),
    .o1(gen_filter_18__u_filter_diff_ctr_d[2]));
 b15nand02as1n03x5 U3636 (.a(net2348),
    .b(n2940),
    .o1(n2937));
 b15aoi012ah1n04x5 U3637 (.a(net2405),
    .b(gen_filter_11__u_filter_diff_ctr_q[0]),
    .c(gen_filter_11__u_filter_diff_ctr_q[1]),
    .o1(n2945));
 b15oaoi13an1n04x5 U3638 (.a(n2945),
    .b(n2937),
    .c(n2939),
    .d(n2938),
    .o1(gen_filter_11__u_filter_diff_ctr_d[2]));
 b15aoai13al1n03x5 U3639 (.a(n2826),
    .b(net2414),
    .c(gen_filter_30__u_filter_diff_ctr_q[1]),
    .d(gen_filter_30__u_filter_diff_ctr_q[0]),
    .o1(n2830));
 b15oab012ar1n02x5 U3640 (.a(n2830),
    .b(net2450),
    .c(n2773),
    .out0(gen_filter_30__u_filter_diff_ctr_d[2]));
 b15aoai13as1n03x5 U3641 (.a(n2848),
    .b(net2385),
    .c(gen_filter_12__u_filter_diff_ctr_q[1]),
    .d(gen_filter_12__u_filter_diff_ctr_q[0]),
    .o1(n2852));
 b15oab012ar1n02x5 U3642 (.a(n2852),
    .b(gen_filter_12__u_filter_diff_ctr_q[3]),
    .c(net2386),
    .out0(gen_filter_12__u_filter_diff_ctr_d[2]));
 b15aoai13al1n06x5 U3643 (.a(n2833),
    .b(gen_filter_22__u_filter_diff_ctr_q[2]),
    .c(gen_filter_22__u_filter_diff_ctr_q[1]),
    .d(gen_filter_22__u_filter_diff_ctr_q[0]),
    .o1(n2837));
 b15oab012ar1n02x5 U3644 (.a(n2837),
    .b(net2553),
    .c(n2775),
    .out0(gen_filter_22__u_filter_diff_ctr_d[2]));
 b15aoai13as1n02x5 U3645 (.a(n2862),
    .b(gen_filter_4__u_filter_diff_ctr_q[2]),
    .c(gen_filter_4__u_filter_diff_ctr_q[1]),
    .d(net2271),
    .o1(n2866));
 b15oab012an1n02x5 U3646 (.a(net2393),
    .b(gen_filter_4__u_filter_diff_ctr_q[3]),
    .c(n2776),
    .out0(gen_filter_4__u_filter_diff_ctr_d[2]));
 b15aoai13ah1n02x5 U3647 (.a(n2855),
    .b(net2369),
    .c(gen_filter_1__u_filter_diff_ctr_q[1]),
    .d(gen_filter_1__u_filter_diff_ctr_q[0]),
    .o1(n2859));
 b15oab012ar1n02x5 U3648 (.a(net2370),
    .b(gen_filter_1__u_filter_diff_ctr_q[3]),
    .c(n2777),
    .out0(gen_filter_1__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3649 (.a(net2279),
    .o1(n2779));
 b15inv000al1n02x5 U3650 (.a(n2808),
    .o1(n2778));
 b15aoai13al1n08x5 U3651 (.a(n2778),
    .b(net2358),
    .c(gen_filter_9__u_filter_diff_ctr_q[1]),
    .d(gen_filter_9__u_filter_diff_ctr_q[0]),
    .o1(n4044));
 b15aoi012ah1n02x5 U3652 (.a(n4044),
    .b(n2780),
    .c(n2779),
    .o1(gen_filter_9__u_filter_diff_ctr_d[2]));
 b15nandp2ah1n02x5 U3653 (.a(net2231),
    .b(n2840),
    .o1(n2845));
 b15aoi012an1n02x5 U3654 (.a(gen_filter_10__u_filter_diff_ctr_q[2]),
    .b(gen_filter_10__u_filter_diff_ctr_q[0]),
    .c(gen_filter_10__u_filter_diff_ctr_q[1]),
    .o1(n2846));
 b15oaoi13as1n02x5 U3655 (.a(n2846),
    .b(net2232),
    .c(n2844),
    .d(n2841),
    .o1(gen_filter_10__u_filter_diff_ctr_d[2]));
 b15nandp2ar1n02x5 U3656 (.a(gen_filter_29__u_filter_diff_ctr_q[3]),
    .b(n2818),
    .o1(n2823));
 b15aoi012al1n02x5 U3657 (.a(net2342),
    .b(net2336),
    .c(gen_filter_29__u_filter_diff_ctr_q[1]),
    .o1(n2824));
 b15oaoi13an1n02x5 U3658 (.a(net2343),
    .b(n2823),
    .c(n2822),
    .d(n2819),
    .o1(gen_filter_29__u_filter_diff_ctr_d[2]));
 b15aoai13ar1n08x5 U3659 (.a(n2781),
    .b(gen_filter_20__u_filter_diff_ctr_q[2]),
    .c(gen_filter_20__u_filter_diff_ctr_q[1]),
    .d(gen_filter_20__u_filter_diff_ctr_q[0]),
    .o1(n4048));
 b15nandp3al1n04x5 U3660 (.a(gen_filter_20__u_filter_diff_ctr_q[2]),
    .b(gen_filter_20__u_filter_diff_ctr_q[1]),
    .c(gen_filter_20__u_filter_diff_ctr_q[3]),
    .o1(n2782));
 b15nor002aq1n08x5 U3661 (.a(n4048),
    .b(n2782),
    .o1(eq_x_81_n25));
 b15aoai13an1n06x5 U3662 (.a(n2783),
    .b(gen_filter_7__u_filter_diff_ctr_q[2]),
    .c(gen_filter_7__u_filter_diff_ctr_q[1]),
    .d(gen_filter_7__u_filter_diff_ctr_q[0]),
    .o1(n4042));
 b15nand03ar1n06x5 U3663 (.a(gen_filter_7__u_filter_diff_ctr_q[2]),
    .b(gen_filter_7__u_filter_diff_ctr_q[1]),
    .c(net2569),
    .o1(n2784));
 b15nor002ah1n06x5 U3664 (.a(n4042),
    .b(n2784),
    .o1(eq_x_146_n25));
 b15inv000al1n02x5 U3665 (.a(gen_filter_19__u_filter_diff_ctr_q[3]),
    .o1(n2787));
 b15aoi012aq1n02x5 U3666 (.a(n2785),
    .b(n2787),
    .c(net2295),
    .o1(gen_filter_19__u_filter_diff_ctr_d[3]));
 b15nonb02an1n02x5 U3667 (.a(gen_filter_19__u_filter_diff_ctr_d[3]),
    .b(n2788),
    .out0(eq_x_86_n25));
 b15inv000ah1n03x5 U3668 (.a(net1976),
    .o1(n2952));
 b15aoi022ah1n02x5 U3669 (.a(net1976),
    .b(net1950),
    .c(n2951),
    .d(n2952),
    .o1(net239));
 b15nor002as1n04x5 U3670 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd),
    .o1(n2792));
 b15inv040ar1n02x5 U3671 (.a(n2792),
    .o1(n2790));
 b15nand03aq1n02x5 U3672 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq),
    .c(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq),
    .o1(n2789));
 b15oai013ar1n08x5 U3673 (.a(n2789),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq),
    .c(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq),
    .d(n2790),
    .o1(n2791));
 b15norp03al1n08x5 U3674 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[0]),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .c(n2791),
    .o1(n2972));
 b15aoi012ah1n12x5 U3675 (.a(n2792),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd),
    .c(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .o1(n2973));
 b15nonb02an1n02x5 U3676 (.a(n2972),
    .b(n2973),
    .out0(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[0]));
 b15nand02ar1n02x5 U3677 (.a(gen_filter_6__u_filter_diff_ctr_q[0]),
    .b(net2570),
    .o1(n2793));
 b15oai012ah1n02x5 U3678 (.a(n2793),
    .b(gen_filter_6__u_filter_diff_ctr_q[0]),
    .c(net2327),
    .o1(n2795));
 b15aoi012al1n04x5 U3679 (.a(n2794),
    .b(n2796),
    .c(n2795),
    .o1(gen_filter_6__u_filter_diff_ctr_d[1]));
 b15nandp3al1n03x5 U3680 (.a(net2456),
    .b(net2354),
    .c(gen_filter_6__u_filter_diff_ctr_q[3]),
    .o1(n2797));
 b15nonb02ah1n04x5 U3681 (.a(gen_filter_6__u_filter_diff_ctr_d[1]),
    .b(n2797),
    .out0(eq_x_151_n25));
 b15nand02ar1n02x5 U3682 (.a(gen_filter_28__u_filter_diff_ctr_q[0]),
    .b(gen_filter_28__u_filter_diff_ctr_q[1]),
    .o1(n2798));
 b15oai012an1n03x5 U3683 (.a(n2798),
    .b(gen_filter_28__u_filter_diff_ctr_q[0]),
    .c(gen_filter_28__u_filter_diff_ctr_q[1]),
    .o1(n2800));
 b15aoi012al1n04x5 U3684 (.a(n2799),
    .b(n2801),
    .c(n2800),
    .o1(gen_filter_28__u_filter_diff_ctr_d[1]));
 b15nand03al1n04x5 U3685 (.a(gen_filter_28__u_filter_diff_ctr_q[1]),
    .b(net2562),
    .c(gen_filter_28__u_filter_diff_ctr_q[3]),
    .o1(n2802));
 b15nonb02al1n04x5 U3686 (.a(gen_filter_28__u_filter_diff_ctr_d[1]),
    .b(n2802),
    .out0(eq_x_41_n25));
 b15nand02ar1n02x5 U3687 (.a(gen_filter_21__u_filter_diff_ctr_q[0]),
    .b(gen_filter_21__u_filter_diff_ctr_q[1]),
    .o1(n2803));
 b15oai012as1n02x5 U3688 (.a(n2803),
    .b(gen_filter_21__u_filter_diff_ctr_q[0]),
    .c(gen_filter_21__u_filter_diff_ctr_q[1]),
    .o1(n2805));
 b15aoi012aq1n06x5 U3689 (.a(n2804),
    .b(n2806),
    .c(n2805),
    .o1(gen_filter_21__u_filter_diff_ctr_d[1]));
 b15nand03ar1n08x5 U3690 (.a(gen_filter_21__u_filter_diff_ctr_q[1]),
    .b(gen_filter_21__u_filter_diff_ctr_q[2]),
    .c(gen_filter_21__u_filter_diff_ctr_q[3]),
    .o1(n2807));
 b15nonb02an1n12x5 U3691 (.a(gen_filter_21__u_filter_diff_ctr_d[1]),
    .b(n2807),
    .out0(eq_x_76_n25));
 b15aoi012ah1n06x5 U3692 (.a(n2808),
    .b(gen_filter_9__u_filter_diff_ctr_q[0]),
    .c(n2809),
    .o1(gen_filter_9__u_filter_diff_ctr_d[0]));
 b15aoi012as1n02x5 U3693 (.a(n2810),
    .b(gen_filter_24__u_filter_diff_ctr_q[0]),
    .c(n2811),
    .o1(gen_filter_24__u_filter_diff_ctr_d[0]));
 b15nandp3an1n03x5 U3694 (.a(gen_filter_24__u_filter_diff_ctr_q[1]),
    .b(net2568),
    .c(gen_filter_24__u_filter_diff_ctr_q[3]),
    .o1(n2812));
 b15nonb02al1n04x5 U3695 (.a(gen_filter_24__u_filter_diff_ctr_d[0]),
    .b(n2812),
    .out0(eq_x_61_n25));
 b15inv020ah1n08x5 U3696 (.a(u_reg_u_reg_if_a_ack),
    .o1(n3864));
 b15aob012aq1n06x5 U3697 (.a(n3864),
    .b(net294),
    .c(net38),
    .out0(u_reg_u_reg_if_N7));
 b15xor002aq1n06x5 U3698 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq),
    .b(n2813),
    .out0(n2976));
 b15qgbxo2an1n10x5 U3699 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq),
    .b(n2814),
    .out0(n2977));
 b15aoi112aq1n06x5 U3700 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .c(n2976),
    .d(n2977),
    .o1(n2975));
 b15aoi022as1n08x5 U3701 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .c(n2814),
    .d(n2813),
    .o1(n2974));
 b15nonb02ar1n02x3 U3702 (.a(n2975),
    .b(n2974),
    .out0(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[0]));
 b15inv000al1n02x5 U3703 (.a(gen_filter_0__u_filter_diff_ctr_q[1]),
    .o1(n2817));
 b15oaoi13ah1n03x5 U3704 (.a(n2815),
    .b(n2816),
    .c(net2304),
    .d(n2817),
    .o1(eq_x_181_n25));
 b15oai012al1n02x5 U3705 (.a(n2818),
    .b(gen_filter_29__u_filter_diff_ctr_q[0]),
    .c(gen_filter_29__u_filter_diff_ctr_q[1]),
    .o1(n2820));
 b15nand03al1n06x5 U3706 (.a(gen_filter_29__u_filter_diff_ctr_q[3]),
    .b(n2819),
    .c(n2818),
    .o1(n2821));
 b15aoai13al1n04x5 U3707 (.a(n2821),
    .b(n2820),
    .c(net2362),
    .d(net2336),
    .o1(gen_filter_29__u_filter_diff_ctr_d[1]));
 b15oai012ah1n04x5 U3708 (.a(n2821),
    .b(net2336),
    .c(n2822),
    .o1(gen_filter_29__u_filter_diff_ctr_d[0]));
 b15norp02ar1n02x5 U3709 (.a(n2824),
    .b(n2823),
    .o1(n2825));
 b15and003as1n03x5 U3710 (.a(n2825),
    .b(gen_filter_29__u_filter_diff_ctr_d[1]),
    .c(gen_filter_29__u_filter_diff_ctr_d[0]),
    .o(eq_x_36_n25));
 b15oai012ar1n04x5 U3711 (.a(n2826),
    .b(gen_filter_30__u_filter_diff_ctr_q[0]),
    .c(gen_filter_30__u_filter_diff_ctr_q[1]),
    .o1(n2827));
 b15nand04aq1n06x5 U3712 (.a(gen_filter_30__u_filter_diff_ctr_q[1]),
    .b(gen_filter_30__u_filter_diff_ctr_q[3]),
    .c(net2414),
    .d(n2826),
    .o1(n2828));
 b15aoai13al1n06x5 U3713 (.a(net2415),
    .b(n2827),
    .c(gen_filter_30__u_filter_diff_ctr_q[1]),
    .d(gen_filter_30__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_30__u_filter_diff_ctr_d[1]));
 b15oai012as1n04x5 U3714 (.a(n2828),
    .b(net2397),
    .c(n2829),
    .o1(gen_filter_30__u_filter_diff_ctr_d[0]));
 b15norp02ar1n02x5 U3715 (.a(n2831),
    .b(n2830),
    .o1(n2832));
 b15and003ah1n03x5 U3716 (.a(n2832),
    .b(gen_filter_30__u_filter_diff_ctr_d[1]),
    .c(gen_filter_30__u_filter_diff_ctr_d[0]),
    .o(eq_x_31_n25));
 b15oai012an1n02x5 U3717 (.a(n2833),
    .b(gen_filter_22__u_filter_diff_ctr_q[0]),
    .c(gen_filter_22__u_filter_diff_ctr_q[1]),
    .o1(n2834));
 b15nand04al1n12x5 U3718 (.a(gen_filter_22__u_filter_diff_ctr_q[1]),
    .b(net2282),
    .c(gen_filter_22__u_filter_diff_ctr_q[2]),
    .d(n2833),
    .o1(n2835));
 b15aoai13ah1n04x5 U3719 (.a(net2283),
    .b(n2834),
    .c(gen_filter_22__u_filter_diff_ctr_q[1]),
    .d(net2565),
    .o1(gen_filter_22__u_filter_diff_ctr_d[1]));
 b15oai012aq1n06x5 U3720 (.a(net2283),
    .b(net2307),
    .c(n2836),
    .o1(gen_filter_22__u_filter_diff_ctr_d[0]));
 b15norp02ah1n03x5 U3721 (.a(n2838),
    .b(n2837),
    .o1(n2839));
 b15and003as1n12x5 U3722 (.a(n2839),
    .b(gen_filter_22__u_filter_diff_ctr_d[1]),
    .c(gen_filter_22__u_filter_diff_ctr_d[0]),
    .o(eq_x_71_n25));
 b15oai012ar1n02x5 U3723 (.a(n2840),
    .b(gen_filter_10__u_filter_diff_ctr_q[0]),
    .c(gen_filter_10__u_filter_diff_ctr_q[1]),
    .o1(n2842));
 b15nand03as1n06x5 U3724 (.a(net2231),
    .b(n2841),
    .c(net2248),
    .o1(n2843));
 b15aoai13as1n03x5 U3725 (.a(net2249),
    .b(n2842),
    .c(gen_filter_10__u_filter_diff_ctr_q[1]),
    .d(gen_filter_10__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_10__u_filter_diff_ctr_d[1]));
 b15oai012al1n08x5 U3726 (.a(net2249),
    .b(net2258),
    .c(n2844),
    .o1(gen_filter_10__u_filter_diff_ctr_d[0]));
 b15norp02ar1n02x5 U3727 (.a(n2846),
    .b(n2845),
    .o1(n2847));
 b15and003al1n04x5 U3728 (.a(n2847),
    .b(gen_filter_10__u_filter_diff_ctr_d[1]),
    .c(gen_filter_10__u_filter_diff_ctr_d[0]),
    .o(eq_x_131_n25));
 b15oai012aq1n02x5 U3729 (.a(n2848),
    .b(gen_filter_12__u_filter_diff_ctr_q[0]),
    .c(gen_filter_12__u_filter_diff_ctr_q[1]),
    .o1(n2849));
 b15nand04ah1n06x5 U3730 (.a(gen_filter_12__u_filter_diff_ctr_q[1]),
    .b(net2407),
    .c(net2385),
    .d(n2848),
    .o1(n2850));
 b15aoai13as1n04x5 U3731 (.a(n2850),
    .b(n2849),
    .c(gen_filter_12__u_filter_diff_ctr_q[1]),
    .d(gen_filter_12__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_12__u_filter_diff_ctr_d[1]));
 b15oai012al1n06x5 U3732 (.a(n2850),
    .b(net2427),
    .c(n2851),
    .o1(gen_filter_12__u_filter_diff_ctr_d[0]));
 b15norp02ar1n02x5 U3733 (.a(n2853),
    .b(n2852),
    .o1(n2854));
 b15and003as1n02x5 U3734 (.a(n2854),
    .b(gen_filter_12__u_filter_diff_ctr_d[1]),
    .c(gen_filter_12__u_filter_diff_ctr_d[0]),
    .o(eq_x_121_n25));
 b15oai012al1n02x5 U3735 (.a(n2855),
    .b(gen_filter_1__u_filter_diff_ctr_q[0]),
    .c(gen_filter_1__u_filter_diff_ctr_q[1]),
    .o1(n2856));
 b15nand04ah1n06x5 U3736 (.a(gen_filter_1__u_filter_diff_ctr_q[1]),
    .b(net2412),
    .c(net2369),
    .d(n2855),
    .o1(n2857));
 b15aoai13al1n04x5 U3737 (.a(n2857),
    .b(n2856),
    .c(gen_filter_1__u_filter_diff_ctr_q[1]),
    .d(gen_filter_1__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_1__u_filter_diff_ctr_d[1]));
 b15oai012ah1n06x5 U3738 (.a(n2857),
    .b(net2387),
    .c(n2858),
    .o1(gen_filter_1__u_filter_diff_ctr_d[0]));
 b15norp02ar1n02x5 U3739 (.a(n2860),
    .b(n2859),
    .o1(n2861));
 b15and003aq1n03x5 U3740 (.a(n2861),
    .b(gen_filter_1__u_filter_diff_ctr_d[1]),
    .c(gen_filter_1__u_filter_diff_ctr_d[0]),
    .o(eq_x_176_n25));
 b15oai012ar1n03x5 U3741 (.a(n2862),
    .b(net2271),
    .c(gen_filter_4__u_filter_diff_ctr_q[1]),
    .o1(n2863));
 b15nand04ar1n12x5 U3742 (.a(gen_filter_4__u_filter_diff_ctr_q[1]),
    .b(gen_filter_4__u_filter_diff_ctr_q[3]),
    .c(gen_filter_4__u_filter_diff_ctr_q[2]),
    .d(n2862),
    .o1(n2864));
 b15aoai13as1n04x5 U3743 (.a(n2864),
    .b(n2863),
    .c(gen_filter_4__u_filter_diff_ctr_q[1]),
    .d(net2271),
    .o1(gen_filter_4__u_filter_diff_ctr_d[1]));
 b15oai012al1n06x5 U3744 (.a(n2864),
    .b(net2271),
    .c(n2865),
    .o1(gen_filter_4__u_filter_diff_ctr_d[0]));
 b15nor002ar1n02x5 U3745 (.a(n2867),
    .b(n2866),
    .o1(n2868));
 b15and003al1n04x5 U3746 (.a(n2868),
    .b(gen_filter_4__u_filter_diff_ctr_d[1]),
    .c(gen_filter_4__u_filter_diff_ctr_d[0]),
    .o(eq_x_161_n25));
 b15aoai13ar1n04x5 U3747 (.a(n2957),
    .b(gen_filter_8__u_filter_diff_ctr_q[2]),
    .c(gen_filter_8__u_filter_diff_ctr_q[0]),
    .d(gen_filter_8__u_filter_diff_ctr_q[1]),
    .o1(n2869));
 b15nonb02an1n03x5 U3748 (.a(gen_filter_8__u_filter_diff_ctr_q[3]),
    .b(n2869),
    .out0(n2962));
 b15oabi12an1n02x5 U3749 (.a(n2962),
    .b(n2958),
    .c(net2299),
    .out0(gen_filter_8__u_filter_diff_ctr_d[2]));
 b15aoai13as1n04x5 U3750 (.a(n2963),
    .b(net687),
    .c(gen_filter_14__u_filter_diff_ctr_q[0]),
    .d(gen_filter_14__u_filter_diff_ctr_q[1]),
    .o1(n2870));
 b15nonb02ah1n03x5 U3751 (.a(gen_filter_14__u_filter_diff_ctr_q[3]),
    .b(n2870),
    .out0(n2968));
 b15oabi12an1n08x5 U3752 (.a(n2968),
    .b(n2964),
    .c(n2870),
    .out0(gen_filter_14__u_filter_diff_ctr_d[2]));
 b15nand02ar1n02x5 U3753 (.a(gen_filter_3__u_filter_diff_ctr_q[0]),
    .b(gen_filter_3__u_filter_diff_ctr_q[1]),
    .o1(n2871));
 b15oai012aq1n03x5 U3754 (.a(n2871),
    .b(gen_filter_3__u_filter_diff_ctr_q[0]),
    .c(gen_filter_3__u_filter_diff_ctr_q[1]),
    .o1(n2872));
 b15oaoi13an1n08x5 U3755 (.a(n2873),
    .b(n2872),
    .c(n2876),
    .d(n2874),
    .o1(gen_filter_3__u_filter_diff_ctr_d[1]));
 b15oaoi13aq1n08x5 U3756 (.a(n2873),
    .b(net2366),
    .c(n2876),
    .d(n2874),
    .o1(gen_filter_3__u_filter_diff_ctr_d[0]));
 b15nandp3ar1n12x5 U3757 (.o1(n2875),
    .a(gen_filter_3__u_filter_diff_ctr_q[2]),
    .b(gen_filter_3__u_filter_diff_ctr_d[1]),
    .c(gen_filter_3__u_filter_diff_ctr_d[0]));
 b15nor002al1n16x5 U3758 (.a(n2876),
    .b(n2875),
    .o1(eq_x_166_n25));
 b15nand02ar1n02x5 U3759 (.a(gen_filter_17__u_filter_diff_ctr_q[0]),
    .b(gen_filter_17__u_filter_diff_ctr_q[1]),
    .o1(n2877));
 b15oai012aq1n02x5 U3760 (.a(n2877),
    .b(gen_filter_17__u_filter_diff_ctr_q[0]),
    .c(gen_filter_17__u_filter_diff_ctr_q[1]),
    .o1(n2878));
 b15oaoi13an1n04x5 U3761 (.a(net2122),
    .b(n2878),
    .c(n2882),
    .d(n2880),
    .o1(gen_filter_17__u_filter_diff_ctr_d[1]));
 b15oaoi13aq1n04x5 U3762 (.a(n2879),
    .b(net2293),
    .c(n2882),
    .d(n2880),
    .o1(gen_filter_17__u_filter_diff_ctr_d[0]));
 b15nand03al1n06x5 U3763 (.a(gen_filter_17__u_filter_diff_ctr_q[2]),
    .b(gen_filter_17__u_filter_diff_ctr_d[1]),
    .c(gen_filter_17__u_filter_diff_ctr_d[0]),
    .o1(n2881));
 b15norp02ah1n04x5 U3764 (.a(n2882),
    .b(n2881),
    .o1(eq_x_96_n25));
 b15nand02ar1n02x5 U3765 (.a(gen_filter_23__u_filter_diff_ctr_q[0]),
    .b(gen_filter_23__u_filter_diff_ctr_q[1]),
    .o1(n2883));
 b15oai012an1n04x5 U3766 (.a(n2883),
    .b(gen_filter_23__u_filter_diff_ctr_q[0]),
    .c(gen_filter_23__u_filter_diff_ctr_q[1]),
    .o1(n2884));
 b15oaoi13al1n04x5 U3767 (.a(net2162),
    .b(n2884),
    .c(n2888),
    .d(n2886),
    .o1(gen_filter_23__u_filter_diff_ctr_d[1]));
 b15oaoi13al1n04x5 U3768 (.a(net2162),
    .b(gen_filter_23__u_filter_diff_ctr_q[0]),
    .c(n2888),
    .d(n2886),
    .o1(gen_filter_23__u_filter_diff_ctr_d[0]));
 b15nand03an1n04x5 U3769 (.a(gen_filter_23__u_filter_diff_ctr_q[2]),
    .b(gen_filter_23__u_filter_diff_ctr_d[1]),
    .c(gen_filter_23__u_filter_diff_ctr_d[0]),
    .o1(n2887));
 b15nor002aq1n04x5 U3770 (.a(n2888),
    .b(n2887),
    .o1(eq_x_66_n25));
 b15nand02ar1n02x5 U3771 (.a(gen_filter_16__u_filter_diff_ctr_q[0]),
    .b(gen_filter_16__u_filter_diff_ctr_q[1]),
    .o1(n2889));
 b15oai012ar1n02x5 U3772 (.a(n2889),
    .b(gen_filter_16__u_filter_diff_ctr_q[0]),
    .c(gen_filter_16__u_filter_diff_ctr_q[1]),
    .o1(n2890));
 b15oaoi13aq1n03x5 U3773 (.a(n2891),
    .b(n2890),
    .c(n2894),
    .d(n2892),
    .o1(gen_filter_16__u_filter_diff_ctr_d[1]));
 b15oaoi13ar1n04x5 U3774 (.a(n2891),
    .b(gen_filter_16__u_filter_diff_ctr_q[0]),
    .c(n2894),
    .d(n2892),
    .o1(gen_filter_16__u_filter_diff_ctr_d[0]));
 b15nandp3ar1n04x5 U3775 (.a(gen_filter_16__u_filter_diff_ctr_q[2]),
    .b(gen_filter_16__u_filter_diff_ctr_d[1]),
    .c(gen_filter_16__u_filter_diff_ctr_d[0]),
    .o1(n2893));
 b15norp02an1n08x5 U3776 (.a(n2894),
    .b(n2893),
    .o1(eq_x_101_n25));
 b15nand02ar1n02x5 U3777 (.a(gen_filter_5__u_filter_diff_ctr_q[0]),
    .b(gen_filter_5__u_filter_diff_ctr_q[1]),
    .o1(n2895));
 b15oai012ar1n04x5 U3778 (.a(n2895),
    .b(gen_filter_5__u_filter_diff_ctr_q[0]),
    .c(gen_filter_5__u_filter_diff_ctr_q[1]),
    .o1(n2896));
 b15oaoi13ar1n04x5 U3779 (.a(n2897),
    .b(n2896),
    .c(n2900),
    .d(n2898),
    .o1(gen_filter_5__u_filter_diff_ctr_d[1]));
 b15oaoi13aq1n03x5 U3780 (.a(n2897),
    .b(net2352),
    .c(n2900),
    .d(n2898),
    .o1(gen_filter_5__u_filter_diff_ctr_d[0]));
 b15nandp3an1n04x5 U3781 (.a(gen_filter_5__u_filter_diff_ctr_q[2]),
    .b(gen_filter_5__u_filter_diff_ctr_d[1]),
    .c(gen_filter_5__u_filter_diff_ctr_d[0]),
    .o1(n2899));
 b15norp02an1n08x5 U3782 (.a(n2900),
    .b(n2899),
    .o1(eq_x_156_n25));
 b15nand02ar1n02x5 U3783 (.a(gen_filter_2__u_filter_diff_ctr_q[0]),
    .b(gen_filter_2__u_filter_diff_ctr_q[1]),
    .o1(n2901));
 b15oai012ar1n04x5 U3784 (.a(n2901),
    .b(gen_filter_2__u_filter_diff_ctr_q[0]),
    .c(gen_filter_2__u_filter_diff_ctr_q[1]),
    .o1(n2902));
 b15oaoi13ar1n04x5 U3785 (.a(n2903),
    .b(n2902),
    .c(n2906),
    .d(n2904),
    .o1(gen_filter_2__u_filter_diff_ctr_d[1]));
 b15oaoi13as1n03x5 U3786 (.a(n2903),
    .b(gen_filter_2__u_filter_diff_ctr_q[0]),
    .c(n2906),
    .d(n2904),
    .o1(gen_filter_2__u_filter_diff_ctr_d[0]));
 b15nand03aq1n04x5 U3787 (.a(net2448),
    .b(gen_filter_2__u_filter_diff_ctr_d[1]),
    .c(gen_filter_2__u_filter_diff_ctr_d[0]),
    .o1(n2905));
 b15nor002an1n06x5 U3788 (.a(n2906),
    .b(n2905),
    .o1(eq_x_171_n25));
 b15nand02ar1n02x5 U3789 (.a(gen_filter_31__u_filter_diff_ctr_q[0]),
    .b(gen_filter_31__u_filter_diff_ctr_q[1]),
    .o1(n2907));
 b15oai012aq1n03x5 U3790 (.a(n2907),
    .b(gen_filter_31__u_filter_diff_ctr_q[0]),
    .c(gen_filter_31__u_filter_diff_ctr_q[1]),
    .o1(n2908));
 b15oaoi13aq1n04x5 U3791 (.a(n2909),
    .b(n2908),
    .c(n2912),
    .d(n2910),
    .o1(gen_filter_31__u_filter_diff_ctr_d[1]));
 b15oaoi13ar1n08x5 U3792 (.a(n2909),
    .b(gen_filter_31__u_filter_diff_ctr_q[0]),
    .c(n2912),
    .d(n2910),
    .o1(gen_filter_31__u_filter_diff_ctr_d[0]));
 b15nandp3ar1n04x5 U3793 (.a(gen_filter_31__u_filter_diff_ctr_q[2]),
    .b(gen_filter_31__u_filter_diff_ctr_d[1]),
    .c(gen_filter_31__u_filter_diff_ctr_d[0]),
    .o1(n2911));
 b15norp02ah1n03x5 U3794 (.a(n2912),
    .b(n2911),
    .o1(eq_x_26_n25));
 b15nand02ar1n02x5 U3795 (.a(gen_filter_15__u_filter_diff_ctr_q[0]),
    .b(gen_filter_15__u_filter_diff_ctr_q[1]),
    .o1(n2913));
 b15oai012ar1n04x5 U3796 (.a(n2913),
    .b(gen_filter_15__u_filter_diff_ctr_q[0]),
    .c(gen_filter_15__u_filter_diff_ctr_q[1]),
    .o1(n2914));
 b15oaoi13ar1n04x5 U3797 (.a(net2181),
    .b(n2914),
    .c(n2918),
    .d(net2203),
    .o1(gen_filter_15__u_filter_diff_ctr_d[1]));
 b15oaoi13ah1n04x5 U3798 (.a(n2915),
    .b(gen_filter_15__u_filter_diff_ctr_q[0]),
    .c(net2153),
    .d(n2916),
    .o1(gen_filter_15__u_filter_diff_ctr_d[0]));
 b15nand03ar1n03x5 U3799 (.a(gen_filter_15__u_filter_diff_ctr_q[2]),
    .b(gen_filter_15__u_filter_diff_ctr_d[1]),
    .c(gen_filter_15__u_filter_diff_ctr_d[0]),
    .o1(n2917));
 b15norp02ah1n02x5 U3800 (.a(n2918),
    .b(n2917),
    .o1(eq_x_106_n25));
 b15nand02ar1n02x5 U3801 (.a(gen_filter_27__u_filter_diff_ctr_q[0]),
    .b(gen_filter_27__u_filter_diff_ctr_q[1]),
    .o1(n2919));
 b15oai012ar1n04x5 U3802 (.a(n2919),
    .b(gen_filter_27__u_filter_diff_ctr_q[0]),
    .c(gen_filter_27__u_filter_diff_ctr_q[1]),
    .o1(n2920));
 b15oaoi13an1n04x5 U3803 (.a(n2921),
    .b(n2920),
    .c(n2924),
    .d(n2922),
    .o1(gen_filter_27__u_filter_diff_ctr_d[1]));
 b15oaoi13al1n08x5 U3804 (.a(n2921),
    .b(gen_filter_27__u_filter_diff_ctr_q[0]),
    .c(n2924),
    .d(n2922),
    .o1(gen_filter_27__u_filter_diff_ctr_d[0]));
 b15nandp3aq1n03x5 U3805 (.a(gen_filter_27__u_filter_diff_ctr_q[2]),
    .b(gen_filter_27__u_filter_diff_ctr_d[1]),
    .c(gen_filter_27__u_filter_diff_ctr_d[0]),
    .o1(n2923));
 b15norp02aq1n04x5 U3806 (.a(n2924),
    .b(n2923),
    .o1(eq_x_46_n25));
 b15oai012aq1n02x5 U3807 (.a(n2925),
    .b(gen_filter_25__u_filter_diff_ctr_q[0]),
    .c(gen_filter_25__u_filter_diff_ctr_q[1]),
    .o1(n2927));
 b15aoi012aq1n04x5 U3808 (.a(n2926),
    .b(n2930),
    .c(n2927),
    .o1(gen_filter_25__u_filter_diff_ctr_d[1]));
 b15inv040aq1n02x5 U3809 (.a(gen_filter_25__u_filter_diff_ctr_d[1]),
    .o1(n2928));
 b15aoi112as1n08x5 U3810 (.a(n2929),
    .b(n2928),
    .c(gen_filter_25__u_filter_diff_ctr_q[0]),
    .d(n2930),
    .o1(eq_x_56_n25));
 b15oai012aq1n02x5 U3811 (.a(n2931),
    .b(gen_filter_13__u_filter_diff_ctr_q[0]),
    .c(gen_filter_13__u_filter_diff_ctr_q[1]),
    .o1(n2933));
 b15aoi012ar1n04x5 U3812 (.a(n2932),
    .b(n2936),
    .c(n2933),
    .o1(gen_filter_13__u_filter_diff_ctr_d[1]));
 b15inv040ar1n02x5 U3813 (.a(gen_filter_13__u_filter_diff_ctr_d[1]),
    .o1(n2934));
 b15aoi112ar1n06x5 U3814 (.a(n2935),
    .b(n2934),
    .c(gen_filter_13__u_filter_diff_ctr_q[0]),
    .d(n2936),
    .o1(eq_x_116_n25));
 b15inv040al1n02x5 U3815 (.a(n2937),
    .o1(n2943));
 b15nand02ah1n04x5 U3816 (.a(n2943),
    .b(n2938),
    .o1(n2941));
 b15oai012aq1n08x5 U3817 (.a(n2941),
    .b(gen_filter_11__u_filter_diff_ctr_q[0]),
    .c(n2939),
    .o1(gen_filter_11__u_filter_diff_ctr_d[0]));
 b15oai012ah1n03x5 U3818 (.a(n2940),
    .b(gen_filter_11__u_filter_diff_ctr_q[0]),
    .c(gen_filter_11__u_filter_diff_ctr_q[1]),
    .o1(n2942));
 b15aoai13an1n08x5 U3819 (.a(n2941),
    .b(n2942),
    .c(gen_filter_11__u_filter_diff_ctr_q[1]),
    .d(gen_filter_11__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_11__u_filter_diff_ctr_d[1]));
 b15nand03an1n04x5 U3820 (.a(n2943),
    .b(gen_filter_11__u_filter_diff_ctr_d[0]),
    .c(gen_filter_11__u_filter_diff_ctr_d[1]),
    .o1(n2944));
 b15nor002as1n04x5 U3821 (.a(n2945),
    .b(n2944),
    .o1(eq_x_126_n25));
 b15nanb02al1n04x5 U3822 (.a(n4046),
    .b(n2946),
    .out0(n2949));
 b15oai012aq1n06x5 U3823 (.a(n2949),
    .b(net2422),
    .c(n2947),
    .o1(gen_filter_18__u_filter_diff_ctr_d[0]));
 b15oai012al1n02x5 U3824 (.a(n2948),
    .b(gen_filter_18__u_filter_diff_ctr_q[0]),
    .c(gen_filter_18__u_filter_diff_ctr_q[1]),
    .o1(n2950));
 b15aoai13ah1n03x5 U3825 (.a(n2949),
    .b(n2950),
    .c(net2356),
    .d(gen_filter_18__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_18__u_filter_diff_ctr_d[1]));
 b15aboi22al1n08x5 U3826 (.a(net1970),
    .b(net1982),
    .c(net1970),
    .d(n2951),
    .out0(net240));
 b15inv000aq1n16x5 U3827 (.a(net2035),
    .o1(net242));
 b15aboi22ar1n08x5 U3828 (.a(net1990),
    .b(n2952),
    .c(net1990),
    .d(net1986),
    .out0(n2955));
 b15aoi022ah1n48x5 U3829 (.a(net674),
    .b(net242),
    .c(net1994),
    .d(n2953),
    .o1(n2954));
 b15xor002aq1n06x5 U3830 (.a(n2955),
    .b(net1995),
    .out0(n2956));
 b15xor002al1n03x5 U3831 (.a(net1996),
    .b(net1983),
    .out0(net298));
 b15xor002al1n03x5 U3832 (.a(net1992),
    .b(n2956),
    .out0(net238));
 b15oai012ar1n02x5 U3833 (.a(n2957),
    .b(gen_filter_8__u_filter_diff_ctr_q[0]),
    .c(gen_filter_8__u_filter_diff_ctr_q[1]),
    .o1(n2959));
 b15nandp2aq1n02x5 U3834 (.a(n2962),
    .b(n2958),
    .o1(n2960));
 b15aoai13ar1n03x5 U3835 (.a(n2960),
    .b(n2959),
    .c(net2328),
    .d(gen_filter_8__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_8__u_filter_diff_ctr_d[1]));
 b15oai012ah1n02x5 U3836 (.a(n2960),
    .b(net2335),
    .c(n2961),
    .o1(gen_filter_8__u_filter_diff_ctr_d[0]));
 b15and003ar1n03x5 U3837 (.a(n2962),
    .b(gen_filter_8__u_filter_diff_ctr_d[1]),
    .c(gen_filter_8__u_filter_diff_ctr_d[0]),
    .o(eq_x_141_n25));
 b15oai012al1n04x5 U3838 (.a(n2963),
    .b(gen_filter_14__u_filter_diff_ctr_q[0]),
    .c(gen_filter_14__u_filter_diff_ctr_q[1]),
    .o1(n2965));
 b15nand02ah1n04x5 U3839 (.a(n2968),
    .b(n2964),
    .o1(n2966));
 b15aoai13ar1n08x5 U3840 (.a(n2966),
    .b(n2965),
    .c(gen_filter_14__u_filter_diff_ctr_q[1]),
    .d(gen_filter_14__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_14__u_filter_diff_ctr_d[1]));
 b15oai012ah1n06x5 U3841 (.a(n2966),
    .b(gen_filter_14__u_filter_diff_ctr_q[0]),
    .c(n2967),
    .o1(gen_filter_14__u_filter_diff_ctr_d[0]));
 b15and003aq1n08x5 U3842 (.a(n2968),
    .b(gen_filter_14__u_filter_diff_ctr_d[1]),
    .c(gen_filter_14__u_filter_diff_ctr_d[0]),
    .o(eq_x_111_n25));
 b15nanb02al1n24x5 U3843 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .b(n2973),
    .out0(n2971));
 b15inv040an1n06x5 U3844 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .o1(n2970));
 b15nandp2ar1n12x5 U3845 (.a(n2971),
    .b(net2455),
    .o1(n2969));
 b15oai012ah1n32x5 U3846 (.a(n2969),
    .b(n2971),
    .c(n2970),
    .o1(gen_alert_tx_0__u_prim_alert_sender_ack_level));
 b15nandp2al1n08x5 U3847 (.a(net2467),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39));
 b15nonb03as1n12x5 U3848 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39),
    .b(n2973),
    .c(n2972),
    .out0(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[1]));
 b15nandp2ah1n05x5 U3849 (.a(net2441),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39));
 b15nonb03al1n12x5 U3850 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39),
    .b(n2975),
    .c(n2974),
    .out0(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[1]));
 b15inv000ah1n10x5 U3851 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .o1(n3355));
 b15nor002ar1n04x5 U3852 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .b(n3355),
    .o1(n2981));
 b15nor002aq1n04x5 U3853 (.a(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .b(gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .o1(n3059));
 b15oabi12aq1n06x5 U3854 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .b(n2977),
    .c(n2976),
    .out0(n2978));
 b15oaoi13as1n08x5 U3855 (.a(gen_alert_tx_0__u_prim_alert_sender_ping_set_q),
    .b(n2978),
    .c(n2980),
    .d(n2979),
    .o1(n3351));
 b15norp02as1n04x5 U3856 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[1]),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[1]),
    .o1(n3867));
 b15inv040as1n05x5 U3857 (.a(n3867),
    .o1(n3361));
 b15aoi112as1n06x5 U3858 (.a(n3351),
    .b(n3361),
    .c(n2981),
    .d(n3059),
    .o1(gen_alert_tx_0__u_prim_alert_sender_ping_set_d));
 b15inv040aq1n05x5 U3859 (.a(net2109),
    .o1(n3018));
 b15aboi22al1n12x5 U3860 (.a(net495),
    .b(n3018),
    .c(net2109),
    .d(net495),
    .out0(n2985));
 b15inv020aq1n28x5 U3861 (.a(net246),
    .o1(n3028));
 b15inv000ar1n16x5 U3862 (.a(net2043),
    .o1(n3071));
 b15aoi022an1n24x5 U3863 (.a(net475),
    .b(n3028),
    .c(net468),
    .d(n3071),
    .o1(n2997));
 b15inv040aq1n12x5 U3864 (.a(net501),
    .o1(n3007));
 b15inv040aq1n05x5 U3865 (.a(net2022),
    .o1(n3000));
 b15aoi022ah1n06x5 U3866 (.a(net2022),
    .b(n3007),
    .c(net501),
    .d(n3000),
    .o1(n2982));
 b15xor002ah1n03x5 U3867 (.a(n2997),
    .b(n2982),
    .out0(n2983));
 b15inv040as1n10x5 U3868 (.a(net470),
    .o1(n2991));
 b15inv020aq1n12x5 U3869 (.a(net2158),
    .o1(n3062));
 b15aoi022ar1n48x5 U3870 (.a(net2136),
    .b(net470),
    .c(n2991),
    .d(net2159),
    .o1(n3055));
 b15xor002as1n03x5 U3871 (.a(n2983),
    .b(n3055),
    .out0(n2984));
 b15xor002ah1n06x5 U3872 (.a(n2985),
    .b(n2984),
    .out0(n2988));
 b15inv040as1n12x5 U3873 (.a(net489),
    .o1(n2992));
 b15inv000ar1n28x5 U3874 (.a(net499),
    .o1(n3031));
 b15aoi022as1n48x5 U3875 (.a(net500),
    .b(net487),
    .c(net454),
    .d(n3031),
    .o1(n3024));
 b15inv040ah1n08x5 U3876 (.a(net457),
    .o1(n3005));
 b15aboi22al1n12x5 U3877 (.a(net2143),
    .b(n3005),
    .c(net456),
    .d(net2143),
    .out0(n2986));
 b15xor002aq1n08x5 U3878 (.a(n3024),
    .b(n2986),
    .out0(n2987));
 b15xor002aq1n08x5 U3879 (.a(net2215),
    .b(n2987),
    .out0(net297));
 b15inv000an1n05x5 U3880 (.a(net469),
    .o1(n3041));
 b15aboi22as1n08x5 U3881 (.a(net254),
    .b(n3041),
    .c(net254),
    .d(net469),
    .out0(n2990));
 b15inv040as1n03x5 U3882 (.a(net2012),
    .o1(n3003));
 b15inv040as1n12x5 U3883 (.a(net459),
    .o1(n3050));
 b15aoi022ah1n12x5 U3884 (.a(net459),
    .b(net2012),
    .c(n3003),
    .d(n3050),
    .o1(n2989));
 b15xor002an1n16x5 U3885 (.a(n2990),
    .b(net2118),
    .out0(n3019));
 b15inv040ah1n28x5 U3886 (.a(net494),
    .o1(n3034));
 b15inv020ah1n40x5 U3887 (.a(net481),
    .o1(n3012));
 b15aoi022as1n48x5 U3888 (.a(net482),
    .b(net491),
    .c(n3034),
    .d(n3012),
    .o1(n2994));
 b15aoi022an1n12x5 U3889 (.a(net471),
    .b(net488),
    .c(n2992),
    .d(n2991),
    .o1(n2993));
 b15xor002ar1n12x5 U3890 (.a(n2994),
    .b(n2993),
    .out0(n2995));
 b15inv040ah1n12x5 U3891 (.a(net474),
    .o1(n3026));
 b15inv000as1n06x5 U3892 (.a(net479),
    .o1(n3008));
 b15aoi022aq1n12x5 U3893 (.a(net479),
    .b(net472),
    .c(net452),
    .d(n3008),
    .o1(n3054));
 b15xor002an1n08x5 U3894 (.a(n2995),
    .b(net404),
    .out0(n2996));
 b15xor002an1n08x5 U3895 (.a(n2997),
    .b(n2996),
    .out0(n2998));
 b15inv040ah1n08x5 U3896 (.a(net466),
    .o1(n3004));
 b15inv000as1n06x5 U3897 (.a(net269),
    .o1(n3045));
 b15aoi022ah1n24x5 U3898 (.a(net269),
    .b(net466),
    .c(n3004),
    .d(n3045),
    .o1(n3064));
 b15xor002ah1n08x5 U3899 (.a(n2998),
    .b(n3064),
    .out0(n2999));
 b15xor002as1n04x5 U3900 (.a(net2119),
    .b(n2999),
    .out0(net296));
 b15inv000aq1n24x5 U3901 (.a(net477),
    .o1(n3015));
 b15inv040as1n24x5 U3902 (.a(net486),
    .o1(n3030));
 b15aoi022ah1n32x5 U3903 (.a(net485),
    .b(net478),
    .c(n3015),
    .d(n3030),
    .o1(n3002));
 b15inv000al1n10x5 U3904 (.a(net2085),
    .o1(n3061));
 b15aoi022as1n16x5 U3905 (.a(net2022),
    .b(n3061),
    .c(net2085),
    .d(n3000),
    .o1(n3001));
 b15xor002ah1n16x5 U3906 (.a(n3002),
    .b(n3001),
    .out0(n3057));
 b15aoi022an1n12x5 U3907 (.a(net2012),
    .b(net2066),
    .c(n3004),
    .d(n3003),
    .o1(n3006));
 b15inv040as1n08x5 U3908 (.a(net2146),
    .o1(n3070));
 b15aoi022al1n32x5 U3909 (.a(net456),
    .b(n3070),
    .c(net2146),
    .d(n3005),
    .o1(n3022));
 b15xor002as1n12x5 U3910 (.a(n3006),
    .b(n3022),
    .out0(n3010));
 b15inv040as1n20x5 U3911 (.a(net460),
    .o1(n3029));
 b15aoi022an1n48x5 U3912 (.a(net461),
    .b(net245),
    .c(n3007),
    .d(net451),
    .o1(n3063));
 b15aboi22al1n16x5 U3913 (.a(net403),
    .b(n3008),
    .c(net479),
    .d(net403),
    .out0(n3009));
 b15xor002ah1n03x5 U3914 (.a(n3010),
    .b(net363),
    .out0(n3011));
 b15xor002aq1n06x5 U3915 (.a(n3057),
    .b(n3011),
    .out0(n3014));
 b15inv020as1n32x5 U3916 (.a(net496),
    .o1(n3016));
 b15aoi022an1n48x5 U3917 (.a(net497),
    .b(net480),
    .c(n3012),
    .d(n3016),
    .o1(n3013));
 b15xor002as1n16x5 U3918 (.a(net2142),
    .b(n3013),
    .out0(n3036));
 b15xor002as1n08x5 U3919 (.a(n3014),
    .b(net2187),
    .out0(net280));
 b15aoi022aq1n32x5 U3920 (.a(net476),
    .b(net498),
    .c(n3016),
    .d(n3015),
    .o1(n3017));
 b15inv040ah1n10x5 U3921 (.a(net504),
    .o1(n3042));
 b15inv000ah1n08x5 U3922 (.a(net464),
    .o1(n3049));
 b15aoi022al1n24x5 U3923 (.a(net464),
    .b(net502),
    .c(net450),
    .d(n3049),
    .o1(n3065));
 b15xor002ah1n03x5 U3924 (.a(n3017),
    .b(net402),
    .out0(n3021));
 b15inv040aq1n05x5 U3925 (.a(net2018),
    .o1(n3027));
 b15aoi022as1n16x5 U3926 (.a(net2109),
    .b(net2018),
    .c(n3027),
    .d(n3018),
    .o1(n3048));
 b15xor002ar1n06x5 U3927 (.a(n3048),
    .b(n3019),
    .out0(n3020));
 b15xor002an1n04x5 U3928 (.a(n3021),
    .b(n3020),
    .out0(n3023));
 b15xor002ah1n04x5 U3929 (.a(n3023),
    .b(n3022),
    .out0(n3025));
 b15xor002aq1n08x5 U3930 (.a(n3025),
    .b(n3024),
    .out0(net290));
 b15aoi022an1n12x5 U3931 (.a(net474),
    .b(net2018),
    .c(n3027),
    .d(n3026),
    .o1(n3040));
 b15aoi022al1n48x5 U3932 (.a(net467),
    .b(net462),
    .c(net451),
    .d(n3028),
    .o1(n3033));
 b15aoi022ah1n24x5 U3933 (.a(net483),
    .b(net255),
    .c(n3031),
    .d(n3030),
    .o1(n3032));
 b15xor002al1n16x5 U3934 (.a(n3033),
    .b(net401),
    .out0(n3038));
 b15inv020as1n06x5 U3935 (.a(net2071),
    .o1(n3046));
 b15aoi022an1n16x5 U3936 (.a(net2071),
    .b(net493),
    .c(n3034),
    .d(n3046),
    .o1(n3035));
 b15xor002as1n16x5 U3937 (.a(net495),
    .b(n3035),
    .out0(n3075));
 b15xor002an1n12x5 U3938 (.a(n3036),
    .b(n3075),
    .out0(n3037));
 b15xor002ah1n12x5 U3939 (.a(n3038),
    .b(n3037),
    .out0(n3039));
 b15xor002as1n12x5 U3940 (.a(n3040),
    .b(n3039),
    .out0(n3044));
 b15aoi022ar1n08x5 U3941 (.a(net469),
    .b(net2024),
    .c(n3042),
    .d(n3041),
    .o1(n3043));
 b15xor002an1n03x5 U3942 (.a(net2113),
    .b(n3043),
    .out0(net259));
 b15aoi022an1n12x5 U3943 (.a(net269),
    .b(net2071),
    .c(n3046),
    .d(n3045),
    .o1(n3047));
 b15xor002as1n06x5 U3944 (.a(n3048),
    .b(n3047),
    .out0(n3052));
 b15aoi022aq1n16x5 U3945 (.a(net465),
    .b(net458),
    .c(net453),
    .d(n3049),
    .o1(n3051));
 b15xor002as1n03x5 U3946 (.a(n3052),
    .b(net400),
    .out0(n3053));
 b15xor002aq1n06x5 U3947 (.a(net404),
    .b(n3053),
    .out0(n3056));
 b15qgbxo2an1n10x5 U3948 (.a(n3056),
    .b(n3055),
    .out0(n3058));
 b15qgbxo2an1n10x5 U3949 (.a(n3058),
    .b(n3057),
    .out0(net270));
 b15oai012an1n12x5 U3950 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .b(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .c(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .o1(n3865));
 b15inv040al1n03x5 U3951 (.a(n3059),
    .o1(n3060));
 b15aoi013ah1n06x5 U3952 (.a(n3361),
    .b(n3865),
    .c(n3355),
    .d(n3060),
    .o1(n3301));
 b15inv040ah1n05x5 U3953 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .o1(n3350));
 b15aoi022ah1n12x5 U3954 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .b(n3350),
    .c(gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .d(n3355),
    .o1(n3442));
 b15nonb02ar1n02x3 U3955 (.a(n3301),
    .b(n3442),
    .out0(gen_alert_tx_0__u_prim_alert_sender_state_d[2]));
 b15aoi022as1n06x5 U3956 (.a(net2085),
    .b(net2136),
    .c(net2159),
    .d(n3061),
    .o1(n3069));
 b15xor002ar1n12x5 U3957 (.a(n3064),
    .b(n3063),
    .out0(n3067));
 b15xor002ah1n16x5 U3958 (.a(net254),
    .b(net402),
    .out0(n3066));
 b15xor002al1n12x5 U3959 (.a(n3067),
    .b(n3066),
    .out0(n3068));
 b15xor002aq1n06x5 U3960 (.a(n3069),
    .b(n3068),
    .out0(n3073));
 b15aoi022an1n16x5 U3961 (.a(net2146),
    .b(net2044),
    .c(n3071),
    .d(n3070),
    .o1(n3072));
 b15xor002an1n12x5 U3962 (.a(n3073),
    .b(n3072),
    .out0(n3074));
 b15xor002an1n16x5 U3963 (.a(n3075),
    .b(n3074),
    .out0(net295));
 b15inv040as1n08x5 U3964 (.a(net92),
    .o1(n3254));
 b15inv040ar1n10x5 U3965 (.a(net91),
    .o1(n3255));
 b15inv000ar1n16x5 U3966 (.a(net93),
    .o1(n3249));
 b15norp03al1n08x5 U3967 (.a(n3254),
    .b(n3255),
    .c(n3249),
    .o1(n3080));
 b15inv040ah1n08x5 U3968 (.a(net90),
    .o1(n3248));
 b15oai112aq1n02x5 U3969 (.a(n3255),
    .b(n3249),
    .c(net95),
    .d(net39),
    .o1(n3076));
 b15oai013as1n03x5 U3970 (.a(n3076),
    .b(net92),
    .c(net90),
    .d(net95),
    .o1(n3077));
 b15obai22aq1n06x5 U3971 (.a(n3080),
    .b(n3248),
    .c(net40),
    .d(n3077),
    .out0(n3299));
 b15norp03an1n08x5 U3972 (.a(net92),
    .b(net93),
    .c(net96),
    .o1(n3288));
 b15inv000al1n12x5 U3973 (.a(net95),
    .o1(n3284));
 b15aoi022ar1n08x5 U3974 (.a(net95),
    .b(net90),
    .c(net91),
    .d(n3284),
    .o1(n3078));
 b15aoi112ah1n04x5 U3975 (.a(net40),
    .b(net39),
    .c(n3288),
    .d(n3078),
    .o1(n3297));
 b15nor002aq1n02x5 U3976 (.a(net93),
    .b(net95),
    .o1(n3079));
 b15inv040as1n05x5 U3977 (.a(net96),
    .o1(n3283));
 b15nor003ar1n06x5 U3978 (.a(net91),
    .b(net90),
    .c(n3283),
    .o1(n3289));
 b15aoai13as1n04x5 U3979 (.a(n3289),
    .b(n3079),
    .c(net95),
    .d(n3254),
    .o1(n3296));
 b15nandp2ah1n32x5 U3980 (.a(net709),
    .b(net98),
    .o1(n3313));
 b15norp03as1n24x5 U3981 (.a(net99),
    .b(net100),
    .c(n3313),
    .o1(n3300));
 b15inv000as1n08x5 U3982 (.a(net43),
    .o1(n3863));
 b15nandp2as1n12x5 U3983 (.a(net672),
    .b(n3863),
    .o1(n3308));
 b15oaoi13aq1n04x5 U3984 (.a(n3308),
    .b(net90),
    .c(n3080),
    .d(n3300),
    .o1(n3295));
 b15inv040as1n04x5 U3985 (.a(net51),
    .o1(n3115));
 b15aoi022an1n16x5 U3986 (.a(net51),
    .b(net96),
    .c(n3283),
    .d(n3115),
    .o1(n3092));
 b15inv040ar1n06x5 U3987 (.a(net53),
    .o1(n3147));
 b15inv040as1n20x5 U3988 (.a(net99),
    .o1(n3311));
 b15aoi022as1n08x5 U3989 (.a(net99),
    .b(net53),
    .c(n3147),
    .d(n3311),
    .o1(n3088));
 b15inv000ah1n05x5 U3990 (.a(net41),
    .o1(n3244));
 b15aboi22aq1n08x5 U3991 (.a(net107),
    .b(n3244),
    .c(net107),
    .d(net41),
    .out0(n3081));
 b15xor002as1n08x5 U3992 (.a(net128),
    .b(n3081),
    .out0(n3256));
 b15xor002ah1n16x5 U3993 (.a(net124),
    .b(net123),
    .out0(n3121));
 b15xor002ar1n12x5 U3994 (.a(n3121),
    .b(net49),
    .out0(n3083));
 b15xor002an1n16x5 U3995 (.a(net101),
    .b(net102),
    .out0(n3242));
 b15xor002ah1n16x5 U3996 (.a(net117),
    .b(net120),
    .out0(n3137));
 b15qgbxo2an1n10x5 U3997 (.a(n3242),
    .b(n3137),
    .out0(n3082));
 b15xor002as1n08x5 U3998 (.a(n3083),
    .b(n3082),
    .out0(n3084));
 b15xor002al1n12x5 U3999 (.a(n3256),
    .b(n3084),
    .out0(n3086));
 b15xor002as1n08x5 U4000 (.a(net112),
    .b(net113),
    .out0(n3085));
 b15xor002aq1n16x5 U4001 (.a(n3086),
    .b(n3085),
    .out0(n3087));
 b15xor002ar1n12x5 U4002 (.a(n3088),
    .b(n3087),
    .out0(n3090));
 b15xor002an1n12x5 U4003 (.a(net122),
    .b(net110),
    .out0(n3089));
 b15xor002al1n12x5 U4004 (.a(n3090),
    .b(n3089),
    .out0(n3091));
 b15qgbxo2an1n10x5 U4005 (.a(n3092),
    .b(n3091),
    .out0(n3114));
 b15qgbin1an1n15x5 U4006 (.a(net50),
    .o1(n3281));
 b15aboi22ah1n16x5 U4007 (.a(net119),
    .b(net50),
    .c(net119),
    .d(n3281),
    .out0(n3113));
 b15nandp2aq1n03x5 U4008 (.a(n3114),
    .b(n3113),
    .o1(n3112));
 b15ztpn00an1n08x5 PHY_64 ();
 b15ztpn00an1n08x5 PHY_63 ();
 b15aoi022ar1n12x5 U4011 (.a(net82),
    .b(n4132),
    .c(net75),
    .d(net694),
    .o1(n3093));
 b15xor002as1n08x5 U4012 (.a(net54),
    .b(n3093),
    .out0(n3094));
 b15xor002as1n12x5 U4013 (.a(n3094),
    .b(net720),
    .out0(n3110));
 b15ztpn00an1n08x5 PHY_62 ();
 b15ztpn00an1n08x5 PHY_61 ();
 b15aoi022ah1n06x5 U4016 (.a(net66),
    .b(n4123),
    .c(net719),
    .d(n4125),
    .o1(n3099));
 b15ztpn00an1n08x5 PHY_60 ();
 b15ztpn00an1n08x5 PHY_59 ();
 b15aoi022ah1n24x5 U4019 (.a(net68),
    .b(net722),
    .c(n4118),
    .d(n4127),
    .o1(n3216));
 b15ztpn00an1n08x5 PHY_58 ();
 b15ztpn00an1n08x5 PHY_57 ();
 b15aoi022ah1n06x5 U4022 (.a(net84),
    .b(net67),
    .c(n4126),
    .d(n4140),
    .o1(n3095));
 b15xor002al1n08x5 U4023 (.a(n3216),
    .b(n3095),
    .out0(n3097));
 b15ztpn00an1n08x5 PHY_56 ();
 b15ztpn00an1n08x5 PHY_55 ();
 b15aoi022ar1n48x5 U4026 (.a(net717),
    .b(net715),
    .c(n4131),
    .d(net701),
    .o1(n3190));
 b15xor002an1n06x5 U4027 (.a(n3190),
    .b(net724),
    .out0(n3096));
 b15xor002al1n08x5 U4028 (.a(n3097),
    .b(n3096),
    .out0(n3098));
 b15xor002as1n06x5 U4029 (.a(n3099),
    .b(n3098),
    .out0(n3100));
 b15inv040as1n60x5 U4030 (.a(net69),
    .o1(n3818));
 b15ztpn00an1n08x5 PHY_54 ();
 b15norp02ah1n48x5 U4032 (.a(n3818),
    .b(net692),
    .o1(n3828));
 b15oabi12as1n24x5 U4033 (.a(n3828),
    .b(net69),
    .c(net87),
    .out0(n3225));
 b15xor002an1n16x5 U4034 (.a(n3100),
    .b(n3225),
    .out0(n3109));
 b15ztpn00an1n08x5 PHY_53 ();
 b15aoi022aq1n16x5 U4036 (.a(net719),
    .b(net723),
    .c(n4117),
    .d(n4123),
    .o1(n3212));
 b15ztpn00an1n08x5 PHY_52 ();
 b15aoi022ar1n32x5 U4038 (.a(net75),
    .b(net714),
    .c(n4133),
    .d(n4132),
    .o1(n3221));
 b15ztpn00an1n08x5 PHY_51 ();
 b15aoi022ar1n24x5 U4040 (.a(net717),
    .b(net88),
    .c(n4144),
    .d(net701),
    .o1(n3101));
 b15xor002al1n16x5 U4041 (.a(n3221),
    .b(n3101),
    .out0(n3103));
 b15ztpn00an1n08x5 PHY_50 ();
 b15ztpn00an1n08x5 PHY_49 ();
 b15aoi022al1n48x5 U4044 (.a(net63),
    .b(net77),
    .c(n4134),
    .d(n4122),
    .o1(n3211));
 b15ztpn00an1n08x5 PHY_48 ();
 b15ztpn00an1n08x5 PHY_47 ();
 b15aoi022aq1n16x5 U4047 (.a(net712),
    .b(net721),
    .c(n4119),
    .d(n4138),
    .o1(n3222));
 b15xor002an1n08x5 U4048 (.a(n3211),
    .b(n3222),
    .out0(n3102));
 b15xor002an1n12x5 U4049 (.a(n3103),
    .b(n3102),
    .out0(n3104));
 b15xor002ar1n12x5 U4050 (.a(n3212),
    .b(n3104),
    .out0(n3105));
 b15ztpn00an1n08x5 PHY_46 ();
 b15aoi022ah1n24x5 U4052 (.a(net67),
    .b(net713),
    .c(n4135),
    .d(n4126),
    .o1(n3176));
 b15xor002an1n12x5 U4053 (.a(n3105),
    .b(n3176),
    .out0(n3108));
 b15ztpn00an1n08x5 PHY_45 ();
 b15ztpn00an1n08x5 PHY_44 ();
 b15oai022ar1n32x5 U4056 (.a(n4120),
    .b(net73),
    .c(n4130),
    .d(net720),
    .o1(n3202));
 b15xnr002aq1n12x5 U4057 (.a(net72),
    .b(n3202),
    .out0(n3107));
 b15oai022al1n08x5 U4058 (.a(n3110),
    .b(n3109),
    .c(n3107),
    .d(n3108),
    .o1(n3106));
 b15aoi122as1n08x5 U4059 (.a(n3106),
    .b(n3110),
    .c(n3109),
    .d(n3108),
    .e(n3107),
    .o1(n3111));
 b15oai112ah1n12x5 U4060 (.a(n3112),
    .b(n3111),
    .c(n3114),
    .d(n3113),
    .o1(n3280));
 b15xor002as1n08x5 U4061 (.a(net106),
    .b(net113),
    .out0(n3118));
 b15inv000ah1n04x5 U4062 (.a(net126),
    .o1(n3149));
 b15aoi022as1n12x5 U4063 (.a(net126),
    .b(net51),
    .c(n3115),
    .d(n3149),
    .o1(n3116));
 b15xor002an1n16x5 U4064 (.a(net129),
    .b(n3116),
    .out0(n3133));
 b15xor002as1n08x5 U4065 (.a(net111),
    .b(n3133),
    .out0(n3117));
 b15xor002as1n16x5 U4066 (.a(n3118),
    .b(n3117),
    .out0(n3257));
 b15inv040an1n12x5 U4067 (.a(net98),
    .o1(n3302));
 b15aboi22an1n08x5 U4068 (.a(net115),
    .b(n3302),
    .c(net98),
    .d(net115),
    .out0(n3128));
 b15inv020ah1n16x5 U4069 (.a(net100),
    .o1(n3303));
 b15aboi22ah1n06x5 U4070 (.a(net120),
    .b(n3303),
    .c(net100),
    .d(net120),
    .out0(n3124));
 b15aoi022ar1n32x5 U4071 (.a(net93),
    .b(net95),
    .c(n3284),
    .d(n3249),
    .o1(n3120));
 b15inv040as1n04x5 U4072 (.a(net52),
    .o1(n3282));
 b15aboi22aq1n08x5 U4073 (.a(net121),
    .b(n3282),
    .c(net52),
    .d(net121),
    .out0(n3119));
 b15xor002ah1n08x5 U4074 (.a(n3120),
    .b(n3119),
    .out0(n3122));
 b15xor002al1n16x5 U4075 (.a(n3122),
    .b(n3121),
    .out0(n3123));
 b15xor002al1n06x5 U4076 (.a(n3124),
    .b(n3123),
    .out0(n3126));
 b15xor002al1n06x5 U4077 (.a(net102),
    .b(net48),
    .out0(n3125));
 b15xor002aq1n06x5 U4078 (.a(n3126),
    .b(n3125),
    .out0(n3127));
 b15xor002as1n08x5 U4079 (.a(n3128),
    .b(n3127),
    .out0(n3130));
 b15xor002ah1n12x5 U4080 (.a(net118),
    .b(net109),
    .out0(n3129));
 b15xor002an1n16x5 U4081 (.a(n3130),
    .b(n3129),
    .out0(n3146));
 b15aboi22as1n24x5 U4082 (.a(net125),
    .b(n3281),
    .c(net125),
    .d(net50),
    .out0(n3258));
 b15xor002ah1n16x5 U4083 (.a(net43),
    .b(n3258),
    .out0(n3162));
 b15inv040as1n02x5 U4084 (.a(net128),
    .o1(n3131));
 b15aboi22aq1n16x5 U4085 (.a(net42),
    .b(n3131),
    .c(net128),
    .d(net42),
    .out0(n3153));
 b15aoi022aq1n06x5 U4086 (.a(net96),
    .b(n3284),
    .c(net95),
    .d(n3283),
    .o1(n3132));
 b15xor002as1n04x5 U4087 (.a(n3153),
    .b(n3132),
    .out0(n3134));
 b15xor002as1n08x5 U4088 (.a(n3134),
    .b(n3133),
    .out0(n3135));
 b15xor002as1n16x5 U4089 (.a(n3162),
    .b(n3135),
    .out0(n3243));
 b15aboi22an1n04x5 U4090 (.a(net104),
    .b(n3248),
    .c(net104),
    .d(net90),
    .out0(n3136));
 b15xor002as1n04x5 U4091 (.a(n3137),
    .b(n3136),
    .out0(n3139));
 b15xor002aq1n16x5 U4092 (.a(net118),
    .b(net119),
    .out0(n3163));
 b15xor002aq1n08x5 U4093 (.a(n3163),
    .b(net106),
    .out0(n3138));
 b15xor002an1n12x5 U4094 (.a(n3139),
    .b(n3138),
    .out0(n3140));
 b15xor002al1n12x5 U4095 (.a(net45),
    .b(n3140),
    .out0(n3143));
 b15xor002ah1n08x5 U4096 (.a(net103),
    .b(net115),
    .out0(n3141));
 b15xor002as1n16x5 U4097 (.a(n3141),
    .b(net114),
    .out0(n3151));
 b15xor002ar1n12x5 U4098 (.a(net107),
    .b(n3151),
    .out0(n3142));
 b15xor002as1n08x5 U4099 (.a(n3143),
    .b(n3142),
    .out0(n3145));
 b15aoi022ah1n06x5 U4100 (.a(n3257),
    .b(n3146),
    .c(n3243),
    .d(n3145),
    .o1(n3144));
 b15oai122as1n16x5 U4101 (.a(n3144),
    .b(n3257),
    .c(n3146),
    .d(n3243),
    .e(n3145),
    .o1(n3279));
 b15aoi022ah1n16x5 U4102 (.a(net53),
    .b(net52),
    .c(n3282),
    .d(n3147),
    .o1(n3267));
 b15xor002ah1n04x5 U4103 (.a(net122),
    .b(n3267),
    .out0(n3148));
 b15xor002an1n08x5 U4104 (.a(n3148),
    .b(net121),
    .out0(n3271));
 b15aoi022an1n12x5 U4105 (.a(net91),
    .b(net126),
    .c(n3149),
    .d(n3255),
    .o1(n3150));
 b15xor002an1n08x5 U4106 (.a(n3151),
    .b(n3150),
    .out0(n3155));
 b15xor002as1n06x5 U4107 (.a(net110),
    .b(net109),
    .out0(n3152));
 b15xor002ah1n12x5 U4108 (.a(n3152),
    .b(net108),
    .out0(n3268));
 b15xor002al1n08x5 U4109 (.a(n3268),
    .b(n3153),
    .out0(n3154));
 b15xor002as1n08x5 U4110 (.a(n3155),
    .b(n3154),
    .out0(n3156));
 b15ztpn00an1n08x5 PHY_43 ();
 b15nor002ar1n16x5 U4112 (.a(n4146),
    .b(net98),
    .o1(n3456));
 b15nand02as1n48x5 U4113 (.a(net98),
    .b(n4146),
    .o1(n3443));
 b15nanb02ah1n24x5 U4114 (.a(n3456),
    .b(n3443),
    .out0(n3319));
 b15xor002as1n06x5 U4115 (.a(n3311),
    .b(n3319),
    .out0(n3253));
 b15xnr002an1n06x5 U4116 (.a(n3156),
    .b(n3253),
    .out0(n3160));
 b15xor002an1n12x5 U4117 (.a(net123),
    .b(net46),
    .out0(n3158));
 b15xor002an1n12x5 U4118 (.a(net125),
    .b(net117),
    .out0(n3157));
 b15xor002an1n16x5 U4119 (.a(n3158),
    .b(n3157),
    .out0(n3159));
 b15xor002al1n08x5 U4120 (.a(n3160),
    .b(n3159),
    .out0(n3241));
 b15aboi22ah1n04x5 U4121 (.a(net129),
    .b(n4146),
    .c(net707),
    .d(net129),
    .out0(n3171));
 b15aboi22ah1n08x5 U4122 (.a(net124),
    .b(n3254),
    .c(net92),
    .d(net124),
    .out0(n3167));
 b15aboi22as1n16x5 U4123 (.a(net101),
    .b(n3303),
    .c(net100),
    .d(net101),
    .out0(n3161));
 b15qgbxo2an1n05x5 U4124 (.a(n3162),
    .b(n3161),
    .out0(n3165));
 b15xor002as1n12x5 U4125 (.a(net104),
    .b(net112),
    .out0(n3259));
 b15xor002al1n08x5 U4126 (.a(n3163),
    .b(n3259),
    .out0(n3164));
 b15xor002an1n08x5 U4127 (.a(n3165),
    .b(n3164),
    .out0(n3166));
 b15xor002an1n12x5 U4128 (.a(n3167),
    .b(n3166),
    .out0(n3169));
 b15xor002ah1n12x5 U4129 (.a(net111),
    .b(net47),
    .out0(n3168));
 b15xor002ah1n16x5 U4130 (.a(n3169),
    .b(n3168),
    .out0(n3170));
 b15xor002aq1n06x5 U4131 (.a(n3171),
    .b(n3170),
    .out0(n3173));
 b15xor002aq1n08x5 U4132 (.a(net114),
    .b(net108),
    .out0(n3172));
 b15xor002an1n12x5 U4133 (.a(n3173),
    .b(n3172),
    .out0(n3270));
 b15ztpn00an1n08x5 PHY_42 ();
 b15inv040as1n36x5 U4135 (.a(net59),
    .o1(n3814));
 b15oai022ah1n16x5 U4136 (.a(n4116),
    .b(n3814),
    .c(net59),
    .d(net724),
    .o1(n3193));
 b15xor002an1n12x5 U4137 (.a(n4138),
    .b(n3193),
    .out0(n3238));
 b15ztpn00an1n08x5 PHY_41 ();
 b15ztpn00an1n08x5 PHY_40 ();
 b15aoi022aq1n12x5 U4140 (.a(net65),
    .b(net711),
    .c(n4142),
    .d(n4124),
    .o1(n3180));
 b15aoi022aq1n06x5 U4141 (.a(net66),
    .b(net73),
    .c(n4130),
    .d(n4125),
    .o1(n3175));
 b15aoi022ar1n12x5 U4142 (.a(net715),
    .b(net87),
    .c(net692),
    .d(n4131),
    .o1(n3174));
 b15xor002ah1n03x5 U4143 (.a(n3175),
    .b(n3174),
    .out0(n3178));
 b15ztpn00an1n08x5 PHY_39 ();
 b15ztpn00an1n08x5 PHY_38 ();
 b15aoi022ar1n16x5 U4146 (.a(net62),
    .b(net718),
    .c(n4128),
    .d(n4121),
    .o1(n3219));
 b15xor002ah1n06x5 U4147 (.a(n3176),
    .b(n3219),
    .out0(n3177));
 b15xor002as1n06x5 U4148 (.a(n3178),
    .b(n3177),
    .out0(n3179));
 b15xor002as1n12x5 U4149 (.a(n3180),
    .b(n3179),
    .out0(n3182));
 b15xor002as1n16x5 U4150 (.a(net63),
    .b(net83),
    .out0(n3181));
 b15xor002as1n06x5 U4151 (.a(n3182),
    .b(n3181),
    .out0(n3237));
 b15norp02as1n48x5 U4152 (.a(n4134),
    .b(net689),
    .o1(n3825));
 b15oabi12an1n06x5 U4153 (.a(n3825),
    .b(net77),
    .c(net59),
    .out0(n3184));
 b15nandp2aq1n02x5 U4154 (.a(n3184),
    .b(net61),
    .o1(n3183));
 b15oai012aq1n08x5 U4155 (.a(n3183),
    .b(net61),
    .c(n3184),
    .o1(n3185));
 b15xor002an1n08x5 U4156 (.a(net62),
    .b(n3185),
    .out0(n3189));
 b15ztpn00an1n08x5 PHY_37 ();
 b15aoi022an1n12x5 U4158 (.a(net80),
    .b(net711),
    .c(n4142),
    .d(n4137),
    .o1(n3187));
 b15aoi022ar1n24x5 U4159 (.a(net82),
    .b(net713),
    .c(n4135),
    .d(net694),
    .o1(n3186));
 b15xor002ah1n12x5 U4160 (.a(n3187),
    .b(n3186),
    .out0(n3188));
 b15qgbxo2an1n05x5 U4161 (.a(n3189),
    .b(n3188),
    .out0(n3208));
 b15ztpn00an1n08x5 PHY_36 ();
 b15aoi022ah1n12x5 U4163 (.a(net88),
    .b(net89),
    .c(n4145),
    .d(n4144),
    .o1(n3198));
 b15ztpn00an1n08x5 PHY_35 ();
 b15aoi022al1n32x5 U4165 (.a(net84),
    .b(net85),
    .c(n4141),
    .d(n4140),
    .o1(n3220));
 b15xor002ah1n06x5 U4166 (.a(n3198),
    .b(n3220),
    .out0(n3192));
 b15xor002as1n08x5 U4167 (.a(n3190),
    .b(net714),
    .out0(n3191));
 b15xor002as1n12x5 U4168 (.a(n3192),
    .b(n3191),
    .out0(n3207));
 b15xor002ah1n03x5 U4169 (.a(net723),
    .b(n3193),
    .out0(n3206));
 b15ztpn00an1n08x5 PHY_34 ();
 b15oai022al1n32x5 U4171 (.a(n4137),
    .b(net79),
    .c(n4136),
    .d(net80),
    .o1(n3218));
 b15aoi022ah1n08x5 U4172 (.a(net68),
    .b(net69),
    .c(n3818),
    .d(n4127),
    .o1(n3197));
 b15norp02ar1n32x5 U4173 (.a(net695),
    .b(n4124),
    .o1(n3822));
 b15oabi12al1n03x5 U4174 (.a(net670),
    .b(net82),
    .c(net65),
    .out0(n3195));
 b15nand02ar1n02x5 U4175 (.a(n3195),
    .b(net94),
    .o1(n3194));
 b15oai012ah1n03x5 U4176 (.a(n3194),
    .b(net94),
    .c(n3195),
    .o1(n3196));
 b15xor002ah1n03x5 U4177 (.a(n3197),
    .b(n3196),
    .out0(n3200));
 b15xor002as1n03x5 U4178 (.a(net721),
    .b(n3198),
    .out0(n3199));
 b15xor002as1n06x5 U4179 (.a(n3200),
    .b(n3199),
    .out0(n3201));
 b15xor002as1n08x5 U4180 (.a(n3218),
    .b(n3201),
    .out0(n3203));
 b15xor002al1n06x5 U4181 (.a(n3203),
    .b(n3202),
    .out0(n3205));
 b15aoi022al1n02x5 U4182 (.a(n3208),
    .b(n3207),
    .c(n3205),
    .d(n3206),
    .o1(n3204));
 b15oai122an1n08x5 U4183 (.a(n3204),
    .b(n3208),
    .c(n3207),
    .d(n3206),
    .e(n3205),
    .o1(n3235));
 b15aoi022ah1n08x5 U4184 (.a(net85),
    .b(n4128),
    .c(net718),
    .d(n4141),
    .o1(n3233));
 b15aoi022aq1n08x5 U4185 (.a(net79),
    .b(net89),
    .c(n4145),
    .d(n4136),
    .o1(n3210));
 b15aoi022ar1n08x5 U4186 (.a(net66),
    .b(net711),
    .c(n4142),
    .d(n4125),
    .o1(n3209));
 b15xor002ah1n03x5 U4187 (.a(n3210),
    .b(n3209),
    .out0(n3214));
 b15xor002an1n03x5 U4188 (.a(n3212),
    .b(n3211),
    .out0(n3213));
 b15xor002as1n03x5 U4189 (.a(n3214),
    .b(n3213),
    .out0(n3215));
 b15xor002ar1n06x5 U4190 (.a(net116),
    .b(n3215),
    .out0(n3217));
 b15xor002as1n04x5 U4191 (.a(n3217),
    .b(n3216),
    .out0(n3232));
 b15xnr002aq1n16x5 U4192 (.a(net105),
    .b(n3218),
    .out0(n3231));
 b15xor002ah1n03x5 U4193 (.a(n3220),
    .b(n3219),
    .out0(n3224));
 b15xor002as1n03x5 U4194 (.a(n3222),
    .b(n3221),
    .out0(n3223));
 b15xor002an1n06x5 U4195 (.a(n3224),
    .b(n3223),
    .out0(n3226));
 b15xor002aq1n08x5 U4196 (.a(n3226),
    .b(n3225),
    .out0(n3228));
 b15aoi022an1n16x5 U4197 (.a(net722),
    .b(net65),
    .c(n4124),
    .d(n4118),
    .o1(n3227));
 b15xor002an1n16x5 U4198 (.a(n3228),
    .b(n3227),
    .out0(n3230));
 b15aoi022an1n06x5 U4199 (.a(n3232),
    .b(n3233),
    .c(n3230),
    .d(n3231),
    .o1(n3229));
 b15oai122aq1n16x5 U4200 (.a(n3229),
    .b(n3233),
    .c(n3232),
    .d(n3231),
    .e(n3230),
    .o1(n3234));
 b15aoi112ar1n06x5 U4201 (.a(n3235),
    .b(n3234),
    .c(n3238),
    .d(n3237),
    .o1(n3236));
 b15oai012aq1n16x5 U4202 (.a(n3236),
    .b(n3238),
    .c(n3237),
    .o1(n3239));
 b15aoi012ah1n02x5 U4203 (.a(n3239),
    .b(n3270),
    .c(n3241),
    .o1(n3240));
 b15oai012aq1n08x5 U4204 (.a(n3240),
    .b(n3271),
    .c(n3241),
    .o1(n3278));
 b15xnr002ah1n02x5 U4205 (.a(n3243),
    .b(n3242),
    .out0(n3246));
 b15xor002an1n04x5 U4206 (.a(n3267),
    .b(n3244),
    .out0(n3245));
 b15xor002as1n02x5 U4207 (.a(n3246),
    .b(n3245),
    .out0(n3247));
 b15xor002aq1n06x5 U4208 (.a(net127),
    .b(n3247),
    .out0(n3251));
 b15aoi022ah1n16x5 U4209 (.a(net90),
    .b(net93),
    .c(n3249),
    .d(n3248),
    .o1(n3263));
 b15xor002aq1n03x5 U4210 (.a(net100),
    .b(n3263),
    .out0(n3250));
 b15xor002ah1n04x5 U4211 (.a(n3251),
    .b(n3250),
    .out0(n3252));
 b15xor002aq1n08x5 U4212 (.a(n3253),
    .b(n3252),
    .out0(n3276));
 b15aoi022ah1n12x5 U4213 (.a(net92),
    .b(net91),
    .c(n3255),
    .d(n3254),
    .o1(n3275));
 b15qgbxo2an1n10x5 U4214 (.a(n3257),
    .b(n3256),
    .out0(n3261));
 b15xor002an1n12x5 U4215 (.a(n3259),
    .b(n3258),
    .out0(n3260));
 b15xor002al1n12x5 U4216 (.a(n3261),
    .b(n3260),
    .out0(n3262));
 b15xor002al1n04x5 U4217 (.a(n3263),
    .b(n3262),
    .out0(n3265));
 b15xor002as1n12x5 U4218 (.a(net103),
    .b(net138),
    .out0(n3264));
 b15xor002al1n03x5 U4219 (.a(n3265),
    .b(n3264),
    .out0(n3266));
 b15xor002al1n03x5 U4220 (.a(n3267),
    .b(n3266),
    .out0(n3269));
 b15xor002as1n03x5 U4221 (.a(n3269),
    .b(n3268),
    .out0(n3274));
 b15nonb02ar1n03x5 U4222 (.a(n3271),
    .b(n3270),
    .out0(n3272));
 b15oaoi13al1n02x5 U4223 (.a(n3272),
    .b(n3274),
    .c(n3276),
    .d(n3275),
    .o1(n3273));
 b15aoai13as1n04x5 U4224 (.a(n3273),
    .b(n3274),
    .c(n3276),
    .d(n3275),
    .o1(n3277));
 b15nor004as1n12x5 U4225 (.a(n3280),
    .b(n3279),
    .c(n3278),
    .d(n3277),
    .o1(n3348));
 b15norp03al1n08x5 U4226 (.a(net51),
    .b(net42),
    .c(n3281),
    .o1(n3293));
 b15nandp2an1n05x5 U4227 (.a(n3282),
    .b(net53),
    .o1(n3291));
 b15inv040aq1n02x5 U4228 (.a(net39),
    .o1(n3287));
 b15nand03ar1n03x5 U4229 (.a(n3287),
    .b(n3284),
    .c(n3283),
    .o1(n3285));
 b15aoai13ah1n02x5 U4230 (.a(n3285),
    .b(net40),
    .c(net39),
    .d(net95),
    .o1(n3286));
 b15oai013aq1n06x5 U4231 (.a(n3286),
    .b(n3289),
    .c(n3288),
    .d(n3287),
    .o1(n3290));
 b15aoi112ah1n03x5 U4232 (.a(n3291),
    .b(n3290),
    .c(net43),
    .d(net41),
    .o1(n3292));
 b15nand04an1n12x5 U4233 (.a(net44),
    .b(n3348),
    .c(n3293),
    .d(n3292),
    .o1(n3294));
 b15aoi112al1n06x5 U4234 (.a(n3295),
    .b(n3294),
    .c(n3297),
    .d(n3296),
    .o1(n3298));
 b15oai013as1n12x5 U4235 (.a(n3298),
    .b(net43),
    .c(net41),
    .d(n3299),
    .o1(u_reg_u_reg_if_N46));
 b15norp03aq1n08x5 U4236 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .b(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .c(n3350),
    .o1(n3349));
 b15norp02al1n32x5 U4237 (.a(n3308),
    .b(u_reg_u_reg_if_N46),
    .o1(n3821));
 b15aoi013aq1n08x5 U4238 (.a(net2301),
    .b(n3300),
    .c(net724),
    .d(n3821),
    .o1(n3352));
 b15aoi012al1n04x5 U4239 (.a(n3352),
    .b(n3349),
    .c(n3301),
    .o1(gen_alert_tx_0__u_prim_alert_sender_alert_test_set_d));
 b15nandp2al1n48x5 U4240 (.a(n4146),
    .b(n3302),
    .o1(n3920));
 b15nor002an1n24x5 U4241 (.a(n3311),
    .b(n3303),
    .o1(n3444));
 b15qgbin1an1n15x5 U4242 (.a(n3444),
    .o1(n3317));
 b15norp02an1n16x5 U4243 (.a(n3920),
    .b(n3317),
    .o1(n3304));
 b15ztpn00an1n08x5 PHY_33 ();
 b15ztpn00an1n08x5 PHY_32 ();
 b15nandp2ah1n48x5 U4246 (.a(net359),
    .b(net399),
    .o1(n3305));
 b15ztpn00an1n08x5 PHY_31 ();
 b15ztpn00an1n08x5 PHY_30 ();
 b15nand02aq1n48x5 U4249 (.a(n3311),
    .b(net100),
    .o1(n3919));
 b15nor002al1n16x5 U4250 (.a(n3313),
    .b(n3919),
    .o1(n3306));
 b15ztpn00an1n08x5 PHY_29 ();
 b15ztpn00an1n08x5 PHY_28 ();
 b15nand02as1n48x5 U4253 (.a(net358),
    .b(net445),
    .o1(n3307));
 b15ztpn00an1n08x5 PHY_27 ();
 b15ztpn00an1n08x5 PHY_26 ();
 b15nonb02as1n16x5 U4256 (.a(n3308),
    .b(u_reg_u_reg_if_N46),
    .out0(n4024));
 b15and002al1n04x5 U4257 (.a(n3456),
    .b(n3444),
    .o(n3415));
 b15ztpn00an1n08x5 PHY_25 ();
 b15inv000ah1n04x5 U4259 (.a(reg2hw_intr_state__q__15_),
    .o1(n3312));
 b15norp03as1n24x5 U4260 (.a(net99),
    .b(net100),
    .c(n3920),
    .o1(n3309));
 b15ztpn00an1n08x5 PHY_24 ();
 b15ztpn00an1n08x5 PHY_23 ();
 b15norp02ah1n32x5 U4263 (.a(n3443),
    .b(n3919),
    .o1(n3908));
 b15nandp2an1n12x5 U4264 (.a(net430),
    .b(net165),
    .o1(n3840));
 b15nor002as1n32x5 U4265 (.a(net100),
    .b(n3311),
    .o1(n3679));
 b15inv000al1n20x5 U4266 (.a(n3679),
    .o1(n3315));
 b15norp02ah1n48x5 U4267 (.a(n3313),
    .b(n3315),
    .o1(n3909));
 b15nand02aq1n24x5 U4268 (.a(net392),
    .b(net197),
    .o1(n3462));
 b15oai112as1n16x5 U4269 (.a(n3840),
    .b(n3462),
    .c(n3312),
    .d(n4174),
    .o1(n3325));
 b15norp02aq1n24x5 U4270 (.a(n3313),
    .b(n3317),
    .o1(n3314));
 b15ztpn00an1n08x5 PHY_22 ();
 b15ztpn00an1n08x5 PHY_21 ();
 b15ztpn00an1n08x5 PHY_20 ();
 b15ztpn00an1n08x5 PHY_19 ();
 b15aoi022ah1n08x5 U4275 (.a(net596),
    .b(net388),
    .c(net557),
    .d(net396),
    .o1(n3323));
 b15norp02aq1n48x5 U4276 (.a(n3920),
    .b(n3315),
    .o1(n3316));
 b15ztpn00an1n08x5 PHY_18 ();
 b15ztpn00an1n08x5 PHY_17 ();
 b15aoi022ah1n08x5 U4279 (.a(reg2hw_intr_ctrl_en_rising__q__15_),
    .b(net446),
    .c(net375),
    .d(u_reg_data_in_qs[15]),
    .o1(n3322));
 b15norp02aq1n48x5 U4280 (.a(n3919),
    .b(net98),
    .o1(n3915));
 b15norp02ah1n16x5 U4281 (.a(net99),
    .b(net100),
    .o1(n3478));
 b15and002as1n24x5 U4282 (.a(n3478),
    .b(n3456),
    .o(n3413));
 b15ztpn00an1n08x5 PHY_16 ();
 b15aoi022as1n16x5 U4284 (.a(net426),
    .b(net147),
    .c(net423),
    .d(reg2hw_intr_enable__q__15_),
    .o1(n3321));
 b15norp02ah1n32x5 U4285 (.a(n3443),
    .b(n3317),
    .o1(n3318));
 b15ztpn00an1n08x5 PHY_15 ();
 b15ztpn00an1n08x5 PHY_14 ();
 b15nandp2ah1n48x5 U4288 (.a(n3679),
    .b(n3319),
    .o1(n3886));
 b15ztpn00an1n08x5 PHY_13 ();
 b15aoi022aq1n48x5 U4290 (.a(net535),
    .b(net371),
    .c(net179),
    .d(n4176),
    .o1(n3320));
 b15nand04as1n16x5 U4291 (.a(n3323),
    .b(n3322),
    .c(n3321),
    .d(n3320),
    .o1(n3324));
 b15aoi112as1n08x5 U4292 (.a(n3325),
    .b(n3324),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__15_),
    .d(net441),
    .o1(n3326));
 b15nandp2an1n24x5 U4293 (.a(net356),
    .b(n3326),
    .o1(u_reg_u_reg_if_N29));
 b15ztpn00an1n08x5 PHY_12 ();
 b15and002al1n32x5 U4295 (.a(n3915),
    .b(net358),
    .o(N113));
 b15nor002ar1n03x5 U4296 (.a(n4144),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[30]));
 b15ztpn00an1n08x5 PHY_11 ();
 b15nor002ah1n02x5 U4299 (.a(n4144),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[30]));
 b15norp02ar1n04x5 U4300 (.a(n4145),
    .b(n3305),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[31]));
 b15nor002ah1n02x5 U4301 (.a(n4141),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[27]));
 b15nor002al1n03x5 U4302 (.a(n4141),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[27]));
 b15norp02aq1n03x5 U4303 (.a(net693),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[26]));
 b15nor002ar1n03x5 U4304 (.a(n4145),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[31]));
 b15norp02aq1n03x5 U4305 (.a(net693),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[26]));
 b15nor002ah1n04x5 U4306 (.a(n4138),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[24]));
 b15norp02an1n03x5 U4307 (.a(n4138),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[24]));
 b15norp02as1n04x5 U4308 (.a(n4142),
    .b(n3307),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[28]));
 b15nor002ar1n02x5 U4309 (.a(n4142),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[28]));
 b15norp02ar1n03x5 U4310 (.a(net691),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[29]));
 b15norp02an1n02x5 U4311 (.a(net691),
    .b(n3307),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[29]));
 b15nor002an1n03x5 U4312 (.a(net697),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[25]));
 b15norp02aq1n04x5 U4313 (.a(net697),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[25]));
 b15ztpn00an1n08x5 PHY_10 ();
 b15nor002al1n04x5 U4315 (.a(n4133),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[19]));
 b15ztpn00an1n08x5 PHY_9 ();
 b15norp02al1n04x5 U4317 (.a(n4133),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[19]));
 b15nor002an1n04x5 U4319 (.a(n4121),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[6]));
 b15ztpn00an1n08x5 PHY_8 ();
 b15nor002as1n04x5 U4321 (.a(n4117),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[1]));
 b15nor002ar1n06x5 U4322 (.a(n4120),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[5]));
 b15norp02aq1n03x5 U4323 (.a(n4120),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[5]));
 b15nor002al1n04x5 U4324 (.a(n4122),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[7]));
 b15norp02aq1n03x5 U4325 (.a(net704),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[1]));
 b15norp02an1n04x5 U4326 (.a(n4119),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[3]));
 b15nor002an1n04x5 U4327 (.a(n4122),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[7]));
 b15norp02an1n04x5 U4328 (.a(n4119),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[3]));
 b15nor002ah1n06x5 U4329 (.a(n4121),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[6]));
 b15norp02as1n03x5 U4330 (.a(n4116),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[0]));
 b15norp02an1n04x5 U4331 (.a(n4136),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[22]));
 b15norp02an1n03x5 U4332 (.a(n4118),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[2]));
 b15nor002an1n03x5 U4333 (.a(net701),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[15]));
 b15norp02as1n03x5 U4334 (.a(n4137),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[23]));
 b15norp02as1n03x5 U4335 (.a(net700),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[15]));
 b15norp02an1n03x5 U4336 (.a(n4130),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[16]));
 b15nor002an1n03x5 U4337 (.a(n4132),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[18]));
 b15nor002aq1n02x5 U4338 (.a(n4127),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[12]));
 b15nor002ar1n06x5 U4339 (.a(n4127),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[12]));
 b15norp02an1n04x5 U4340 (.a(n4123),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[8]));
 b15nor002aq1n03x5 U4341 (.a(net706),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[0]));
 b15nor002al1n06x5 U4342 (.a(n4123),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[8]));
 b15nor002al1n04x5 U4343 (.a(n4132),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[18]));
 b15norp02aq1n04x5 U4344 (.a(n4137),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[23]));
 b15nor002an1n03x5 U4345 (.a(net702),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[14]));
 b15norp02as1n03x5 U4346 (.a(n4118),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[2]));
 b15nor002as1n02x5 U4347 (.a(n4136),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[22]));
 b15norp02as1n03x5 U4348 (.a(n4126),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[11]));
 b15qgbno2an1n05x5 U4349 (.o1(u_reg_u_intr_ctrl_en_rising_wr_data[16]),
    .a(n4130),
    .b(net346));
 b15nor002as1n04x5 U4350 (.a(n4128),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[14]));
 b15nor002ah1n02x5 U4351 (.a(n4126),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[11]));
 b15norp02as1n04x5 U4352 (.a(n4135),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[21]));
 b15nor002aq1n06x5 U4353 (.a(n4135),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[21]));
 b15norp02al1n02x5 U4354 (.a(net689),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[4]));
 b15nor002ar1n04x5 U4355 (.a(n3814),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[4]));
 b15nor002an1n03x5 U4356 (.a(n3818),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[13]));
 b15norp02al1n04x5 U4357 (.a(n3818),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[13]));
 b15norp02al1n04x5 U4358 (.a(n4125),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[10]));
 b15nor002as1n02x5 U4359 (.a(n4125),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[10]));
 b15nor002ah1n02x5 U4360 (.a(n4131),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[17]));
 b15norp02aq1n03x5 U4361 (.a(n4131),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[17]));
 b15nandp2ar1n24x5 U4363 (.a(net358),
    .b(net439),
    .o1(n3344));
 b15ztpn00an1n08x5 PHY_7 ();
 b15ztpn00an1n08x5 PHY_6 ();
 b15norp02an1n03x5 U4366 (.a(n4133),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[19]));
 b15norp02as1n04x5 U4367 (.a(n4124),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[9]));
 b15norp02aq1n03x5 U4368 (.a(n4124),
    .b(net344),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[9]));
 b15ztpn00an1n08x5 PHY_5 ();
 b15nandp2ah1n48x5 U4370 (.a(net358),
    .b(net420),
    .o1(n3343));
 b15ztpn00an1n08x5 PHY_4 ();
 b15ztpn00an1n08x5 PHY_3 ();
 b15norp02as1n03x5 U4373 (.a(n4133),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[19]));
 b15ztpn00an1n08x5 PHY_2 ();
 b15ztpn00an1n08x5 PHY_1 ();
 b15norp02al1n04x5 U4376 (.a(n4119),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[3]));
 b15ztpn00an1n08x5 PHY_0 ();
 b15norp02an1n04x5 U4379 (.a(n4120),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[5]));
 b15nor002an1n04x5 U4380 (.a(n4120),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[5]));
 b15nor002al1n04x5 U4381 (.a(n4121),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[6]));
 b15nor002ar1n08x5 U4382 (.a(net704),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[1]));
 b15nor002ah1n02x5 U4383 (.a(n4119),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[3]));
 b15nor002ah1n03x5 U4384 (.a(n4122),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[7]));
 b15nor002aq1n03x5 U4385 (.a(n4122),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[7]));
 b15nor002as1n04x5 U4386 (.a(net704),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[1]));
 b15norp02as1n04x5 U4387 (.a(n4121),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[6]));
 b15nor002aq1n03x5 U4388 (.a(net706),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[0]));
 b15norp02al1n03x5 U4389 (.a(net702),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[14]));
 b15qgbno2an1n05x5 U4390 (.o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[8]),
    .a(n4123),
    .b(net338));
 b15nor002an1n03x5 U4391 (.a(net705),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[0]));
 b15norp02ah1n04x5 U4392 (.a(n4126),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[11]));
 b15norp02al1n04x5 U4393 (.a(net701),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[15]));
 b15nor002an1n02x5 U4394 (.a(n4130),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[16]));
 b15nor002al1n03x5 U4395 (.a(n4123),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[8]));
 b15norp02as1n03x5 U4396 (.a(n4127),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[12]));
 b15nor002aq1n03x5 U4397 (.a(n4118),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[2]));
 b15norp02ar1n04x5 U4398 (.a(n4132),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[18]));
 b15norp02ar1n04x5 U4399 (.a(n4127),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[12]));
 b15nor002an1n06x5 U4400 (.a(net699),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[20]));
 b15nor002ar1n04x5 U4401 (.a(n4136),
    .b(n3343),
    .o1(u_reg_u_intr_enable_wr_data[22]));
 b15norp02an1n04x5 U4402 (.a(n4137),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[23]));
 b15nor002ar1n08x5 U4403 (.a(n4130),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[16]));
 b15nor002ah1n02x5 U4404 (.a(n4137),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[23]));
 b15nor002ah1n02x5 U4405 (.a(net703),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[14]));
 b15norp02as1n03x5 U4406 (.a(n4126),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[11]));
 b15nor002an1n03x5 U4407 (.a(n4118),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[2]));
 b15norp02al1n04x5 U4408 (.a(n4132),
    .b(n3344),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[18]));
 b15nor002ah1n02x5 U4409 (.a(n4129),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[15]));
 b15nor002aq1n04x5 U4410 (.a(net698),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[20]));
 b15norp02an1n04x5 U4411 (.a(n4135),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[21]));
 b15norp02ar1n08x5 U4412 (.a(n4136),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[22]));
 b15norp02ah1n03x5 U4413 (.a(n4135),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[21]));
 b15norp02as1n03x5 U4414 (.a(n4125),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[10]));
 b15nor002ar1n06x5 U4415 (.a(net688),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[4]));
 b15norp02as1n03x5 U4416 (.a(n3818),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[13]));
 b15norp02an1n04x5 U4417 (.a(net688),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[4]));
 b15nor002ar1n04x5 U4418 (.a(n4125),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[10]));
 b15norp02aq1n03x5 U4419 (.a(n3818),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[13]));
 b15nor002aq1n02x5 U4420 (.a(n4131),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[17]));
 b15norp02as1n03x5 U4421 (.a(n4131),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[17]));
 b15norp02an1n03x5 U4422 (.a(n4124),
    .b(net337),
    .o1(u_reg_u_intr_enable_wr_data[9]));
 b15nor002ah1n03x5 U4423 (.a(n4124),
    .b(net338),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[9]));
 b15nor002al1n04x5 U4424 (.a(net699),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[20]));
 b15nor002an1n06x5 U4425 (.a(net699),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[20]));
 b15nor002aq1n03x5 U4428 (.a(n4144),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[30]));
 b15nor002ah1n02x5 U4431 (.a(n4144),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[30]));
 b15nor002al1n04x5 U4432 (.a(net693),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[26]));
 b15qgbno2an1n05x5 U4433 (.o1(u_reg_u_intr_enable_wr_data[27]),
    .a(n4141),
    .b(net336));
 b15nor002as1n02x5 U4434 (.a(n4141),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[27]));
 b15norp02aq1n03x5 U4435 (.a(n4145),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[31]));
 b15norp02as1n03x5 U4436 (.a(n4145),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[31]));
 b15norp02as1n03x5 U4437 (.a(net693),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[26]));
 b15nor002aq1n03x5 U4438 (.a(n4138),
    .b(n3344),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[24]));
 b15nor002ah1n04x5 U4439 (.a(n4138),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[24]));
 b15nor002ar1n04x5 U4440 (.a(n4142),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[28]));
 b15nor002as1n03x5 U4441 (.a(n4142),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[28]));
 b15nor002an1n03x5 U4442 (.a(net691),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[29]));
 b15nor002ah1n02x5 U4443 (.a(net690),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[29]));
 b15nor002aq1n03x5 U4444 (.a(net697),
    .b(net339),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[25]));
 b15norp02an1n08x5 U4445 (.a(net697),
    .b(net336),
    .o1(u_reg_u_intr_enable_wr_data[25]));
 b15oabi12as1n16x5 U4446 (.a(net2472),
    .b(n3348),
    .c(n3347),
    .out0(n1439));
 b15orn002aq1n04x5 U4447 (.a(net2238),
    .b(n1439),
    .o(gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger));
 b15oaoi13aq1n08x5 U4448 (.a(n3349),
    .b(n3350),
    .c(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .d(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .o1(n3357));
 b15nor002as1n02x5 U4449 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .b(n3351),
    .o1(n3358));
 b15nonb02al1n12x5 U4450 (.a(n3352),
    .b(gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger),
    .out0(n3360));
 b15aoi013ar1n02x5 U4451 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .b(n3355),
    .c(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .d(gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .o1(n3353));
 b15inv000al1n02x5 U4452 (.a(n3353),
    .o1(n3354));
 b15aoi013ah1n03x5 U4453 (.a(n3354),
    .b(n3358),
    .c(n3360),
    .d(n3355),
    .o1(n3356));
 b15aoi112ar1n06x5 U4454 (.a(n3356),
    .b(n3361),
    .c(gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .d(n3357),
    .o1(gen_alert_tx_0__u_prim_alert_sender_state_d[1]));
 b15nor002an1n02x5 U4455 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .b(n3358),
    .o1(n3359));
 b15oaoi13aq1n08x5 U4456 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .b(n3359),
    .c(gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .d(n3360),
    .o1(n3866));
 b15aoi012an1n02x5 U4457 (.a(n3361),
    .b(n3866),
    .c(n3865),
    .o1(gen_alert_tx_0__u_prim_alert_sender_alert_nd));
 b15aoi022al1n04x5 U4459 (.a(reg2hw_ctrl_en_input_filter__q__11_),
    .b(net386),
    .c(net549),
    .d(net437),
    .o1(n3369));
 b15aoi022as1n08x5 U4461 (.a(net418),
    .b(reg2hw_intr_enable__q__11_),
    .c(net376),
    .d(net2139),
    .o1(n3368));
 b15inv000al1n20x5 U4463 (.a(net638),
    .o1(n3690));
 b15aoi022al1n48x5 U4465 (.a(net435),
    .b(net514),
    .c(net428),
    .d(net661),
    .o1(n3362));
 b15oai012ah1n08x5 U4466 (.a(n3362),
    .b(n3690),
    .c(n3886),
    .o1(n3365));
 b15aoi022aq1n24x5 U4467 (.a(reg2hw_intr_ctrl_en_lvllow__q__11_),
    .b(net372),
    .c(reg2hw_intr_ctrl_en_falling__q__11_),
    .d(net399),
    .o1(n3363));
 b15qgbna2an1n10x5 U4468 (.a(net431),
    .b(net160),
    .o1(n3834));
 b15nandp2an1n08x5 U4469 (.a(net394),
    .b(net192),
    .o1(n3460));
 b15nand04as1n16x5 U4470 (.a(n4024),
    .b(n3363),
    .c(n3834),
    .d(n3460),
    .o1(n3364));
 b15aoi112as1n08x5 U4471 (.a(n3365),
    .b(n3364),
    .c(reg2hw_intr_ctrl_en_rising__q__11_),
    .d(net444),
    .o1(n3367));
 b15nand03as1n06x5 U4472 (.a(n3369),
    .b(net2140),
    .c(n3367),
    .o1(u_reg_u_reg_if_N25));
 b15aoi022ah1n08x5 U4474 (.a(reg2hw_intr_ctrl_en_rising__q__6_),
    .b(net445),
    .c(net381),
    .d(net2103),
    .o1(n3377));
 b15aoi022ar1n32x5 U4475 (.a(reg2hw_intr_ctrl_en_falling__q__6_),
    .b(net399),
    .c(net435),
    .d(net505),
    .o1(n3376));
 b15inv000al1n16x5 U4476 (.a(net614),
    .o1(n3694));
 b15aoi022aq1n32x5 U4477 (.a(net532),
    .b(net368),
    .c(net425),
    .d(net169),
    .o1(n3371));
 b15oai012ar1n12x5 U4478 (.a(n3371),
    .b(n3694),
    .c(n3886),
    .o1(n3374));
 b15aoi022al1n16x5 U4479 (.a(net542),
    .b(net437),
    .c(net419),
    .d(reg2hw_intr_enable__q__6_),
    .o1(n3372));
 b15qgbna2an1n10x5 U4480 (.a(net431),
    .b(net2558),
    .o1(n3848));
 b15nand02as1n08x5 U4481 (.a(net390),
    .b(net2419),
    .o1(n3458));
 b15nand04as1n08x5 U4482 (.a(n4024),
    .b(n3372),
    .c(n3848),
    .d(n3458),
    .o1(n3373));
 b15aoi112aq1n08x5 U4483 (.a(n3374),
    .b(n3373),
    .c(net567),
    .d(net382),
    .o1(n3375));
 b15nandp3aq1n24x5 U4484 (.a(net2104),
    .b(n3376),
    .c(n3375),
    .o1(u_reg_u_reg_if_N20));
 b15aoi022ar1n24x5 U4485 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__8_),
    .b(net437),
    .c(net433),
    .d(reg2hw_intr_state__q__8_),
    .o1(n3384));
 b15aoi022ar1n16x5 U4486 (.a(reg2hw_intr_ctrl_en_rising__q__8_),
    .b(net443),
    .c(reg2hw_intr_ctrl_en_lvllow__q__8_),
    .d(net370),
    .o1(n3383));
 b15inv000ah1n20x5 U4487 (.a(net203),
    .o1(n3804));
 b15aoi022ah1n06x5 U4488 (.a(net418),
    .b(reg2hw_intr_enable__q__8_),
    .c(net376),
    .d(net2275),
    .o1(n3378));
 b15oai012ah1n12x5 U4489 (.a(n3378),
    .b(n3804),
    .c(net366),
    .o1(n3381));
 b15aoi022an1n48x5 U4490 (.a(net564),
    .b(net386),
    .c(net427),
    .d(net171),
    .o1(n3379));
 b15nand02aq1n16x5 U4491 (.a(net431),
    .b(net650),
    .o1(n3850));
 b15nand02aq1n48x5 U4492 (.a(net393),
    .b(net622),
    .o1(n3466));
 b15nand04as1n16x5 U4493 (.a(net357),
    .b(n3379),
    .c(n3850),
    .d(n3466),
    .o1(n3380));
 b15aoi112aq1n08x5 U4494 (.a(n3381),
    .b(n3380),
    .c(reg2hw_intr_ctrl_en_falling__q__8_),
    .d(net396),
    .o1(n3382));
 b15nandp3as1n24x5 U4495 (.a(n3384),
    .b(n3383),
    .c(n3382),
    .o1(u_reg_u_reg_if_N22));
 b15aoi022as1n06x5 U4496 (.a(reg2hw_intr_ctrl_en_rising__q__3_),
    .b(net443),
    .c(net376),
    .d(net2229),
    .o1(n3391));
 b15aoi022an1n12x5 U4497 (.a(net433),
    .b(net509),
    .c(net427),
    .d(net166),
    .o1(n3390));
 b15inv040an1n16x5 U4499 (.a(net198),
    .o1(n3685));
 b15aoi022an1n06x5 U4501 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__3_),
    .b(net437),
    .c(reg2hw_intr_ctrl_en_lvllow__q__3_),
    .d(net371),
    .o1(n3385));
 b15oai012ah1n04x5 U4502 (.a(n3385),
    .b(n3685),
    .c(net366),
    .o1(n3388));
 b15aoi022ah1n08x5 U4503 (.a(net553),
    .b(net396),
    .c(net420),
    .d(reg2hw_intr_enable__q__3_),
    .o1(n3386));
 b15nandp2al1n24x5 U4504 (.a(net430),
    .b(net151),
    .o1(n3836));
 b15nand02an1n32x5 U4505 (.a(net392),
    .b(net630),
    .o1(n3470));
 b15nand04as1n16x5 U4506 (.a(net357),
    .b(n3386),
    .c(n3836),
    .d(n3470),
    .o1(n3387));
 b15aoi112al1n06x5 U4507 (.a(n3388),
    .b(n3387),
    .c(net576),
    .d(net386),
    .o1(n3389));
 b15nand03aq1n16x5 U4508 (.a(n3391),
    .b(n3390),
    .c(n3389),
    .o1(u_reg_u_reg_if_N17));
 b15aoi022ar1n32x5 U4509 (.a(net526),
    .b(net446),
    .c(net426),
    .d(net146),
    .o1(n3398));
 b15aoi022al1n16x5 U4510 (.a(net599),
    .b(net386),
    .c(net423),
    .d(reg2hw_intr_enable__q__14_),
    .o1(n3397));
 b15inv000ar1n20x5 U4511 (.a(net633),
    .o1(n3802));
 b15aoi022as1n02x5 U4512 (.a(reg2hw_intr_ctrl_en_falling__q__14_),
    .b(net396),
    .c(net433),
    .d(reg2hw_intr_state__q__14_),
    .o1(n3392));
 b15oai012al1n08x5 U4513 (.a(n3392),
    .b(n3802),
    .c(net367),
    .o1(n3395));
 b15aoi022al1n24x5 U4514 (.a(net537),
    .b(net370),
    .c(net379),
    .d(u_reg_data_in_qs[14]),
    .o1(n3393));
 b15nandp2an1n08x5 U4515 (.a(net430),
    .b(net164),
    .o1(n3852));
 b15nandp2as1n12x5 U4516 (.a(net392),
    .b(net196),
    .o1(n3468));
 b15nand04as1n16x5 U4517 (.a(net355),
    .b(n3393),
    .c(n3852),
    .d(n3468),
    .o1(n3394));
 b15aoi112as1n08x5 U4518 (.a(n3395),
    .b(n3394),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__14_),
    .d(net439),
    .o1(n3396));
 b15nandp3an1n24x5 U4519 (.a(n3398),
    .b(n3397),
    .c(n3396),
    .o1(u_reg_u_reg_if_N28));
 b15aoi022an1n12x5 U4520 (.a(net603),
    .b(net388),
    .c(net559),
    .d(net396),
    .o1(n3405));
 b15aoi022an1n12x5 U4521 (.a(reg2hw_intr_ctrl_en_rising__q__12_),
    .b(net447),
    .c(reg2hw_intr_ctrl_en_lvllow__q__12_),
    .d(net370),
    .o1(n3404));
 b15inv040al1n12x5 U4522 (.a(net637),
    .o1(n3688));
 b15aoi022al1n32x5 U4523 (.a(net433),
    .b(net513),
    .c(net426),
    .d(net144),
    .o1(n3399));
 b15oai012ah1n06x5 U4524 (.a(n3399),
    .b(n3688),
    .c(net367),
    .o1(n3402));
 b15aoi022ah1n06x5 U4525 (.a(net422),
    .b(net524),
    .c(net374),
    .d(net2100),
    .o1(n3400));
 b15nandp2ah1n16x5 U4526 (.a(net430),
    .b(net161),
    .o1(n3838));
 b15nandp2ar1n24x5 U4527 (.a(net392),
    .b(net193),
    .o1(n3464));
 b15nand04ah1n12x5 U4528 (.a(net355),
    .b(net2101),
    .c(n3838),
    .d(n3464),
    .o1(n3401));
 b15aoi112ah1n08x5 U4529 (.a(n3402),
    .b(n3401),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__12_),
    .d(net441),
    .o1(n3403));
 b15nandp3as1n24x5 U4530 (.a(n3405),
    .b(n3404),
    .c(n3403),
    .o1(u_reg_u_reg_if_N26));
 b15aoi022aq1n12x5 U4531 (.a(net565),
    .b(net385),
    .c(net373),
    .d(net2073),
    .o1(n3412));
 b15aoi022as1n08x5 U4532 (.a(reg2hw_intr_ctrl_en_rising__q__7_),
    .b(net446),
    .c(net436),
    .d(reg2hw_intr_state__q__7_),
    .o1(n3411));
 b15inv000al1n20x5 U4533 (.a(net613),
    .o1(n3806));
 b15aoi022ar1n06x5 U4534 (.a(reg2hw_intr_ctrl_en_falling__q__7_),
    .b(net399),
    .c(net419),
    .d(reg2hw_intr_enable__q__7_),
    .o1(n3406));
 b15oai012aq1n08x5 U4535 (.a(n3406),
    .b(n3806),
    .c(net366),
    .o1(n3409));
 b15aoi022as1n48x5 U4536 (.a(net530),
    .b(net368),
    .c(net425),
    .d(net639),
    .o1(n3407));
 b15nandp2ah1n08x5 U4537 (.a(net431),
    .b(net2050),
    .o1(n3844));
 b15nand02as1n08x5 U4538 (.a(net390),
    .b(net2559),
    .o1(n3472));
 b15nand04as1n16x5 U4539 (.a(net357),
    .b(n3407),
    .c(n3844),
    .d(n3472),
    .o1(n3408));
 b15aoi112an1n08x5 U4540 (.a(n3409),
    .b(n3408),
    .c(net541),
    .d(net437),
    .o1(n3410));
 b15nandp3aq1n24x5 U4541 (.a(net2074),
    .b(n3411),
    .c(n3410),
    .o1(u_reg_u_reg_if_N21));
 b15aoi022aq1n12x5 U4543 (.a(net610),
    .b(net386),
    .c(net418),
    .d(reg2hw_intr_enable__q__1_),
    .o1(n3423));
 b15aoi022al1n24x5 U4544 (.a(net529),
    .b(net443),
    .c(net427),
    .d(net664),
    .o1(n3422));
 b15inv000al1n20x5 U4546 (.a(net184),
    .o1(n3809));
 b15aoi022ar1n04x5 U4547 (.a(reg2hw_intr_ctrl_en_lvllow__q__1_),
    .b(net371),
    .c(net436),
    .d(net517),
    .o1(n3416));
 b15oai012ah1n06x5 U4548 (.a(n3416),
    .b(n3809),
    .c(net366),
    .o1(n3419));
 b15aoi022ah1n08x5 U4549 (.a(net560),
    .b(net396),
    .c(net375),
    .d(net2431),
    .o1(n3417));
 b15nand02al1n16x5 U4550 (.a(net430),
    .b(net149),
    .o1(n3856));
 b15nandp2as1n16x5 U4551 (.a(net392),
    .b(net181),
    .o1(n3756));
 b15nand04as1n16x5 U4552 (.a(net355),
    .b(n3417),
    .c(n3856),
    .d(n3756),
    .o1(n3418));
 b15aoi112ar1n08x5 U4553 (.a(n3419),
    .b(n3418),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__1_),
    .d(net437),
    .o1(n3421));
 b15nand03an1n12x5 U4554 (.a(n3423),
    .b(n3422),
    .c(n3421),
    .o1(u_reg_u_reg_if_N15));
 b15aoi022an1n16x5 U4555 (.a(reg2hw_intr_ctrl_en_rising__q__10_),
    .b(net444),
    .c(reg2hw_intr_ctrl_en_falling__q__10_),
    .d(net399),
    .o1(n3430));
 b15aoi022an1n48x5 U4556 (.a(net539),
    .b(net372),
    .c(net428),
    .d(net142),
    .o1(n3429));
 b15qbfin1bn1n16x5 U4558 (.a(net174),
    .o1(n3697));
 b15aoi022ar1n32x5 U4559 (.a(net419),
    .b(reg2hw_intr_enable__q__10_),
    .c(net376),
    .d(net2315),
    .o1(n3424));
 b15oai012al1n16x5 U4560 (.a(n3424),
    .b(n3697),
    .c(n3886),
    .o1(n3427));
 b15aoi022ar1n32x5 U4561 (.a(reg2hw_ctrl_en_input_filter__q__10_),
    .b(net386),
    .c(net550),
    .d(net437),
    .o1(n3425));
 b15nandp2aq1n24x5 U4562 (.a(net432),
    .b(net647),
    .o1(n3846));
 b15nandp2al1n16x5 U4563 (.a(net390),
    .b(net620),
    .o1(n3751));
 b15nand04as1n06x5 U4564 (.a(n4024),
    .b(n3425),
    .c(n3846),
    .d(n3751),
    .o1(n3426));
 b15aoi112as1n08x5 U4565 (.a(n3427),
    .b(n3426),
    .c(net435),
    .d(net516),
    .o1(n3428));
 b15nandp3aq1n24x5 U4566 (.a(n3430),
    .b(n3429),
    .c(net2316),
    .o1(u_reg_u_reg_if_N24));
 b15aoi022ah1n12x5 U4567 (.a(net569),
    .b(net385),
    .c(reg2hw_intr_ctrl_en_lvllow__q__5_),
    .d(net372),
    .o1(n3439));
 b15aoi022ar1n48x5 U4568 (.a(net435),
    .b(net506),
    .c(net425),
    .d(net641),
    .o1(n3438));
 b15inv040as1n08x5 U4570 (.a(net200),
    .o1(n3692));
 b15aoi022an1n16x5 U4571 (.a(net419),
    .b(net518),
    .c(net376),
    .d(net2191),
    .o1(n3432));
 b15oai012aq1n16x5 U4572 (.a(net2192),
    .b(n3692),
    .c(n3886),
    .o1(n3435));
 b15aoi022aq1n16x5 U4573 (.a(net543),
    .b(net437),
    .c(reg2hw_intr_ctrl_en_rising__q__5_),
    .d(net444),
    .o1(n3433));
 b15nandp2ar1n24x5 U4574 (.a(n3908),
    .b(net154),
    .o1(n3832));
 b15nand02as1n08x5 U4575 (.a(net394),
    .b(net2554),
    .o1(n3474));
 b15nand04as1n16x5 U4576 (.a(net357),
    .b(n3433),
    .c(n3832),
    .d(n3474),
    .o1(n3434));
 b15aoi112as1n08x5 U4577 (.a(n3435),
    .b(n3434),
    .c(reg2hw_intr_ctrl_en_falling__q__5_),
    .d(net399),
    .o1(n3437));
 b15nandp3ah1n12x5 U4578 (.o1(u_reg_u_reg_if_N19),
    .a(n3439),
    .b(n3438),
    .c(net2193));
 b15inv040ar1n02x5 U4579 (.a(n3866),
    .o1(n3441));
 b15nand02an1n02x5 U4580 (.a(n3867),
    .b(n3865),
    .o1(n3440));
 b15oaoi13al1n04x5 U4581 (.a(n3440),
    .b(n3441),
    .c(n3442),
    .d(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .o1(gen_alert_tx_0__u_prim_alert_sender_state_d[0]));
 b15norp02as1n32x5 U4584 (.a(n3443),
    .b(net349),
    .o1(n3680));
 b15nand02ah1n48x5 U4585 (.a(n3680),
    .b(n3444),
    .o1(n3448));
 b15nor002an1n03x5 U4588 (.a(n4133),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[19]));
 b15nor002ar1n03x5 U4591 (.a(n4117),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[1]));
 b15norp02as1n03x5 U4592 (.a(n4119),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[3]));
 b15nor002an1n04x5 U4593 (.a(n4122),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[7]));
 b15nor002ah1n04x5 U4594 (.a(n4120),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[5]));
 b15nor002aq1n04x5 U4595 (.a(n4121),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[6]));
 b15nor002as1n03x5 U4596 (.a(net703),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[14]));
 b15norp02aq1n04x5 U4597 (.a(net706),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[0]));
 b15nor002ar1n06x5 U4598 (.a(n4136),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[22]));
 b15nor002as1n03x5 U4599 (.a(n4123),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[8]));
 b15norp02ah1n04x5 U4600 (.a(n4126),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[11]));
 b15nor002aq1n04x5 U4601 (.a(n4135),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[21]));
 b15nor002aq1n02x5 U4602 (.a(n4130),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[16]));
 b15norp02aq1n03x5 U4603 (.a(n4127),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[12]));
 b15norp02ar1n08x5 U4604 (.a(n4137),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[23]));
 b15nor002ah1n02x5 U4605 (.a(n4132),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[18]));
 b15nor002as1n03x5 U4606 (.a(n4118),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[2]));
 b15nor002as1n03x5 U4607 (.a(net700),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[15]));
 b15norp02aq1n03x5 U4608 (.a(n3818),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[13]));
 b15nor002aq1n04x5 U4609 (.a(net688),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[4]));
 b15nor002as1n03x5 U4610 (.a(n4125),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[10]));
 b15norp02an1n03x5 U4611 (.a(n4131),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[17]));
 b15norp02as1n03x5 U4612 (.a(n4124),
    .b(net313),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[9]));
 b15nor002ah1n02x5 U4615 (.a(n4144),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[30]));
 b15norp02al1n04x5 U4616 (.a(n4145),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[31]));
 b15nor002as1n03x5 U4617 (.a(net698),
    .b(n3448),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[20]));
 b15nor002ah1n02x5 U4618 (.a(n4141),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[27]));
 b15nor002ar1n03x5 U4619 (.a(net693),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[26]));
 b15norp02al1n03x5 U4620 (.a(n4138),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[24]));
 b15norp02ah1n04x5 U4621 (.a(n4142),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[28]));
 b15norp02aq1n48x5 U4622 (.a(net349),
    .b(n4177),
    .o1(u_reg_reg_we_check_15_));
 b15nor002an1n04x5 U4625 (.a(n4144),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[30]));
 b15nor002al1n04x5 U4626 (.a(n4145),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[31]));
 b15nor002aq1n03x5 U4627 (.a(n4141),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[27]));
 b15norp02as1n03x5 U4628 (.a(n4140),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[26]));
 b15norp02ah1n04x5 U4629 (.a(net690),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[29]));
 b15norp02as1n03x5 U4630 (.a(n4138),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[24]));
 b15norp02al1n03x5 U4631 (.a(net697),
    .b(net312),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[25]));
 b15norp02an1n04x5 U4632 (.a(n4142),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[28]));
 b15norp02al1n04x5 U4634 (.a(n4133),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[19]));
 b15norp02as1n03x5 U4636 (.a(n4121),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[6]));
 b15nor002aq1n03x5 U4637 (.a(n4117),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[1]));
 b15nor002aq1n03x5 U4638 (.a(net690),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[29]));
 b15nor002al1n04x5 U4639 (.a(n4120),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[5]));
 b15nor002ah1n03x5 U4640 (.a(n4122),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[7]));
 b15nor002ar1n06x5 U4641 (.a(n4119),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[3]));
 b15nor002aq1n03x5 U4642 (.a(n4139),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[25]));
 b15norp02aq1n04x5 U4643 (.a(net706),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[0]));
 b15nor002al1n06x5 U4644 (.a(n4118),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[2]));
 b15nor002al1n04x5 U4645 (.a(n4126),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[11]));
 b15norp02al1n04x5 U4646 (.a(net700),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[15]));
 b15norp02aq1n04x5 U4647 (.a(n4123),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[8]));
 b15norp02as1n03x5 U4648 (.a(n4128),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[14]));
 b15nor002ar1n04x5 U4649 (.a(n4130),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[16]));
 b15nor002ah1n06x5 U4650 (.a(n4135),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[21]));
 b15nor002as1n03x5 U4651 (.a(n4132),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[18]));
 b15nor002an1n03x5 U4652 (.a(n4137),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[23]));
 b15norp02an1n04x5 U4653 (.a(n4136),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[22]));
 b15nor002ah1n03x5 U4654 (.a(n4127),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[12]));
 b15norp02an1n04x5 U4655 (.a(n4125),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[10]));
 b15norp02as1n03x5 U4656 (.a(net688),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[4]));
 b15nor002aq1n03x5 U4657 (.a(n3818),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[13]));
 b15norp02as1n03x5 U4658 (.a(n4131),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[17]));
 b15nor002ah1n03x5 U4659 (.a(n4124),
    .b(net319),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[9]));
 b15nor002an1n06x5 U4660 (.a(net698),
    .b(net320),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[20]));
 b15nandp2aq1n32x5 U4661 (.a(net358),
    .b(net394),
    .o1(n3749));
 b15nandp2ah1n04x5 U4663 (.a(n3456),
    .b(n3679),
    .o1(n3935));
 b15nor002al1n16x5 U4664 (.a(net349),
    .b(net416),
    .o1(n3754));
 b15aoai13as1n02x5 U4665 (.a(net79),
    .b(net328),
    .c(net331),
    .d(net62),
    .o1(n3457));
 b15oai013ah1n04x5 U4666 (.a(n3457),
    .b(net79),
    .c(net349),
    .d(n3458),
    .o1(N62));
 b15aoai13an1n02x5 U4667 (.a(net85),
    .b(net326),
    .c(net67),
    .d(net331),
    .o1(n3459));
 b15oai013as1n02x5 U4668 (.a(n3459),
    .b(net85),
    .c(net349),
    .d(n3460),
    .o1(N67));
 b15aoai13ah1n02x5 U4669 (.a(net89),
    .b(net329),
    .c(net717),
    .d(n4181),
    .o1(n3461));
 b15oai013aq1n06x5 U4670 (.a(n3461),
    .b(net89),
    .c(net351),
    .d(n3462),
    .o1(N71));
 b15aoai13al1n02x5 U4671 (.a(net86),
    .b(net327),
    .c(net68),
    .d(n4181),
    .o1(n3463));
 b15oai013an1n03x5 U4672 (.a(n3463),
    .b(net86),
    .c(net351),
    .d(n3464),
    .o1(N68));
 b15aoai13an1n06x5 U4673 (.a(net712),
    .b(net329),
    .c(net331),
    .d(net719),
    .o1(n3465));
 b15oai013as1n12x5 U4674 (.a(n3465),
    .b(net712),
    .c(net349),
    .d(n3466),
    .o1(N64));
 b15aoai13al1n02x5 U4675 (.a(net88),
    .b(net327),
    .c(n4181),
    .d(net70),
    .o1(n3467));
 b15oai013ar1n04x5 U4676 (.a(n3467),
    .b(net88),
    .c(net351),
    .d(n3468),
    .o1(N70));
 b15aoai13as1n06x5 U4677 (.a(net714),
    .b(net326),
    .c(net721),
    .d(net331),
    .o1(n3469));
 b15oai013as1n12x5 U4678 (.a(n3469),
    .b(net714),
    .c(net349),
    .d(n3470),
    .o1(N59));
 b15aoai13al1n03x5 U4679 (.a(net80),
    .b(net328),
    .c(net63),
    .d(net331),
    .o1(n3471));
 b15oai013aq1n06x5 U4680 (.a(n3471),
    .b(net80),
    .c(net349),
    .d(n3472),
    .o1(N63));
 b15aoai13ar1n04x5 U4681 (.a(net713),
    .b(net326),
    .c(net720),
    .d(net331),
    .o1(n3473));
 b15oai013ah1n03x5 U4682 (.a(n3473),
    .b(net713),
    .c(net349),
    .d(n3474),
    .o1(N61));
 b15inv040as1n20x5 U4683 (.a(net632),
    .o1(n3934));
 b15aoai13as1n06x5 U4684 (.a(net75),
    .b(net329),
    .c(net722),
    .d(n4181),
    .o1(n3475));
 b15oai013as1n12x5 U4685 (.a(n3475),
    .b(net75),
    .c(n3749),
    .d(net415),
    .o1(N58));
 b15inv040al1n04x5 U4686 (.a(net686),
    .o1(n3477));
 b15nandp2an1n05x5 U4687 (.a(net588),
    .b(gen_filter_19__u_filter_stored_value_q),
    .o1(n3476));
 b15oai012an1n24x5 U4688 (.a(n3476),
    .b(net588),
    .c(n3477),
    .o1(u_reg_u_data_in_wr_data[19]));
 b15nand02ar1n24x5 U4689 (.a(net358),
    .b(net433),
    .o1(n3513));
 b15nonb02ah1n03x5 U4691 (.a(reg2hw_intr_ctrl_en_rising__q__19_),
    .b(net2254),
    .out0(n3481));
 b15aoi012aq1n02x5 U4692 (.a(reg2hw_intr_ctrl_en_lvllow__q__19_),
    .b(net2254),
    .c(reg2hw_intr_ctrl_en_falling__q__19_),
    .o1(n3479));
 b15nandp2aq1n48x5 U4693 (.a(n3478),
    .b(n3680),
    .o1(n3494));
 b15oai022ah1n04x5 U4695 (.a(n3479),
    .b(u_reg_u_data_in_wr_data[19]),
    .c(n4133),
    .d(net307),
    .o1(n3480));
 b15oaoi13as1n08x5 U4696 (.a(n3480),
    .b(u_reg_u_data_in_wr_data[19]),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__19_),
    .d(n3481),
    .o1(n3771));
 b15aboi22ah1n04x5 U4697 (.a(reg2hw_intr_state__q__19_),
    .b(net2255),
    .c(net714),
    .d(n4180),
    .out0(u_reg_u_intr_state_wr_data[19]));
 b15nandp2an1n12x5 U4698 (.a(net575),
    .b(gen_filter_30__u_filter_stored_value_q),
    .o1(n3482));
 b15oai012as1n48x5 U4699 (.a(n3482),
    .b(net574),
    .c(n3483),
    .o1(u_reg_u_data_in_wr_data[30]));
 b15nonb02al1n04x5 U4700 (.a(reg2hw_intr_ctrl_en_rising__q__30_),
    .b(data_in_q[30]),
    .out0(n3486));
 b15aoi012al1n02x5 U4701 (.a(reg2hw_intr_ctrl_en_lvllow__q__30_),
    .b(data_in_q[30]),
    .c(reg2hw_intr_ctrl_en_falling__q__30_),
    .o1(n3484));
 b15oai022ah1n04x5 U4702 (.a(n3484),
    .b(u_reg_u_data_in_wr_data[30]),
    .c(n4144),
    .d(net310),
    .o1(n3485));
 b15oaoi13as1n08x5 U4703 (.a(n3485),
    .b(u_reg_u_data_in_wr_data[30]),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__30_),
    .d(n3486),
    .o1(n3772));
 b15aboi22ar1n12x5 U4704 (.a(reg2hw_intr_state__q__30_),
    .b(n3772),
    .c(net88),
    .d(n4180),
    .out0(u_reg_u_intr_state_wr_data[30]));
 b15aoai13aq1n03x5 U4706 (.a(net331),
    .b(n3825),
    .c(net185),
    .d(net699),
    .o1(n3487));
 b15oai012aq1n03x5 U4707 (.a(n3487),
    .b(n4186),
    .c(net698),
    .o1(N60));
 b15aoai13as1n08x5 U4708 (.a(net330),
    .b(net670),
    .c(net190),
    .d(net696),
    .o1(n3488));
 b15oai012ar1n32x5 U4709 (.a(net306),
    .b(net321),
    .c(net695),
    .o1(N65));
 b15aoai13as1n06x5 U4710 (.a(n4181),
    .b(n3828),
    .c(net616),
    .d(n4143),
    .o1(n3490));
 b15oai012an1n04x5 U4711 (.a(n3490),
    .b(net322),
    .c(n4143),
    .o1(N69));
 b15nandp2aq1n08x5 U4712 (.a(net563),
    .b(net2367),
    .o1(n3491));
 b15oai012as1n32x5 U4713 (.a(n3491),
    .b(net563),
    .c(n3492),
    .o1(u_reg_u_data_in_wr_data[8]));
 b15inv040ar1n02x5 U4717 (.a(data_in_q[8]),
    .o1(n3495));
 b15aoai13as1n04x5 U4718 (.a(u_reg_u_data_in_wr_data[8]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__8_),
    .c(reg2hw_intr_ctrl_en_rising__q__8_),
    .d(n3495),
    .o1(n3498));
 b15inv000al1n02x5 U4719 (.a(u_reg_u_data_in_wr_data[8]),
    .o1(n3496));
 b15aoai13an1n08x5 U4720 (.a(n3496),
    .b(reg2hw_intr_ctrl_en_lvllow__q__8_),
    .c(reg2hw_intr_ctrl_en_falling__q__8_),
    .d(data_in_q[8]),
    .o1(n3497));
 b15oai112as1n16x5 U4721 (.a(n3498),
    .b(n3497),
    .c(net308),
    .d(n4123),
    .o1(n3773));
 b15oa0022al1n03x5 U4722 (.a(n4123),
    .b(net335),
    .c(n3773),
    .d(reg2hw_intr_state__q__8_),
    .o(u_reg_u_intr_state_wr_data[8]));
 b15inv000al1n06x5 U4723 (.a(net679),
    .o1(n3500));
 b15nand02an1n08x5 U4724 (.a(net567),
    .b(net2430),
    .o1(n3499));
 b15oai012ah1n24x5 U4725 (.a(n3499),
    .b(net567),
    .c(n3500),
    .o1(u_reg_u_data_in_wr_data[6]));
 b15inv000an1n02x5 U4726 (.a(data_in_q[6]),
    .o1(n3501));
 b15aoai13an1n06x5 U4727 (.a(u_reg_u_data_in_wr_data[6]),
    .b(net542),
    .c(reg2hw_intr_ctrl_en_rising__q__6_),
    .d(n3501),
    .o1(n3504));
 b15inv000al1n02x5 U4728 (.a(u_reg_u_data_in_wr_data[6]),
    .o1(n3502));
 b15aoai13ar1n08x5 U4729 (.a(n3502),
    .b(net533),
    .c(reg2hw_intr_ctrl_en_falling__q__6_),
    .d(data_in_q[6]),
    .o1(n3503));
 b15oai112as1n16x5 U4730 (.a(n3504),
    .b(n3503),
    .c(net309),
    .d(n4121),
    .o1(n3757));
 b15oa0022al1n04x5 U4731 (.a(n4121),
    .b(net335),
    .c(n3757),
    .d(net2434),
    .o(u_reg_u_intr_state_wr_data[6]));
 b15qbfna2bn1n16x5 U4732 (.a(net606),
    .b(gen_filter_11__u_filter_stored_value_q),
    .o1(n3505));
 b15oai012as1n48x5 U4733 (.a(n3505),
    .b(net606),
    .c(n3506),
    .o1(u_reg_u_data_in_wr_data[11]));
 b15inv000al1n02x5 U4734 (.a(data_in_q[11]),
    .o1(n3507));
 b15aoai13as1n04x5 U4735 (.a(u_reg_u_data_in_wr_data[11]),
    .b(net549),
    .c(reg2hw_intr_ctrl_en_rising__q__11_),
    .d(n3507),
    .o1(n3510));
 b15inv000al1n02x5 U4736 (.a(u_reg_u_data_in_wr_data[11]),
    .o1(n3508));
 b15aoai13ah1n06x5 U4737 (.a(n3508),
    .b(reg2hw_intr_ctrl_en_lvllow__q__11_),
    .c(reg2hw_intr_ctrl_en_falling__q__11_),
    .d(data_in_q[11]),
    .o1(n3509));
 b15oai112as1n16x5 U4738 (.a(n3510),
    .b(n3509),
    .c(net309),
    .d(n4126),
    .o1(n3758));
 b15oa0022ar1n04x5 U4739 (.a(n4126),
    .b(net335),
    .c(n3758),
    .d(reg2hw_intr_state__q__11_),
    .o(u_reg_u_intr_state_wr_data[11]));
 b15inv000aq1n06x5 U4740 (.a(gen_filter_13__u_filter_filter_synced),
    .o1(n3512));
 b15nand02an1n12x5 U4741 (.a(net601),
    .b(gen_filter_13__u_filter_stored_value_q),
    .o1(n3511));
 b15oai012as1n32x5 U4742 (.a(n3511),
    .b(net601),
    .c(n3512),
    .o1(u_reg_u_data_in_wr_data[13]));
 b15inv000as1n02x5 U4745 (.a(data_in_q[13]),
    .o1(n3515));
 b15aoai13ar1n08x5 U4746 (.a(u_reg_u_data_in_wr_data[13]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__13_),
    .c(net528),
    .d(n3515),
    .o1(n3518));
 b15inv000al1n02x5 U4747 (.a(u_reg_u_data_in_wr_data[13]),
    .o1(n3516));
 b15aoai13as1n04x5 U4748 (.a(n3516),
    .b(net538),
    .c(net558),
    .d(net2243),
    .o1(n3517));
 b15oai112as1n12x5 U4749 (.a(n3518),
    .b(n3517),
    .c(net308),
    .d(n3818),
    .o1(n3785));
 b15oa0022al1n02x5 U4750 (.a(n3818),
    .b(net335),
    .c(net2244),
    .d(reg2hw_intr_state__q__13_),
    .o(u_reg_u_intr_state_wr_data[13]));
 b15nand02al1n12x5 U4751 (.a(net608),
    .b(gen_filter_10__u_filter_stored_value_q),
    .o1(n3519));
 b15oai012an1n32x5 U4752 (.a(n3519),
    .b(net608),
    .c(n3520),
    .o1(u_reg_u_data_in_wr_data[10]));
 b15inv020ar1n04x5 U4753 (.a(data_in_q[10]),
    .o1(n3521));
 b15aoai13al1n08x5 U4754 (.a(u_reg_u_data_in_wr_data[10]),
    .b(net550),
    .c(reg2hw_intr_ctrl_en_rising__q__10_),
    .d(n3521),
    .o1(n3524));
 b15inv040ar1n02x5 U4755 (.a(u_reg_u_data_in_wr_data[10]),
    .o1(n3522));
 b15aoai13ah1n06x5 U4756 (.a(n3522),
    .b(reg2hw_intr_ctrl_en_lvllow__q__10_),
    .c(reg2hw_intr_ctrl_en_falling__q__10_),
    .d(data_in_q[10]),
    .o1(n3523));
 b15oai112as1n16x5 U4757 (.a(n3524),
    .b(n3523),
    .c(net309),
    .d(n4125),
    .o1(n3761));
 b15oa0022ah1n02x5 U4758 (.a(n4125),
    .b(net335),
    .c(n3761),
    .d(net2438),
    .o(u_reg_u_intr_state_wr_data[10]));
 b15nand02aq1n12x5 U4759 (.a(net598),
    .b(gen_filter_14__u_filter_stored_value_q),
    .o1(n3525));
 b15oai012ar1n48x5 U4760 (.a(n3525),
    .b(net598),
    .c(n3526),
    .o1(u_reg_u_data_in_wr_data[14]));
 b15inv000al1n02x5 U4761 (.a(net2331),
    .o1(n3527));
 b15aoai13ah1n03x5 U4762 (.a(u_reg_u_data_in_wr_data[14]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__14_),
    .c(reg2hw_intr_ctrl_en_rising__q__14_),
    .d(n3527),
    .o1(n3530));
 b15inv000al1n02x5 U4763 (.a(u_reg_u_data_in_wr_data[14]),
    .o1(n3528));
 b15aoai13an1n04x5 U4764 (.a(n3528),
    .b(net537),
    .c(reg2hw_intr_ctrl_en_falling__q__14_),
    .d(net2331),
    .o1(n3529));
 b15oai112an1n16x5 U4765 (.a(n3530),
    .b(n3529),
    .c(net308),
    .d(net702),
    .o1(n3782));
 b15oa0022al1n03x5 U4766 (.a(net702),
    .b(net335),
    .c(n3782),
    .d(reg2hw_intr_state__q__14_),
    .o(u_reg_u_intr_state_wr_data[14]));
 b15inv040aq1n05x5 U4767 (.a(net681),
    .o1(n3532));
 b15nand02ar1n16x5 U4768 (.a(net568),
    .b(gen_filter_5__u_filter_stored_value_q),
    .o1(n3531));
 b15oai012ah1n32x5 U4769 (.a(n3531),
    .b(net568),
    .c(n3532),
    .o1(u_reg_u_data_in_wr_data[5]));
 b15inv020aq1n03x5 U4770 (.a(data_in_q[5]),
    .o1(n3533));
 b15aoai13ah1n06x5 U4771 (.a(u_reg_u_data_in_wr_data[5]),
    .b(net543),
    .c(reg2hw_intr_ctrl_en_rising__q__5_),
    .d(n3533),
    .o1(n3536));
 b15inv040al1n02x5 U4772 (.a(u_reg_u_data_in_wr_data[5]),
    .o1(n3534));
 b15aoai13al1n08x5 U4773 (.a(n3534),
    .b(reg2hw_intr_ctrl_en_lvllow__q__5_),
    .c(reg2hw_intr_ctrl_en_falling__q__5_),
    .d(data_in_q[5]),
    .o1(n3535));
 b15oai112as1n16x5 U4774 (.a(n3536),
    .b(n3535),
    .c(net309),
    .d(n4120),
    .o1(n3778));
 b15oa0022ah1n04x5 U4775 (.a(n4120),
    .b(net334),
    .c(n3778),
    .d(net2464),
    .o(u_reg_u_intr_state_wr_data[5]));
 b15inv000as1n03x5 U4776 (.a(gen_filter_21__u_filter_filter_synced),
    .o1(n3538));
 b15nandp2an1n05x5 U4777 (.a(net587),
    .b(net2234),
    .o1(n3537));
 b15oai012ah1n16x5 U4778 (.a(n3537),
    .b(net587),
    .c(n3538),
    .o1(u_reg_u_data_in_wr_data[21]));
 b15inv020ah1n03x5 U4779 (.a(data_in_q[21]),
    .o1(n3539));
 b15aoai13as1n08x5 U4780 (.a(u_reg_u_data_in_wr_data[21]),
    .b(net546),
    .c(reg2hw_intr_ctrl_en_rising__q__21_),
    .d(n3539),
    .o1(n3542));
 b15inv000an1n02x5 U4781 (.a(u_reg_u_data_in_wr_data[21]),
    .o1(n3540));
 b15aoai13as1n08x5 U4782 (.a(n3540),
    .b(reg2hw_intr_ctrl_en_lvllow__q__21_),
    .c(reg2hw_intr_ctrl_en_falling__q__21_),
    .d(data_in_q[21]),
    .o1(n3541));
 b15oai112as1n16x5 U4783 (.a(n3542),
    .b(n3541),
    .c(net307),
    .d(n4135),
    .o1(n3765));
 b15oa0022an1n03x5 U4784 (.a(n4135),
    .b(net334),
    .c(n3765),
    .d(reg2hw_intr_state__q__21_),
    .o(u_reg_u_intr_state_wr_data[21]));
 b15inv020ah1n06x5 U4785 (.a(gen_filter_15__u_filter_filter_synced),
    .o1(n3544));
 b15nand02aq1n08x5 U4786 (.a(net597),
    .b(net2449),
    .o1(n3543));
 b15oai012an1n32x5 U4787 (.a(n3543),
    .b(net597),
    .c(n3544),
    .o1(u_reg_u_data_in_wr_data[15]));
 b15inv000al1n02x5 U4788 (.a(net2223),
    .o1(n3545));
 b15aoai13as1n04x5 U4789 (.a(u_reg_u_data_in_wr_data[15]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__15_),
    .c(reg2hw_intr_ctrl_en_rising__q__15_),
    .d(n3545),
    .o1(n3548));
 b15inv000al1n02x5 U4790 (.a(u_reg_u_data_in_wr_data[15]),
    .o1(n3546));
 b15aoai13as1n06x5 U4791 (.a(n3546),
    .b(net536),
    .c(net557),
    .d(net2223),
    .o1(n3547));
 b15oai112aq1n16x5 U4792 (.a(n3548),
    .b(n3547),
    .c(net308),
    .d(n4129),
    .o1(n3774));
 b15oa0022ah1n02x5 U4793 (.a(n4129),
    .b(net335),
    .c(n3774),
    .d(reg2hw_intr_state__q__15_),
    .o(u_reg_u_intr_state_wr_data[15]));
 b15inv040ah1n04x5 U4794 (.a(gen_filter_0__u_filter_filter_synced),
    .o1(n3550));
 b15nandp2aq1n02x5 U4795 (.a(reg2hw_ctrl_en_input_filter__q__0_),
    .b(gen_filter_0__u_filter_stored_value_q),
    .o1(n3549));
 b15oai012al1n06x5 U4796 (.a(n3549),
    .b(reg2hw_ctrl_en_input_filter__q__0_),
    .c(n3550),
    .o1(u_reg_u_data_in_wr_data[0]));
 b15inv000as1n03x5 U4797 (.a(data_in_q[0]),
    .o1(n3551));
 b15aoai13as1n08x5 U4798 (.a(net365),
    .b(net551),
    .c(reg2hw_intr_ctrl_en_rising__q__0_),
    .d(n3551),
    .o1(n3554));
 b15inv000aq1n02x5 U4799 (.a(net365),
    .o1(n3552));
 b15aoai13as1n08x5 U4800 (.a(n3552),
    .b(reg2hw_intr_ctrl_en_lvllow__q__0_),
    .c(net562),
    .d(data_in_q[0]),
    .o1(n3553));
 b15oai112as1n16x5 U4801 (.a(n3554),
    .b(n3553),
    .c(net308),
    .d(net705),
    .o1(n3781));
 b15oa0022ar1n03x5 U4802 (.a(net705),
    .b(net335),
    .c(n3781),
    .d(reg2hw_intr_state__q__0_),
    .o(u_reg_u_intr_state_wr_data[0]));
 b15nand02al1n06x5 U4803 (.a(net590),
    .b(net2246),
    .o1(n3555));
 b15oai012al1n16x5 U4804 (.a(n3555),
    .b(net590),
    .c(n3556),
    .o1(u_reg_u_data_in_wr_data[18]));
 b15inv000as1n02x5 U4805 (.a(data_in_q[18]),
    .o1(n3557));
 b15aoai13as1n06x5 U4806 (.a(u_reg_u_data_in_wr_data[18]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__18_),
    .c(reg2hw_intr_ctrl_en_rising__q__18_),
    .d(n3557),
    .o1(n3560));
 b15inv000al1n02x5 U4807 (.a(u_reg_u_data_in_wr_data[18]),
    .o1(n3558));
 b15aoai13al1n08x5 U4808 (.a(n3558),
    .b(reg2hw_intr_ctrl_en_lvllow__q__18_),
    .c(net556),
    .d(net2284),
    .o1(n3559));
 b15oai112as1n16x5 U4809 (.a(n3560),
    .b(n3559),
    .c(net307),
    .d(n4132),
    .o1(n3786));
 b15oa0022ah1n02x5 U4810 (.a(n4132),
    .b(net334),
    .c(net2285),
    .d(reg2hw_intr_state__q__18_),
    .o(u_reg_u_intr_state_wr_data[18]));
 b15inv000an1n05x5 U4811 (.a(gen_filter_16__u_filter_filter_synced),
    .o1(n3562));
 b15nandp2as1n04x5 U4812 (.a(net594),
    .b(net2264),
    .o1(n3561));
 b15oai012an1n24x5 U4813 (.a(n3561),
    .b(net594),
    .c(n3562),
    .o1(u_reg_u_data_in_wr_data[16]));
 b15inv040ar1n02x5 U4814 (.a(data_in_q[16]),
    .o1(n3563));
 b15aoai13an1n06x5 U4815 (.a(u_reg_u_data_in_wr_data[16]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__16_),
    .c(reg2hw_intr_ctrl_en_rising__q__16_),
    .d(n3563),
    .o1(n3566));
 b15inv000al1n02x5 U4816 (.a(u_reg_u_data_in_wr_data[16]),
    .o1(n3564));
 b15aoai13ah1n04x5 U4817 (.a(n3564),
    .b(reg2hw_intr_ctrl_en_lvllow__q__16_),
    .c(reg2hw_intr_ctrl_en_falling__q__16_),
    .d(net2475),
    .o1(n3565));
 b15oai112as1n16x5 U4818 (.a(n3566),
    .b(n3565),
    .c(net307),
    .d(n4130),
    .o1(n3762));
 b15oa0022an1n02x5 U4819 (.a(n4130),
    .b(net334),
    .c(n3762),
    .d(reg2hw_intr_state__q__16_),
    .o(u_reg_u_intr_state_wr_data[16]));
 b15nandp2aq1n02x5 U4820 (.a(net566),
    .b(gen_filter_7__u_filter_stored_value_q),
    .o1(n3567));
 b15oai012al1n06x5 U4821 (.a(n3567),
    .b(net566),
    .c(n3568),
    .o1(u_reg_u_data_in_wr_data[7]));
 b15inv040al1n02x5 U4822 (.a(data_in_q[7]),
    .o1(n3569));
 b15aoai13as1n06x5 U4823 (.a(net364),
    .b(net541),
    .c(reg2hw_intr_ctrl_en_rising__q__7_),
    .d(n3569),
    .o1(n3572));
 b15inv040al1n02x5 U4824 (.a(net364),
    .o1(n3570));
 b15aoai13as1n08x5 U4825 (.a(n3570),
    .b(reg2hw_intr_ctrl_en_lvllow__q__7_),
    .c(reg2hw_intr_ctrl_en_falling__q__7_),
    .d(data_in_q[7]),
    .o1(n3571));
 b15oai112as1n16x5 U4826 (.a(n3572),
    .b(n3571),
    .c(net311),
    .d(n4122),
    .o1(n3787));
 b15oa0022as1n02x5 U4827 (.a(n4122),
    .b(net334),
    .c(n3787),
    .d(reg2hw_intr_state__q__7_),
    .o(u_reg_u_intr_state_wr_data[7]));
 b15inv040as1n02x5 U4828 (.a(gen_filter_28__u_filter_filter_synced),
    .o1(n3574));
 b15nandp2an1n04x5 U4829 (.a(net579),
    .b(net2465),
    .o1(n3573));
 b15oai012ah1n12x5 U4830 (.a(n3573),
    .b(net579),
    .c(n3574),
    .o1(u_reg_u_data_in_wr_data[28]));
 b15inv000ar1n03x5 U4832 (.a(data_in_q[28]),
    .o1(n3576));
 b15aoai13as1n06x5 U4833 (.a(u_reg_u_data_in_wr_data[28]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__28_),
    .c(reg2hw_intr_ctrl_en_rising__q__28_),
    .d(n3576),
    .o1(n3579));
 b15inv000al1n02x5 U4834 (.a(u_reg_u_data_in_wr_data[28]),
    .o1(n3577));
 b15aoai13al1n08x5 U4835 (.a(n3577),
    .b(reg2hw_intr_ctrl_en_lvllow__q__28_),
    .c(reg2hw_intr_ctrl_en_falling__q__28_),
    .d(data_in_q[28]),
    .o1(n3578));
 b15oai112as1n16x5 U4836 (.a(n3579),
    .b(n3578),
    .c(net310),
    .d(n4142),
    .o1(n3766));
 b15oa0022aq1n02x5 U4837 (.a(n4142),
    .b(n3513),
    .c(n3766),
    .d(reg2hw_intr_state__q__28_),
    .o(u_reg_u_intr_state_wr_data[28]));
 b15inv020as1n08x5 U4838 (.a(gen_filter_3__u_filter_filter_synced),
    .o1(n3581));
 b15nandp2al1n12x5 U4839 (.a(net577),
    .b(gen_filter_3__u_filter_stored_value_q),
    .o1(n3580));
 b15oai012an1n48x5 U4840 (.a(n3580),
    .b(net577),
    .c(n3581),
    .o1(u_reg_u_data_in_wr_data[3]));
 b15inv040ar1n03x5 U4841 (.a(data_in_q[3]),
    .o1(n3582));
 b15aoai13al1n08x5 U4842 (.a(u_reg_u_data_in_wr_data[3]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__3_),
    .c(reg2hw_intr_ctrl_en_rising__q__3_),
    .d(n3582),
    .o1(n3585));
 b15inv000al1n02x5 U4843 (.a(u_reg_u_data_in_wr_data[3]),
    .o1(n3583));
 b15aoai13al1n08x5 U4844 (.a(n3583),
    .b(reg2hw_intr_ctrl_en_lvllow__q__3_),
    .c(net553),
    .d(data_in_q[3]),
    .o1(n3584));
 b15oai112as1n16x5 U4845 (.a(n3585),
    .b(n3584),
    .c(net308),
    .d(n4119),
    .o1(n3783));
 b15oa0022as1n02x5 U4846 (.a(n4119),
    .b(net335),
    .c(n3783),
    .d(net509),
    .o(u_reg_u_intr_state_wr_data[3]));
 b15inv020ah1n16x5 U4847 (.a(reg2hw_ctrl_en_input_filter__q__2_),
    .o1(n3884));
 b15nand02ah1n06x5 U4848 (.a(reg2hw_ctrl_en_input_filter__q__2_),
    .b(net2481),
    .o1(n3586));
 b15aob012as1n24x5 U4849 (.a(n3586),
    .b(n3884),
    .c(gen_filter_2__u_filter_filter_synced),
    .out0(u_reg_u_data_in_wr_data[2]));
 b15inv000ah1n02x5 U4850 (.a(data_in_q[2]),
    .o1(n3587));
 b15aoai13ar1n08x5 U4851 (.a(u_reg_u_data_in_wr_data[2]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__2_),
    .c(reg2hw_intr_ctrl_en_rising__q__2_),
    .d(n3587),
    .o1(n3590));
 b15inv020an1n03x5 U4852 (.a(u_reg_u_data_in_wr_data[2]),
    .o1(n3588));
 b15aoai13ah1n08x5 U4853 (.a(n3588),
    .b(reg2hw_intr_ctrl_en_lvllow__q__2_),
    .c(net554),
    .d(data_in_q[2]),
    .o1(n3589));
 b15oai112as1n16x5 U4854 (.a(n3590),
    .b(n3589),
    .c(net311),
    .d(n4118),
    .o1(n3767));
 b15oa0022al1n03x5 U4855 (.a(n4118),
    .b(net335),
    .c(n3767),
    .d(reg2hw_intr_state__q__2_),
    .o(u_reg_u_intr_state_wr_data[2]));
 b15nand02aq1n16x5 U4856 (.a(reg2hw_ctrl_en_input_filter__q__1_),
    .b(gen_filter_1__u_filter_stored_value_q),
    .o1(n3591));
 b15oai012ah1n48x5 U4857 (.a(n3591),
    .b(net609),
    .c(n3592),
    .o1(u_reg_u_data_in_wr_data[1]));
 b15inv040aq1n02x5 U4858 (.a(data_in_q[1]),
    .o1(n3593));
 b15aoai13an1n08x5 U4859 (.a(u_reg_u_data_in_wr_data[1]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__1_),
    .c(net529),
    .d(n3593),
    .o1(n3596));
 b15inv000al1n02x5 U4860 (.a(u_reg_u_data_in_wr_data[1]),
    .o1(n3594));
 b15aoai13as1n06x5 U4861 (.a(n3594),
    .b(reg2hw_intr_ctrl_en_lvllow__q__1_),
    .c(net561),
    .d(data_in_q[1]),
    .o1(n3595));
 b15oai112as1n16x5 U4862 (.a(n3596),
    .b(n3595),
    .c(net308),
    .d(net704),
    .o1(n3779));
 b15oa0022ah1n03x5 U4863 (.a(net704),
    .b(net335),
    .c(n3779),
    .d(net2391),
    .o(u_reg_u_intr_state_wr_data[1]));
 b15qgbna2an1n10x5 U4864 (.a(net572),
    .b(gen_filter_4__u_filter_stored_value_q),
    .o1(n3597));
 b15oai012ah1n32x5 U4865 (.a(n3597),
    .b(net572),
    .c(n3598),
    .o1(u_reg_u_data_in_wr_data[4]));
 b15inv000as1n03x5 U4866 (.a(data_in_q[4]),
    .o1(n3599));
 b15aoai13ah1n06x5 U4867 (.a(u_reg_u_data_in_wr_data[4]),
    .b(net544),
    .c(reg2hw_intr_ctrl_en_rising__q__4_),
    .d(n3599),
    .o1(n3602));
 b15inv000aq1n02x5 U4868 (.a(u_reg_u_data_in_wr_data[4]),
    .o1(n3600));
 b15aoai13aq1n08x5 U4869 (.a(n3600),
    .b(reg2hw_intr_ctrl_en_lvllow__q__4_),
    .c(reg2hw_intr_ctrl_en_falling__q__4_),
    .d(data_in_q[4]),
    .o1(n3601));
 b15oai112as1n16x5 U4870 (.a(n3602),
    .b(n3601),
    .c(net309),
    .d(net689),
    .o1(n3795));
 b15oa0022ar1n06x5 U4871 (.a(net689),
    .b(net334),
    .c(n3795),
    .d(reg2hw_intr_state__q__4_),
    .o(u_reg_u_intr_state_wr_data[4]));
 b15inv000an1n04x5 U4872 (.a(gen_filter_27__u_filter_filter_synced),
    .o1(n3604));
 b15qgbna2an1n05x5 U4873 (.o1(n3603),
    .a(reg2hw_ctrl_en_input_filter__q__27_),
    .b(net2268));
 b15oai012ah1n16x5 U4874 (.a(n3603),
    .b(reg2hw_ctrl_en_input_filter__q__27_),
    .c(n3604),
    .o1(u_reg_u_data_in_wr_data[27]));
 b15inv000al1n02x5 U4875 (.a(data_in_q[27]),
    .o1(n3605));
 b15aoai13as1n04x5 U4876 (.a(u_reg_u_data_in_wr_data[27]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__27_),
    .c(net525),
    .d(n3605),
    .o1(n3608));
 b15inv000al1n02x5 U4877 (.a(u_reg_u_data_in_wr_data[27]),
    .o1(n3606));
 b15aoai13as1n04x5 U4878 (.a(n3606),
    .b(reg2hw_intr_ctrl_en_lvllow__q__27_),
    .c(net555),
    .d(data_in_q[27]),
    .o1(n3607));
 b15oai112as1n16x5 U4879 (.a(n3608),
    .b(n3607),
    .c(net311),
    .d(n4141),
    .o1(n3763));
 b15oa0022aq1n03x5 U4880 (.a(n4141),
    .b(net334),
    .c(n3763),
    .d(reg2hw_intr_state__q__27_),
    .o(u_reg_u_intr_state_wr_data[27]));
 b15inv040aq1n03x5 U4881 (.a(gen_filter_23__u_filter_filter_synced),
    .o1(n3610));
 b15nand02an1n06x5 U4882 (.a(net584),
    .b(net2230),
    .o1(n3609));
 b15oai012as1n16x5 U4883 (.a(n3609),
    .b(net584),
    .c(n3610),
    .o1(u_reg_u_data_in_wr_data[23]));
 b15inv040ar1n03x5 U4884 (.a(data_in_q[23]),
    .o1(n3611));
 b15aoai13al1n08x5 U4885 (.a(u_reg_u_data_in_wr_data[23]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__23_),
    .c(reg2hw_intr_ctrl_en_rising__q__23_),
    .d(n3611),
    .o1(n3614));
 b15inv000al1n02x5 U4886 (.a(u_reg_u_data_in_wr_data[23]),
    .o1(n3612));
 b15aoai13ar1n08x5 U4887 (.a(n3612),
    .b(reg2hw_intr_ctrl_en_lvllow__q__23_),
    .c(reg2hw_intr_ctrl_en_falling__q__23_),
    .d(data_in_q[23]),
    .o1(n3613));
 b15oai112as1n16x5 U4888 (.a(n3614),
    .b(n3613),
    .c(n3494),
    .d(n4137),
    .o1(n3759));
 b15oa0022aq1n02x5 U4889 (.a(n4137),
    .b(net335),
    .c(n3759),
    .d(reg2hw_intr_state__q__23_),
    .o(u_reg_u_intr_state_wr_data[23]));
 b15inv000al1n12x5 U4890 (.a(gen_filter_31__u_filter_filter_synced),
    .o1(n3616));
 b15nandp2ar1n12x5 U4891 (.a(reg2hw_ctrl_en_input_filter__q__31_),
    .b(gen_filter_31__u_filter_stored_value_q),
    .o1(n3615));
 b15oai012as1n32x5 U4892 (.a(n3615),
    .b(reg2hw_ctrl_en_input_filter__q__31_),
    .c(n3616),
    .o1(u_reg_u_data_in_wr_data[31]));
 b15inv000al1n02x5 U4893 (.a(data_in_q[31]),
    .o1(n3617));
 b15aoai13as1n04x5 U4894 (.a(u_reg_u_data_in_wr_data[31]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__31_),
    .c(reg2hw_intr_ctrl_en_rising__q__31_),
    .d(n3617),
    .o1(n3620));
 b15inv000al1n02x5 U4895 (.a(u_reg_u_data_in_wr_data[31]),
    .o1(n3618));
 b15aoai13an1n06x5 U4896 (.a(n3618),
    .b(reg2hw_intr_ctrl_en_lvllow__q__31_),
    .c(reg2hw_intr_ctrl_en_falling__q__31_),
    .d(data_in_q[31]),
    .o1(n3619));
 b15oai112as1n16x5 U4897 (.a(n3620),
    .b(n3619),
    .c(net310),
    .d(n4145),
    .o1(n3780));
 b15oa0022an1n02x5 U4898 (.a(n4145),
    .b(net334),
    .c(n3780),
    .d(reg2hw_intr_state__q__31_),
    .o(u_reg_u_intr_state_wr_data[31]));
 b15inv020an1n06x5 U4899 (.a(gen_filter_17__u_filter_filter_synced),
    .o1(n3622));
 b15nand02aq1n04x5 U4900 (.a(net592),
    .b(gen_filter_17__u_filter_stored_value_q),
    .o1(n3621));
 b15oai012al1n16x5 U4901 (.a(n3621),
    .b(net592),
    .c(n3622),
    .o1(u_reg_u_data_in_wr_data[17]));
 b15inv000al1n02x5 U4902 (.a(data_in_q[17]),
    .o1(n3623));
 b15aoai13aq1n04x5 U4903 (.a(u_reg_u_data_in_wr_data[17]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__17_),
    .c(reg2hw_intr_ctrl_en_rising__q__17_),
    .d(n3623),
    .o1(n3626));
 b15inv000al1n02x5 U4904 (.a(u_reg_u_data_in_wr_data[17]),
    .o1(n3624));
 b15aoai13an1n06x5 U4905 (.a(n3624),
    .b(reg2hw_intr_ctrl_en_lvllow__q__17_),
    .c(reg2hw_intr_ctrl_en_falling__q__17_),
    .d(data_in_q[17]),
    .o1(n3625));
 b15oai112aq1n16x5 U4906 (.a(n3626),
    .b(n3625),
    .c(net308),
    .d(n4131),
    .o1(n3775));
 b15oa0022ar1n04x5 U4907 (.a(n4131),
    .b(net335),
    .c(n3775),
    .d(reg2hw_intr_state__q__17_),
    .o(u_reg_u_intr_state_wr_data[17]));
 b15nand02ar1n16x5 U4908 (.a(net604),
    .b(gen_filter_12__u_filter_stored_value_q),
    .o1(n3627));
 b15oai012ar1n48x5 U4909 (.a(n3627),
    .b(net604),
    .c(n3628),
    .o1(u_reg_u_data_in_wr_data[12]));
 b15inv000aq1n02x5 U4910 (.a(net2263),
    .o1(n3629));
 b15aoai13ah1n06x5 U4911 (.a(u_reg_u_data_in_wr_data[12]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__12_),
    .c(reg2hw_intr_ctrl_en_rising__q__12_),
    .d(n3629),
    .o1(n3632));
 b15inv000al1n02x5 U4912 (.a(u_reg_u_data_in_wr_data[12]),
    .o1(n3630));
 b15aoai13ah1n04x5 U4913 (.a(n3630),
    .b(reg2hw_intr_ctrl_en_lvllow__q__12_),
    .c(net559),
    .d(net2263),
    .o1(n3631));
 b15oai112an1n12x5 U4914 (.a(n3632),
    .b(n3631),
    .c(net308),
    .d(n4127),
    .o1(n3768));
 b15oa0022an1n02x5 U4915 (.a(n4127),
    .b(net335),
    .c(n3768),
    .d(reg2hw_intr_state__q__12_),
    .o(u_reg_u_intr_state_wr_data[12]));
 b15nand02aq1n12x5 U4916 (.a(reg2hw_ctrl_en_input_filter__q__20_),
    .b(net2460),
    .o1(n3633));
 b15oai012as1n12x5 U4917 (.a(n3633),
    .b(reg2hw_ctrl_en_input_filter__q__20_),
    .c(n3634),
    .o1(u_reg_u_data_in_wr_data[20]));
 b15inv020ah1n03x5 U4918 (.a(data_in_q[20]),
    .o1(n3635));
 b15aoai13as1n08x5 U4919 (.a(u_reg_u_data_in_wr_data[20]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__20_),
    .c(reg2hw_intr_ctrl_en_rising__q__20_),
    .d(n3635),
    .o1(n3638));
 b15inv000ah1n02x5 U4920 (.a(u_reg_u_data_in_wr_data[20]),
    .o1(n3636));
 b15aoai13ah1n08x5 U4921 (.a(n3636),
    .b(reg2hw_intr_ctrl_en_lvllow__q__20_),
    .c(reg2hw_intr_ctrl_en_falling__q__20_),
    .d(data_in_q[20]),
    .o1(n3637));
 b15oai112as1n16x5 U4922 (.a(n3638),
    .b(n3637),
    .c(net307),
    .d(net698),
    .o1(n3777));
 b15oa0022al1n03x5 U4923 (.a(net699),
    .b(net334),
    .c(n3777),
    .d(reg2hw_intr_state__q__20_),
    .o(u_reg_u_intr_state_wr_data[20]));
 b15inv020as1n10x5 U4924 (.a(net684),
    .o1(n3640));
 b15nand02aq1n16x5 U4925 (.a(net581),
    .b(net2313),
    .o1(n3639));
 b15oai012ah1n48x5 U4926 (.a(n3639),
    .b(net580),
    .c(n3640),
    .o1(u_reg_u_data_in_wr_data[26]));
 b15inv000al1n02x5 U4927 (.a(data_in_q[26]),
    .o1(n3641));
 b15aoai13ah1n04x5 U4928 (.a(u_reg_u_data_in_wr_data[26]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__26_),
    .c(reg2hw_intr_ctrl_en_rising__q__26_),
    .d(n3641),
    .o1(n3644));
 b15inv000al1n02x5 U4929 (.a(u_reg_u_data_in_wr_data[26]),
    .o1(n3642));
 b15aoai13aq1n06x5 U4930 (.a(n3642),
    .b(reg2hw_intr_ctrl_en_lvllow__q__26_),
    .c(reg2hw_intr_ctrl_en_falling__q__26_),
    .d(data_in_q[26]),
    .o1(n3643));
 b15oai112as1n16x5 U4931 (.a(n3644),
    .b(n3643),
    .c(net307),
    .d(net693),
    .o1(n3796));
 b15oa0022an1n02x5 U4932 (.a(net693),
    .b(net334),
    .c(n3796),
    .d(reg2hw_intr_state__q__26_),
    .o(u_reg_u_intr_state_wr_data[26]));
 b15inv040ar1n03x5 U4933 (.a(gen_filter_9__u_filter_filter_synced),
    .o1(n3646));
 b15nandp2aq1n04x5 U4934 (.a(reg2hw_ctrl_en_input_filter__q__9_),
    .b(net2480),
    .o1(n3645));
 b15oai012aq1n16x5 U4935 (.a(n3645),
    .b(reg2hw_ctrl_en_input_filter__q__9_),
    .c(n3646),
    .o1(u_reg_u_data_in_wr_data[9]));
 b15inv020ar1n04x5 U4936 (.a(data_in_q[9]),
    .o1(n3647));
 b15aoai13ar1n08x5 U4937 (.a(u_reg_u_data_in_wr_data[9]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__9_),
    .c(reg2hw_intr_ctrl_en_rising__q__9_),
    .d(n3647),
    .o1(n3650));
 b15inv000al1n02x5 U4938 (.a(u_reg_u_data_in_wr_data[9]),
    .o1(n3648));
 b15aoai13ar1n08x5 U4939 (.a(n3648),
    .b(reg2hw_intr_ctrl_en_lvllow__q__9_),
    .c(reg2hw_intr_ctrl_en_falling__q__9_),
    .d(data_in_q[9]),
    .o1(n3649));
 b15oai112as1n16x5 U4940 (.a(n3650),
    .b(n3649),
    .c(net311),
    .d(n4124),
    .o1(n3760));
 b15oa0022as1n02x5 U4941 (.a(n4124),
    .b(net335),
    .c(n3760),
    .d(reg2hw_intr_state__q__9_),
    .o(u_reg_u_intr_state_wr_data[9]));
 b15nand02al1n12x5 U4942 (.a(net585),
    .b(net2451),
    .o1(n3653));
 b15oai012aq1n32x5 U4943 (.a(n3653),
    .b(net585),
    .c(n3654),
    .o1(u_reg_u_data_in_wr_data[22]));
 b15inv000aq1n02x5 U4944 (.a(data_in_q[22]),
    .o1(n3655));
 b15aoai13as1n06x5 U4945 (.a(u_reg_u_data_in_wr_data[22]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__22_),
    .c(reg2hw_intr_ctrl_en_rising__q__22_),
    .d(n3655),
    .o1(n3658));
 b15inv000al1n02x5 U4946 (.a(u_reg_u_data_in_wr_data[22]),
    .o1(n3656));
 b15aoai13as1n04x5 U4947 (.a(n3656),
    .b(reg2hw_intr_ctrl_en_lvllow__q__22_),
    .c(reg2hw_intr_ctrl_en_falling__q__22_),
    .d(data_in_q[22]),
    .o1(n3657));
 b15oai112as1n16x5 U4948 (.a(n3658),
    .b(n3657),
    .c(net310),
    .d(n4136),
    .o1(n3776));
 b15oa0022ar1n04x5 U4949 (.a(n4136),
    .b(net334),
    .c(n3776),
    .d(reg2hw_intr_state__q__22_),
    .o(u_reg_u_intr_state_wr_data[22]));
 b15nand02aq1n04x5 U4950 (.a(net578),
    .b(net2446),
    .o1(n3659));
 b15oai012aq1n16x5 U4951 (.a(n3659),
    .b(net578),
    .c(n3660),
    .o1(u_reg_u_data_in_wr_data[29]));
 b15inv040al1n03x5 U4952 (.a(data_in_q[29]),
    .o1(n3661));
 b15aoai13al1n08x5 U4953 (.a(u_reg_u_data_in_wr_data[29]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__29_),
    .c(reg2hw_intr_ctrl_en_rising__q__29_),
    .d(n3661),
    .o1(n3664));
 b15inv000al1n02x5 U4954 (.a(u_reg_u_data_in_wr_data[29]),
    .o1(n3662));
 b15aoai13an1n08x5 U4955 (.a(n3662),
    .b(reg2hw_intr_ctrl_en_lvllow__q__29_),
    .c(reg2hw_intr_ctrl_en_falling__q__29_),
    .d(data_in_q[29]),
    .o1(n3663));
 b15oai112as1n16x5 U4956 (.a(n3664),
    .b(n3663),
    .c(net310),
    .d(net691),
    .o1(n3784));
 b15oa0022al1n03x5 U4957 (.a(net690),
    .b(net334),
    .c(n3784),
    .d(net2453),
    .o(u_reg_u_intr_state_wr_data[29]));
 b15inv040ah1n04x5 U4958 (.a(gen_filter_25__u_filter_filter_synced),
    .o1(n3666));
 b15nand02an1n08x5 U4959 (.a(reg2hw_ctrl_en_input_filter__q__25_),
    .b(net2466),
    .o1(n3665));
 b15oai012ah1n24x5 U4960 (.a(n3665),
    .b(reg2hw_ctrl_en_input_filter__q__25_),
    .c(n3666),
    .o1(u_reg_u_data_in_wr_data[25]));
 b15inv020ar1n04x5 U4961 (.a(data_in_q[25]),
    .o1(n3667));
 b15aoai13aq1n08x5 U4962 (.a(u_reg_u_data_in_wr_data[25]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__25_),
    .c(reg2hw_intr_ctrl_en_rising__q__25_),
    .d(n3667),
    .o1(n3670));
 b15inv020ar1n04x5 U4963 (.a(u_reg_u_data_in_wr_data[25]),
    .o1(n3668));
 b15aoai13as1n08x5 U4964 (.a(n3668),
    .b(reg2hw_intr_ctrl_en_lvllow__q__25_),
    .c(reg2hw_intr_ctrl_en_falling__q__25_),
    .d(data_in_q[25]),
    .o1(n3669));
 b15oai112as1n16x5 U4965 (.a(n3670),
    .b(n3669),
    .c(net307),
    .d(net696),
    .o1(n3788));
 b15oa0022ah1n02x5 U4966 (.a(net696),
    .b(net334),
    .c(n3788),
    .d(reg2hw_intr_state__q__25_),
    .o(u_reg_u_intr_state_wr_data[25]));
 b15inv040ah1n06x5 U4967 (.a(gen_filter_24__u_filter_filter_synced),
    .o1(n3672));
 b15nand02ah1n12x5 U4968 (.a(net582),
    .b(gen_filter_24__u_filter_stored_value_q),
    .o1(n3671));
 b15oai012aq1n48x5 U4969 (.a(n3671),
    .b(net582),
    .c(n3672),
    .o1(u_reg_u_data_in_wr_data[24]));
 b15inv000as1n02x5 U4970 (.a(data_in_q[24]),
    .o1(n3673));
 b15aoai13al1n08x5 U4971 (.a(u_reg_u_data_in_wr_data[24]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__24_),
    .c(reg2hw_intr_ctrl_en_rising__q__24_),
    .d(n3673),
    .o1(n3676));
 b15inv000al1n02x5 U4972 (.a(u_reg_u_data_in_wr_data[24]),
    .o1(n3674));
 b15aoai13as1n06x5 U4973 (.a(n3674),
    .b(reg2hw_intr_ctrl_en_lvllow__q__24_),
    .c(reg2hw_intr_ctrl_en_falling__q__24_),
    .d(data_in_q[24]),
    .o1(n3675));
 b15oai112as1n16x5 U4974 (.a(n3676),
    .b(n3675),
    .c(n4138),
    .d(net310),
    .o1(n3764));
 b15oa0022an1n03x5 U4975 (.a(n4138),
    .b(net334),
    .c(n3764),
    .d(reg2hw_intr_state__q__24_),
    .o(u_reg_u_intr_state_wr_data[24]));
 b15nandp2ah1n48x5 U4976 (.a(n3680),
    .b(n3679),
    .o1(n3812));
 b15aoai13ah1n02x5 U4978 (.a(n4189),
    .b(n3825),
    .c(net199),
    .d(n4134),
    .o1(n3681));
 b15oai012aq1n08x5 U4979 (.a(n3681),
    .b(n4186),
    .c(net689),
    .o1(N43));
 b15aoai13an1n03x5 U4980 (.a(n4189),
    .b(n3822),
    .c(net204),
    .d(net695),
    .o1(n3682));
 b15oai012ar1n02x5 U4981 (.a(n3682),
    .b(net321),
    .c(n4124),
    .o1(N48));
 b15aoai13an1n08x5 U4982 (.a(n4189),
    .b(n3828),
    .c(net636),
    .d(net692),
    .o1(n3683));
 b15oai012an1n24x5 U4983 (.a(n3683),
    .b(net322),
    .c(n3818),
    .o1(N52));
 b15aoai13as1n08x5 U4984 (.a(net721),
    .b(net326),
    .c(n4189),
    .d(net714),
    .o1(n3684));
 b15oai013as1n12x5 U4985 (.a(n3684),
    .b(net714),
    .c(net305),
    .d(n3685),
    .o1(N42));
 b15inv000ah1n16x5 U4986 (.a(net195),
    .o1(n3887));
 b15aoai13as1n08x5 U4987 (.a(net722),
    .b(net326),
    .c(n4189),
    .d(net75),
    .o1(n3686));
 b15oai013as1n12x5 U4988 (.a(n3686),
    .b(net75),
    .c(net305),
    .d(n3887),
    .o1(N41));
 b15aoai13aq1n08x5 U4989 (.a(net68),
    .b(net327),
    .c(n4189),
    .d(net86),
    .o1(n3687));
 b15oai013as1n12x5 U4990 (.a(n3687),
    .b(net86),
    .c(net304),
    .d(n3688),
    .o1(N51));
 b15aoai13an1n06x5 U4991 (.a(net67),
    .b(net328),
    .c(n4189),
    .d(net85),
    .o1(n3689));
 b15oai013as1n12x5 U4992 (.a(n3689),
    .b(net85),
    .c(n3812),
    .d(n3690),
    .o1(N50));
 b15aoai13ah1n04x5 U4993 (.a(net720),
    .b(net328),
    .c(n4189),
    .d(net78),
    .o1(n3691));
 b15oai013as1n12x5 U4994 (.a(n3691),
    .b(net78),
    .c(n3812),
    .d(n3692),
    .o1(N44));
 b15aoai13an1n06x5 U4995 (.a(net62),
    .b(net328),
    .c(net79),
    .d(n4189),
    .o1(n3693));
 b15oai013as1n12x5 U4996 (.a(n3693),
    .b(net79),
    .c(n3812),
    .d(n3694),
    .o1(N45));
 b15aoai13ah1n04x5 U4997 (.a(net66),
    .b(net328),
    .c(net84),
    .d(n4189),
    .o1(n3696));
 b15oai013as1n12x5 U4998 (.a(n3696),
    .b(net84),
    .c(n3812),
    .d(n3697),
    .o1(N49));
 b15nand02an1n08x5 U5001 (.a(net708),
    .b(n4142),
    .o1(n3701));
 b15oai012as1n48x5 U5002 (.a(net342),
    .b(net660),
    .c(net669),
    .o1(n3700));
 b15aoi012an1n32x5 U5003 (.a(n3700),
    .b(n4127),
    .c(net669),
    .o1(N126));
 b15nand02an1n32x5 U5004 (.a(net708),
    .b(n4145),
    .o1(n3705));
 b15oai012aq1n03x5 U5005 (.a(net343),
    .b(net147),
    .c(n3705),
    .o1(n3704));
 b15aoi012ar1n04x5 U5006 (.a(n3704),
    .b(n4129),
    .c(n3705),
    .o1(N129));
 b15nandp2al1n48x5 U5007 (.a(net709),
    .b(n4135),
    .o1(n3709));
 b15oai012al1n48x5 U5008 (.a(net340),
    .b(net168),
    .c(n3709),
    .o1(n3708));
 b15aoi012ah1n16x5 U5009 (.a(n3708),
    .b(n4120),
    .c(n3709),
    .o1(N119));
 b15nandp2as1n24x5 U5010 (.a(net709),
    .b(n4130),
    .o1(n3713));
 b15oai012ar1n08x5 U5011 (.a(net343),
    .b(net666),
    .c(n3713),
    .o1(n3712));
 b15aoi012ah1n08x5 U5012 (.a(n3712),
    .b(net706),
    .c(n3713),
    .o1(N114));
 b15nand02ah1n24x5 U5013 (.a(net708),
    .b(n4137),
    .o1(n3716));
 b15oai012an1n24x5 U5014 (.a(net340),
    .b(net170),
    .c(net668),
    .o1(n3715));
 b15aoi012as1n12x5 U5015 (.a(net325),
    .b(n4122),
    .c(n3716),
    .o1(N121));
 b15nandp2as1n24x5 U5016 (.a(net708),
    .b(n4133),
    .o1(n3720));
 b15oai012ah1n02x5 U5017 (.a(net343),
    .b(net166),
    .c(n3720),
    .o1(n3719));
 b15aoi012ar1n04x5 U5018 (.a(n3719),
    .b(n4119),
    .c(n3720),
    .o1(N117));
 b15nand02ah1n24x5 U5019 (.a(net708),
    .b(n4132),
    .o1(n3724));
 b15oai012ar1n03x5 U5020 (.a(net343),
    .b(net163),
    .c(n3724),
    .o1(n3723));
 b15aoi012an1n02x5 U5021 (.a(n3723),
    .b(n4118),
    .c(n3724),
    .o1(N116));
 b15nand02as1n48x5 U5022 (.a(net709),
    .b(n4141),
    .o1(n3728));
 b15oai012as1n32x5 U5023 (.a(net340),
    .b(net143),
    .c(n3728),
    .o1(n3727));
 b15aoi012as1n16x5 U5024 (.a(n3727),
    .b(n4126),
    .c(n3728),
    .o1(N125));
 b15nandp2aq1n04x5 U5025 (.a(net708),
    .b(n4136),
    .o1(n3732));
 b15oai012as1n48x5 U5026 (.a(net340),
    .b(net640),
    .c(net667),
    .o1(n3731));
 b15aoi012aq1n32x5 U5027 (.a(n3731),
    .b(n4121),
    .c(net667),
    .o1(N120));
 b15nand02ah1n32x5 U5028 (.a(net708),
    .b(n4144),
    .o1(n3736));
 b15oai012ah1n03x5 U5029 (.a(net343),
    .b(net146),
    .c(n3736),
    .o1(n3735));
 b15aoi012ah1n04x5 U5030 (.a(n3735),
    .b(net703),
    .c(n3736),
    .o1(N128));
 b15nand02as1n48x5 U5031 (.a(net708),
    .b(n4140),
    .o1(n3740));
 b15oai012al1n48x5 U5032 (.a(net340),
    .b(net662),
    .c(n3740),
    .o1(n3739));
 b15aoi012ah1n16x5 U5033 (.a(n3739),
    .b(n4125),
    .c(n3740),
    .o1(N124));
 b15nandp2ar1n32x5 U5034 (.a(net708),
    .b(n4131),
    .o1(n3743));
 b15oai012ah1n03x5 U5035 (.a(net343),
    .b(net664),
    .c(n3743),
    .o1(n3742));
 b15aoi012ah1n04x5 U5036 (.a(n3742),
    .b(net704),
    .c(n3743),
    .o1(N115));
 b15nand02ah1n24x5 U5037 (.a(net708),
    .b(n4138),
    .o1(n3747));
 b15oai012ah1n02x5 U5038 (.a(net343),
    .b(net171),
    .c(n3747),
    .o1(n3746));
 b15aoi012ah1n02x5 U5039 (.a(n3746),
    .b(n4123),
    .c(n3747),
    .o1(N122));
 b15nandp2an1n32x5 U5040 (.a(net322),
    .b(n3749),
    .o1(N55));
 b15oai112al1n06x5 U5042 (.a(net84),
    .b(N55),
    .c(net66),
    .d(net408),
    .o1(n3750));
 b15oai013al1n08x5 U5043 (.a(n3750),
    .b(net84),
    .c(net349),
    .d(n3751),
    .o1(N66));
 b15nandp2al1n08x5 U5044 (.a(net392),
    .b(net180),
    .o1(n3869));
 b15oai112al1n12x5 U5045 (.a(net73),
    .b(N55),
    .c(net724),
    .d(net408),
    .o1(n3752));
 b15oai013as1n12x5 U5046 (.a(n3752),
    .b(net73),
    .c(net349),
    .d(net362),
    .o1(N56));
 b15nand02as1n16x5 U5047 (.a(net358),
    .b(n4131),
    .o1(n3857));
 b15oai112as1n16x5 U5048 (.a(net715),
    .b(N55),
    .c(net723),
    .d(net327),
    .o1(n3755));
 b15oai012aq1n16x5 U5049 (.a(n3755),
    .b(n3756),
    .c(n3857),
    .o1(N57));
 b15nor004ah1n08x5 U5050 (.a(n3760),
    .b(n3759),
    .c(n3758),
    .d(n3757),
    .o1(n3799));
 b15nor004an1n08x5 U5051 (.a(n3764),
    .b(n3763),
    .c(n3762),
    .d(n3761),
    .o1(n3798));
 b15nor004aq1n04x5 U5052 (.a(n3768),
    .b(n3767),
    .c(n3766),
    .d(n3765),
    .o1(n3770));
 b15nand04aq1n08x5 U5053 (.a(n3772),
    .b(n3771),
    .c(n3770),
    .d(net334),
    .o1(n3794));
 b15nor004al1n06x5 U5054 (.a(n3776),
    .b(n3775),
    .c(n3774),
    .d(n3773),
    .o1(n3792));
 b15nor004aq1n08x5 U5055 (.a(n3780),
    .b(n3779),
    .c(n3778),
    .d(n3777),
    .o1(n3791));
 b15nor004ah1n12x5 U5056 (.a(n3784),
    .b(n3783),
    .c(n3782),
    .d(n3781),
    .o1(n3790));
 b15nor004an1n03x5 U5057 (.a(n3788),
    .b(n3787),
    .c(n3786),
    .d(n3785),
    .o1(n3789));
 b15nand04aq1n08x5 U5058 (.a(n3792),
    .b(n3791),
    .c(n3790),
    .d(n3789),
    .o1(n3793));
 b15nor004aq1n06x5 U5059 (.a(n3796),
    .b(n3795),
    .c(n3794),
    .d(n3793),
    .o1(n3797));
 b15nand03ar1n16x5 U5060 (.a(n3799),
    .b(n3798),
    .c(n3797),
    .o1(u_reg_u_intr_state_n1));
 b15nandp2ar1n24x5 U5061 (.a(net322),
    .b(net304),
    .o1(N38));
 b15oai112an1n08x5 U5062 (.a(net718),
    .b(N38),
    .c(net88),
    .d(net406),
    .o1(n3801));
 b15oai013as1n12x5 U5063 (.a(n3801),
    .b(net88),
    .c(net304),
    .d(n3802),
    .o1(N53));
 b15oai112ah1n08x5 U5064 (.a(net719),
    .b(net300),
    .c(net712),
    .d(net411),
    .o1(n3803));
 b15oai013as1n12x5 U5065 (.a(n3803),
    .b(net712),
    .c(net305),
    .d(n3804),
    .o1(N47));
 b15oai112as1n02x5 U5066 (.a(net63),
    .b(net300),
    .c(net80),
    .d(net407),
    .o1(n3805));
 b15oai013aq1n08x5 U5067 (.a(n3805),
    .b(net80),
    .c(n3812),
    .d(n3806),
    .o1(N46));
 b15inv000as1n16x5 U5068 (.a(net173),
    .o1(n3874));
 b15oai112al1n12x5 U5069 (.a(net724),
    .b(net300),
    .c(net73),
    .d(net408),
    .o1(n3807));
 b15oai013as1n12x5 U5070 (.a(n3807),
    .b(net73),
    .c(net305),
    .d(n3874),
    .o1(N39));
 b15oai112as1n16x5 U5071 (.a(net723),
    .b(net300),
    .c(net715),
    .d(net408),
    .o1(n3808));
 b15oai013as1n12x5 U5072 (.a(n3808),
    .b(net715),
    .c(net305),
    .d(n3809),
    .o1(N40));
 b15inv000ah1n20x5 U5073 (.a(net179),
    .o1(n3811));
 b15oai112as1n16x5 U5074 (.a(net717),
    .b(N38),
    .c(net89),
    .d(net406),
    .o1(n3810));
 b15oai013as1n12x5 U5075 (.a(n3810),
    .b(net89),
    .c(net304),
    .d(n3811),
    .o1(N54));
 b15aoi012as1n32x5 U5076 (.a(n3825),
    .b(net167),
    .c(n4134),
    .o1(n3815));
 b15nandp2aq1n48x5 U5077 (.a(net710),
    .b(N113),
    .o1(n3819));
 b15nand02an1n48x5 U5078 (.a(net341),
    .b(n4146),
    .o1(n3861));
 b15oai022ah1n48x5 U5079 (.a(n3815),
    .b(n3819),
    .c(net688),
    .d(net324),
    .o1(N118));
 b15aoi012ar1n12x5 U5080 (.a(n3822),
    .b(net172),
    .c(net695),
    .o1(n3817));
 b15oai022an1n08x5 U5081 (.a(n3817),
    .b(n3819),
    .c(n4124),
    .d(net324),
    .o1(N123));
 b15aoi012as1n32x5 U5082 (.a(n3828),
    .b(net145),
    .c(n4143),
    .o1(n3820));
 b15oai022ah1n48x5 U5083 (.a(n3820),
    .b(n3819),
    .c(n3818),
    .d(net323),
    .o1(N127));
 b15and002aq1n12x5 U5084 (.a(net432),
    .b(net359),
    .o(n3859));
 b15aoai13al1n08x5 U5085 (.a(net333),
    .b(net670),
    .c(net158),
    .d(net696),
    .o1(n3823));
 b15oai012an1n04x5 U5086 (.a(n3823),
    .b(n3861),
    .c(net694),
    .o1(N140));
 b15aoai13ar1n03x5 U5087 (.a(net333),
    .b(n3825),
    .c(net153),
    .d(net698),
    .o1(n3826));
 b15oai012aq1n06x5 U5088 (.a(n3826),
    .b(n3861),
    .c(net698),
    .o1(N135));
 b15aoai13an1n08x5 U5089 (.a(net332),
    .b(n3828),
    .c(net162),
    .d(n4143),
    .o1(n3829));
 b15oai012aq1n06x5 U5090 (.a(n3829),
    .b(net323),
    .c(net692),
    .o1(N144));
 b15aoai13al1n06x5 U5092 (.a(net713),
    .b(n4188),
    .c(net720),
    .d(net333),
    .o1(n3831));
 b15oai013aq1n12x5 U5093 (.a(n3831),
    .b(net713),
    .c(net350),
    .d(n3832),
    .o1(N136));
 b15aoai13ar1n02x5 U5094 (.a(net85),
    .b(n4188),
    .c(net67),
    .d(n3859),
    .o1(n3833));
 b15oai013an1n02x5 U5095 (.a(n3833),
    .b(net85),
    .c(net349),
    .d(n3834),
    .o1(N142));
 b15aoai13al1n02x5 U5096 (.a(net76),
    .b(net318),
    .c(net721),
    .d(net332),
    .o1(n3835));
 b15oai013ar1n02x5 U5097 (.a(n3835),
    .b(net76),
    .c(net351),
    .d(n3836),
    .o1(N134));
 b15aoai13as1n02x5 U5098 (.a(net86),
    .b(net318),
    .c(net68),
    .d(net332),
    .o1(n3837));
 b15oai013as1n06x5 U5099 (.a(n3837),
    .b(net86),
    .c(net351),
    .d(n3838),
    .o1(N143));
 b15aoai13aq1n02x5 U5100 (.a(net89),
    .b(net318),
    .c(net717),
    .d(net332),
    .o1(n3839));
 b15oai013as1n02x5 U5101 (.a(n3839),
    .b(net89),
    .c(net351),
    .d(n3840),
    .o1(N146));
 b15nandp2as1n24x5 U5102 (.a(net430),
    .b(net658),
    .o1(n3881));
 b15aoai13al1n02x5 U5103 (.a(net75),
    .b(net318),
    .c(net722),
    .d(net332),
    .o1(n3842));
 b15oai013aq1n04x5 U5104 (.a(n3842),
    .b(net75),
    .c(net351),
    .d(n3881),
    .o1(N133));
 b15aoai13as1n04x5 U5105 (.a(net80),
    .b(n4188),
    .c(net63),
    .d(n3859),
    .o1(n3843));
 b15oai013as1n03x5 U5106 (.a(n3843),
    .b(net80),
    .c(net349),
    .d(n3844),
    .o1(N138));
 b15aoai13an1n02x5 U5107 (.a(net84),
    .b(n4188),
    .c(n3859),
    .d(net66),
    .o1(n3845));
 b15oai013ah1n04x5 U5108 (.a(n3845),
    .b(net84),
    .c(net349),
    .d(n3846),
    .o1(N141));
 b15aoai13ar1n06x5 U5109 (.a(net79),
    .b(n4188),
    .c(n3859),
    .d(net62),
    .o1(n3847));
 b15oai013aq1n06x5 U5110 (.a(n3847),
    .b(net79),
    .c(net349),
    .d(n3848),
    .o1(N137));
 b15aoai13aq1n03x5 U5111 (.a(net712),
    .b(n4188),
    .c(net333),
    .d(net719),
    .o1(n3849));
 b15oai013aq1n12x5 U5112 (.a(n3849),
    .b(net712),
    .c(net349),
    .d(n3850),
    .o1(N139));
 b15aoai13ar1n02x5 U5113 (.a(net88),
    .b(net318),
    .c(net332),
    .d(net718),
    .o1(n3851));
 b15oai013an1n02x5 U5114 (.a(n3851),
    .b(net88),
    .c(net351),
    .d(n3852),
    .o1(N145));
 b15oai012aq1n08x5 U5115 (.a(net715),
    .b(net723),
    .c(net318),
    .o1(n3855));
 b15nor002as1n08x5 U5116 (.a(net332),
    .b(net318),
    .o1(n3858));
 b15oaoi13as1n08x5 U5117 (.a(n3858),
    .b(n3855),
    .c(n3857),
    .d(n3856),
    .o1(N132));
 b15inv000ah1n08x5 U5118 (.a(n3858),
    .o1(N130));
 b15aoai13an1n06x5 U5119 (.a(N130),
    .b(net716),
    .c(net332),
    .d(net148),
    .o1(n3860));
 b15aoi013aq1n03x5 U5120 (.a(n3860),
    .b(net716),
    .c(net705),
    .d(net323),
    .o1(N131));
 b15nor004ar1n08x5 U5121 (.a(net41),
    .b(net42),
    .c(n3864),
    .d(n3863),
    .o1(u_reg_u_reg_if_rd_req));
 b15and003ar1n08x5 U5122 (.a(n3867),
    .b(n3866),
    .c(n3865),
    .o(gen_alert_tx_0__u_prim_alert_sender_alert_pd));
 b15aoi022ah1n06x5 U5123 (.a(net551),
    .b(net437),
    .c(net562),
    .d(net396),
    .o1(n3879));
 b15aoi022as1n48x5 U5124 (.a(net430),
    .b(net659),
    .c(net379),
    .d(net678),
    .o1(n3878));
 b15inv040as1n02x5 U5125 (.a(reg2hw_intr_state__q__0_),
    .o1(n3872));
 b15aoi022ar1n48x5 U5127 (.a(net540),
    .b(net371),
    .c(net427),
    .d(net665),
    .o1(n3870));
 b15oai112al1n16x5 U5128 (.a(n3870),
    .b(net362),
    .c(n3872),
    .d(n4174),
    .o1(n3876));
 b15aoi022an1n12x5 U5129 (.a(reg2hw_intr_ctrl_en_rising__q__0_),
    .b(net443),
    .c(net419),
    .d(reg2hw_intr_enable__q__0_),
    .o1(n3873));
 b15oai012al1n08x5 U5130 (.a(n3873),
    .b(n3874),
    .c(net367),
    .o1(n3875));
 b15aoi112as1n08x5 U5131 (.a(n3876),
    .b(n3875),
    .c(net611),
    .d(net388),
    .o1(n3877));
 b15nand04as1n16x5 U5132 (.a(net357),
    .b(n3879),
    .c(n3878),
    .d(n3877),
    .o1(u_reg_u_reg_if_N14));
 b15aoi022ar1n32x5 U5133 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__2_),
    .b(net437),
    .c(net391),
    .d(net182),
    .o1(n3892));
 b15aoi022ah1n12x5 U5134 (.a(net554),
    .b(net396),
    .c(net433),
    .d(reg2hw_intr_state__q__2_),
    .o1(n3891));
 b15aoi022as1n04x5 U5136 (.a(reg2hw_intr_ctrl_en_rising__q__2_),
    .b(net444),
    .c(reg2hw_intr_ctrl_en_lvllow__q__2_),
    .d(net369),
    .o1(n3882));
 b15oai112as1n16x5 U5137 (.a(n3882),
    .b(n3881),
    .c(n3884),
    .d(n4177),
    .o1(n3889));
 b15aoi022as1n08x5 U5138 (.a(net418),
    .b(reg2hw_intr_enable__q__2_),
    .c(net376),
    .d(u_reg_data_in_qs[2]),
    .o1(n3885));
 b15oai012al1n08x5 U5139 (.a(n3885),
    .b(n3887),
    .c(net366),
    .o1(n3888));
 b15aoi112as1n08x5 U5140 (.a(n3889),
    .b(n3888),
    .c(net427),
    .d(net163),
    .o1(n3890));
 b15nand04as1n16x5 U5141 (.a(net357),
    .b(n3892),
    .c(n3891),
    .d(n3890),
    .o1(u_reg_u_reg_if_N16));
 b15aoi022an1n48x5 U5143 (.a(net552),
    .b(net399),
    .c(net425),
    .d(net642),
    .o1(n3896));
 b15aoi022aq1n08x5 U5144 (.a(reg2hw_intr_ctrl_en_rising__q__4_),
    .b(net444),
    .c(net420),
    .d(reg2hw_intr_enable__q__4_),
    .o1(n3895));
 b15aoi022ar1n32x5 U5145 (.a(net570),
    .b(net384),
    .c(net431),
    .d(net657),
    .o1(n3894));
 b15aoi022as1n12x5 U5146 (.a(reg2hw_intr_ctrl_en_lvllow__q__4_),
    .b(net372),
    .c(net199),
    .d(n4176),
    .o1(n3893));
 b15nand04ah1n12x5 U5147 (.a(n3896),
    .b(n3895),
    .c(n3894),
    .d(n3893),
    .o1(n3899));
 b15aoi022as1n16x5 U5148 (.a(net544),
    .b(net437),
    .c(net373),
    .d(u_reg_data_in_qs[4]),
    .o1(n3898));
 b15aoi022as1n12x5 U5149 (.a(net436),
    .b(net508),
    .c(net394),
    .d(net185),
    .o1(n3897));
 b15nona23as1n24x5 U5150 (.a(net352),
    .b(n3899),
    .c(n3898),
    .d(n3897),
    .out0(u_reg_u_reg_if_N18));
 b15aoi022ah1n08x5 U5151 (.a(reg2hw_intr_ctrl_en_falling__q__9_),
    .b(net396),
    .c(net375),
    .d(net2256),
    .o1(n3904));
 b15aoi022ah1n06x5 U5152 (.a(reg2hw_intr_ctrl_en_rising__q__9_),
    .b(net443),
    .c(net418),
    .d(reg2hw_intr_enable__q__9_),
    .o1(n3903));
 b15aoi022ah1n08x5 U5153 (.a(reg2hw_ctrl_en_input_filter__q__9_),
    .b(net386),
    .c(net436),
    .d(reg2hw_intr_state__q__9_),
    .o1(n3902));
 b15aoi022an1n32x5 U5154 (.a(net427),
    .b(net172),
    .c(net204),
    .d(n4176),
    .o1(n3901));
 b15nand04as1n16x5 U5155 (.a(n3904),
    .b(n3903),
    .c(n3902),
    .d(n3901),
    .o1(n3907));
 b15aoi022ah1n48x5 U5156 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__9_),
    .b(net437),
    .c(reg2hw_intr_ctrl_en_lvllow__q__9_),
    .d(net371),
    .o1(n3906));
 b15aoi022ah1n24x5 U5157 (.a(net429),
    .b(net648),
    .c(n3909),
    .d(net621),
    .o1(n3905));
 b15nona23as1n08x5 U5158 (.a(net354),
    .b(n3907),
    .c(n3906),
    .d(n3905),
    .out0(u_reg_u_reg_if_N23));
 b15aoi022al1n24x5 U5159 (.a(net548),
    .b(net439),
    .c(net430),
    .d(net162),
    .o1(n3914));
 b15aoi022al1n24x5 U5160 (.a(net558),
    .b(net396),
    .c(net422),
    .d(net523),
    .o1(n3913));
 b15aoi022al1n24x5 U5161 (.a(net527),
    .b(net447),
    .c(net392),
    .d(net616),
    .o1(n3912));
 b15aoi022ar1n32x5 U5162 (.a(net636),
    .b(n4176),
    .c(net379),
    .d(u_reg_data_in_qs[13]),
    .o1(n3911));
 b15nand04as1n16x5 U5163 (.a(n3914),
    .b(n3913),
    .c(n3912),
    .d(n3911),
    .o1(n3918));
 b15aoi022as1n16x5 U5164 (.a(net600),
    .b(net388),
    .c(net538),
    .d(net370),
    .o1(n3917));
 b15aoi022as1n32x5 U5165 (.a(net433),
    .b(net512),
    .c(net426),
    .d(net145),
    .o1(n3916));
 b15nona23as1n32x5 U5166 (.a(n4178),
    .b(n3918),
    .c(n3917),
    .d(n3916),
    .out0(u_reg_u_reg_if_N27));
 b15aoi022aq1n32x5 U5167 (.a(net547),
    .b(net439),
    .c(net410),
    .d(net180),
    .o1(n3926));
 b15aoi022as1n06x5 U5168 (.a(reg2hw_intr_ctrl_en_lvllow__q__16_),
    .b(net370),
    .c(net374),
    .d(net2126),
    .o1(n3925));
 b15norp02al1n32x5 U5169 (.a(n3920),
    .b(n3919),
    .o1(n4026));
 b15aoi022ar1n48x5 U5170 (.a(net148),
    .b(net412),
    .c(net422),
    .d(net522),
    .o1(n3924));
 b15aoi022ar1n02x5 U5171 (.a(reg2hw_intr_ctrl_en_rising__q__16_),
    .b(net447),
    .c(reg2hw_intr_ctrl_en_falling__q__16_),
    .d(net397),
    .o1(n3921));
 b15aob012al1n06x5 U5172 (.a(n3921),
    .b(net433),
    .c(reg2hw_intr_state__q__16_),
    .out0(n3922));
 b15aoi112aq1n06x5 U5173 (.a(net353),
    .b(n3922),
    .c(net594),
    .d(net383),
    .o1(n3923));
 b15nand04ah1n08x5 U5174 (.a(n3926),
    .b(net2127),
    .c(n3924),
    .d(n3923),
    .o1(u_reg_u_reg_if_N30));
 b15aoi022aq1n08x5 U5175 (.a(net2376),
    .b(net439),
    .c(reg2hw_intr_ctrl_en_lvllow__q__17_),
    .d(net368),
    .o1(n3932));
 b15aoi022an1n08x5 U5176 (.a(reg2hw_intr_ctrl_en_rising__q__17_),
    .b(net447),
    .c(net422),
    .d(reg2hw_intr_enable__q__17_),
    .o1(n3931));
 b15aoi022ah1n32x5 U5177 (.a(net410),
    .b(net181),
    .c(net374),
    .d(u_reg_data_in_qs[17]),
    .o1(n3930));
 b15aoi022an1n02x5 U5178 (.a(reg2hw_intr_ctrl_en_falling__q__17_),
    .b(net397),
    .c(net149),
    .d(net412),
    .o1(n3927));
 b15aob012aq1n04x5 U5179 (.a(n3927),
    .b(net433),
    .c(reg2hw_intr_state__q__17_),
    .out0(n3928));
 b15aoi112al1n08x5 U5180 (.a(net353),
    .b(n3928),
    .c(net592),
    .d(net383),
    .o1(n3929));
 b15nand04as1n16x5 U5181 (.a(n3932),
    .b(n3931),
    .c(n3930),
    .d(n3929),
    .o1(u_reg_u_reg_if_N31));
 b15aoi022aq1n08x5 U5182 (.a(reg2hw_intr_ctrl_en_rising__q__18_),
    .b(net447),
    .c(net422),
    .d(reg2hw_intr_enable__q__18_),
    .o1(n3940));
 b15aoi022ah1n06x5 U5183 (.a(net590),
    .b(net383),
    .c(net556),
    .d(net397),
    .o1(n3939));
 b15aoi022ah1n08x5 U5184 (.a(net433),
    .b(reg2hw_intr_state__q__18_),
    .c(net658),
    .d(net412),
    .o1(n3938));
 b15aoi022an1n02x5 U5185 (.a(reg2hw_intr_ctrl_en_lvllow__q__18_),
    .b(net368),
    .c(net374),
    .d(net2014),
    .o1(n3933));
 b15oai012as1n03x5 U5186 (.a(net2015),
    .b(net416),
    .c(net415),
    .o1(n3936));
 b15aoi112ar1n08x5 U5187 (.a(net353),
    .b(n3936),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__18_),
    .d(net439),
    .o1(n3937));
 b15nand04ah1n16x5 U5188 (.a(n3940),
    .b(n3939),
    .c(n3938),
    .d(net2016),
    .o1(u_reg_u_reg_if_N32));
 b15aoi022as1n04x5 U5189 (.a(net588),
    .b(net383),
    .c(net2552),
    .d(net440),
    .o1(n3946));
 b15aoi022ar1n08x5 U5190 (.a(reg2hw_intr_ctrl_en_falling__q__19_),
    .b(net398),
    .c(net422),
    .d(reg2hw_intr_enable__q__19_),
    .o1(n3945));
 b15aoi022ar1n02x3 U5191 (.a(net433),
    .b(reg2hw_intr_state__q__19_),
    .c(net410),
    .d(net629),
    .o1(n3943));
 b15aoi022ar1n02x3 U5192 (.a(reg2hw_intr_ctrl_en_rising__q__19_),
    .b(net447),
    .c(net151),
    .d(net412),
    .o1(n3942));
 b15aoi022ar1n02x5 U5193 (.a(reg2hw_intr_ctrl_en_lvllow__q__19_),
    .b(net368),
    .c(net374),
    .d(net2005),
    .o1(n3941));
 b15and003as1n02x5 U5194 (.a(n3943),
    .b(n3942),
    .c(net2006),
    .o(n3944));
 b15nand04as1n12x5 U5195 (.a(net355),
    .b(n3946),
    .c(n3945),
    .d(n3944),
    .o1(u_reg_u_reg_if_N33));
 b15aoi022ah1n06x5 U5196 (.a(reg2hw_ctrl_en_input_filter__q__20_),
    .b(net384),
    .c(net417),
    .d(reg2hw_intr_enable__q__20_),
    .o1(n3952));
 b15aoi022as1n08x5 U5197 (.a(reg2hw_intr_ctrl_en_lvllow__q__20_),
    .b(n3318),
    .c(reg2hw_intr_ctrl_en_falling__q__20_),
    .d(net398),
    .o1(n3951));
 b15aoi022ah1n08x5 U5198 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__20_),
    .b(net438),
    .c(n3316),
    .d(net2056),
    .o1(n3950));
 b15aoi022aq1n16x5 U5199 (.a(net407),
    .b(net628),
    .c(net656),
    .d(n4026),
    .o1(n3947));
 b15aob012ar1n08x5 U5200 (.a(net361),
    .b(net434),
    .c(reg2hw_intr_state__q__20_),
    .out0(n3948));
 b15aoi112al1n08x5 U5201 (.a(net354),
    .b(n3948),
    .c(reg2hw_intr_ctrl_en_rising__q__20_),
    .d(net442),
    .o1(n3949));
 b15nand04ah1n16x5 U5202 (.a(n3952),
    .b(n3951),
    .c(net2057),
    .d(n3949),
    .o1(u_reg_u_reg_if_N34));
 b15aoi022ar1n12x5 U5203 (.a(net546),
    .b(net437),
    .c(net409),
    .d(net627),
    .o1(n3958));
 b15aoi022ar1n12x5 U5204 (.a(net587),
    .b(net384),
    .c(net380),
    .d(net2087),
    .o1(n3957));
 b15aoi022as1n04x5 U5205 (.a(reg2hw_intr_ctrl_en_lvllow__q__21_),
    .b(net368),
    .c(n3413),
    .d(reg2hw_intr_enable__q__21_),
    .o1(n3956));
 b15aoi022al1n08x5 U5206 (.a(reg2hw_intr_ctrl_en_falling__q__21_),
    .b(net398),
    .c(net154),
    .d(net413),
    .o1(n3953));
 b15aob012ar1n08x5 U5207 (.a(n3953),
    .b(net434),
    .c(reg2hw_intr_state__q__21_),
    .out0(n3954));
 b15aoi112aq1n06x5 U5208 (.a(net354),
    .b(n3954),
    .c(reg2hw_intr_ctrl_en_rising__q__21_),
    .d(net442),
    .o1(n3955));
 b15nand04aq1n16x5 U5209 (.a(n3958),
    .b(net2088),
    .c(n3956),
    .d(n3955),
    .o1(u_reg_u_reg_if_N35));
 b15aoi022ah1n08x5 U5210 (.a(reg2hw_intr_ctrl_en_rising__q__22_),
    .b(net448),
    .c(net424),
    .d(reg2hw_intr_enable__q__22_),
    .o1(n3964));
 b15aoi022an1n32x5 U5211 (.a(net406),
    .b(net625),
    .c(net378),
    .d(net2205),
    .o1(n3963));
 b15aoi022as1n08x5 U5212 (.a(net586),
    .b(net383),
    .c(reg2hw_intr_ctrl_en_falling__q__22_),
    .d(net398),
    .o1(n3962));
 b15aoi022ar1n12x5 U5213 (.a(reg2hw_intr_ctrl_en_lvllow__q__22_),
    .b(net368),
    .c(net654),
    .d(net413),
    .o1(n3959));
 b15aob012as1n04x5 U5214 (.a(n3959),
    .b(net433),
    .c(reg2hw_intr_state__q__22_),
    .out0(n3960));
 b15aoi112al1n08x5 U5215 (.a(net353),
    .b(n3960),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__22_),
    .d(net440),
    .o1(n3961));
 b15nand04as1n16x5 U5216 (.a(n3964),
    .b(net2206),
    .c(n3962),
    .d(n3961),
    .o1(u_reg_u_reg_if_N36));
 b15aoi022as1n48x5 U5217 (.a(net408),
    .b(net624),
    .c(net651),
    .d(net414),
    .o1(n3971));
 b15aoi022an1n08x5 U5218 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__23_),
    .b(net440),
    .c(reg2hw_intr_ctrl_en_falling__q__23_),
    .d(net398),
    .o1(n3970));
 b15aoi022al1n12x5 U5219 (.a(reg2hw_intr_ctrl_en_rising__q__23_),
    .b(net448),
    .c(net378),
    .d(net2195),
    .o1(n3969));
 b15aoi022ar1n02x5 U5220 (.a(reg2hw_intr_ctrl_en_lvllow__q__23_),
    .b(net368),
    .c(net424),
    .d(reg2hw_intr_enable__q__23_),
    .o1(n3966));
 b15aob012ah1n04x5 U5221 (.a(n3966),
    .b(n3309),
    .c(reg2hw_intr_state__q__23_),
    .out0(n3967));
 b15aoi112an1n06x5 U5222 (.a(net353),
    .b(n3967),
    .c(net584),
    .d(net383),
    .o1(n3968));
 b15nand04as1n16x5 U5223 (.a(n3971),
    .b(n3970),
    .c(net2196),
    .d(n3968),
    .o1(u_reg_u_reg_if_N37));
 b15aoi022al1n32x5 U5225 (.a(n4175),
    .b(net189),
    .c(net380),
    .d(u_reg_data_in_qs[24]),
    .o1(n3979));
 b15aoi022aq1n08x5 U5226 (.a(reg2hw_intr_ctrl_en_falling__q__24_),
    .b(net395),
    .c(net421),
    .d(net521),
    .o1(n3978));
 b15aoi022aq1n08x5 U5227 (.a(reg2hw_intr_ctrl_en_rising__q__24_),
    .b(net442),
    .c(net157),
    .d(net413),
    .o1(n3977));
 b15aoi022ar1n12x5 U5228 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__24_),
    .b(net437),
    .c(reg2hw_intr_ctrl_en_lvllow__q__24_),
    .d(net368),
    .o1(n3973));
 b15aob012as1n06x5 U5229 (.a(n3973),
    .b(net434),
    .c(reg2hw_intr_state__q__24_),
    .out0(n3974));
 b15aoi112aq1n08x5 U5230 (.a(net354),
    .b(n3974),
    .c(reg2hw_ctrl_en_input_filter__q__24_),
    .d(net384),
    .o1(n3976));
 b15nand04as1n16x5 U5231 (.a(n3979),
    .b(net2221),
    .c(n3977),
    .d(n3976),
    .o1(u_reg_u_reg_if_N38));
 b15aoi022ar1n24x5 U5232 (.a(net158),
    .b(net413),
    .c(net417),
    .d(net520),
    .o1(n3986));
 b15aoi022al1n12x5 U5233 (.a(reg2hw_ctrl_en_input_filter__q__25_),
    .b(net384),
    .c(net380),
    .d(net2045),
    .o1(n3985));
 b15aoi022aq1n08x5 U5234 (.a(reg2hw_intr_ctrl_en_rising__q__25_),
    .b(net442),
    .c(reg2hw_intr_ctrl_en_falling__q__25_),
    .d(net398),
    .o1(n3984));
 b15aoi022al1n32x5 U5235 (.a(net534),
    .b(net368),
    .c(net409),
    .d(net190),
    .o1(n3980));
 b15aob012as1n03x5 U5236 (.a(n3980),
    .b(net434),
    .c(reg2hw_intr_state__q__25_),
    .out0(n3981));
 b15aoi112as1n04x5 U5237 (.a(net354),
    .b(n3981),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__25_),
    .d(net438),
    .o1(n3983));
 b15nand04as1n16x5 U5238 (.a(n3986),
    .b(net2046),
    .c(n3984),
    .d(n3983),
    .o1(u_reg_u_reg_if_N39));
 b15aoi022an1n16x5 U5239 (.a(net2400),
    .b(net437),
    .c(n3413),
    .d(reg2hw_intr_enable__q__26_),
    .o1(n3992));
 b15aoi022as1n32x5 U5240 (.a(net408),
    .b(net191),
    .c(net159),
    .d(net414),
    .o1(n3991));
 b15aoi022al1n12x5 U5241 (.a(reg2hw_intr_ctrl_en_lvllow__q__26_),
    .b(net368),
    .c(net380),
    .d(u_reg_data_in_qs[26]),
    .o1(n3990));
 b15aoi022al1n06x5 U5242 (.a(reg2hw_intr_ctrl_en_rising__q__26_),
    .b(net442),
    .c(reg2hw_intr_ctrl_en_falling__q__26_),
    .d(net395),
    .o1(n3987));
 b15aob012an1n12x5 U5243 (.a(n3987),
    .b(net434),
    .c(reg2hw_intr_state__q__26_),
    .out0(n3988));
 b15aoi112ah1n06x5 U5244 (.a(net354),
    .b(n3988),
    .c(reg2hw_ctrl_en_input_filter__q__26_),
    .d(net384),
    .o1(n3989));
 b15nand04as1n16x5 U5245 (.a(n3992),
    .b(n3991),
    .c(n3990),
    .d(n3989),
    .o1(u_reg_u_reg_if_N40));
 b15aoi022aq1n08x5 U5246 (.a(reg2hw_ctrl_en_input_filter__q__27_),
    .b(net384),
    .c(net417),
    .d(net519),
    .o1(n3998));
 b15aoi022an1n24x5 U5247 (.a(net405),
    .b(net192),
    .c(net377),
    .d(u_reg_data_in_qs[27]),
    .o1(n3997));
 b15aoi022ah1n06x5 U5248 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__27_),
    .b(net437),
    .c(net525),
    .d(net444),
    .o1(n3996));
 b15aoi022an1n12x5 U5249 (.a(net555),
    .b(net399),
    .c(net160),
    .d(net414),
    .o1(n3993));
 b15aob012as1n03x5 U5250 (.a(n3993),
    .b(net436),
    .c(reg2hw_intr_state__q__27_),
    .out0(n3994));
 b15aoi112ar1n08x5 U5251 (.a(net354),
    .b(n3994),
    .c(reg2hw_intr_ctrl_en_lvllow__q__27_),
    .d(net368),
    .o1(n3995));
 b15nand04as1n16x5 U5252 (.a(n3998),
    .b(n3997),
    .c(n3996),
    .d(n3995),
    .o1(u_reg_u_reg_if_N41));
 b15aoi022aq1n08x5 U5253 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__28_),
    .b(net440),
    .c(net424),
    .d(reg2hw_intr_enable__q__28_),
    .o1(n4005));
 b15aoi022aq1n12x5 U5254 (.a(net579),
    .b(net389),
    .c(net378),
    .d(net2062),
    .o1(n4004));
 b15aoi022as1n48x5 U5255 (.a(net410),
    .b(net617),
    .c(net645),
    .d(net412),
    .o1(n4003));
 b15aoi022ar1n02x3 U5256 (.a(reg2hw_intr_ctrl_en_lvllow__q__28_),
    .b(net368),
    .c(reg2hw_intr_ctrl_en_falling__q__28_),
    .d(net398),
    .o1(n3999));
 b15aob012an1n03x5 U5257 (.a(n3999),
    .b(net434),
    .c(reg2hw_intr_state__q__28_),
    .out0(n4000));
 b15aoi112an1n06x5 U5258 (.a(net353),
    .b(n4000),
    .c(reg2hw_intr_ctrl_en_rising__q__28_),
    .d(net448),
    .o1(n4002));
 b15nand04as1n16x5 U5259 (.a(n4005),
    .b(net2063),
    .c(n4003),
    .d(n4002),
    .o1(u_reg_u_reg_if_N42));
 b15aoi022aq1n48x5 U5260 (.a(net410),
    .b(net194),
    .c(net644),
    .d(net412),
    .o1(n4013));
 b15aoi022as1n06x5 U5261 (.a(reg2hw_intr_ctrl_en_rising__q__29_),
    .b(net449),
    .c(net424),
    .d(net2134),
    .o1(n4012));
 b15aoi022aq1n08x5 U5262 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__29_),
    .b(net440),
    .c(reg2hw_intr_ctrl_en_lvllow__q__29_),
    .d(net368),
    .o1(n4011));
 b15aoi022al1n04x5 U5263 (.a(reg2hw_intr_ctrl_en_falling__q__29_),
    .b(net398),
    .c(net378),
    .d(net2563),
    .o1(n4008));
 b15aob012ah1n03x5 U5264 (.a(n4008),
    .b(net433),
    .c(net510),
    .out0(n4009));
 b15aoi112aq1n08x5 U5265 (.a(net353),
    .b(n4009),
    .c(net578),
    .d(net387),
    .o1(n4010));
 b15nand04as1n16x5 U5266 (.a(n4013),
    .b(n4012),
    .c(n4011),
    .d(n4010),
    .o1(u_reg_u_reg_if_N43));
 b15aoi022ah1n08x5 U5267 (.a(net575),
    .b(net383),
    .c(net2269),
    .d(net398),
    .o1(n4023));
 b15aoi022an1n16x5 U5268 (.a(reg2hw_intr_ctrl_en_rising__q__30_),
    .b(net448),
    .c(net378),
    .d(net673),
    .o1(n4022));
 b15aoi022an1n06x5 U5269 (.a(net433),
    .b(reg2hw_intr_state__q__30_),
    .c(net424),
    .d(reg2hw_intr_enable__q__30_),
    .o1(n4020));
 b15aoi022as1n08x5 U5270 (.a(reg2hw_intr_ctrl_en_lvllow__q__30_),
    .b(net368),
    .c(net406),
    .d(net196),
    .o1(n4019));
 b15aoi022ar1n06x5 U5271 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__30_),
    .b(net440),
    .c(net164),
    .d(net413),
    .o1(n4018));
 b15and003ar1n08x5 U5272 (.a(n4020),
    .b(n4019),
    .c(n4018),
    .o(n4021));
 b15nand04as1n16x5 U5273 (.a(net356),
    .b(n4023),
    .c(n4022),
    .d(n4021),
    .o1(u_reg_u_reg_if_N44));
 b15aoi022as1n08x5 U5274 (.a(net643),
    .b(net413),
    .c(net424),
    .d(reg2hw_intr_enable__q__31_),
    .o1(n4041));
 b15aoi022as1n06x5 U5275 (.a(reg2hw_intr_ctrl_en_rising__q__31_),
    .b(net449),
    .c(reg2hw_intr_ctrl_en_falling__q__31_),
    .d(net395),
    .o1(n4040));
 b15aoi022ar1n16x5 U5276 (.a(reg2hw_intr_ctrl_en_lvllow__q__31_),
    .b(net368),
    .c(net379),
    .d(net2252),
    .o1(n4039));
 b15aoi022ah1n24x5 U5277 (.a(net545),
    .b(net440),
    .c(net406),
    .d(net197),
    .o1(n4033));
 b15aob012aq1n04x5 U5278 (.a(n4033),
    .b(net433),
    .c(reg2hw_intr_state__q__31_),
    .out0(n4035));
 b15aoi112ar1n08x5 U5279 (.a(net354),
    .b(n4035),
    .c(net573),
    .d(net383),
    .o1(n4038));
 b15nand04as1n16x5 U5280 (.a(n4041),
    .b(n4040),
    .c(n4039),
    .d(n4038),
    .o1(u_reg_u_reg_if_N45));
 b15oab012ar1n02x5 U5282 (.a(n4042),
    .b(net2560),
    .c(n4043),
    .out0(gen_filter_7__u_filter_diff_ctr_d[2]));
 b15nano23al1n08x5 U5283 (.a(net2279),
    .b(gen_filter_9__u_filter_diff_ctr_d[0]),
    .c(n4045),
    .d(n4044),
    .out0(eq_x_136_n25));
 b15nano23an1n12x5 U5284 (.a(gen_filter_18__u_filter_diff_ctr_d[1]),
    .b(gen_filter_18__u_filter_diff_ctr_d[0]),
    .c(n4047),
    .d(n4046),
    .out0(eq_x_91_n25));
 b15oab012ar1n02x5 U5285 (.a(n4048),
    .b(gen_filter_20__u_filter_diff_ctr_q[3]),
    .c(n4049),
    .out0(gen_filter_20__u_filter_diff_ctr_d[2]));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_0__cio_gpio_en_q_reg_1_ (.rb(net742),
    .clk(clknet_1_1__leaf_net2075),
    .d1(N114),
    .d2(N115),
    .o1(net141),
    .o2(net152),
    .si1(net761),
    .si2(net762),
    .ssb(net1500));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_10__cio_gpio_en_q_reg_11_ (.rb(net727),
    .clk(clknet_1_0__leaf_net2075),
    .d1(N124),
    .d2(N125),
    .o1(net142),
    .o2(net143),
    .si1(net763),
    .si2(net764),
    .ssb(net1501));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_12__cio_gpio_en_q_reg_13_ (.rb(net747),
    .clk(clknet_1_1__leaf_net2075),
    .d1(N126),
    .d2(N127),
    .o1(net144),
    .o2(net145),
    .si1(net765),
    .si2(net766),
    .ssb(net1502));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_14__cio_gpio_en_q_reg_15_ (.rb(net742),
    .clk(clknet_1_1__leaf_net2075),
    .d1(N128),
    .d2(N129),
    .o1(net146),
    .o2(net147),
    .si1(net767),
    .si2(net768),
    .ssb(net1503));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_16__cio_gpio_en_q_reg_17_ (.rb(net747),
    .clk(clknet_1_1__leaf_net2070),
    .d1(N131),
    .d2(N132),
    .o1(net148),
    .o2(net149),
    .si1(net769),
    .si2(net770),
    .ssb(net1504));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_18__cio_gpio_en_q_reg_19_ (.rb(net747),
    .clk(clknet_1_1__leaf_net2070),
    .d1(N133),
    .d2(N134),
    .o1(net150),
    .o2(net151),
    .si1(net771),
    .si2(net772),
    .ssb(net1505));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_20__cio_gpio_en_q_reg_21_ (.rb(net749),
    .clk(clknet_1_0__leaf_net2070),
    .d1(N135),
    .d2(N136),
    .o1(net153),
    .o2(net154),
    .si1(net773),
    .si2(net774),
    .ssb(net1506));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_22__cio_gpio_en_q_reg_23_ (.rb(net739),
    .clk(clknet_1_0__leaf_net2070),
    .d1(N137),
    .d2(N138),
    .o1(net155),
    .o2(net156),
    .si1(net775),
    .si2(net776),
    .ssb(net1507));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_24__cio_gpio_en_q_reg_25_ (.rb(net738),
    .clk(clknet_1_0__leaf_net2070),
    .d1(N139),
    .d2(N140),
    .o1(net157),
    .o2(net158),
    .si1(net777),
    .si2(net778),
    .ssb(net1508));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_26__cio_gpio_en_q_reg_27_ (.rb(net739),
    .clk(clknet_1_0__leaf_net2070),
    .d1(N141),
    .d2(N142),
    .o1(net159),
    .o2(net160),
    .si1(net779),
    .si2(net780),
    .ssb(net1509));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_28__cio_gpio_en_q_reg_29_ (.rb(net747),
    .clk(clknet_1_1__leaf_net2070),
    .d1(N143),
    .d2(N144),
    .o1(net161),
    .o2(net162),
    .si1(net781),
    .si2(net782),
    .ssb(net1510));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_2__cio_gpio_en_q_reg_3_ (.rb(net742),
    .clk(clknet_1_1__leaf_net2075),
    .d1(N116),
    .d2(N117),
    .o1(net163),
    .o2(net166),
    .si1(net783),
    .si2(net784),
    .ssb(net1511));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_30__cio_gpio_en_q_reg_31_ (.rb(net753),
    .clk(clknet_1_1__leaf_net2070),
    .d1(N145),
    .d2(N146),
    .o1(net164),
    .o2(net165),
    .si1(net785),
    .si2(net786),
    .ssb(net1512));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_4__cio_gpio_en_q_reg_5_ (.rb(net727),
    .clk(clknet_1_0__leaf_net2075),
    .d1(N118),
    .d2(N119),
    .o1(net167),
    .o2(net168),
    .si1(net787),
    .si2(net788),
    .ssb(net1513));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_6__cio_gpio_en_q_reg_7_ (.rb(net734),
    .clk(clknet_1_0__leaf_net2075),
    .d1(N120),
    .d2(net303),
    .o1(net169),
    .o2(net170),
    .si1(net789),
    .si2(net790),
    .ssb(net1514));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_8__cio_gpio_en_q_reg_9_ (.rb(net742),
    .clk(clknet_1_0__leaf_net2075),
    .d1(N122),
    .d2(N123),
    .o1(net171),
    .o2(net172),
    .si1(net791),
    .si2(net792),
    .ssb(net1515));
 b15fqy203ar1n02x5 cio_gpio_q_reg_0__cio_gpio_q_reg_1_ (.rb(net728),
    .clk(clknet_1_0__leaf_net2065),
    .d1(N39),
    .d2(N40),
    .o1(net173),
    .o2(net184),
    .si1(net793),
    .si2(net794),
    .ssb(net1516));
 b15fqy203ar1n02x5 cio_gpio_q_reg_10__cio_gpio_q_reg_11_ (.rb(net726),
    .clk(clknet_1_1__leaf_net2065),
    .d1(N49),
    .d2(N50),
    .o1(net174),
    .o2(net175),
    .si1(net795),
    .si2(net796),
    .ssb(net1517));
 b15fqy203ar1n02x5 cio_gpio_q_reg_12__cio_gpio_q_reg_13_ (.rb(net744),
    .clk(clknet_1_1__leaf_net2065),
    .d1(N51),
    .d2(N52),
    .o1(net176),
    .o2(net177),
    .si1(net797),
    .si2(net798),
    .ssb(net1518));
 b15fqy203ar1n02x5 cio_gpio_q_reg_14__cio_gpio_q_reg_15_ (.rb(net742),
    .clk(clknet_1_0__leaf_net2065),
    .d1(net299),
    .d2(N54),
    .o1(net178),
    .o2(net179),
    .si1(net799),
    .si2(net800),
    .ssb(net1519));
 b15fqy203ar1n02x5 cio_gpio_q_reg_16__cio_gpio_q_reg_17_ (.rb(net747),
    .clk(clknet_1_0__leaf_net2059),
    .d1(N56),
    .d2(N57),
    .o1(net180),
    .o2(net181),
    .si1(net801),
    .si2(net802),
    .ssb(net1520));
 b15fqy203ar1n02x5 cio_gpio_q_reg_18__cio_gpio_q_reg_19_ (.rb(net728),
    .clk(clknet_1_1__leaf_net2059),
    .d1(N58),
    .d2(N59),
    .o1(net182),
    .o2(net183),
    .si1(net803),
    .si2(net804),
    .ssb(net1521));
 b15fqy203ar1n02x5 cio_gpio_q_reg_20__cio_gpio_q_reg_21_ (.rb(net739),
    .clk(clknet_1_0__leaf_net2059),
    .d1(N60),
    .d2(N61),
    .o1(net185),
    .o2(net186),
    .si1(net805),
    .si2(net806),
    .ssb(net1522));
 b15fqy203ar1n02x5 cio_gpio_q_reg_22__cio_gpio_q_reg_23_ (.rb(net739),
    .clk(clknet_1_1__leaf_net2059),
    .d1(N62),
    .d2(N63),
    .o1(net187),
    .o2(net188),
    .si1(net807),
    .si2(net808),
    .ssb(net1523));
 b15fqy203ar1n02x5 cio_gpio_q_reg_24__cio_gpio_q_reg_25_ (.rb(net736),
    .clk(clknet_1_1__leaf_net2059),
    .d1(N64),
    .d2(net301),
    .o1(net189),
    .o2(net190),
    .si1(net809),
    .si2(net810),
    .ssb(net1524));
 b15fqy203ar1n02x5 cio_gpio_q_reg_26__cio_gpio_q_reg_27_ (.rb(net739),
    .clk(clknet_1_1__leaf_net2059),
    .d1(N66),
    .d2(N67),
    .o1(net191),
    .o2(net192),
    .si1(net811),
    .si2(net812),
    .ssb(net1525));
 b15fqy203ar1n02x5 cio_gpio_q_reg_28__cio_gpio_q_reg_29_ (.rb(net747),
    .clk(clknet_1_0__leaf_net2059),
    .d1(N68),
    .d2(N69),
    .o1(net193),
    .o2(net194),
    .si1(net813),
    .si2(net814),
    .ssb(net1526));
 b15fqy203ar1n02x5 cio_gpio_q_reg_2__cio_gpio_q_reg_3_ (.rb(net742),
    .clk(clknet_1_0__leaf_net2065),
    .d1(N41),
    .d2(N42),
    .o1(net195),
    .o2(net198),
    .si1(net815),
    .si2(net816),
    .ssb(net1527));
 b15fqy203ar1n02x5 cio_gpio_q_reg_30__cio_gpio_q_reg_31_ (.rb(net753),
    .clk(clknet_1_0__leaf_net2059),
    .d1(N70),
    .d2(N71),
    .o1(net196),
    .o2(net197),
    .si1(net817),
    .si2(net818),
    .ssb(net1528));
 b15fqy203ar1n02x5 cio_gpio_q_reg_4__cio_gpio_q_reg_5_ (.rb(net726),
    .clk(clknet_1_1__leaf_net2065),
    .d1(N43),
    .d2(N44),
    .o1(net199),
    .o2(net200),
    .si1(net819),
    .si2(net820),
    .ssb(net1529));
 b15fqy203ar1n02x5 cio_gpio_q_reg_6__cio_gpio_q_reg_7_ (.rb(net726),
    .clk(clknet_1_1__leaf_net2065),
    .d1(N45),
    .d2(N46),
    .o1(net201),
    .o2(net202),
    .si1(net821),
    .si2(net822),
    .ssb(net1530));
 b15fqy203ar1n02x5 cio_gpio_q_reg_8__cio_gpio_q_reg_9_ (.rb(net742),
    .clk(clknet_1_0__leaf_net2065),
    .d1(N47),
    .d2(N48),
    .o1(net203),
    .o2(net204),
    .si1(net823),
    .si2(net824),
    .ssb(net1531));
 b15cilb05ah1n02x3 clk_gate_cio_gpio_en_q_reg_0_latch (.clk(clknet_leaf_11_clk_i),
    .clkout(net2075),
    .en(net343),
    .te(net825));
 b15cilb05ah1n02x3 clk_gate_cio_gpio_en_q_reg_latch (.clk(clknet_leaf_7_clk_i),
    .clkout(net2070),
    .en(N130),
    .te(net826));
 b15cilb05ah1n02x3 clk_gate_cio_gpio_q_reg_0_latch (.clk(clknet_leaf_12_clk_i),
    .clkout(net2065),
    .en(net300),
    .te(net827));
 b15cilb05ah1n02x3 clk_gate_cio_gpio_q_reg_latch (.clk(clknet_leaf_1_clk_i),
    .clkout(net2059),
    .en(N55),
    .te(net828));
 b15fpy200ar1n02x5 data_in_q_reg_0__data_in_q_reg_1_ (.clk(clknet_leaf_11_clk_i),
    .d1(net365),
    .d2(u_reg_u_data_in_wr_data[1]),
    .o1(data_in_q[0]),
    .o2(data_in_q[1]),
    .si1(net829),
    .si2(net830),
    .ssb(net1532));
 b15fpy200ar1n02x5 data_in_q_reg_10__data_in_q_reg_11_ (.clk(clknet_leaf_0_clk_i),
    .d1(u_reg_u_data_in_wr_data[10]),
    .d2(u_reg_u_data_in_wr_data[11]),
    .o1(data_in_q[10]),
    .o2(data_in_q[11]),
    .si1(net831),
    .si2(net832),
    .ssb(net1533));
 b15fpy200ar1n02x5 data_in_q_reg_12__data_in_q_reg_13_ (.clk(clknet_leaf_8_clk_i),
    .d1(u_reg_u_data_in_wr_data[12]),
    .d2(u_reg_u_data_in_wr_data[13]),
    .o1(data_in_q[12]),
    .o2(data_in_q[13]),
    .si1(net833),
    .si2(net834),
    .ssb(net1534));
 b15fpy200ar1n02x5 data_in_q_reg_14__data_in_q_reg_15_ (.clk(clknet_leaf_8_clk_i),
    .d1(u_reg_u_data_in_wr_data[14]),
    .d2(u_reg_u_data_in_wr_data[15]),
    .o1(data_in_q[14]),
    .o2(data_in_q[15]),
    .si1(net835),
    .si2(net836),
    .ssb(net1535));
 b15fpy200ar1n02x5 data_in_q_reg_16__data_in_q_reg_17_ (.clk(clknet_leaf_9_clk_i),
    .d1(u_reg_u_data_in_wr_data[16]),
    .d2(u_reg_u_data_in_wr_data[17]),
    .o1(data_in_q[16]),
    .o2(data_in_q[17]),
    .si1(net837),
    .si2(net838),
    .ssb(net1536));
 b15fpy200ar1n02x5 data_in_q_reg_18__data_in_q_reg_19_ (.clk(clknet_leaf_7_clk_i),
    .d1(u_reg_u_data_in_wr_data[18]),
    .d2(u_reg_u_data_in_wr_data[19]),
    .o1(data_in_q[18]),
    .o2(data_in_q[19]),
    .si1(net839),
    .si2(net840),
    .ssb(net1537));
 b15fpy200ar1n02x5 data_in_q_reg_20__data_in_q_reg_21_ (.clk(clknet_leaf_4_clk_i),
    .d1(u_reg_u_data_in_wr_data[20]),
    .d2(u_reg_u_data_in_wr_data[21]),
    .o1(data_in_q[20]),
    .o2(data_in_q[21]),
    .si1(net841),
    .si2(net842),
    .ssb(net1538));
 b15fpy200ar1n02x5 data_in_q_reg_22__data_in_q_reg_23_ (.clk(clknet_leaf_6_clk_i),
    .d1(u_reg_u_data_in_wr_data[22]),
    .d2(u_reg_u_data_in_wr_data[23]),
    .o1(data_in_q[22]),
    .o2(data_in_q[23]),
    .si1(net843),
    .si2(net844),
    .ssb(net1539));
 b15fpy200ar1n02x5 data_in_q_reg_24__data_in_q_reg_25_ (.clk(clknet_leaf_4_clk_i),
    .d1(u_reg_u_data_in_wr_data[24]),
    .d2(u_reg_u_data_in_wr_data[25]),
    .o1(data_in_q[24]),
    .o2(data_in_q[25]),
    .si1(net845),
    .si2(net846),
    .ssb(net1540));
 b15fpy200ar1n02x5 data_in_q_reg_26__data_in_q_reg_27_ (.clk(clknet_leaf_3_clk_i),
    .d1(u_reg_u_data_in_wr_data[26]),
    .d2(u_reg_u_data_in_wr_data[27]),
    .o1(data_in_q[26]),
    .o2(data_in_q[27]),
    .si1(net847),
    .si2(net848),
    .ssb(net1541));
 b15fpy200ar1n02x5 data_in_q_reg_28__data_in_q_reg_29_ (.clk(clknet_leaf_6_clk_i),
    .d1(u_reg_u_data_in_wr_data[28]),
    .d2(u_reg_u_data_in_wr_data[29]),
    .o1(data_in_q[28]),
    .o2(data_in_q[29]),
    .si1(net849),
    .si2(net850),
    .ssb(net1542));
 b15fpy200ar1n02x5 data_in_q_reg_2__data_in_q_reg_3_ (.clk(clknet_leaf_11_clk_i),
    .d1(u_reg_u_data_in_wr_data[2]),
    .d2(u_reg_u_data_in_wr_data[3]),
    .o1(data_in_q[2]),
    .o2(data_in_q[3]),
    .si1(net851),
    .si2(net852),
    .ssb(net1543));
 b15fpy200ar1n02x5 data_in_q_reg_30__data_in_q_reg_31_ (.clk(clknet_leaf_4_clk_i),
    .d1(u_reg_u_data_in_wr_data[30]),
    .d2(u_reg_u_data_in_wr_data[31]),
    .o1(data_in_q[30]),
    .o2(data_in_q[31]),
    .si1(net853),
    .si2(net854),
    .ssb(net1544));
 b15fpy200ar1n02x5 data_in_q_reg_4__data_in_q_reg_5_ (.clk(clknet_leaf_0_clk_i),
    .d1(u_reg_u_data_in_wr_data[4]),
    .d2(u_reg_u_data_in_wr_data[5]),
    .o1(data_in_q[4]),
    .o2(data_in_q[5]),
    .si1(net855),
    .si2(net856),
    .ssb(net1545));
 b15fpy200ar1n02x5 data_in_q_reg_6__data_in_q_reg_7_ (.clk(clknet_leaf_0_clk_i),
    .d1(u_reg_u_data_in_wr_data[6]),
    .d2(net364),
    .o1(data_in_q[6]),
    .o2(data_in_q[7]),
    .si1(net857),
    .si2(net858),
    .ssb(net1546));
 b15fpy200ar1n02x5 data_in_q_reg_8__data_in_q_reg_9_ (.clk(clknet_leaf_11_clk_i),
    .d1(u_reg_u_data_in_wr_data[8]),
    .d2(u_reg_u_data_in_wr_data[9]),
    .o1(data_in_q[8]),
    .o2(data_in_q[9]),
    .si1(net859),
    .si2(net860),
    .ssb(net1547));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg (.rb(net726),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger),
    .d2(gen_alert_tx_0__u_prim_alert_sender_alert_test_set_d),
    .o1(gen_alert_tx_0__u_prim_alert_sender_n1),
    .o2(gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q),
    .si1(net861),
    .si2(net862),
    .ssb(net1548));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg (.rb(net734),
    .clk(clknet_leaf_1_clk_i),
    .d1(gen_alert_tx_0__u_prim_alert_sender_ping_set_d),
    .d2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .o1(gen_alert_tx_0__u_prim_alert_sender_ping_set_q),
    .o2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq),
    .si1(net863),
    .si2(net864),
    .ssb(net1549));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0__gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1_ (.rb(net727),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_alert_tx_0__u_prim_alert_sender_state_d[0]),
    .d2(gen_alert_tx_0__u_prim_alert_sender_state_d[1]),
    .o1(gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .o2(gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .si1(net865),
    .si2(net866),
    .ssb(net1550));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net727),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_alert_tx_0__u_prim_alert_sender_state_d[2]),
    .d2(net2),
    .o1(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .o2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_intq_0_),
    .si1(net867),
    .si2(net868),
    .ssb(net1551));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq_reg (.clk(clknet_leaf_1_clk_i),
    .d(net2377),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq),
    .psb(net734),
    .si(net869),
    .ssb(net1552));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_1_clk_i),
    .d(net1),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_intq_0_),
    .psb(net734),
    .si(net870),
    .ssb(net1553));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_1_clk_i),
    .d(net2212),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd),
    .psb(net734),
    .si(net871),
    .ssb(net1554));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg (.rb(net734),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2149),
    .d2(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .o2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q),
    .si1(net872),
    .si2(net873),
    .ssb(net1555));
 b15fqy043ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_0_ (.clk(clknet_leaf_1_clk_i),
    .d(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[0]),
    .den(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[0]),
    .rb(net734),
    .si(net874),
    .ssb(net1556));
 b15fqy043ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_1_ (.clk(clknet_leaf_1_clk_i),
    .d(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[1]),
    .den(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .rb(net734),
    .si(net875),
    .ssb(net1557));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq_reg (.clk(clknet_leaf_14_clk_i),
    .d(net2479),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq),
    .psb(net727),
    .si(net876),
    .ssb(net1558));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net727),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2440),
    .d2(net4),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq),
    .o2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_intq_0_),
    .si1(net877),
    .si2(net878),
    .ssb(net1559));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_0_clk_i),
    .d(net3),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_intq_0_),
    .psb(net726),
    .si(net879),
    .ssb(net1560));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_14_clk_i),
    .d(net2125),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .psb(net726),
    .si(net880),
    .ssb(net1561));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg (.rb(net727),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2198),
    .d2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_n3),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .o2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q),
    .si1(net881),
    .si2(net882),
    .ssb(net1562));
 b15fqy043ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_0_ (.clk(clknet_leaf_14_clk_i),
    .d(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[0]),
    .den(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .rb(net727),
    .si(net883),
    .ssb(net1563));
 b15fqy043ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_1_ (.clk(clknet_leaf_14_clk_i),
    .d(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[1]),
    .den(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .rb(net727),
    .si(net884),
    .ssb(net1564));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net727),
    .clk(clknet_leaf_14_clk_i),
    .d1(gen_alert_tx_0__u_prim_alert_sender_alert_pd),
    .d2(net32),
    .o1(net140),
    .o2(gen_filter_5__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net885),
    .si2(net886),
    .ssb(net1565));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_1_ (.clk(clknet_leaf_0_clk_i),
    .d(gen_alert_tx_0__u_prim_alert_sender_alert_nd),
    .o(net139),
    .psb(net727),
    .si(net887),
    .ssb(net1566));
 b15fqy203ar1n02x5 gen_filter_0__u_filter_diff_ctr_q_reg_0__gen_filter_0__u_filter_diff_ctr_q_reg_1_ (.rb(net725),
    .clk(clknet_leaf_13_clk_i),
    .d1(net2305),
    .d2(gen_filter_0__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_0__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_0__u_filter_diff_ctr_q[1]),
    .si1(net888),
    .si2(net889),
    .ssb(net1567));
 b15fqy203ar1n02x5 gen_filter_0__u_filter_diff_ctr_q_reg_2__gen_filter_0__u_filter_diff_ctr_q_reg_3_ (.rb(net725),
    .clk(clknet_leaf_13_clk_i),
    .d1(net2404),
    .d2(net2303),
    .o1(gen_filter_0__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_0__u_filter_diff_ctr_q[3]),
    .si1(net890),
    .si2(net891),
    .ssb(net1568));
 b15fqy203ar1n02x5 gen_filter_0__u_filter_filter_q_reg_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net725),
    .clk(clknet_leaf_13_clk_i),
    .d1(gen_filter_0__u_filter_filter_synced),
    .d2(net5),
    .o1(gen_filter_0__u_filter_filter_q),
    .o2(gen_filter_0__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net892),
    .si2(net893),
    .ssb(net1569));
 b15fqy203ar1n02x5 gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_1__u_filter_diff_ctr_q_reg_0_ (.rb(net725),
    .clk(clknet_leaf_13_clk_i),
    .d1(net2210),
    .d2(net2388),
    .o1(gen_filter_0__u_filter_filter_synced),
    .o2(gen_filter_1__u_filter_diff_ctr_q[0]),
    .si1(net894),
    .si2(net895),
    .ssb(net1570));
 b15fqy043ar1n02x5 gen_filter_0__u_filter_stored_value_q_reg (.clk(clknet_leaf_13_clk_i),
    .d(gen_filter_0__u_filter_filter_synced),
    .den(eq_x_181_n25),
    .o(gen_filter_0__u_filter_stored_value_q),
    .rb(net725),
    .si(net896),
    .ssb(net1571));
 b15fqy203ar1n02x5 gen_filter_10__u_filter_diff_ctr_q_reg_1__gen_filter_10__u_filter_diff_ctr_q_reg_2_ (.rb(net725),
    .clk(clknet_leaf_13_clk_i),
    .d1(net2250),
    .d2(net2233),
    .o1(gen_filter_10__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_10__u_filter_diff_ctr_q[2]),
    .si1(net897),
    .si2(net898),
    .ssb(net1572));
 b15fqy203ar1n02x5 gen_filter_10__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_filter_q_reg (.rb(net725),
    .clk(clknet_leaf_14_clk_i),
    .d1(gen_filter_10__u_filter_diff_ctr_d[3]),
    .d2(net2273),
    .o1(gen_filter_10__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_10__u_filter_filter_q),
    .si1(net899),
    .si2(net900),
    .ssb(net1573));
 b15fqy203ar1n02x5 gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net725),
    .clk(clknet_leaf_14_clk_i),
    .d1(net6),
    .d2(net2166),
    .o1(gen_filter_10__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_10__u_filter_filter_synced),
    .si1(net901),
    .si2(net902),
    .ssb(net1574));
 b15fqy043ar1n02x5 gen_filter_10__u_filter_stored_value_q_reg (.clk(clknet_leaf_14_clk_i),
    .d(net2273),
    .den(eq_x_131_n25),
    .o(gen_filter_10__u_filter_stored_value_q),
    .rb(net725),
    .si(net903),
    .ssb(net1575));
 b15fqy203ar1n02x5 gen_filter_11__u_filter_diff_ctr_q_reg_0__gen_filter_12__u_filter_diff_ctr_q_reg_0_ (.rb(net742),
    .clk(clknet_leaf_10_clk_i),
    .d1(gen_filter_11__u_filter_diff_ctr_d[0]),
    .d2(net2428),
    .o1(gen_filter_11__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_12__u_filter_diff_ctr_q[0]),
    .si1(net904),
    .si2(net905),
    .ssb(net1576));
 b15fqy203ar1n02x5 gen_filter_11__u_filter_diff_ctr_q_reg_2__gen_filter_11__u_filter_diff_ctr_q_reg_3_ (.rb(net742),
    .clk(clknet_leaf_10_clk_i),
    .d1(net2406),
    .d2(net2349),
    .o1(gen_filter_11__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_11__u_filter_diff_ctr_q[3]),
    .si1(net906),
    .si2(net907),
    .ssb(net1577));
 b15fqy203ar1n02x5 gen_filter_11__u_filter_filter_q_reg_gen_filter_12__u_filter_filter_q_reg (.rb(net743),
    .clk(clknet_leaf_10_clk_i),
    .d1(gen_filter_11__u_filter_filter_synced),
    .d2(gen_filter_12__u_filter_filter_synced),
    .o1(gen_filter_11__u_filter_filter_q),
    .o2(gen_filter_12__u_filter_filter_q),
    .si1(net908),
    .si2(net909),
    .ssb(net1578));
 b15fqy203ar1n02x5 gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_3_ (.rb(net742),
    .clk(clknet_leaf_11_clk_i),
    .d1(net2297),
    .d2(net2443),
    .o1(gen_filter_11__u_filter_filter_synced),
    .o2(gen_filter_14__u_filter_diff_ctr_q[3]),
    .si1(net910),
    .si2(net911),
    .ssb(net1579));
 b15fqy043ar1n02x5 gen_filter_11__u_filter_stored_value_q_reg (.clk(clknet_leaf_11_clk_i),
    .d(gen_filter_11__u_filter_filter_synced),
    .den(eq_x_126_n25),
    .o(gen_filter_11__u_filter_stored_value_q),
    .rb(net742),
    .si(net912),
    .ssb(net1580));
 b15fqy203ar1n02x5 gen_filter_12__u_filter_diff_ctr_q_reg_1__gen_filter_12__u_filter_diff_ctr_q_reg_2_ (.rb(net746),
    .clk(clknet_leaf_10_clk_i),
    .d1(net2361),
    .d2(net2408),
    .o1(gen_filter_12__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_12__u_filter_diff_ctr_q[2]),
    .si1(net913),
    .si2(net914),
    .ssb(net1581));
 b15fqy203ar1n02x5 gen_filter_12__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_diff_ctr_q_reg_0_ (.rb(net746),
    .clk(clknet_leaf_10_clk_i),
    .d1(gen_filter_12__u_filter_diff_ctr_d[3]),
    .d2(net2365),
    .o1(gen_filter_12__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_13__u_filter_diff_ctr_q[0]),
    .si1(net915),
    .si2(net916),
    .ssb(net1582));
 b15fqy203ar1n02x5 gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net743),
    .clk(clknet_leaf_10_clk_i),
    .d1(net8),
    .d2(net2167),
    .o1(gen_filter_12__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_12__u_filter_filter_synced),
    .si1(net917),
    .si2(net918),
    .ssb(net1583));
 b15fqy043ar1n02x5 gen_filter_12__u_filter_stored_value_q_reg (.clk(clknet_leaf_10_clk_i),
    .d(gen_filter_12__u_filter_filter_synced),
    .den(eq_x_121_n25),
    .o(gen_filter_12__u_filter_stored_value_q),
    .rb(net743),
    .si(net919),
    .ssb(net1584));
 b15fqy203ar1n02x5 gen_filter_13__u_filter_diff_ctr_q_reg_1__gen_filter_13__u_filter_diff_ctr_q_reg_2_ (.rb(net746),
    .clk(clknet_leaf_10_clk_i),
    .d1(net2325),
    .d2(gen_filter_13__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_13__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_13__u_filter_diff_ctr_q[2]),
    .si1(net920),
    .si2(net921),
    .ssb(net1585));
 b15fqy203ar1n02x5 gen_filter_13__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_filter_q_reg (.rb(net746),
    .clk(clknet_leaf_10_clk_i),
    .d1(gen_filter_13__u_filter_diff_ctr_d[3]),
    .d2(net2471),
    .o1(gen_filter_13__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_13__u_filter_filter_q),
    .si1(net922),
    .si2(net923),
    .ssb(net1586));
 b15fqy203ar1n02x5 gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net743),
    .clk(clknet_leaf_10_clk_i),
    .d1(net9),
    .d2(net2169),
    .o1(gen_filter_13__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_13__u_filter_filter_synced),
    .si1(net924),
    .si2(net925),
    .ssb(net1587));
 b15fqy043ar1n02x5 gen_filter_13__u_filter_stored_value_q_reg (.clk(clknet_leaf_10_clk_i),
    .d(gen_filter_13__u_filter_filter_synced),
    .den(eq_x_116_n25),
    .o(gen_filter_13__u_filter_stored_value_q),
    .rb(net746),
    .si(net926),
    .ssb(net1588));
 b15fqy203ar1n02x5 gen_filter_14__u_filter_diff_ctr_q_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_1_ (.rb(net728),
    .clk(clknet_leaf_12_clk_i),
    .d1(gen_filter_14__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_14__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_14__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_14__u_filter_diff_ctr_q[1]),
    .si1(net927),
    .si2(net928),
    .ssb(net1589));
 b15fqy203ar1n02x5 gen_filter_14__u_filter_diff_ctr_q_reg_2__gen_filter_26__u_filter_diff_ctr_q_reg_0_ (.rb(net726),
    .clk(clknet_leaf_0_clk_i),
    .d1(net360),
    .d2(gen_filter_26__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_14__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_26__u_filter_diff_ctr_q[0]),
    .si1(net929),
    .si2(net930),
    .ssb(net1590));
 b15fqy203ar1n02x5 gen_filter_14__u_filter_filter_q_reg_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net743),
    .clk(clknet_leaf_11_clk_i),
    .d1(net2380),
    .d2(net10),
    .o1(gen_filter_14__u_filter_filter_q),
    .o2(gen_filter_14__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net931),
    .si2(net932),
    .ssb(net1591));
 b15fqy203ar1n02x5 gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_diff_ctr_q_reg_0_ (.rb(net743),
    .clk(clknet_leaf_10_clk_i),
    .d1(net2145),
    .d2(net2154),
    .o1(gen_filter_14__u_filter_filter_synced),
    .o2(gen_filter_15__u_filter_diff_ctr_q[0]),
    .si1(net933),
    .si2(net934),
    .ssb(net1592));
 b15fqy043ar1n02x5 gen_filter_14__u_filter_stored_value_q_reg (.clk(clknet_leaf_11_clk_i),
    .d(gen_filter_14__u_filter_filter_synced),
    .den(eq_x_111_n25),
    .o(gen_filter_14__u_filter_stored_value_q),
    .rb(net743),
    .si(net935),
    .ssb(net1593));
 b15fqy203ar1n02x5 gen_filter_15__u_filter_diff_ctr_q_reg_1__gen_filter_15__u_filter_diff_ctr_q_reg_2_ (.rb(net746),
    .clk(clknet_leaf_10_clk_i),
    .d1(net2204),
    .d2(net2182),
    .o1(gen_filter_15__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_15__u_filter_diff_ctr_q[2]),
    .si1(net936),
    .si2(net937),
    .ssb(net1594));
 b15fqy203ar1n02x5 gen_filter_15__u_filter_filter_q_reg_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net746),
    .clk(clknet_leaf_10_clk_i),
    .d1(net2278),
    .d2(net11),
    .o1(gen_filter_15__u_filter_filter_q),
    .o2(gen_filter_15__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net938),
    .si2(net939),
    .ssb(net1595));
 b15fqy203ar1n02x5 gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_diff_ctr_q_reg_0_ (.rb(net746),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2457),
    .d2(net2277),
    .o1(gen_filter_15__u_filter_filter_synced),
    .o2(gen_filter_19__u_filter_diff_ctr_q[0]),
    .si1(net940),
    .si2(net941),
    .ssb(net1596));
 b15fqy043ar1n02x5 gen_filter_15__u_filter_stored_value_q_reg (.clk(clknet_leaf_10_clk_i),
    .d(net2278),
    .den(eq_x_106_n25),
    .o(gen_filter_15__u_filter_stored_value_q),
    .rb(net743),
    .si(net942),
    .ssb(net1597));
 b15fqy203ar1n02x5 gen_filter_16__u_filter_diff_ctr_q_reg_0__gen_filter_16__u_filter_diff_ctr_q_reg_1_ (.rb(net747),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2322),
    .d2(net2347),
    .o1(gen_filter_16__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_16__u_filter_diff_ctr_q[1]),
    .si1(net943),
    .si2(net944),
    .ssb(net1598));
 b15fqy203ar1n02x5 gen_filter_16__u_filter_diff_ctr_q_reg_2__gen_filter_16__u_filter_diff_ctr_q_reg_3_ (.rb(net748),
    .clk(clknet_leaf_9_clk_i),
    .d1(gen_filter_16__u_filter_diff_ctr_d[2]),
    .d2(net2334),
    .o1(gen_filter_16__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_16__u_filter_diff_ctr_q[3]),
    .si1(net945),
    .si2(net946),
    .ssb(net1599));
 b15fqy203ar1n02x5 gen_filter_16__u_filter_filter_q_reg_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net748),
    .clk(clknet_leaf_9_clk_i),
    .d1(gen_filter_16__u_filter_filter_synced),
    .d2(net12),
    .o1(gen_filter_16__u_filter_filter_q),
    .o2(gen_filter_16__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net947),
    .si2(net948),
    .ssb(net1600));
 b15fqy203ar1n02x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net748),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2190),
    .d2(net13),
    .o1(gen_filter_16__u_filter_filter_synced),
    .o2(gen_filter_17__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net949),
    .si2(net950),
    .ssb(net1601));
 b15fqy043ar1n02x5 gen_filter_16__u_filter_stored_value_q_reg (.clk(clknet_leaf_9_clk_i),
    .d(gen_filter_16__u_filter_filter_synced),
    .den(eq_x_101_n25),
    .o(gen_filter_16__u_filter_stored_value_q),
    .rb(net747),
    .si(net951),
    .ssb(net1602));
 b15fqy203ar1n02x5 gen_filter_17__u_filter_diff_ctr_q_reg_1__gen_filter_17__u_filter_diff_ctr_q_reg_2_ (.rb(net746),
    .clk(clknet_leaf_10_clk_i),
    .d1(net2123),
    .d2(net2156),
    .o1(gen_filter_17__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_17__u_filter_diff_ctr_q[2]),
    .si1(net952),
    .si2(net953),
    .ssb(net1603));
 b15fqy203ar1n02x5 gen_filter_17__u_filter_diff_ctr_q_reg_3__gen_filter_17__u_filter_filter_q_reg (.rb(net746),
    .clk(clknet_leaf_9_clk_i),
    .d1(gen_filter_17__u_filter_diff_ctr_d[3]),
    .d2(gen_filter_17__u_filter_filter_synced),
    .o1(gen_filter_17__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_17__u_filter_filter_q),
    .si1(net954),
    .si2(net955),
    .ssb(net1604));
 b15fqy203ar1n02x5 gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_18__u_filter_diff_ctr_q_reg_0_ (.rb(net748),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2292),
    .d2(net2423),
    .o1(gen_filter_17__u_filter_filter_synced),
    .o2(gen_filter_18__u_filter_diff_ctr_q[0]),
    .si1(net956),
    .si2(net957),
    .ssb(net1605));
 b15fqy043ar1n02x5 gen_filter_17__u_filter_stored_value_q_reg (.clk(clknet_leaf_9_clk_i),
    .d(gen_filter_17__u_filter_filter_synced),
    .den(eq_x_96_n25),
    .o(gen_filter_17__u_filter_stored_value_q),
    .rb(net746),
    .si(net958),
    .ssb(net1606));
 b15fqy203ar1n02x5 gen_filter_18__u_filter_diff_ctr_q_reg_1__gen_filter_18__u_filter_diff_ctr_q_reg_2_ (.rb(net748),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2357),
    .d2(net2309),
    .o1(gen_filter_18__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_18__u_filter_diff_ctr_q[2]),
    .si1(net959),
    .si2(net960),
    .ssb(net1607));
 b15fqy203ar1n02x5 gen_filter_18__u_filter_diff_ctr_q_reg_3__gen_filter_18__u_filter_filter_q_reg (.rb(net748),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2418),
    .d2(gen_filter_18__u_filter_filter_synced),
    .o1(gen_filter_18__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_18__u_filter_filter_q),
    .si1(net961),
    .si2(net962),
    .ssb(net1608));
 b15fqy203ar1n02x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net755),
    .clk(clknet_leaf_5_clk_i),
    .d1(net14),
    .d2(net28),
    .o1(gen_filter_18__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_30__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net963),
    .si2(net964),
    .ssb(net1609));
 b15fqy203ar1n02x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net753),
    .clk(clknet_leaf_6_clk_i),
    .d1(gen_filter_18__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .d2(net2226),
    .o1(gen_filter_18__u_filter_filter_synced),
    .o2(gen_filter_19__u_filter_filter_synced),
    .si1(net965),
    .si2(net966),
    .ssb(net1610));
 b15fqy043ar1n02x5 gen_filter_18__u_filter_stored_value_q_reg (.clk(clknet_leaf_7_clk_i),
    .d(gen_filter_18__u_filter_filter_synced),
    .den(eq_x_91_n25),
    .o(gen_filter_18__u_filter_stored_value_q),
    .rb(net753),
    .si(net967),
    .ssb(net1611));
 b15fqy203ar1n02x5 gen_filter_19__u_filter_diff_ctr_q_reg_1__gen_filter_19__u_filter_diff_ctr_q_reg_2_ (.rb(net747),
    .clk(clknet_leaf_9_clk_i),
    .d1(gen_filter_19__u_filter_diff_ctr_d[1]),
    .d2(gen_filter_19__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_19__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_19__u_filter_diff_ctr_q[2]),
    .si1(net968),
    .si2(net969),
    .ssb(net1612));
 b15fqy203ar1n02x5 gen_filter_19__u_filter_diff_ctr_q_reg_3__gen_filter_19__u_filter_filter_q_reg (.rb(net747),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2296),
    .d2(net686),
    .o1(gen_filter_19__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_19__u_filter_filter_q),
    .si1(net970),
    .si2(net971),
    .ssb(net1613));
 b15fqy203ar1n02x5 gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net755),
    .clk(clknet_leaf_6_clk_i),
    .d1(net15),
    .d2(net17),
    .o1(gen_filter_19__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_20__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net972),
    .si2(net973),
    .ssb(net1614));
 b15fqy043ar1n02x5 gen_filter_19__u_filter_stored_value_q_reg (.clk(clknet_leaf_9_clk_i),
    .d(net686),
    .den(eq_x_86_n25),
    .o(gen_filter_19__u_filter_stored_value_q),
    .rb(net747),
    .si(net974),
    .ssb(net1615));
 b15fqy203ar1n02x5 gen_filter_1__u_filter_diff_ctr_q_reg_1__gen_filter_1__u_filter_diff_ctr_q_reg_2_ (.rb(net728),
    .clk(clknet_leaf_13_clk_i),
    .d1(net2413),
    .d2(net2371),
    .o1(gen_filter_1__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_1__u_filter_diff_ctr_q[2]),
    .si1(net975),
    .si2(net976),
    .ssb(net1616));
 b15fqy203ar1n02x5 gen_filter_1__u_filter_diff_ctr_q_reg_3__gen_filter_1__u_filter_filter_q_reg (.rb(net728),
    .clk(clknet_leaf_13_clk_i),
    .d1(gen_filter_1__u_filter_diff_ctr_d[3]),
    .d2(net2468),
    .o1(gen_filter_1__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_1__u_filter_filter_q),
    .si1(net977),
    .si2(net978),
    .ssb(net1617));
 b15fqy203ar1n02x5 gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net728),
    .clk(clknet_leaf_13_clk_i),
    .d1(net16),
    .d2(net2168),
    .o1(gen_filter_1__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_1__u_filter_filter_synced),
    .si1(net979),
    .si2(net980),
    .ssb(net1618));
 b15fqy043ar1n02x5 gen_filter_1__u_filter_stored_value_q_reg (.clk(clknet_leaf_13_clk_i),
    .d(gen_filter_1__u_filter_filter_synced),
    .den(eq_x_176_n25),
    .o(gen_filter_1__u_filter_stored_value_q),
    .rb(net728),
    .si(net981),
    .ssb(net1619));
 b15fqy203ar1n02x5 gen_filter_20__u_filter_diff_ctr_q_reg_0__gen_filter_20__u_filter_diff_ctr_q_reg_1_ (.rb(net737),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_20__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_20__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_20__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_20__u_filter_diff_ctr_q[1]),
    .si1(net982),
    .si2(net983),
    .ssb(net1620));
 b15fqy203ar1n02x5 gen_filter_20__u_filter_diff_ctr_q_reg_2__gen_filter_20__u_filter_diff_ctr_q_reg_3_ (.rb(net737),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_20__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_20__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_20__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_20__u_filter_diff_ctr_q[3]),
    .si1(net984),
    .si2(net985),
    .ssb(net1621));
 b15fqy203ar1n02x5 gen_filter_20__u_filter_filter_q_reg_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net751),
    .clk(clknet_leaf_4_clk_i),
    .d1(gen_filter_20__u_filter_filter_synced),
    .d2(net685),
    .o1(gen_filter_20__u_filter_filter_q),
    .o2(gen_filter_20__u_filter_filter_synced),
    .si1(net986),
    .si2(net987),
    .ssb(net1622));
 b15fqy043ar1n02x5 gen_filter_20__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(gen_filter_20__u_filter_filter_synced),
    .den(eq_x_81_n25),
    .o(gen_filter_20__u_filter_stored_value_q),
    .rb(net736),
    .si(net988),
    .ssb(net1623));
 b15fqy203ar1n02x5 gen_filter_21__u_filter_diff_ctr_q_reg_0__gen_filter_21__u_filter_diff_ctr_q_reg_1_ (.rb(net736),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_filter_21__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_21__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_21__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_21__u_filter_diff_ctr_q[1]),
    .si1(net989),
    .si2(net990),
    .ssb(net1624));
 b15fqy203ar1n02x5 gen_filter_21__u_filter_diff_ctr_q_reg_2__gen_filter_21__u_filter_diff_ctr_q_reg_3_ (.rb(net736),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_filter_21__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_21__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_21__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_21__u_filter_diff_ctr_q[3]),
    .si1(net991),
    .si2(net992),
    .ssb(net1625));
 b15fqy203ar1n02x5 gen_filter_21__u_filter_filter_q_reg_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net751),
    .clk(clknet_leaf_5_clk_i),
    .d1(gen_filter_21__u_filter_filter_synced),
    .d2(net18),
    .o1(gen_filter_21__u_filter_filter_q),
    .o2(gen_filter_21__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net993),
    .si2(net994),
    .ssb(net1626));
 b15fqy203ar1n02x5 gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_diff_ctr_q_reg_0_ (.rb(net751),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2239),
    .d2(net2340),
    .o1(gen_filter_21__u_filter_filter_synced),
    .o2(gen_filter_28__u_filter_diff_ctr_q[0]),
    .si1(net995),
    .si2(net996),
    .ssb(net1627));
 b15fqy043ar1n02x5 gen_filter_21__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(gen_filter_21__u_filter_filter_synced),
    .den(eq_x_76_n25),
    .o(gen_filter_21__u_filter_stored_value_q),
    .rb(net751),
    .si(net997),
    .ssb(net1628));
 b15fqy203ar1n02x5 gen_filter_22__u_filter_diff_ctr_q_reg_0__gen_filter_22__u_filter_diff_ctr_q_reg_1_ (.rb(net736),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_filter_22__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_22__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_22__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_22__u_filter_diff_ctr_q[1]),
    .si1(net998),
    .si2(net999),
    .ssb(net1629));
 b15fqy203ar1n02x5 gen_filter_22__u_filter_diff_ctr_q_reg_2__gen_filter_22__u_filter_diff_ctr_q_reg_3_ (.rb(net751),
    .clk(clknet_leaf_4_clk_i),
    .d1(gen_filter_22__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_22__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_22__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_22__u_filter_diff_ctr_q[3]),
    .si1(net1000),
    .si2(net1001),
    .ssb(net1630));
 b15fqy203ar1n02x5 gen_filter_22__u_filter_filter_q_reg_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net755),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2429),
    .d2(net19),
    .o1(gen_filter_22__u_filter_filter_q),
    .o2(gen_filter_22__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1002),
    .si2(net1003),
    .ssb(net1631));
 b15fqy203ar1n02x5 gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_diff_ctr_q_reg_0_ (.rb(net755),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2199),
    .d2(net2178),
    .o1(gen_filter_22__u_filter_filter_synced),
    .o2(gen_filter_23__u_filter_diff_ctr_q[0]),
    .si1(net1004),
    .si2(net1005),
    .ssb(net1632));
 b15fqy043ar1n02x5 gen_filter_22__u_filter_stored_value_q_reg (.clk(clknet_leaf_6_clk_i),
    .d(gen_filter_22__u_filter_filter_synced),
    .den(eq_x_71_n25),
    .o(gen_filter_22__u_filter_stored_value_q),
    .rb(net754),
    .si(net1006),
    .ssb(net1633));
 b15fqy203ar1n02x5 gen_filter_23__u_filter_diff_ctr_q_reg_1__gen_filter_23__u_filter_diff_ctr_q_reg_2_ (.rb(net755),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2163),
    .d2(gen_filter_23__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_23__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_23__u_filter_diff_ctr_q[2]),
    .si1(net1007),
    .si2(net1008),
    .ssb(net1634));
 b15fqy203ar1n02x5 gen_filter_23__u_filter_diff_ctr_q_reg_3__gen_filter_23__u_filter_filter_q_reg (.rb(net755),
    .clk(clknet_leaf_6_clk_i),
    .d1(gen_filter_23__u_filter_diff_ctr_d[3]),
    .d2(gen_filter_23__u_filter_filter_synced),
    .o1(gen_filter_23__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_23__u_filter_filter_q),
    .si1(net1009),
    .si2(net1010),
    .ssb(net1635));
 b15fqy203ar1n02x5 gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net753),
    .clk(clknet_leaf_6_clk_i),
    .d1(net20),
    .d2(net2164),
    .o1(gen_filter_23__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_23__u_filter_filter_synced),
    .si1(net1011),
    .si2(net1012),
    .ssb(net1636));
 b15fqy043ar1n02x5 gen_filter_23__u_filter_stored_value_q_reg (.clk(clknet_leaf_6_clk_i),
    .d(gen_filter_23__u_filter_filter_synced),
    .den(eq_x_66_n25),
    .o(gen_filter_23__u_filter_stored_value_q),
    .rb(net757),
    .si(net1013),
    .ssb(net1637));
 b15fqy203ar1n02x5 gen_filter_24__u_filter_diff_ctr_q_reg_0__gen_filter_24__u_filter_diff_ctr_q_reg_1_ (.rb(net735),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2242),
    .d2(gen_filter_24__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_24__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_24__u_filter_diff_ctr_q[1]),
    .si1(net1014),
    .si2(net1015),
    .ssb(net1638));
 b15fqy203ar1n02x5 gen_filter_24__u_filter_diff_ctr_q_reg_2__gen_filter_24__u_filter_diff_ctr_q_reg_3_ (.rb(net735),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2262),
    .d2(gen_filter_24__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_24__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_24__u_filter_diff_ctr_q[3]),
    .si1(net1016),
    .si2(net1017),
    .ssb(net1639));
 b15fqy203ar1n02x5 gen_filter_24__u_filter_filter_q_reg_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net735),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_24__u_filter_filter_synced),
    .d2(net21),
    .o1(gen_filter_24__u_filter_filter_q),
    .o2(gen_filter_24__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1018),
    .si2(net1019),
    .ssb(net1640));
 b15fqy203ar1n02x5 gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_25__u_filter_diff_ctr_q_reg_0_ (.rb(net735),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2189),
    .d2(gen_filter_25__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_24__u_filter_filter_synced),
    .o2(gen_filter_25__u_filter_diff_ctr_q[0]),
    .si1(net1020),
    .si2(net1021),
    .ssb(net1641));
 b15fqy043ar1n02x5 gen_filter_24__u_filter_stored_value_q_reg (.clk(clknet_leaf_2_clk_i),
    .d(gen_filter_24__u_filter_filter_synced),
    .den(eq_x_61_n25),
    .o(gen_filter_24__u_filter_stored_value_q),
    .rb(net735),
    .si(net1022),
    .ssb(net1642));
 b15fqy203ar1n02x5 gen_filter_25__u_filter_diff_ctr_q_reg_1__gen_filter_25__u_filter_diff_ctr_q_reg_2_ (.rb(net735),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2373),
    .d2(net2320),
    .o1(gen_filter_25__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_25__u_filter_diff_ctr_q[2]),
    .si1(net1023),
    .si2(net1024),
    .ssb(net1643));
 b15fqy203ar1n02x5 gen_filter_25__u_filter_diff_ctr_q_reg_3__gen_filter_25__u_filter_filter_q_reg (.rb(net735),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_25__u_filter_diff_ctr_d[3]),
    .d2(gen_filter_25__u_filter_filter_synced),
    .o1(gen_filter_25__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_25__u_filter_filter_q),
    .si1(net1025),
    .si2(net1026),
    .ssb(net1644));
 b15fqy203ar1n02x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_0_ (.rb(net737),
    .clk(clknet_leaf_3_clk_i),
    .d1(net22),
    .d2(intr_hw_N32),
    .o1(gen_filter_25__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(net205),
    .si1(net1027),
    .si2(net1028),
    .ssb(net1645));
 b15fqy203ar1n02x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_27__u_filter_diff_ctr_q_reg_0_ (.rb(net737),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2165),
    .d2(gen_filter_27__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_25__u_filter_filter_synced),
    .o2(gen_filter_27__u_filter_diff_ctr_q[0]),
    .si1(net1029),
    .si2(net1030),
    .ssb(net1646));
 b15fqy043ar1n02x5 gen_filter_25__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(gen_filter_25__u_filter_filter_synced),
    .den(eq_x_56_n25),
    .o(gen_filter_25__u_filter_stored_value_q),
    .rb(net737),
    .si(net1031),
    .ssb(net1647));
 b15fqy203ar1n02x5 gen_filter_26__u_filter_diff_ctr_q_reg_1__gen_filter_26__u_filter_diff_ctr_q_reg_2_ (.rb(net734),
    .clk(clknet_leaf_1_clk_i),
    .d1(gen_filter_26__u_filter_diff_ctr_d[1]),
    .d2(gen_filter_26__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_26__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_26__u_filter_diff_ctr_q[2]),
    .si1(net1032),
    .si2(net1033),
    .ssb(net1648));
 b15fqy203ar1n02x5 gen_filter_26__u_filter_diff_ctr_q_reg_3__gen_filter_26__u_filter_filter_q_reg (.rb(net734),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2426),
    .d2(net683),
    .o1(gen_filter_26__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_26__u_filter_filter_q),
    .si1(net1034),
    .si2(net1035),
    .ssb(net1649));
 b15fqy203ar1n02x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net729),
    .clk(clknet_leaf_12_clk_i),
    .d1(net23),
    .d2(net2172),
    .o1(gen_filter_26__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_26__u_filter_filter_synced),
    .si1(net1036),
    .si2(net1037),
    .ssb(net1650));
 b15fqy043ar1n02x5 gen_filter_26__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(net684),
    .den(eq_x_51_n25),
    .o(gen_filter_26__u_filter_stored_value_q),
    .rb(net739),
    .si(net1038),
    .ssb(net1651));
 b15fqy203ar1n02x5 gen_filter_27__u_filter_diff_ctr_q_reg_1__gen_filter_27__u_filter_diff_ctr_q_reg_2_ (.rb(net737),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_27__u_filter_diff_ctr_d[1]),
    .d2(gen_filter_27__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_27__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_27__u_filter_diff_ctr_q[2]),
    .si1(net1039),
    .si2(net1040),
    .ssb(net1652));
 b15fqy203ar1n02x5 gen_filter_27__u_filter_diff_ctr_q_reg_3__gen_filter_27__u_filter_filter_q_reg (.rb(net737),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2375),
    .d2(net2330),
    .o1(gen_filter_27__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_27__u_filter_filter_q),
    .si1(net1041),
    .si2(net1042),
    .ssb(net1653));
 b15fqy203ar1n02x5 gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net736),
    .clk(clknet_leaf_3_clk_i),
    .d1(net24),
    .d2(net2170),
    .o1(gen_filter_27__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_27__u_filter_filter_synced),
    .si1(net1043),
    .si2(net1044),
    .ssb(net1654));
 b15fqy043ar1n02x5 gen_filter_27__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(gen_filter_27__u_filter_filter_synced),
    .den(eq_x_46_n25),
    .o(gen_filter_27__u_filter_stored_value_q),
    .rb(net737),
    .si(net1045),
    .ssb(net1655));
 b15fqy203ar1n02x5 gen_filter_28__u_filter_diff_ctr_q_reg_1__gen_filter_28__u_filter_diff_ctr_q_reg_2_ (.rb(net754),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2462),
    .d2(net2421),
    .o1(gen_filter_28__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_28__u_filter_diff_ctr_q[2]),
    .si1(net1046),
    .si2(net1047),
    .ssb(net1656));
 b15fqy203ar1n02x5 gen_filter_28__u_filter_diff_ctr_q_reg_3__gen_filter_28__u_filter_filter_q_reg (.rb(net754),
    .clk(clknet_leaf_5_clk_i),
    .d1(gen_filter_28__u_filter_diff_ctr_d[3]),
    .d2(gen_filter_28__u_filter_filter_synced),
    .o1(gen_filter_28__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_28__u_filter_filter_q),
    .si1(net1048),
    .si2(net1049),
    .ssb(net1657));
 b15fqy203ar1n02x5 gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net754),
    .clk(clknet_leaf_5_clk_i),
    .d1(net25),
    .d2(net2176),
    .o1(gen_filter_28__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_28__u_filter_filter_synced),
    .si1(net1050),
    .si2(net1051),
    .ssb(net1658));
 b15fqy043ar1n02x5 gen_filter_28__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(gen_filter_28__u_filter_filter_synced),
    .den(eq_x_41_n25),
    .o(gen_filter_28__u_filter_stored_value_q),
    .rb(net754),
    .si(net1052),
    .ssb(net1659));
 b15fqy203ar1n02x5 gen_filter_29__u_filter_diff_ctr_q_reg_0__gen_filter_29__u_filter_diff_ctr_q_reg_1_ (.rb(net755),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2337),
    .d2(net2363),
    .o1(gen_filter_29__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_29__u_filter_diff_ctr_q[1]),
    .si1(net1053),
    .si2(net1054),
    .ssb(net1660));
 b15fqy203ar1n02x5 gen_filter_29__u_filter_diff_ctr_q_reg_2__gen_filter_29__u_filter_diff_ctr_q_reg_3_ (.rb(net755),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2344),
    .d2(gen_filter_29__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_29__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_29__u_filter_diff_ctr_q[3]),
    .si1(net1055),
    .si2(net1056),
    .ssb(net1661));
 b15fqy203ar1n02x5 gen_filter_29__u_filter_filter_q_reg_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net755),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2259),
    .d2(net26),
    .o1(gen_filter_29__u_filter_filter_q),
    .o2(gen_filter_29__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1057),
    .si2(net1058),
    .ssb(net1662));
 b15fqy003ar1n02x5 gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net755),
    .clk(clknet_leaf_5_clk_i),
    .d(net2157),
    .o(gen_filter_29__u_filter_filter_synced),
    .si(net1059),
    .ssb(net1663));
 b15fqy043ar1n02x5 gen_filter_29__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(net2259),
    .den(eq_x_36_n25),
    .o(gen_filter_29__u_filter_stored_value_q),
    .rb(net755),
    .si(net1060),
    .ssb(net1664));
 b15fqy203ar1n02x5 gen_filter_2__u_filter_diff_ctr_q_reg_0__gen_filter_2__u_filter_diff_ctr_q_reg_1_ (.rb(net727),
    .clk(clknet_leaf_14_clk_i),
    .d1(net2312),
    .d2(gen_filter_2__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_2__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_2__u_filter_diff_ctr_q[1]),
    .si1(net1061),
    .si2(net1062),
    .ssb(net1665));
 b15fqy203ar1n02x5 gen_filter_2__u_filter_diff_ctr_q_reg_2__gen_filter_2__u_filter_diff_ctr_q_reg_3_ (.rb(net725),
    .clk(clknet_leaf_14_clk_i),
    .d1(gen_filter_2__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_2__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_2__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_2__u_filter_diff_ctr_q[3]),
    .si1(net1063),
    .si2(net1064),
    .ssb(net1666));
 b15fqy203ar1n02x5 gen_filter_2__u_filter_filter_q_reg_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net725),
    .clk(clknet_leaf_14_clk_i),
    .d1(gen_filter_2__u_filter_filter_synced),
    .d2(net2447),
    .o1(gen_filter_2__u_filter_filter_q),
    .o2(gen_filter_2__u_filter_filter_synced),
    .si1(net1065),
    .si2(net1066),
    .ssb(net1667));
 b15fqy203ar1n02x5 gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net725),
    .clk(clknet_leaf_13_clk_i),
    .d1(net27),
    .d2(net2225),
    .o1(gen_filter_2__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_3__u_filter_filter_synced),
    .si1(net1067),
    .si2(net1068),
    .ssb(net1668));
 b15fqy043ar1n02x5 gen_filter_2__u_filter_stored_value_q_reg (.clk(clknet_leaf_14_clk_i),
    .d(gen_filter_2__u_filter_filter_synced),
    .den(eq_x_171_n25),
    .o(gen_filter_2__u_filter_stored_value_q),
    .rb(net725),
    .si(net1069),
    .ssb(net1669));
 b15fqy203ar1n02x5 gen_filter_30__u_filter_diff_ctr_q_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_1_ (.rb(net751),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2398),
    .d2(net2416),
    .o1(gen_filter_30__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_30__u_filter_diff_ctr_q[1]),
    .si1(net1070),
    .si2(net1071),
    .ssb(net1670));
 b15fqy203ar1n02x5 gen_filter_30__u_filter_diff_ctr_q_reg_2__gen_filter_30__u_filter_diff_ctr_q_reg_3_ (.rb(net751),
    .clk(clknet_leaf_5_clk_i),
    .d1(gen_filter_30__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_30__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_30__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_30__u_filter_diff_ctr_q[3]),
    .si1(net1072),
    .si2(net1073),
    .ssb(net1671));
 b15fqy203ar1n02x5 gen_filter_30__u_filter_filter_q_reg_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net754),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2476),
    .d2(net2389),
    .o1(gen_filter_30__u_filter_filter_q),
    .o2(gen_filter_30__u_filter_filter_synced),
    .si1(net1074),
    .si2(net1075),
    .ssb(net1672));
 b15fqy043ar1n02x5 gen_filter_30__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(gen_filter_30__u_filter_filter_synced),
    .den(eq_x_31_n25),
    .o(gen_filter_30__u_filter_stored_value_q),
    .rb(net751),
    .si(net1076),
    .ssb(net1673));
 b15fqy203ar1n02x5 gen_filter_31__u_filter_diff_ctr_q_reg_0__gen_filter_31__u_filter_diff_ctr_q_reg_1_ (.rb(net737),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_filter_31__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_31__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_31__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_31__u_filter_diff_ctr_q[1]),
    .si1(net1077),
    .si2(net1078),
    .ssb(net1674));
 b15fqy203ar1n02x5 gen_filter_31__u_filter_diff_ctr_q_reg_2__gen_filter_31__u_filter_diff_ctr_q_reg_3_ (.rb(net737),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2289),
    .d2(net2287),
    .o1(gen_filter_31__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_31__u_filter_diff_ctr_q[3]),
    .si1(net1079),
    .si2(net1080),
    .ssb(net1675));
 b15fqy203ar1n02x5 gen_filter_31__u_filter_filter_q_reg_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net736),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_filter_31__u_filter_filter_synced),
    .d2(net29),
    .o1(gen_filter_31__u_filter_filter_q),
    .o2(gen_filter_31__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1081),
    .si2(net1082),
    .ssb(net1676));
 b15fqy203ar1n02x5 gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_3_ (.rb(net751),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2435),
    .d2(intr_hw_N29),
    .o1(gen_filter_31__u_filter_filter_synced),
    .o2(net230),
    .si1(net1083),
    .si2(net1084),
    .ssb(net1677));
 b15fqy043ar1n02x5 gen_filter_31__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(gen_filter_31__u_filter_filter_synced),
    .den(eq_x_26_n25),
    .o(gen_filter_31__u_filter_stored_value_q),
    .rb(net737),
    .si(net1085),
    .ssb(net1678));
 b15fqy203ar1n02x5 gen_filter_3__u_filter_diff_ctr_q_reg_0__gen_filter_3__u_filter_diff_ctr_q_reg_1_ (.rb(net734),
    .clk(clknet_leaf_1_clk_i),
    .d1(gen_filter_3__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_3__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_3__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_3__u_filter_diff_ctr_q[1]),
    .si1(net1086),
    .si2(net1087),
    .ssb(net1679));
 b15fqy203ar1n02x5 gen_filter_3__u_filter_diff_ctr_q_reg_2__gen_filter_3__u_filter_diff_ctr_q_reg_3_ (.rb(net734),
    .clk(clknet_leaf_1_clk_i),
    .d1(gen_filter_3__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_3__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_3__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_3__u_filter_diff_ctr_q[3]),
    .si1(net1088),
    .si2(net1089),
    .ssb(net1680));
 b15fqy203ar1n02x5 gen_filter_3__u_filter_filter_q_reg_gen_filter_4__u_filter_diff_ctr_q_reg_0_ (.rb(net725),
    .clk(clknet_leaf_14_clk_i),
    .d1(net682),
    .d2(gen_filter_4__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_3__u_filter_filter_q),
    .o2(gen_filter_4__u_filter_diff_ctr_q[0]),
    .si1(net1090),
    .si2(net1091),
    .ssb(net1681));
 b15fqy203ar1n02x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net725),
    .clk(clknet_leaf_13_clk_i),
    .d1(net30),
    .d2(net31),
    .o1(gen_filter_3__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_4__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1092),
    .si2(net1093),
    .ssb(net1682));
 b15fqy043ar1n02x5 gen_filter_3__u_filter_stored_value_q_reg (.clk(clknet_leaf_14_clk_i),
    .d(net682),
    .den(eq_x_166_n25),
    .o(gen_filter_3__u_filter_stored_value_q),
    .rb(net726),
    .si(net1094),
    .ssb(net1683));
 b15fqy203ar1n02x5 gen_filter_4__u_filter_diff_ctr_q_reg_1__gen_filter_4__u_filter_diff_ctr_q_reg_2_ (.rb(net732),
    .clk(clknet_leaf_13_clk_i),
    .d1(net2272),
    .d2(net2394),
    .o1(gen_filter_4__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_4__u_filter_diff_ctr_q[2]),
    .si1(net1095),
    .si2(net1096),
    .ssb(net1684));
 b15fqy203ar1n02x5 gen_filter_4__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_diff_ctr_q_reg_0_ (.rb(net725),
    .clk(clknet_leaf_13_clk_i),
    .d1(gen_filter_4__u_filter_diff_ctr_d[3]),
    .d2(gen_filter_10__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_4__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_10__u_filter_diff_ctr_q[0]),
    .si1(net1097),
    .si2(net1098),
    .ssb(net1685));
 b15fqy203ar1n02x5 gen_filter_4__u_filter_filter_q_reg_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net732),
    .clk(clknet_leaf_13_clk_i),
    .d1(net2290),
    .d2(net2310),
    .o1(gen_filter_4__u_filter_filter_q),
    .o2(gen_filter_4__u_filter_filter_synced),
    .si1(net1099),
    .si2(net1100),
    .ssb(net1686));
 b15fqy043ar1n02x5 gen_filter_4__u_filter_stored_value_q_reg (.clk(clknet_leaf_13_clk_i),
    .d(net2290),
    .den(eq_x_161_n25),
    .o(gen_filter_4__u_filter_stored_value_q),
    .rb(net732),
    .si(net1101),
    .ssb(net1687));
 b15fqy203ar1n02x5 gen_filter_5__u_filter_diff_ctr_q_reg_0__gen_filter_5__u_filter_diff_ctr_q_reg_1_ (.rb(net735),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2353),
    .d2(gen_filter_5__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_5__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_5__u_filter_diff_ctr_q[1]),
    .si1(net1102),
    .si2(net1103),
    .ssb(net1688));
 b15fqy203ar1n02x5 gen_filter_5__u_filter_diff_ctr_q_reg_2__gen_filter_5__u_filter_filter_q_reg (.rb(net734),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2411),
    .d2(net680),
    .o1(gen_filter_5__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_5__u_filter_filter_q),
    .si1(net1104),
    .si2(net1105),
    .ssb(net1689));
 b15fqy203ar1n02x5 gen_filter_5__u_filter_diff_ctr_q_reg_3__gen_filter_6__u_filter_diff_ctr_q_reg_0_ (.rb(net737),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_5__u_filter_diff_ctr_d[3]),
    .d2(net2266),
    .o1(gen_filter_5__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_6__u_filter_diff_ctr_q[0]),
    .si1(net1106),
    .si2(net1107),
    .ssb(net1690));
 b15fqy203ar1n02x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_diff_ctr_q_reg_0_ (.rb(net728),
    .clk(clknet_leaf_12_clk_i),
    .d1(gen_filter_5__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .d2(gen_filter_9__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_5__u_filter_filter_synced),
    .o2(gen_filter_9__u_filter_diff_ctr_q[0]),
    .si1(net1108),
    .si2(net1109),
    .ssb(net1691));
 b15fqy043ar1n02x5 gen_filter_5__u_filter_stored_value_q_reg (.clk(clknet_leaf_1_clk_i),
    .d(net680),
    .den(eq_x_156_n25),
    .o(gen_filter_5__u_filter_stored_value_q),
    .rb(net739),
    .si(net1110),
    .ssb(net1692));
 b15fqy203ar1n02x5 gen_filter_6__u_filter_diff_ctr_q_reg_1__gen_filter_6__u_filter_diff_ctr_q_reg_2_ (.rb(net737),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_filter_6__u_filter_diff_ctr_d[1]),
    .d2(gen_filter_6__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_6__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_6__u_filter_diff_ctr_q[2]),
    .si1(net1111),
    .si2(net1112),
    .ssb(net1693));
 b15fqy203ar1n02x5 gen_filter_6__u_filter_diff_ctr_q_reg_3__gen_filter_6__u_filter_filter_q_reg (.rb(net734),
    .clk(clknet_leaf_1_clk_i),
    .d1(gen_filter_6__u_filter_diff_ctr_d[3]),
    .d2(net679),
    .o1(gen_filter_6__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_6__u_filter_filter_q),
    .si1(net1113),
    .si2(net1114),
    .ssb(net1694));
 b15fqy203ar1n02x5 gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net726),
    .clk(clknet_leaf_0_clk_i),
    .d1(net33),
    .d2(net2171),
    .o1(gen_filter_6__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_6__u_filter_filter_synced),
    .si1(net1115),
    .si2(net1116),
    .ssb(net1695));
 b15fqy043ar1n02x5 gen_filter_6__u_filter_stored_value_q_reg (.clk(clknet_leaf_1_clk_i),
    .d(net679),
    .den(eq_x_151_n25),
    .o(gen_filter_6__u_filter_stored_value_q),
    .rb(net734),
    .si(net1117),
    .ssb(net1696));
 b15fqy203ar1n02x5 gen_filter_7__u_filter_diff_ctr_q_reg_0__gen_filter_7__u_filter_diff_ctr_q_reg_1_ (.rb(net746),
    .clk(clknet_leaf_9_clk_i),
    .d1(gen_filter_7__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_7__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_7__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_7__u_filter_diff_ctr_q[1]),
    .si1(net1118),
    .si2(net1119),
    .ssb(net1697));
 b15fqy203ar1n02x5 gen_filter_7__u_filter_diff_ctr_q_reg_2__gen_filter_7__u_filter_diff_ctr_q_reg_3_ (.rb(net748),
    .clk(clknet_leaf_9_clk_i),
    .d1(gen_filter_7__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_7__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_7__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_7__u_filter_diff_ctr_q[3]),
    .si1(net1120),
    .si2(net1121),
    .ssb(net1698));
 b15fqy203ar1n02x5 gen_filter_7__u_filter_filter_q_reg_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net747),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2341),
    .d2(net34),
    .o1(gen_filter_7__u_filter_filter_q),
    .o2(gen_filter_7__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1122),
    .si2(net1123),
    .ssb(net1699));
 b15fqy203ar1n02x5 gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_diff_ctr_q_reg_3_ (.rb(net746),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2224),
    .d2(gen_filter_15__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_7__u_filter_filter_synced),
    .o2(gen_filter_15__u_filter_diff_ctr_q[3]),
    .si1(net1124),
    .si2(net1125),
    .ssb(net1700));
 b15fqy043ar1n02x5 gen_filter_7__u_filter_stored_value_q_reg (.clk(clknet_leaf_9_clk_i),
    .d(net2341),
    .den(eq_x_146_n25),
    .o(gen_filter_7__u_filter_stored_value_q),
    .rb(net744),
    .si(net1126),
    .ssb(net1701));
 b15fqy203ar1n02x5 gen_filter_8__u_filter_diff_ctr_q_reg_0__gen_filter_8__u_filter_diff_ctr_q_reg_1_ (.rb(net748),
    .clk(clknet_leaf_10_clk_i),
    .d1(gen_filter_8__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_8__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_8__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_8__u_filter_diff_ctr_q[1]),
    .si1(net1127),
    .si2(net1128),
    .ssb(net1702));
 b15fqy203ar1n02x5 gen_filter_8__u_filter_diff_ctr_q_reg_2__gen_filter_8__u_filter_diff_ctr_q_reg_3_ (.rb(net748),
    .clk(clknet_leaf_10_clk_i),
    .d1(net2300),
    .d2(gen_filter_8__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_8__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_8__u_filter_diff_ctr_q[3]),
    .si1(net1129),
    .si2(net1130),
    .ssb(net1703));
 b15fqy203ar1n02x5 gen_filter_8__u_filter_filter_q_reg_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net746),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2216),
    .d2(net35),
    .o1(gen_filter_8__u_filter_filter_q),
    .o2(gen_filter_8__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1131),
    .si2(net1132),
    .ssb(net1704));
 b15fqy203ar1n02x5 gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_diff_ctr_q_reg_0_ (.rb(net746),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2179),
    .d2(gen_filter_17__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_8__u_filter_filter_synced),
    .o2(gen_filter_17__u_filter_diff_ctr_q[0]),
    .si1(net1133),
    .si2(net1134),
    .ssb(net1705));
 b15fqy043ar1n02x5 gen_filter_8__u_filter_stored_value_q_reg (.clk(clknet_leaf_10_clk_i),
    .d(net2216),
    .den(eq_x_141_n25),
    .o(gen_filter_8__u_filter_stored_value_q),
    .rb(net746),
    .si(net1135),
    .ssb(net1706));
 b15fqy203ar1n02x5 gen_filter_9__u_filter_diff_ctr_q_reg_1__gen_filter_9__u_filter_diff_ctr_q_reg_2_ (.rb(net729),
    .clk(clknet_leaf_12_clk_i),
    .d1(gen_filter_9__u_filter_diff_ctr_d[1]),
    .d2(gen_filter_9__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_9__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_9__u_filter_diff_ctr_q[2]),
    .si1(net1136),
    .si2(net1137),
    .ssb(net1707));
 b15fqy203ar1n02x5 gen_filter_9__u_filter_diff_ctr_q_reg_3__gen_filter_9__u_filter_filter_q_reg (.rb(net729),
    .clk(clknet_leaf_12_clk_i),
    .d1(gen_filter_9__u_filter_diff_ctr_d[3]),
    .d2(gen_filter_9__u_filter_filter_synced),
    .o1(gen_filter_9__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_9__u_filter_filter_q),
    .si1(net1138),
    .si2(net1139),
    .ssb(net1708));
 b15fqy203ar1n02x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_1_ (.rb(net742),
    .clk(clknet_leaf_11_clk_i),
    .d1(net36),
    .d2(gen_filter_11__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_9__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_11__u_filter_diff_ctr_q[1]),
    .si1(net1140),
    .si2(net1141),
    .ssb(net1709));
 b15fqy203ar1n02x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net742),
    .clk(clknet_leaf_11_clk_i),
    .d1(net2213),
    .d2(net7),
    .o1(gen_filter_9__u_filter_filter_synced),
    .o2(gen_filter_11__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1142),
    .si2(net1143),
    .ssb(net1710));
 b15fqy043ar1n02x5 gen_filter_9__u_filter_stored_value_q_reg (.clk(clknet_leaf_11_clk_i),
    .d(gen_filter_9__u_filter_filter_synced),
    .den(net2280),
    .o(gen_filter_9__u_filter_stored_value_q),
    .rb(net742),
    .si(net1144),
    .ssb(net1711));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_10__intr_hw_intr_o_reg_11_ (.rb(net726),
    .clk(clknet_leaf_14_clk_i),
    .d1(intr_hw_N22),
    .d2(intr_hw_N21),
    .o1(net206),
    .o2(net207),
    .si1(net1145),
    .si2(net1146),
    .ssb(net1712));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_12__intr_hw_intr_o_reg_13_ (.rb(net747),
    .clk(clknet_leaf_9_clk_i),
    .d1(intr_hw_N20),
    .d2(intr_hw_N19),
    .o1(net208),
    .o2(net209),
    .si1(net1147),
    .si2(net1148),
    .ssb(net1713));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_14__intr_hw_intr_o_reg_15_ (.rb(net743),
    .clk(clknet_leaf_10_clk_i),
    .d1(intr_hw_N18),
    .d2(intr_hw_N17),
    .o1(net210),
    .o2(net211),
    .si1(net1149),
    .si2(net1150),
    .ssb(net1714));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_16__intr_hw_intr_o_reg_17_ (.rb(net757),
    .clk(clknet_leaf_7_clk_i),
    .d1(intr_hw_N16),
    .d2(intr_hw_N15),
    .o1(net212),
    .o2(net213),
    .si1(net1151),
    .si2(net1152),
    .ssb(net1715));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_19__intr_hw_intr_o_reg_20_ (.rb(net754),
    .clk(clknet_leaf_5_clk_i),
    .d1(intr_hw_N13),
    .d2(intr_hw_N12),
    .o1(net215),
    .o2(net217),
    .si1(net1153),
    .si2(net1154),
    .ssb(net1716));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_1__intr_hw_intr_o_reg_2_ (.rb(net729),
    .clk(clknet_leaf_12_clk_i),
    .d1(intr_hw_N31),
    .d2(intr_hw_N30),
    .o1(net216),
    .o2(net227),
    .si1(net1155),
    .si2(net1156),
    .ssb(net1717));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_21__intr_hw_intr_o_reg_30_ (.rb(net751),
    .clk(clknet_leaf_5_clk_i),
    .d1(intr_hw_N11),
    .d2(intr_hw_N2),
    .o1(net218),
    .o2(net228),
    .si1(net1157),
    .si2(net1158),
    .ssb(net1718));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_22__intr_hw_intr_o_reg_23_ (.rb(net757),
    .clk(clknet_leaf_6_clk_i),
    .d1(intr_hw_N10),
    .d2(intr_hw_N9),
    .o1(net219),
    .o2(net220),
    .si1(net1159),
    .si2(net1160),
    .ssb(net1719));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_24__intr_hw_intr_o_reg_25_ (.rb(net736),
    .clk(clknet_leaf_3_clk_i),
    .d1(intr_hw_N8),
    .d2(intr_hw_N7),
    .o1(net221),
    .o2(net222),
    .si1(net1161),
    .si2(net1162),
    .ssb(net1720));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_26__intr_hw_intr_o_reg_27_ (.rb(net737),
    .clk(clknet_leaf_3_clk_i),
    .d1(intr_hw_N6),
    .d2(intr_hw_N5),
    .o1(net223),
    .o2(net224),
    .si1(net1163),
    .si2(net1164),
    .ssb(net1721));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_28__intr_hw_intr_o_reg_29_ (.rb(net755),
    .clk(clknet_leaf_6_clk_i),
    .d1(intr_hw_N4),
    .d2(intr_hw_N3),
    .o1(net225),
    .o2(net226),
    .si1(net1165),
    .si2(net1166),
    .ssb(net1722));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_31__u_reg_u_data_in_q_reg_3_ (.rb(net742),
    .clk(clknet_leaf_11_clk_i),
    .d1(intr_hw_N1),
    .d2(u_reg_u_data_in_wr_data[3]),
    .o1(net229),
    .o2(u_reg_data_in_qs[3]),
    .si1(net1167),
    .si2(net1168),
    .ssb(net1723));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_4__intr_hw_intr_o_reg_5_ (.rb(net726),
    .clk(clknet_leaf_0_clk_i),
    .d1(intr_hw_N28),
    .d2(intr_hw_N27),
    .o1(net231),
    .o2(net232),
    .si1(net1169),
    .si2(net1170),
    .ssb(net1724));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_6__intr_hw_intr_o_reg_7_ (.rb(net739),
    .clk(clknet_leaf_1_clk_i),
    .d1(intr_hw_N26),
    .d2(intr_hw_N25),
    .o1(net233),
    .o2(net234),
    .si1(net1171),
    .si2(net1172),
    .ssb(net1725));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_8__intr_hw_intr_o_reg_18_ (.rb(net747),
    .clk(clknet_leaf_9_clk_i),
    .d1(intr_hw_N24),
    .d2(intr_hw_N14),
    .o1(net235),
    .o2(net214),
    .si1(net1173),
    .si2(net1174),
    .ssb(net1726));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_9__u_reg_u_data_in_q_reg_5_ (.rb(net726),
    .clk(clknet_leaf_14_clk_i),
    .d1(intr_hw_N23),
    .d2(u_reg_u_data_in_wr_data[5]),
    .o1(net236),
    .o2(u_reg_data_in_qs[5]),
    .si1(net1175),
    .si2(net1176),
    .ssb(net1727));
 b15fqy203ar1n02x5 u_reg_err_q_reg_u_reg_u_data_in_q_reg_6_ (.rb(net734),
    .clk(clknet_leaf_1_clk_i),
    .d1(n1439),
    .d2(u_reg_u_data_in_wr_data[6]),
    .o1(u_reg_err_q),
    .o2(u_reg_data_in_qs[6]),
    .si1(net1177),
    .si2(net1178),
    .ssb(net1728));
 b15cilb05ah1n02x3 u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_0_latch (.clk(clknet_leaf_3_clk_i),
    .clkout(u_reg_u_ctrl_en_input_filter_net2098),
    .en(u_reg_reg_we_check_15_),
    .te(net1179));
 b15cilb05ah1n02x3 u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_latch (.clk(clknet_leaf_13_clk_i),
    .clkout(u_reg_u_ctrl_en_input_filter_net2092),
    .en(u_reg_reg_we_check_15_),
    .te(net1180));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_0__u_reg_u_ctrl_en_input_filter_q_reg_1_ (.rb(net728),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2092),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[0]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[1]),
    .o1(reg2hw_ctrl_en_input_filter__q__0_),
    .o2(reg2hw_ctrl_en_input_filter__q__1_),
    .si1(net1181),
    .si2(net1182),
    .ssb(net1729));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_10__u_reg_u_ctrl_en_input_filter_q_reg_11_ (.rb(net728),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2092),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[10]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[11]),
    .o1(reg2hw_ctrl_en_input_filter__q__10_),
    .o2(reg2hw_ctrl_en_input_filter__q__11_),
    .si1(net1183),
    .si2(net1184),
    .ssb(net1730));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_12__u_reg_u_ctrl_en_input_filter_q_reg_13_ (.rb(net728),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2092),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[12]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[13]),
    .o1(reg2hw_ctrl_en_input_filter__q__12_),
    .o2(reg2hw_ctrl_en_input_filter__q__13_),
    .si1(net1185),
    .si2(net1186),
    .ssb(net1731));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_14__u_reg_u_ctrl_en_input_filter_q_reg_15_ (.rb(net728),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2092),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[14]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[15]),
    .o1(reg2hw_ctrl_en_input_filter__q__14_),
    .o2(reg2hw_ctrl_en_input_filter__q__15_),
    .si1(net1187),
    .si2(net1188),
    .ssb(net1732));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_16__u_reg_u_ctrl_en_input_filter_q_reg_17_ (.rb(net739),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2098),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[16]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[17]),
    .o1(reg2hw_ctrl_en_input_filter__q__16_),
    .o2(reg2hw_ctrl_en_input_filter__q__17_),
    .si1(net1189),
    .si2(net1190),
    .ssb(net1733));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_18__u_reg_u_ctrl_en_input_filter_q_reg_19_ (.rb(net738),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2098),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[18]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[19]),
    .o1(reg2hw_ctrl_en_input_filter__q__18_),
    .o2(reg2hw_ctrl_en_input_filter__q__19_),
    .si1(net1191),
    .si2(net1192),
    .ssb(net1734));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_20__u_reg_u_ctrl_en_input_filter_q_reg_21_ (.rb(net736),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2098),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[20]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[21]),
    .o1(reg2hw_ctrl_en_input_filter__q__20_),
    .o2(reg2hw_ctrl_en_input_filter__q__21_),
    .si1(net1193),
    .si2(net1194),
    .ssb(net1735));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_22__u_reg_u_ctrl_en_input_filter_q_reg_23_ (.rb(net739),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2098),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[22]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[23]),
    .o1(reg2hw_ctrl_en_input_filter__q__22_),
    .o2(reg2hw_ctrl_en_input_filter__q__23_),
    .si1(net1195),
    .si2(net1196),
    .ssb(net1736));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_24__u_reg_u_ctrl_en_input_filter_q_reg_25_ (.rb(net736),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2098),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[24]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[25]),
    .o1(reg2hw_ctrl_en_input_filter__q__24_),
    .o2(reg2hw_ctrl_en_input_filter__q__25_),
    .si1(net1197),
    .si2(net1198),
    .ssb(net1737));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_26__u_reg_u_ctrl_en_input_filter_q_reg_27_ (.rb(net739),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2098),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[26]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[27]),
    .o1(reg2hw_ctrl_en_input_filter__q__26_),
    .o2(reg2hw_ctrl_en_input_filter__q__27_),
    .si1(net1199),
    .si2(net1200),
    .ssb(net1738));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_28__u_reg_u_ctrl_en_input_filter_q_reg_29_ (.rb(net736),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2098),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[28]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[29]),
    .o1(reg2hw_ctrl_en_input_filter__q__28_),
    .o2(reg2hw_ctrl_en_input_filter__q__29_),
    .si1(net1201),
    .si2(net1202),
    .ssb(net1739));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_2__u_reg_u_ctrl_en_input_filter_q_reg_3_ (.rb(net728),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2092),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[2]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[3]),
    .o1(reg2hw_ctrl_en_input_filter__q__2_),
    .o2(reg2hw_ctrl_en_input_filter__q__3_),
    .si1(net1203),
    .si2(net1204),
    .ssb(net1740));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_30__u_reg_u_ctrl_en_input_filter_q_reg_31_ (.rb(net736),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2098),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[30]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[31]),
    .o1(reg2hw_ctrl_en_input_filter__q__30_),
    .o2(reg2hw_ctrl_en_input_filter__q__31_),
    .si1(net1205),
    .si2(net1206),
    .ssb(net1741));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_4__u_reg_u_ctrl_en_input_filter_q_reg_5_ (.rb(net728),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2092),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[4]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[5]),
    .o1(reg2hw_ctrl_en_input_filter__q__4_),
    .o2(reg2hw_ctrl_en_input_filter__q__5_),
    .si1(net1207),
    .si2(net1208),
    .ssb(net1742));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_6__u_reg_u_ctrl_en_input_filter_q_reg_7_ (.rb(net728),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2092),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[6]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[7]),
    .o1(reg2hw_ctrl_en_input_filter__q__6_),
    .o2(reg2hw_ctrl_en_input_filter__q__7_),
    .si1(net1209),
    .si2(net1210),
    .ssb(net1743));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_8__u_reg_u_ctrl_en_input_filter_q_reg_9_ (.rb(net728),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2092),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[8]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[9]),
    .o1(reg2hw_ctrl_en_input_filter__q__8_),
    .o2(reg2hw_ctrl_en_input_filter__q__9_),
    .si1(net1211),
    .si2(net1212),
    .ssb(net1744));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_0__u_reg_u_data_in_q_reg_1_ (.rb(net744),
    .clk(clknet_leaf_9_clk_i),
    .d1(net365),
    .d2(u_reg_u_data_in_wr_data[1]),
    .o1(u_reg_data_in_qs[0]),
    .o2(u_reg_data_in_qs[1]),
    .si1(net1213),
    .si2(net1214),
    .ssb(net1745));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_11__u_reg_u_data_in_q_reg_16_ (.rb(net744),
    .clk(clknet_leaf_8_clk_i),
    .d1(u_reg_u_data_in_wr_data[11]),
    .d2(u_reg_u_data_in_wr_data[16]),
    .o1(u_reg_data_in_qs[11]),
    .o2(u_reg_data_in_qs[16]),
    .si1(net1215),
    .si2(net1216),
    .ssb(net1746));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_12__u_reg_u_data_in_q_reg_17_ (.rb(net747),
    .clk(clknet_leaf_9_clk_i),
    .d1(u_reg_u_data_in_wr_data[12]),
    .d2(u_reg_u_data_in_wr_data[17]),
    .o1(u_reg_data_in_qs[12]),
    .o2(u_reg_data_in_qs[17]),
    .si1(net1217),
    .si2(net1218),
    .ssb(net1747));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_13__u_reg_u_data_in_q_reg_14_ (.rb(net747),
    .clk(clknet_leaf_9_clk_i),
    .d1(u_reg_u_data_in_wr_data[13]),
    .d2(u_reg_u_data_in_wr_data[14]),
    .o1(u_reg_data_in_qs[13]),
    .o2(u_reg_data_in_qs[14]),
    .si1(net1219),
    .si2(net1220),
    .ssb(net1748));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_18__u_reg_u_data_in_q_reg_19_ (.rb(net753),
    .clk(clknet_leaf_7_clk_i),
    .d1(u_reg_u_data_in_wr_data[18]),
    .d2(u_reg_u_data_in_wr_data[19]),
    .o1(u_reg_data_in_qs[18]),
    .o2(u_reg_data_in_qs[19]),
    .si1(net1221),
    .si2(net1222),
    .ssb(net1749));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_20__u_reg_u_data_in_q_reg_21_ (.rb(net751),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_reg_u_data_in_wr_data[20]),
    .d2(u_reg_u_data_in_wr_data[21]),
    .o1(u_reg_data_in_qs[20]),
    .o2(u_reg_data_in_qs[21]),
    .si1(net1223),
    .si2(net1224),
    .ssb(net1750));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_22__u_reg_u_data_in_q_reg_23_ (.rb(net757),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_reg_u_data_in_wr_data[22]),
    .d2(u_reg_u_data_in_wr_data[23]),
    .o1(u_reg_data_in_qs[22]),
    .o2(u_reg_data_in_qs[23]),
    .si1(net1225),
    .si2(net1226),
    .ssb(net1751));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_24__u_reg_u_data_in_q_reg_25_ (.rb(net751),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_reg_u_data_in_wr_data[24]),
    .d2(u_reg_u_data_in_wr_data[25]),
    .o1(u_reg_data_in_qs[24]),
    .o2(u_reg_data_in_qs[25]),
    .si1(net1227),
    .si2(net1228),
    .ssb(net1752));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_26__u_reg_u_reg_if_rspop_q_reg_1_ (.rb(net737),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_reg_u_data_in_wr_data[26]),
    .d2(n1429),
    .o1(u_reg_data_in_qs[26]),
    .o2(net292),
    .si1(net1229),
    .si2(net1230),
    .ssb(net1753));
 b15fqy003ar1n02x5 u_reg_u_data_in_q_reg_27_ (.rb(net739),
    .clk(clknet_leaf_3_clk_i),
    .d(u_reg_u_data_in_wr_data[27]),
    .o(u_reg_data_in_qs[27]),
    .si(net1231),
    .ssb(net1754));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_28__u_reg_u_data_in_q_reg_29_ (.rb(net754),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_reg_u_data_in_wr_data[28]),
    .d2(u_reg_u_data_in_wr_data[29]),
    .o1(u_reg_data_in_qs[28]),
    .o2(u_reg_data_in_qs[29]),
    .si1(net1232),
    .si2(net1233),
    .ssb(net1755));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_2__u_reg_u_data_in_q_reg_8_ (.rb(net742),
    .clk(clknet_leaf_11_clk_i),
    .d1(u_reg_u_data_in_wr_data[2]),
    .d2(u_reg_u_data_in_wr_data[8]),
    .o1(u_reg_data_in_qs[2]),
    .o2(u_reg_data_in_qs[8]),
    .si1(net1234),
    .si2(net1235),
    .ssb(net1756));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_30__u_reg_u_reg_if_rspop_q_reg_2_ (.rb(net737),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_reg_u_data_in_wr_data[30]),
    .d2(n1432),
    .o1(u_reg_data_in_qs[30]),
    .o2(net293),
    .si1(net1236),
    .si2(net1237),
    .ssb(net1757));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_4__u_reg_u_data_in_q_reg_10_ (.rb(net726),
    .clk(clknet_leaf_14_clk_i),
    .d1(u_reg_u_data_in_wr_data[4]),
    .d2(u_reg_u_data_in_wr_data[10]),
    .o1(u_reg_data_in_qs[4]),
    .o2(u_reg_data_in_qs[10]),
    .si1(net1238),
    .si2(net1239),
    .ssb(net1758));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_7__u_reg_u_data_in_q_reg_31_ (.rb(net749),
    .clk(clknet_leaf_8_clk_i),
    .d1(net364),
    .d2(u_reg_u_data_in_wr_data[31]),
    .o1(u_reg_data_in_qs[7]),
    .o2(u_reg_data_in_qs[31]),
    .si1(net1240),
    .si2(net1241),
    .ssb(net1759));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_9__u_reg_u_data_in_q_reg_15_ (.rb(net744),
    .clk(clknet_leaf_11_clk_i),
    .d1(u_reg_u_data_in_wr_data[9]),
    .d2(u_reg_u_data_in_wr_data[15]),
    .o1(u_reg_data_in_qs[9]),
    .o2(u_reg_data_in_qs[15]),
    .si1(net1242),
    .si2(net1243),
    .ssb(net1760));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_0_latch (.clk(clknet_leaf_4_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_falling_net2098),
    .en(n4185),
    .te(net1244));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_latch (.clk(clknet_leaf_0_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_falling_net2092),
    .en(n4185),
    .te(net1245));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_0__u_reg_u_intr_ctrl_en_falling_q_reg_1_ (.rb(net726),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2092),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[0]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[1]),
    .o1(reg2hw_intr_ctrl_en_falling__q__0_),
    .o2(reg2hw_intr_ctrl_en_falling__q__1_),
    .si1(net1246),
    .si2(net1247),
    .ssb(net1761));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_10__u_reg_u_intr_ctrl_en_falling_q_reg_11_ (.rb(net726),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2092),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[10]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[11]),
    .o1(reg2hw_intr_ctrl_en_falling__q__10_),
    .o2(reg2hw_intr_ctrl_en_falling__q__11_),
    .si1(net1248),
    .si2(net1249),
    .ssb(net1762));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_12__u_reg_u_intr_ctrl_en_falling_q_reg_13_ (.rb(net730),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2092),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[12]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[13]),
    .o1(reg2hw_intr_ctrl_en_falling__q__12_),
    .o2(reg2hw_intr_ctrl_en_falling__q__13_),
    .si1(net1250),
    .si2(net1251),
    .ssb(net1763));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_14__u_reg_u_intr_ctrl_en_falling_q_reg_15_ (.rb(net730),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2092),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[14]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[15]),
    .o1(reg2hw_intr_ctrl_en_falling__q__14_),
    .o2(reg2hw_intr_ctrl_en_falling__q__15_),
    .si1(net1252),
    .si2(net1253),
    .ssb(net1764));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_16__u_reg_u_intr_ctrl_en_falling_q_reg_17_ (.rb(net749),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2098),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[16]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[17]),
    .o1(reg2hw_intr_ctrl_en_falling__q__16_),
    .o2(reg2hw_intr_ctrl_en_falling__q__17_),
    .si1(net1254),
    .si2(net1255),
    .ssb(net1765));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_18__u_reg_u_intr_ctrl_en_falling_q_reg_19_ (.rb(net751),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2098),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[18]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[19]),
    .o1(reg2hw_intr_ctrl_en_falling__q__18_),
    .o2(reg2hw_intr_ctrl_en_falling__q__19_),
    .si1(net1256),
    .si2(net1257),
    .ssb(net1766));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_20__u_reg_u_intr_ctrl_en_falling_q_reg_21_ (.rb(net752),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2098),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[20]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[21]),
    .o1(reg2hw_intr_ctrl_en_falling__q__20_),
    .o2(reg2hw_intr_ctrl_en_falling__q__21_),
    .si1(net1258),
    .si2(net1259),
    .ssb(net1767));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_22__u_reg_u_intr_ctrl_en_falling_q_reg_23_ (.rb(net749),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2098),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[22]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[23]),
    .o1(reg2hw_intr_ctrl_en_falling__q__22_),
    .o2(reg2hw_intr_ctrl_en_falling__q__23_),
    .si1(net1260),
    .si2(net1261),
    .ssb(net1768));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_24__u_reg_u_intr_ctrl_en_falling_q_reg_25_ (.rb(net752),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2098),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[24]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[25]),
    .o1(reg2hw_intr_ctrl_en_falling__q__24_),
    .o2(reg2hw_intr_ctrl_en_falling__q__25_),
    .si1(net1262),
    .si2(net1263),
    .ssb(net1769));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_26__u_reg_u_intr_ctrl_en_falling_q_reg_27_ (.rb(net749),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2098),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[26]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[27]),
    .o1(reg2hw_intr_ctrl_en_falling__q__26_),
    .o2(reg2hw_intr_ctrl_en_falling__q__27_),
    .si1(net1264),
    .si2(net1265),
    .ssb(net1770));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_28__u_reg_u_intr_ctrl_en_falling_q_reg_29_ (.rb(net752),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2098),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[28]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[29]),
    .o1(reg2hw_intr_ctrl_en_falling__q__28_),
    .o2(reg2hw_intr_ctrl_en_falling__q__29_),
    .si1(net1266),
    .si2(net1267),
    .ssb(net1771));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_2__u_reg_u_intr_ctrl_en_falling_q_reg_3_ (.rb(net730),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2092),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[2]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[3]),
    .o1(reg2hw_intr_ctrl_en_falling__q__2_),
    .o2(reg2hw_intr_ctrl_en_falling__q__3_),
    .si1(net1268),
    .si2(net1269),
    .ssb(net1772));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_30__u_reg_u_intr_ctrl_en_falling_q_reg_31_ (.rb(net750),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2098),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[30]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[31]),
    .o1(reg2hw_intr_ctrl_en_falling__q__30_),
    .o2(reg2hw_intr_ctrl_en_falling__q__31_),
    .si1(net1270),
    .si2(net1271),
    .ssb(net1773));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_4__u_reg_u_intr_ctrl_en_falling_q_reg_5_ (.rb(net726),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2092),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[4]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[5]),
    .o1(reg2hw_intr_ctrl_en_falling__q__4_),
    .o2(reg2hw_intr_ctrl_en_falling__q__5_),
    .si1(net1272),
    .si2(net1273),
    .ssb(net1774));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_6__u_reg_u_intr_ctrl_en_falling_q_reg_7_ (.rb(net727),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2092),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[6]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[7]),
    .o1(reg2hw_intr_ctrl_en_falling__q__6_),
    .o2(reg2hw_intr_ctrl_en_falling__q__7_),
    .si1(net1274),
    .si2(net1275),
    .ssb(net1775));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_8__u_reg_u_intr_ctrl_en_falling_q_reg_9_ (.rb(net730),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2092),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[8]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[9]),
    .o1(reg2hw_intr_ctrl_en_falling__q__8_),
    .o2(reg2hw_intr_ctrl_en_falling__q__9_),
    .si1(net1276),
    .si2(net1277),
    .ssb(net1776));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_0_latch (.clk(clknet_leaf_7_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .en(n4183),
    .te(net1278));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_latch (.clk(clknet_leaf_11_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .en(n4183),
    .te(net1279));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1_ (.rb(net744),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[0]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[1]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__0_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__1_),
    .si1(net1280),
    .si2(net1281),
    .ssb(net1777));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11_ (.rb(net744),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[10]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[11]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__10_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__11_),
    .si1(net1282),
    .si2(net1283),
    .ssb(net1778));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13_ (.rb(net744),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[12]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[13]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__12_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__13_),
    .si1(net1284),
    .si2(net1285),
    .ssb(net1779));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15_ (.rb(net744),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[14]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[15]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__14_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__15_),
    .si1(net1286),
    .si2(net1287),
    .ssb(net1780));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17_ (.rb(net750),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[16]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[17]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__16_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__17_),
    .si1(net1288),
    .si2(net1289),
    .ssb(net1781));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19_ (.rb(net753),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[18]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[19]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__18_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__19_),
    .si1(net1290),
    .si2(net1291),
    .ssb(net1782));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21_ (.rb(net750),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[20]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[21]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__20_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__21_),
    .si1(net1292),
    .si2(net1293),
    .ssb(net1783));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23_ (.rb(net753),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[22]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[23]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__22_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__23_),
    .si1(net1294),
    .si2(net1295),
    .ssb(net1784));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25_ (.rb(net750),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[24]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[25]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__24_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__25_),
    .si1(net1296),
    .si2(net1297),
    .ssb(net1785));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27_ (.rb(net750),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[26]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[27]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__26_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__27_),
    .si1(net1298),
    .si2(net1299),
    .ssb(net1786));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29_ (.rb(net753),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[28]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[29]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__28_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__29_),
    .si1(net1300),
    .si2(net1301),
    .ssb(net1787));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3_ (.rb(net744),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[2]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[3]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__2_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__3_),
    .si1(net1302),
    .si2(net1303),
    .ssb(net1788));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31_ (.rb(net753),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[30]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[31]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__30_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__31_),
    .si1(net1304),
    .si2(net1305),
    .ssb(net1789));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5_ (.rb(net744),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[4]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[5]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__4_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__5_),
    .si1(net1306),
    .si2(net1307),
    .ssb(net1790));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7_ (.rb(net744),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[6]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[7]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__6_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__7_),
    .si1(net1308),
    .si2(net1309),
    .ssb(net1791));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9_ (.rb(net745),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[8]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[9]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__8_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__9_),
    .si1(net1310),
    .si2(net1311),
    .ssb(net1792));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_0_latch (.clk(clknet_leaf_4_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_lvllow_net2098),
    .en(n4190),
    .te(net1312));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_latch (.clk(clknet_leaf_12_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_lvllow_net2092),
    .en(n4190),
    .te(net1313));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_reg_u_intr_ctrl_en_lvllow_q_reg_1_ (.rb(net730),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[0]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[1]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__0_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__1_),
    .si1(net1314),
    .si2(net1315),
    .ssb(net1793));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_reg_u_intr_ctrl_en_lvllow_q_reg_11_ (.rb(net730),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[10]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[11]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__10_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__11_),
    .si1(net1316),
    .si2(net1317),
    .ssb(net1794));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_reg_u_intr_ctrl_en_lvllow_q_reg_13_ (.rb(net730),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[12]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[13]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__12_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__13_),
    .si1(net1318),
    .si2(net1319),
    .ssb(net1795));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_reg_u_intr_ctrl_en_lvllow_q_reg_15_ (.rb(net730),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[14]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[15]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__14_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__15_),
    .si1(net1320),
    .si2(net1321),
    .ssb(net1796));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_reg_u_intr_ctrl_en_lvllow_q_reg_17_ (.rb(net749),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[16]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[17]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__16_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__17_),
    .si1(net1322),
    .si2(net1323),
    .ssb(net1797));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_reg_u_intr_ctrl_en_lvllow_q_reg_19_ (.rb(net749),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[18]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[19]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__18_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__19_),
    .si1(net1324),
    .si2(net1325),
    .ssb(net1798));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_reg_u_intr_ctrl_en_lvllow_q_reg_21_ (.rb(net749),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[20]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[21]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__20_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__21_),
    .si1(net1326),
    .si2(net1327),
    .ssb(net1799));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_reg_u_intr_ctrl_en_lvllow_q_reg_23_ (.rb(net749),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[22]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[23]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__22_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__23_),
    .si1(net1328),
    .si2(net1329),
    .ssb(net1800));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_reg_u_intr_ctrl_en_lvllow_q_reg_25_ (.rb(net749),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[24]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[25]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__24_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__25_),
    .si1(net1330),
    .si2(net1331),
    .ssb(net1801));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_reg_u_intr_ctrl_en_lvllow_q_reg_27_ (.rb(net749),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[26]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[27]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__26_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__27_),
    .si1(net1332),
    .si2(net1333),
    .ssb(net1802));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_reg_u_intr_ctrl_en_lvllow_q_reg_29_ (.rb(net749),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[28]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[29]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__28_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__29_),
    .si1(net1334),
    .si2(net1335),
    .ssb(net1803));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_reg_u_intr_ctrl_en_lvllow_q_reg_3_ (.rb(net730),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[2]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[3]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__2_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__3_),
    .si1(net1336),
    .si2(net1337),
    .ssb(net1804));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_reg_u_intr_ctrl_en_lvllow_q_reg_31_ (.rb(net749),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[30]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[31]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__30_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__31_),
    .si1(net1338),
    .si2(net1339),
    .ssb(net1805));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_reg_u_intr_ctrl_en_lvllow_q_reg_5_ (.rb(net730),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[4]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[5]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__4_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__5_),
    .si1(net1340),
    .si2(net1341),
    .ssb(net1806));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_reg_u_intr_ctrl_en_lvllow_q_reg_7_ (.rb(net730),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[6]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[7]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__6_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__7_),
    .si1(net1342),
    .si2(net1343),
    .ssb(net1807));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_reg_u_intr_ctrl_en_lvllow_q_reg_9_ (.rb(net730),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[8]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[9]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__8_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__9_),
    .si1(net1344),
    .si2(net1345),
    .ssb(net1808));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_0_latch (.clk(clknet_leaf_5_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_rising_net2098),
    .en(n4184),
    .te(net1346));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_latch (.clk(clknet_leaf_12_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_rising_net2092),
    .en(n4184),
    .te(net1347));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_0__u_reg_u_intr_ctrl_en_rising_q_reg_1_ (.rb(net730),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2092),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[0]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[1]),
    .o1(reg2hw_intr_ctrl_en_rising__q__0_),
    .o2(reg2hw_intr_ctrl_en_rising__q__1_),
    .si1(net1348),
    .si2(net1349),
    .ssb(net1809));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_10__u_reg_u_intr_ctrl_en_rising_q_reg_11_ (.rb(net730),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2092),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[10]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[11]),
    .o1(reg2hw_intr_ctrl_en_rising__q__10_),
    .o2(reg2hw_intr_ctrl_en_rising__q__11_),
    .si1(net1350),
    .si2(net1351),
    .ssb(net1810));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_12__u_reg_u_intr_ctrl_en_rising_q_reg_13_ (.rb(net730),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2092),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[12]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[13]),
    .o1(reg2hw_intr_ctrl_en_rising__q__12_),
    .o2(reg2hw_intr_ctrl_en_rising__q__13_),
    .si1(net1352),
    .si2(net1353),
    .ssb(net1811));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_14__u_reg_u_intr_ctrl_en_rising_q_reg_15_ (.rb(net730),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2092),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[14]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[15]),
    .o1(reg2hw_intr_ctrl_en_rising__q__14_),
    .o2(reg2hw_intr_ctrl_en_rising__q__15_),
    .si1(net1354),
    .si2(net1355),
    .ssb(net1812));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_16__u_reg_u_intr_ctrl_en_rising_q_reg_17_ (.rb(net754),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2098),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[16]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[17]),
    .o1(reg2hw_intr_ctrl_en_rising__q__16_),
    .o2(reg2hw_intr_ctrl_en_rising__q__17_),
    .si1(net1356),
    .si2(net1357),
    .ssb(net1813));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_18__u_reg_u_intr_ctrl_en_rising_q_reg_19_ (.rb(net754),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2098),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[18]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[19]),
    .o1(reg2hw_intr_ctrl_en_rising__q__18_),
    .o2(reg2hw_intr_ctrl_en_rising__q__19_),
    .si1(net1358),
    .si2(net1359),
    .ssb(net1814));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_20__u_reg_u_intr_ctrl_en_rising_q_reg_21_ (.rb(net754),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2098),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[20]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[21]),
    .o1(reg2hw_intr_ctrl_en_rising__q__20_),
    .o2(reg2hw_intr_ctrl_en_rising__q__21_),
    .si1(net1360),
    .si2(net1361),
    .ssb(net1815));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_22__u_reg_u_intr_ctrl_en_rising_q_reg_23_ (.rb(net754),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2098),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[22]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[23]),
    .o1(reg2hw_intr_ctrl_en_rising__q__22_),
    .o2(reg2hw_intr_ctrl_en_rising__q__23_),
    .si1(net1362),
    .si2(net1363),
    .ssb(net1816));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_24__u_reg_u_intr_ctrl_en_rising_q_reg_25_ (.rb(net754),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2098),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[24]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[25]),
    .o1(reg2hw_intr_ctrl_en_rising__q__24_),
    .o2(reg2hw_intr_ctrl_en_rising__q__25_),
    .si1(net1364),
    .si2(net1365),
    .ssb(net1817));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_26__u_reg_u_intr_ctrl_en_rising_q_reg_27_ (.rb(net754),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2098),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[26]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[27]),
    .o1(reg2hw_intr_ctrl_en_rising__q__26_),
    .o2(reg2hw_intr_ctrl_en_rising__q__27_),
    .si1(net1366),
    .si2(net1367),
    .ssb(net1818));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_28__u_reg_u_intr_ctrl_en_rising_q_reg_29_ (.rb(net754),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2098),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[28]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[29]),
    .o1(reg2hw_intr_ctrl_en_rising__q__28_),
    .o2(reg2hw_intr_ctrl_en_rising__q__29_),
    .si1(net1368),
    .si2(net1369),
    .ssb(net1819));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_2__u_reg_u_intr_ctrl_en_rising_q_reg_3_ (.rb(net733),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2092),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[2]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[3]),
    .o1(reg2hw_intr_ctrl_en_rising__q__2_),
    .o2(reg2hw_intr_ctrl_en_rising__q__3_),
    .si1(net1370),
    .si2(net1371),
    .ssb(net1820));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_30__u_reg_u_intr_ctrl_en_rising_q_reg_31_ (.rb(net754),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2098),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[30]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[31]),
    .o1(reg2hw_intr_ctrl_en_rising__q__30_),
    .o2(reg2hw_intr_ctrl_en_rising__q__31_),
    .si1(net1372),
    .si2(net1373),
    .ssb(net1821));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_4__u_reg_u_intr_ctrl_en_rising_q_reg_5_ (.rb(net733),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2092),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[4]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[5]),
    .o1(reg2hw_intr_ctrl_en_rising__q__4_),
    .o2(reg2hw_intr_ctrl_en_rising__q__5_),
    .si1(net1374),
    .si2(net1375),
    .ssb(net1822));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_6__u_reg_u_intr_ctrl_en_rising_q_reg_7_ (.rb(net733),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2092),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[6]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[7]),
    .o1(reg2hw_intr_ctrl_en_rising__q__6_),
    .o2(reg2hw_intr_ctrl_en_rising__q__7_),
    .si1(net1376),
    .si2(net1377),
    .ssb(net1823));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_8__u_reg_u_intr_ctrl_en_rising_q_reg_9_ (.rb(net733),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2092),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[8]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[9]),
    .o1(reg2hw_intr_ctrl_en_rising__q__8_),
    .o2(reg2hw_intr_ctrl_en_rising__q__9_),
    .si1(net1378),
    .si2(net1379),
    .ssb(net1824));
 b15cilb05ah1n02x3 u_reg_u_intr_enable_clk_gate_q_reg_0_latch (.clk(clknet_leaf_7_clk_i),
    .clkout(u_reg_u_intr_enable_net2098),
    .en(n4182),
    .te(net1380));
 b15cilb05ah1n02x3 u_reg_u_intr_enable_clk_gate_q_reg_latch (.clk(clknet_leaf_12_clk_i),
    .clkout(u_reg_u_intr_enable_net2092),
    .en(n4182),
    .te(net1381));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_0__u_reg_u_intr_enable_q_reg_1_ (.rb(net729),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2092),
    .d1(u_reg_u_intr_enable_wr_data[0]),
    .d2(u_reg_u_intr_enable_wr_data[1]),
    .o1(reg2hw_intr_enable__q__0_),
    .o2(reg2hw_intr_enable__q__1_),
    .si1(net1382),
    .si2(net1383),
    .ssb(net1825));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_10__u_reg_u_intr_enable_q_reg_11_ (.rb(net729),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2092),
    .d1(u_reg_u_intr_enable_wr_data[10]),
    .d2(u_reg_u_intr_enable_wr_data[11]),
    .o1(reg2hw_intr_enable__q__10_),
    .o2(reg2hw_intr_enable__q__11_),
    .si1(net1384),
    .si2(net1385),
    .ssb(net1826));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_12__u_reg_u_intr_enable_q_reg_13_ (.rb(net729),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2092),
    .d1(u_reg_u_intr_enable_wr_data[12]),
    .d2(u_reg_u_intr_enable_wr_data[13]),
    .o1(reg2hw_intr_enable__q__12_),
    .o2(reg2hw_intr_enable__q__13_),
    .si1(net1386),
    .si2(net1387),
    .ssb(net1827));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_14__u_reg_u_intr_enable_q_reg_15_ (.rb(net729),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2092),
    .d1(u_reg_u_intr_enable_wr_data[14]),
    .d2(u_reg_u_intr_enable_wr_data[15]),
    .o1(reg2hw_intr_enable__q__14_),
    .o2(reg2hw_intr_enable__q__15_),
    .si1(net1388),
    .si2(net1389),
    .ssb(net1828));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_16__u_reg_u_intr_enable_q_reg_17_ (.rb(net757),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2098),
    .d1(u_reg_u_intr_enable_wr_data[16]),
    .d2(u_reg_u_intr_enable_wr_data[17]),
    .o1(reg2hw_intr_enable__q__16_),
    .o2(reg2hw_intr_enable__q__17_),
    .si1(net1390),
    .si2(net1391),
    .ssb(net1829));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_18__u_reg_u_intr_enable_q_reg_19_ (.rb(net753),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2098),
    .d1(u_reg_u_intr_enable_wr_data[18]),
    .d2(u_reg_u_intr_enable_wr_data[19]),
    .o1(reg2hw_intr_enable__q__18_),
    .o2(reg2hw_intr_enable__q__19_),
    .si1(net1392),
    .si2(net1393),
    .ssb(net1830));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_20__u_reg_u_intr_enable_q_reg_21_ (.rb(net753),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2098),
    .d1(u_reg_u_intr_enable_wr_data[20]),
    .d2(u_reg_u_intr_enable_wr_data[21]),
    .o1(reg2hw_intr_enable__q__20_),
    .o2(reg2hw_intr_enable__q__21_),
    .si1(net1394),
    .si2(net1395),
    .ssb(net1831));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_22__u_reg_u_intr_enable_q_reg_23_ (.rb(net757),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2098),
    .d1(u_reg_u_intr_enable_wr_data[22]),
    .d2(u_reg_u_intr_enable_wr_data[23]),
    .o1(reg2hw_intr_enable__q__22_),
    .o2(reg2hw_intr_enable__q__23_),
    .si1(net1396),
    .si2(net1397),
    .ssb(net1832));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_24__u_reg_u_intr_enable_q_reg_25_ (.rb(net753),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2098),
    .d1(u_reg_u_intr_enable_wr_data[24]),
    .d2(u_reg_u_intr_enable_wr_data[25]),
    .o1(reg2hw_intr_enable__q__24_),
    .o2(reg2hw_intr_enable__q__25_),
    .si1(net1398),
    .si2(net1399),
    .ssb(net1833));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_26__u_reg_u_intr_enable_q_reg_27_ (.rb(net753),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2098),
    .d1(u_reg_u_intr_enable_wr_data[26]),
    .d2(u_reg_u_intr_enable_wr_data[27]),
    .o1(reg2hw_intr_enable__q__26_),
    .o2(reg2hw_intr_enable__q__27_),
    .si1(net1400),
    .si2(net1401),
    .ssb(net1834));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_28__u_reg_u_intr_enable_q_reg_29_ (.rb(net757),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2098),
    .d1(u_reg_u_intr_enable_wr_data[28]),
    .d2(u_reg_u_intr_enable_wr_data[29]),
    .o1(reg2hw_intr_enable__q__28_),
    .o2(reg2hw_intr_enable__q__29_),
    .si1(net1402),
    .si2(net1403),
    .ssb(net1835));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_2__u_reg_u_intr_enable_q_reg_3_ (.rb(net729),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2092),
    .d1(u_reg_u_intr_enable_wr_data[2]),
    .d2(u_reg_u_intr_enable_wr_data[3]),
    .o1(reg2hw_intr_enable__q__2_),
    .o2(reg2hw_intr_enable__q__3_),
    .si1(net1404),
    .si2(net1405),
    .ssb(net1836));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_30__u_reg_u_intr_enable_q_reg_31_ (.rb(net753),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2098),
    .d1(u_reg_u_intr_enable_wr_data[30]),
    .d2(u_reg_u_intr_enable_wr_data[31]),
    .o1(reg2hw_intr_enable__q__30_),
    .o2(reg2hw_intr_enable__q__31_),
    .si1(net1406),
    .si2(net1407),
    .ssb(net1837));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_4__u_reg_u_intr_enable_q_reg_5_ (.rb(net729),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2092),
    .d1(u_reg_u_intr_enable_wr_data[4]),
    .d2(u_reg_u_intr_enable_wr_data[5]),
    .o1(reg2hw_intr_enable__q__4_),
    .o2(reg2hw_intr_enable__q__5_),
    .si1(net1408),
    .si2(net1409),
    .ssb(net1838));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_6__u_reg_u_intr_enable_q_reg_7_ (.rb(net729),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2092),
    .d1(u_reg_u_intr_enable_wr_data[6]),
    .d2(u_reg_u_intr_enable_wr_data[7]),
    .o1(reg2hw_intr_enable__q__6_),
    .o2(reg2hw_intr_enable__q__7_),
    .si1(net1410),
    .si2(net1411),
    .ssb(net1839));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_8__u_reg_u_intr_enable_q_reg_9_ (.rb(net729),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2092),
    .d1(u_reg_u_intr_enable_wr_data[8]),
    .d2(u_reg_u_intr_enable_wr_data[9]),
    .o1(reg2hw_intr_enable__q__8_),
    .o2(reg2hw_intr_enable__q__9_),
    .si1(net1412),
    .si2(net1413),
    .ssb(net1840));
 b15cilb05ah1n02x3 u_reg_u_intr_state_clk_gate_q_reg_0_latch (.clk(clknet_leaf_7_clk_i),
    .clkout(u_reg_u_intr_state_net2121),
    .en(u_reg_u_intr_state_n1),
    .te(net1414));
 b15cilb05ah1n02x3 u_reg_u_intr_state_clk_gate_q_reg_latch (.clk(clknet_leaf_8_clk_i),
    .clkout(u_reg_u_intr_state_net2115),
    .en(u_reg_u_intr_state_n1),
    .te(net1415));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_0__u_reg_u_intr_state_q_reg_1_ (.rb(net745),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2115),
    .d1(u_reg_u_intr_state_wr_data[0]),
    .d2(u_reg_u_intr_state_wr_data[1]),
    .o1(reg2hw_intr_state__q__0_),
    .o2(reg2hw_intr_state__q__1_),
    .si1(net1416),
    .si2(net1417),
    .ssb(net1841));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_10__u_reg_u_intr_state_q_reg_11_ (.rb(net744),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2115),
    .d1(u_reg_u_intr_state_wr_data[10]),
    .d2(u_reg_u_intr_state_wr_data[11]),
    .o1(reg2hw_intr_state__q__10_),
    .o2(reg2hw_intr_state__q__11_),
    .si1(net1418),
    .si2(net1419),
    .ssb(net1842));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_12__u_reg_u_intr_state_q_reg_13_ (.rb(net745),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2115),
    .d1(u_reg_u_intr_state_wr_data[12]),
    .d2(u_reg_u_intr_state_wr_data[13]),
    .o1(reg2hw_intr_state__q__12_),
    .o2(reg2hw_intr_state__q__13_),
    .si1(net1420),
    .si2(net1421),
    .ssb(net1843));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_14__u_reg_u_intr_state_q_reg_15_ (.rb(net745),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2115),
    .d1(u_reg_u_intr_state_wr_data[14]),
    .d2(u_reg_u_intr_state_wr_data[15]),
    .o1(reg2hw_intr_state__q__14_),
    .o2(reg2hw_intr_state__q__15_),
    .si1(net1422),
    .si2(net1423),
    .ssb(net1844));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_16__u_reg_u_intr_state_q_reg_17_ (.rb(net750),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2121),
    .d1(u_reg_u_intr_state_wr_data[16]),
    .d2(u_reg_u_intr_state_wr_data[17]),
    .o1(reg2hw_intr_state__q__16_),
    .o2(reg2hw_intr_state__q__17_),
    .si1(net1424),
    .si2(net1425),
    .ssb(net1845));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_18__u_reg_u_intr_state_q_reg_19_ (.rb(net750),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2121),
    .d1(u_reg_u_intr_state_wr_data[18]),
    .d2(u_reg_u_intr_state_wr_data[19]),
    .o1(reg2hw_intr_state__q__18_),
    .o2(reg2hw_intr_state__q__19_),
    .si1(net1426),
    .si2(net1427),
    .ssb(net1846));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_20__u_reg_u_intr_state_q_reg_21_ (.rb(net750),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2121),
    .d1(u_reg_u_intr_state_wr_data[20]),
    .d2(u_reg_u_intr_state_wr_data[21]),
    .o1(reg2hw_intr_state__q__20_),
    .o2(reg2hw_intr_state__q__21_),
    .si1(net1428),
    .si2(net1429),
    .ssb(net1847));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_22__u_reg_u_intr_state_q_reg_23_ (.rb(net750),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2121),
    .d1(u_reg_u_intr_state_wr_data[22]),
    .d2(u_reg_u_intr_state_wr_data[23]),
    .o1(reg2hw_intr_state__q__22_),
    .o2(reg2hw_intr_state__q__23_),
    .si1(net1430),
    .si2(net1431),
    .ssb(net1848));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_24__u_reg_u_intr_state_q_reg_25_ (.rb(net749),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2121),
    .d1(u_reg_u_intr_state_wr_data[24]),
    .d2(u_reg_u_intr_state_wr_data[25]),
    .o1(reg2hw_intr_state__q__24_),
    .o2(reg2hw_intr_state__q__25_),
    .si1(net1432),
    .si2(net1433),
    .ssb(net1849));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_26__u_reg_u_intr_state_q_reg_27_ (.rb(net749),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2121),
    .d1(u_reg_u_intr_state_wr_data[26]),
    .d2(u_reg_u_intr_state_wr_data[27]),
    .o1(reg2hw_intr_state__q__26_),
    .o2(reg2hw_intr_state__q__27_),
    .si1(net1434),
    .si2(net1435),
    .ssb(net1850));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_28__u_reg_u_intr_state_q_reg_29_ (.rb(net750),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2121),
    .d1(u_reg_u_intr_state_wr_data[28]),
    .d2(u_reg_u_intr_state_wr_data[29]),
    .o1(reg2hw_intr_state__q__28_),
    .o2(reg2hw_intr_state__q__29_),
    .si1(net1436),
    .si2(net1437),
    .ssb(net1851));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_2__u_reg_u_intr_state_q_reg_3_ (.rb(net744),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2115),
    .d1(u_reg_u_intr_state_wr_data[2]),
    .d2(u_reg_u_intr_state_wr_data[3]),
    .o1(reg2hw_intr_state__q__2_),
    .o2(reg2hw_intr_state__q__3_),
    .si1(net1438),
    .si2(net1439),
    .ssb(net1852));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_30__u_reg_u_intr_state_q_reg_31_ (.rb(net749),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2121),
    .d1(u_reg_u_intr_state_wr_data[30]),
    .d2(u_reg_u_intr_state_wr_data[31]),
    .o1(reg2hw_intr_state__q__30_),
    .o2(reg2hw_intr_state__q__31_),
    .si1(net1440),
    .si2(net1441),
    .ssb(net1853));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_4__u_reg_u_intr_state_q_reg_5_ (.rb(net745),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2115),
    .d1(u_reg_u_intr_state_wr_data[4]),
    .d2(u_reg_u_intr_state_wr_data[5]),
    .o1(reg2hw_intr_state__q__4_),
    .o2(reg2hw_intr_state__q__5_),
    .si1(net1442),
    .si2(net1443),
    .ssb(net1854));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_6__u_reg_u_intr_state_q_reg_7_ (.rb(net744),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2115),
    .d1(u_reg_u_intr_state_wr_data[6]),
    .d2(u_reg_u_intr_state_wr_data[7]),
    .o1(reg2hw_intr_state__q__6_),
    .o2(reg2hw_intr_state__q__7_),
    .si1(net1444),
    .si2(net1445),
    .ssb(net1855));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_8__u_reg_u_intr_state_q_reg_9_ (.rb(net744),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2115),
    .d1(u_reg_u_intr_state_wr_data[8]),
    .d2(u_reg_u_intr_state_wr_data[9]),
    .o1(reg2hw_intr_state__q__8_),
    .o2(reg2hw_intr_state__q__9_),
    .si1(net1446),
    .si2(net1447),
    .ssb(net1856));
 b15cilb05ah1n02x3 u_reg_u_reg_if_clk_gate_rdata_q_reg_0_latch (.clk(clknet_leaf_5_clk_i),
    .clkout(u_reg_u_reg_if_net2149),
    .en(net671),
    .te(net1448));
 b15cilb05ah1n02x3 u_reg_u_reg_if_clk_gate_rdata_q_reg_latch (.clk(clknet_leaf_2_clk_i),
    .clkout(u_reg_u_reg_if_net2144),
    .en(net672),
    .te(net1449));
 b15cilb05ah1n02x3 u_reg_u_reg_if_clk_gate_reqid_q_reg_latch (.clk(clknet_leaf_2_clk_i),
    .clkout(u_reg_u_reg_if_net2138),
    .en(net672),
    .te(net1450));
 b15fqy043ar1n02x5 u_reg_u_reg_if_error_q_reg (.clk(clknet_leaf_2_clk_i),
    .d(u_reg_u_reg_if_N46),
    .den(net671),
    .o(net248),
    .rb(net735),
    .si(net1451),
    .ssb(net1857));
 b15fqy043ar1n02x5 u_reg_u_reg_if_outstanding_q_reg (.clk(clknet_leaf_2_clk_i),
    .d(u_reg_u_reg_if_a_ack),
    .den(u_reg_u_reg_if_N7),
    .o(net294),
    .rb(net735),
    .si(net1452),
    .ssb(net1858));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_0__u_reg_u_reg_if_rdata_q_reg_1_ (.rb(net736),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2144),
    .d1(u_reg_u_reg_if_N14),
    .d2(net314),
    .o1(net244),
    .o2(net245),
    .si1(net1453),
    .si2(net1454),
    .ssb(net1859));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_10__u_reg_u_reg_if_rdata_q_reg_11_ (.rb(net741),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2144),
    .d1(net2317),
    .d2(net317),
    .o1(net255),
    .o2(net256),
    .si1(net1455),
    .si2(net1456),
    .ssb(net1860));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_12__u_reg_u_reg_if_rdata_q_reg_13_ (.rb(net736),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2144),
    .d1(net2102),
    .d2(net2351),
    .o1(net257),
    .o2(net258),
    .si1(net1457),
    .si2(net1458),
    .ssb(net1861));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_14__u_reg_u_reg_if_rdata_q_reg_15_ (.rb(net736),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2144),
    .d1(net315),
    .d2(u_reg_u_reg_if_N29),
    .o1(net260),
    .o2(net261),
    .si1(net1459),
    .si2(net1460),
    .ssb(net1862));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_16__u_reg_u_reg_if_rdata_q_reg_17_ (.rb(net752),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2149),
    .d1(net302),
    .d2(u_reg_u_reg_if_N31),
    .o1(net262),
    .o2(net263),
    .si1(net1461),
    .si2(net1462),
    .ssb(net1863));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_18__u_reg_u_reg_if_rdata_q_reg_19_ (.rb(net753),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2149),
    .d1(net2017),
    .d2(net2007),
    .o1(net264),
    .o2(net265),
    .si1(net1463),
    .si2(net1464),
    .ssb(net1864));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_20__u_reg_u_reg_if_rdata_q_reg_21_ (.rb(net751),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2149),
    .d1(net2058),
    .d2(net2089),
    .o1(net266),
    .o2(net267),
    .si1(net1465),
    .si2(net1466),
    .ssb(net1865));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_22__u_reg_u_reg_if_rdata_q_reg_23_ (.rb(net755),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2149),
    .d1(net2207),
    .d2(net2197),
    .o1(net268),
    .o2(net269),
    .si1(net1467),
    .si2(net1468),
    .ssb(net1866));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_24__u_reg_u_reg_if_rdata_q_reg_25_ (.rb(net751),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2149),
    .d1(net2222),
    .d2(net2047),
    .o1(net271),
    .o2(net272),
    .si1(net1469),
    .si2(net1470),
    .ssb(net1867));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_26__u_reg_u_reg_if_rdata_q_reg_27_ (.rb(net751),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2149),
    .d1(net2401),
    .d2(net2228),
    .o1(net273),
    .o2(net274),
    .si1(net1471),
    .si2(net1472),
    .ssb(net1868));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_28__u_reg_u_reg_if_rdata_q_reg_29_ (.rb(net752),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2149),
    .d1(net2064),
    .d2(net2135),
    .o1(net275),
    .o2(net276),
    .si1(net1473),
    .si2(net1474),
    .ssb(net1869));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_2__u_reg_u_reg_if_rdata_q_reg_3_ (.rb(net736),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2144),
    .d1(u_reg_u_reg_if_N16),
    .d2(net316),
    .o1(net246),
    .o2(net247),
    .si1(net1475),
    .si2(net1476),
    .ssb(net1870));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_30__u_reg_u_reg_if_rdata_q_reg_31_ (.rb(net752),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2149),
    .d1(net2270),
    .d2(net2253),
    .o1(net277),
    .o2(net278),
    .si1(net1477),
    .si2(net1478),
    .ssb(net1871));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_4__u_reg_u_reg_if_rdata_q_reg_5_ (.rb(net741),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2144),
    .d1(net2237),
    .d2(net2194),
    .o1(net249),
    .o2(net250),
    .si1(net1479),
    .si2(net1480),
    .ssb(net1872));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_6__u_reg_u_reg_if_rdata_q_reg_7_ (.rb(net738),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2144),
    .d1(net2105),
    .d2(net2076),
    .o1(net251),
    .o2(net252),
    .si1(net1481),
    .si2(net1482),
    .ssb(net1873));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_q_reg_8__u_reg_u_reg_if_rdata_q_reg_9_ (.rb(net740),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2144),
    .d1(u_reg_u_reg_if_N22),
    .d2(u_reg_u_reg_if_N23),
    .o1(net253),
    .o2(net254),
    .si1(net1483),
    .si2(net1484),
    .ssb(net1874));
 b15fqy203ar1n02x5 u_reg_u_reg_if_reqid_q_reg_0__u_reg_u_reg_if_reqid_q_reg_1_ (.rb(net735),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2138),
    .d1(net130),
    .d2(net131),
    .o1(net279),
    .o2(net281),
    .si1(net1485),
    .si2(net1486),
    .ssb(net1875));
 b15fqy203ar1n02x5 u_reg_u_reg_if_reqid_q_reg_2__u_reg_u_reg_if_reqid_q_reg_3_ (.rb(net735),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2138),
    .d1(net132),
    .d2(net133),
    .o1(net282),
    .o2(net283),
    .si1(net1487),
    .si2(net1488),
    .ssb(net1876));
 b15fqy203ar1n02x5 u_reg_u_reg_if_reqid_q_reg_4__u_reg_u_reg_if_reqid_q_reg_5_ (.rb(net735),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2138),
    .d1(net134),
    .d2(net135),
    .o1(net284),
    .o2(net285),
    .si1(net1489),
    .si2(net1490),
    .ssb(net1877));
 b15fqy203ar1n02x5 u_reg_u_reg_if_reqid_q_reg_6__u_reg_u_reg_if_reqid_q_reg_7_ (.rb(net735),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2138),
    .d1(net136),
    .d2(net137),
    .o1(net286),
    .o2(net287),
    .si1(net1491),
    .si2(net1492),
    .ssb(net1878));
 b15fqy043ar1n02x5 u_reg_u_reg_if_reqsz_q_reg_0_ (.clk(clknet_leaf_2_clk_i),
    .d(net39),
    .den(net672),
    .o(net288),
    .rb(net735),
    .si(net1493),
    .ssb(net1879));
 b15fqy043ar1n02x5 u_reg_u_reg_if_reqsz_q_reg_1_ (.clk(clknet_leaf_2_clk_i),
    .d(net40),
    .den(net672),
    .o(net289),
    .rb(net740),
    .si(net1494),
    .ssb(net1880));
 b15fqy043ar1n02x5 u_reg_u_reg_if_rspop_q_reg_0_ (.clk(clknet_leaf_2_clk_i),
    .d(u_reg_u_reg_if_rd_req),
    .den(u_reg_u_reg_if_a_ack),
    .o(net291),
    .rb(net735),
    .si(net1495),
    .ssb(net1881));
 b15tihi00an1n03x5 U3339_1496 (.o(net1496));
 b15cbf000an1n16x5 clkbuf_leaf_0_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_0_clk_i));
 b15ztpn00an1n08x5 PHY_92 ();
 b15ztpn00an1n08x5 PHY_93 ();
 b15ztpn00an1n08x5 PHY_94 ();
 b15ztpn00an1n08x5 PHY_95 ();
 b15ztpn00an1n08x5 PHY_96 ();
 b15ztpn00an1n08x5 PHY_97 ();
 b15ztpn00an1n08x5 PHY_98 ();
 b15ztpn00an1n08x5 PHY_99 ();
 b15ztpn00an1n08x5 PHY_100 ();
 b15ztpn00an1n08x5 PHY_101 ();
 b15ztpn00an1n08x5 PHY_102 ();
 b15ztpn00an1n08x5 PHY_103 ();
 b15ztpn00an1n08x5 PHY_104 ();
 b15ztpn00an1n08x5 PHY_105 ();
 b15ztpn00an1n08x5 PHY_106 ();
 b15ztpn00an1n08x5 PHY_107 ();
 b15ztpn00an1n08x5 PHY_108 ();
 b15ztpn00an1n08x5 PHY_109 ();
 b15ztpn00an1n08x5 PHY_110 ();
 b15ztpn00an1n08x5 PHY_111 ();
 b15ztpn00an1n08x5 PHY_112 ();
 b15ztpn00an1n08x5 PHY_113 ();
 b15ztpn00an1n08x5 PHY_114 ();
 b15ztpn00an1n08x5 PHY_115 ();
 b15ztpn00an1n08x5 PHY_116 ();
 b15ztpn00an1n08x5 PHY_117 ();
 b15ztpn00an1n08x5 PHY_118 ();
 b15ztpn00an1n08x5 PHY_119 ();
 b15ztpn00an1n08x5 PHY_120 ();
 b15ztpn00an1n08x5 PHY_121 ();
 b15ztpn00an1n08x5 PHY_122 ();
 b15ztpn00an1n08x5 PHY_123 ();
 b15ztpn00an1n08x5 PHY_124 ();
 b15ztpn00an1n08x5 PHY_125 ();
 b15ztpn00an1n08x5 PHY_126 ();
 b15ztpn00an1n08x5 PHY_127 ();
 b15ztpn00an1n08x5 PHY_128 ();
 b15ztpn00an1n08x5 PHY_129 ();
 b15ztpn00an1n08x5 PHY_130 ();
 b15ztpn00an1n08x5 PHY_131 ();
 b15ztpn00an1n08x5 PHY_132 ();
 b15ztpn00an1n08x5 PHY_133 ();
 b15ztpn00an1n08x5 PHY_134 ();
 b15ztpn00an1n08x5 PHY_135 ();
 b15ztpn00an1n08x5 PHY_136 ();
 b15ztpn00an1n08x5 PHY_137 ();
 b15ztpn00an1n08x5 PHY_138 ();
 b15ztpn00an1n08x5 PHY_139 ();
 b15ztpn00an1n08x5 PHY_140 ();
 b15ztpn00an1n08x5 PHY_141 ();
 b15ztpn00an1n08x5 PHY_142 ();
 b15ztpn00an1n08x5 PHY_143 ();
 b15ztpn00an1n08x5 PHY_144 ();
 b15ztpn00an1n08x5 PHY_145 ();
 b15ztpn00an1n08x5 PHY_146 ();
 b15ztpn00an1n08x5 PHY_147 ();
 b15ztpn00an1n08x5 PHY_148 ();
 b15ztpn00an1n08x5 PHY_149 ();
 b15ztpn00an1n08x5 PHY_150 ();
 b15ztpn00an1n08x5 PHY_151 ();
 b15ztpn00an1n08x5 PHY_152 ();
 b15ztpn00an1n08x5 PHY_153 ();
 b15ztpn00an1n08x5 PHY_154 ();
 b15ztpn00an1n08x5 PHY_155 ();
 b15ztpn00an1n08x5 PHY_156 ();
 b15ztpn00an1n08x5 PHY_157 ();
 b15ztpn00an1n08x5 PHY_158 ();
 b15ztpn00an1n08x5 PHY_159 ();
 b15ztpn00an1n08x5 PHY_160 ();
 b15ztpn00an1n08x5 PHY_161 ();
 b15ztpn00an1n08x5 PHY_162 ();
 b15ztpn00an1n08x5 PHY_163 ();
 b15ztpn00an1n08x5 PHY_164 ();
 b15ztpn00an1n08x5 PHY_165 ();
 b15ztpn00an1n08x5 PHY_166 ();
 b15ztpn00an1n08x5 PHY_167 ();
 b15ztpn00an1n08x5 PHY_168 ();
 b15ztpn00an1n08x5 PHY_169 ();
 b15ztpn00an1n08x5 PHY_170 ();
 b15ztpn00an1n08x5 PHY_171 ();
 b15ztpn00an1n08x5 PHY_172 ();
 b15ztpn00an1n08x5 PHY_173 ();
 b15ztpn00an1n08x5 PHY_174 ();
 b15ztpn00an1n08x5 PHY_175 ();
 b15ztpn00an1n08x5 PHY_176 ();
 b15ztpn00an1n08x5 PHY_177 ();
 b15ztpn00an1n08x5 PHY_178 ();
 b15ztpn00an1n08x5 PHY_179 ();
 b15ztpn00an1n08x5 PHY_180 ();
 b15ztpn00an1n08x5 PHY_181 ();
 b15ztpn00an1n08x5 PHY_182 ();
 b15ztpn00an1n08x5 PHY_183 ();
 b15ztpn00an1n08x5 PHY_184 ();
 b15ztpn00an1n08x5 PHY_185 ();
 b15ztpn00an1n08x5 PHY_186 ();
 b15ztpn00an1n08x5 PHY_187 ();
 b15ztpn00an1n08x5 PHY_188 ();
 b15ztpn00an1n08x5 PHY_189 ();
 b15ztpn00an1n08x5 PHY_190 ();
 b15ztpn00an1n08x5 PHY_191 ();
 b15ztpn00an1n08x5 PHY_192 ();
 b15ztpn00an1n08x5 PHY_193 ();
 b15ztpn00an1n08x5 PHY_194 ();
 b15ztpn00an1n08x5 PHY_195 ();
 b15ztpn00an1n08x5 PHY_196 ();
 b15ztpn00an1n08x5 PHY_197 ();
 b15ztpn00an1n08x5 PHY_198 ();
 b15ztpn00an1n08x5 PHY_199 ();
 b15ztpn00an1n08x5 PHY_200 ();
 b15ztpn00an1n08x5 PHY_201 ();
 b15ztpn00an1n08x5 PHY_202 ();
 b15ztpn00an1n08x5 PHY_203 ();
 b15ztpn00an1n08x5 PHY_204 ();
 b15ztpn00an1n08x5 PHY_205 ();
 b15ztpn00an1n08x5 PHY_206 ();
 b15ztpn00an1n08x5 PHY_207 ();
 b15ztpn00an1n08x5 PHY_208 ();
 b15ztpn00an1n08x5 PHY_209 ();
 b15ztpn00an1n08x5 PHY_210 ();
 b15ztpn00an1n08x5 PHY_211 ();
 b15ztpn00an1n08x5 PHY_212 ();
 b15ztpn00an1n08x5 PHY_213 ();
 b15ztpn00an1n08x5 PHY_214 ();
 b15ztpn00an1n08x5 PHY_215 ();
 b15ztpn00an1n08x5 PHY_216 ();
 b15ztpn00an1n08x5 PHY_217 ();
 b15ztpn00an1n08x5 PHY_218 ();
 b15ztpn00an1n08x5 PHY_219 ();
 b15ztpn00an1n08x5 PHY_220 ();
 b15ztpn00an1n08x5 PHY_221 ();
 b15ztpn00an1n08x5 PHY_222 ();
 b15ztpn00an1n08x5 PHY_223 ();
 b15ztpn00an1n08x5 PHY_224 ();
 b15ztpn00an1n08x5 PHY_225 ();
 b15ztpn00an1n08x5 PHY_226 ();
 b15ztpn00an1n08x5 PHY_227 ();
 b15ztpn00an1n08x5 PHY_228 ();
 b15ztpn00an1n08x5 PHY_229 ();
 b15ztpn00an1n08x5 PHY_230 ();
 b15ztpn00an1n08x5 PHY_231 ();
 b15ztpn00an1n08x5 PHY_232 ();
 b15ztpn00an1n08x5 PHY_233 ();
 b15ztpn00an1n08x5 PHY_234 ();
 b15ztpn00an1n08x5 PHY_235 ();
 b15ztpn00an1n08x5 PHY_236 ();
 b15ztpn00an1n08x5 PHY_237 ();
 b15ztpn00an1n08x5 PHY_238 ();
 b15ztpn00an1n08x5 PHY_239 ();
 b15ztpn00an1n08x5 PHY_240 ();
 b15ztpn00an1n08x5 PHY_241 ();
 b15ztpn00an1n08x5 PHY_242 ();
 b15ztpn00an1n08x5 PHY_243 ();
 b15ztpn00an1n08x5 PHY_244 ();
 b15ztpn00an1n08x5 PHY_245 ();
 b15ztpn00an1n08x5 PHY_246 ();
 b15ztpn00an1n08x5 PHY_247 ();
 b15ztpn00an1n08x5 PHY_248 ();
 b15ztpn00an1n08x5 PHY_249 ();
 b15ztpn00an1n08x5 PHY_250 ();
 b15ztpn00an1n08x5 PHY_251 ();
 b15ztpn00an1n08x5 PHY_252 ();
 b15ztpn00an1n08x5 PHY_253 ();
 b15ztpn00an1n08x5 PHY_254 ();
 b15ztpn00an1n08x5 PHY_255 ();
 b15ztpn00an1n08x5 PHY_256 ();
 b15ztpn00an1n08x5 PHY_257 ();
 b15ztpn00an1n08x5 PHY_258 ();
 b15ztpn00an1n08x5 PHY_259 ();
 b15ztpn00an1n08x5 PHY_260 ();
 b15ztpn00an1n08x5 PHY_261 ();
 b15ztpn00an1n08x5 PHY_262 ();
 b15ztpn00an1n08x5 PHY_263 ();
 b15ztpn00an1n08x5 PHY_264 ();
 b15ztpn00an1n08x5 PHY_265 ();
 b15ztpn00an1n08x5 PHY_266 ();
 b15ztpn00an1n08x5 PHY_267 ();
 b15ztpn00an1n08x5 PHY_268 ();
 b15ztpn00an1n08x5 PHY_269 ();
 b15ztpn00an1n08x5 PHY_270 ();
 b15ztpn00an1n08x5 PHY_271 ();
 b15ztpn00an1n08x5 PHY_272 ();
 b15ztpn00an1n08x5 PHY_273 ();
 b15ztpn00an1n08x5 PHY_274 ();
 b15ztpn00an1n08x5 PHY_275 ();
 b15ztpn00an1n08x5 PHY_276 ();
 b15ztpn00an1n08x5 PHY_277 ();
 b15ztpn00an1n08x5 PHY_278 ();
 b15ztpn00an1n08x5 PHY_279 ();
 b15ztpn00an1n08x5 PHY_280 ();
 b15ztpn00an1n08x5 PHY_281 ();
 b15ztpn00an1n08x5 PHY_282 ();
 b15ztpn00an1n08x5 PHY_283 ();
 b15ztpn00an1n08x5 PHY_284 ();
 b15ztpn00an1n08x5 PHY_285 ();
 b15ztpn00an1n08x5 PHY_286 ();
 b15ztpn00an1n08x5 PHY_287 ();
 b15ztpn00an1n08x5 PHY_288 ();
 b15ztpn00an1n08x5 PHY_289 ();
 b15ztpn00an1n08x5 PHY_290 ();
 b15ztpn00an1n08x5 PHY_291 ();
 b15ztpn00an1n08x5 PHY_292 ();
 b15ztpn00an1n08x5 PHY_293 ();
 b15ztpn00an1n08x5 PHY_294 ();
 b15ztpn00an1n08x5 PHY_295 ();
 b15ztpn00an1n08x5 PHY_296 ();
 b15ztpn00an1n08x5 PHY_297 ();
 b15ztpn00an1n08x5 PHY_298 ();
 b15ztpn00an1n08x5 PHY_299 ();
 b15ztpn00an1n08x5 PHY_300 ();
 b15ztpn00an1n08x5 PHY_301 ();
 b15ztpn00an1n08x5 PHY_302 ();
 b15ztpn00an1n08x5 PHY_303 ();
 b15ztpn00an1n08x5 PHY_304 ();
 b15ztpn00an1n08x5 PHY_305 ();
 b15ztpn00an1n08x5 PHY_306 ();
 b15ztpn00an1n08x5 PHY_307 ();
 b15ztpn00an1n08x5 PHY_308 ();
 b15ztpn00an1n08x5 PHY_309 ();
 b15ztpn00an1n08x5 PHY_310 ();
 b15ztpn00an1n08x5 PHY_311 ();
 b15ztpn00an1n08x5 PHY_312 ();
 b15ztpn00an1n08x5 PHY_313 ();
 b15ztpn00an1n08x5 PHY_314 ();
 b15ztpn00an1n08x5 PHY_315 ();
 b15ztpn00an1n08x5 PHY_316 ();
 b15ztpn00an1n08x5 PHY_317 ();
 b15ztpn00an1n08x5 PHY_318 ();
 b15ztpn00an1n08x5 PHY_319 ();
 b15ztpn00an1n08x5 PHY_320 ();
 b15ztpn00an1n08x5 PHY_321 ();
 b15ztpn00an1n08x5 PHY_322 ();
 b15ztpn00an1n08x5 PHY_323 ();
 b15ztpn00an1n08x5 PHY_324 ();
 b15ztpn00an1n08x5 PHY_325 ();
 b15ztpn00an1n08x5 PHY_326 ();
 b15ztpn00an1n08x5 PHY_327 ();
 b15ztpn00an1n08x5 PHY_328 ();
 b15ztpn00an1n08x5 PHY_329 ();
 b15ztpn00an1n08x5 PHY_330 ();
 b15ztpn00an1n08x5 PHY_331 ();
 b15ztpn00an1n08x5 PHY_332 ();
 b15ztpn00an1n08x5 PHY_333 ();
 b15ztpn00an1n08x5 PHY_334 ();
 b15ztpn00an1n08x5 PHY_335 ();
 b15ztpn00an1n08x5 PHY_336 ();
 b15ztpn00an1n08x5 PHY_337 ();
 b15ztpn00an1n08x5 PHY_338 ();
 b15ztpn00an1n08x5 PHY_339 ();
 b15ztpn00an1n08x5 PHY_340 ();
 b15ztpn00an1n08x5 PHY_341 ();
 b15ztpn00an1n08x5 PHY_342 ();
 b15ztpn00an1n08x5 PHY_343 ();
 b15ztpn00an1n08x5 PHY_344 ();
 b15ztpn00an1n08x5 PHY_345 ();
 b15ztpn00an1n08x5 PHY_346 ();
 b15ztpn00an1n08x5 PHY_347 ();
 b15ztpn00an1n08x5 PHY_348 ();
 b15ztpn00an1n08x5 PHY_349 ();
 b15ztpn00an1n08x5 PHY_350 ();
 b15ztpn00an1n08x5 PHY_351 ();
 b15ztpn00an1n08x5 PHY_352 ();
 b15ztpn00an1n08x5 PHY_353 ();
 b15ztpn00an1n08x5 PHY_354 ();
 b15ztpn00an1n08x5 PHY_355 ();
 b15ztpn00an1n08x5 PHY_356 ();
 b15ztpn00an1n08x5 PHY_357 ();
 b15ztpn00an1n08x5 PHY_358 ();
 b15ztpn00an1n08x5 PHY_359 ();
 b15ztpn00an1n08x5 PHY_360 ();
 b15ztpn00an1n08x5 PHY_361 ();
 b15ztpn00an1n08x5 PHY_362 ();
 b15ztpn00an1n08x5 PHY_363 ();
 b15ztpn00an1n08x5 PHY_364 ();
 b15ztpn00an1n08x5 PHY_365 ();
 b15ztpn00an1n08x5 PHY_366 ();
 b15ztpn00an1n08x5 PHY_367 ();
 b15ztpn00an1n08x5 PHY_368 ();
 b15ztpn00an1n08x5 PHY_369 ();
 b15ztpn00an1n08x5 PHY_370 ();
 b15ztpn00an1n08x5 PHY_371 ();
 b15ztpn00an1n08x5 PHY_372 ();
 b15ztpn00an1n08x5 PHY_373 ();
 b15ztpn00an1n08x5 PHY_374 ();
 b15ztpn00an1n08x5 PHY_375 ();
 b15ztpn00an1n08x5 PHY_376 ();
 b15ztpn00an1n08x5 PHY_377 ();
 b15ztpn00an1n08x5 PHY_378 ();
 b15ztpn00an1n08x5 PHY_379 ();
 b15ztpn00an1n08x5 PHY_380 ();
 b15ztpn00an1n08x5 PHY_381 ();
 b15ztpn00an1n08x5 PHY_382 ();
 b15ztpn00an1n08x5 PHY_383 ();
 b15ztpn00an1n08x5 PHY_384 ();
 b15ztpn00an1n08x5 PHY_385 ();
 b15ztpn00an1n08x5 PHY_386 ();
 b15ztpn00an1n08x5 PHY_387 ();
 b15ztpn00an1n08x5 PHY_388 ();
 b15ztpn00an1n08x5 PHY_389 ();
 b15ztpn00an1n08x5 TAP_390 ();
 b15ztpn00an1n08x5 TAP_391 ();
 b15ztpn00an1n08x5 TAP_392 ();
 b15ztpn00an1n08x5 TAP_393 ();
 b15ztpn00an1n08x5 TAP_394 ();
 b15ztpn00an1n08x5 TAP_395 ();
 b15ztpn00an1n08x5 TAP_396 ();
 b15ztpn00an1n08x5 TAP_397 ();
 b15ztpn00an1n08x5 TAP_398 ();
 b15ztpn00an1n08x5 TAP_399 ();
 b15ztpn00an1n08x5 TAP_400 ();
 b15ztpn00an1n08x5 TAP_401 ();
 b15ztpn00an1n08x5 TAP_402 ();
 b15ztpn00an1n08x5 TAP_403 ();
 b15ztpn00an1n08x5 TAP_404 ();
 b15ztpn00an1n08x5 TAP_405 ();
 b15ztpn00an1n08x5 TAP_406 ();
 b15ztpn00an1n08x5 TAP_407 ();
 b15ztpn00an1n08x5 TAP_408 ();
 b15ztpn00an1n08x5 TAP_409 ();
 b15ztpn00an1n08x5 TAP_410 ();
 b15ztpn00an1n08x5 TAP_411 ();
 b15ztpn00an1n08x5 TAP_412 ();
 b15ztpn00an1n08x5 TAP_413 ();
 b15ztpn00an1n08x5 TAP_414 ();
 b15ztpn00an1n08x5 TAP_415 ();
 b15ztpn00an1n08x5 TAP_416 ();
 b15ztpn00an1n08x5 TAP_417 ();
 b15ztpn00an1n08x5 TAP_418 ();
 b15ztpn00an1n08x5 TAP_419 ();
 b15ztpn00an1n08x5 TAP_420 ();
 b15ztpn00an1n08x5 TAP_421 ();
 b15ztpn00an1n08x5 TAP_422 ();
 b15ztpn00an1n08x5 TAP_423 ();
 b15ztpn00an1n08x5 TAP_424 ();
 b15ztpn00an1n08x5 TAP_425 ();
 b15ztpn00an1n08x5 TAP_426 ();
 b15ztpn00an1n08x5 TAP_427 ();
 b15ztpn00an1n08x5 TAP_428 ();
 b15ztpn00an1n08x5 TAP_429 ();
 b15ztpn00an1n08x5 TAP_430 ();
 b15ztpn00an1n08x5 TAP_431 ();
 b15ztpn00an1n08x5 TAP_432 ();
 b15ztpn00an1n08x5 TAP_433 ();
 b15ztpn00an1n08x5 TAP_434 ();
 b15ztpn00an1n08x5 TAP_435 ();
 b15ztpn00an1n08x5 TAP_436 ();
 b15ztpn00an1n08x5 TAP_437 ();
 b15ztpn00an1n08x5 TAP_438 ();
 b15ztpn00an1n08x5 TAP_439 ();
 b15ztpn00an1n08x5 TAP_440 ();
 b15ztpn00an1n08x5 TAP_441 ();
 b15ztpn00an1n08x5 TAP_442 ();
 b15ztpn00an1n08x5 TAP_443 ();
 b15ztpn00an1n08x5 TAP_444 ();
 b15ztpn00an1n08x5 TAP_445 ();
 b15ztpn00an1n08x5 TAP_446 ();
 b15ztpn00an1n08x5 TAP_447 ();
 b15ztpn00an1n08x5 TAP_448 ();
 b15ztpn00an1n08x5 TAP_449 ();
 b15ztpn00an1n08x5 TAP_450 ();
 b15ztpn00an1n08x5 TAP_451 ();
 b15ztpn00an1n08x5 TAP_452 ();
 b15ztpn00an1n08x5 TAP_453 ();
 b15ztpn00an1n08x5 TAP_454 ();
 b15ztpn00an1n08x5 TAP_455 ();
 b15ztpn00an1n08x5 TAP_456 ();
 b15ztpn00an1n08x5 TAP_457 ();
 b15ztpn00an1n08x5 TAP_458 ();
 b15ztpn00an1n08x5 TAP_459 ();
 b15ztpn00an1n08x5 TAP_460 ();
 b15ztpn00an1n08x5 TAP_461 ();
 b15ztpn00an1n08x5 TAP_462 ();
 b15ztpn00an1n08x5 TAP_463 ();
 b15ztpn00an1n08x5 TAP_464 ();
 b15ztpn00an1n08x5 TAP_465 ();
 b15ztpn00an1n08x5 TAP_466 ();
 b15ztpn00an1n08x5 TAP_467 ();
 b15ztpn00an1n08x5 TAP_468 ();
 b15ztpn00an1n08x5 TAP_469 ();
 b15ztpn00an1n08x5 TAP_470 ();
 b15ztpn00an1n08x5 TAP_471 ();
 b15ztpn00an1n08x5 TAP_472 ();
 b15ztpn00an1n08x5 TAP_473 ();
 b15ztpn00an1n08x5 TAP_474 ();
 b15ztpn00an1n08x5 TAP_475 ();
 b15ztpn00an1n08x5 TAP_476 ();
 b15ztpn00an1n08x5 TAP_477 ();
 b15ztpn00an1n08x5 TAP_478 ();
 b15ztpn00an1n08x5 TAP_479 ();
 b15ztpn00an1n08x5 TAP_480 ();
 b15ztpn00an1n08x5 TAP_481 ();
 b15ztpn00an1n08x5 TAP_482 ();
 b15ztpn00an1n08x5 TAP_483 ();
 b15ztpn00an1n08x5 TAP_484 ();
 b15ztpn00an1n08x5 TAP_485 ();
 b15ztpn00an1n08x5 TAP_486 ();
 b15ztpn00an1n08x5 TAP_487 ();
 b15ztpn00an1n08x5 TAP_488 ();
 b15ztpn00an1n08x5 TAP_489 ();
 b15ztpn00an1n08x5 TAP_490 ();
 b15ztpn00an1n08x5 TAP_491 ();
 b15ztpn00an1n08x5 TAP_492 ();
 b15ztpn00an1n08x5 TAP_493 ();
 b15ztpn00an1n08x5 TAP_494 ();
 b15ztpn00an1n08x5 TAP_495 ();
 b15ztpn00an1n08x5 TAP_496 ();
 b15ztpn00an1n08x5 TAP_497 ();
 b15ztpn00an1n08x5 TAP_498 ();
 b15ztpn00an1n08x5 TAP_499 ();
 b15ztpn00an1n08x5 TAP_500 ();
 b15ztpn00an1n08x5 TAP_501 ();
 b15ztpn00an1n08x5 TAP_502 ();
 b15ztpn00an1n08x5 TAP_503 ();
 b15ztpn00an1n08x5 TAP_504 ();
 b15ztpn00an1n08x5 TAP_505 ();
 b15ztpn00an1n08x5 TAP_506 ();
 b15ztpn00an1n08x5 TAP_507 ();
 b15ztpn00an1n08x5 TAP_508 ();
 b15ztpn00an1n08x5 TAP_509 ();
 b15ztpn00an1n08x5 TAP_510 ();
 b15ztpn00an1n08x5 TAP_511 ();
 b15ztpn00an1n08x5 TAP_512 ();
 b15ztpn00an1n08x5 TAP_513 ();
 b15ztpn00an1n08x5 TAP_514 ();
 b15ztpn00an1n08x5 TAP_515 ();
 b15ztpn00an1n08x5 TAP_516 ();
 b15ztpn00an1n08x5 TAP_517 ();
 b15ztpn00an1n08x5 TAP_518 ();
 b15ztpn00an1n08x5 TAP_519 ();
 b15ztpn00an1n08x5 TAP_520 ();
 b15ztpn00an1n08x5 TAP_521 ();
 b15ztpn00an1n08x5 TAP_522 ();
 b15ztpn00an1n08x5 TAP_523 ();
 b15ztpn00an1n08x5 TAP_524 ();
 b15ztpn00an1n08x5 TAP_525 ();
 b15ztpn00an1n08x5 TAP_526 ();
 b15ztpn00an1n08x5 TAP_527 ();
 b15ztpn00an1n08x5 TAP_528 ();
 b15ztpn00an1n08x5 TAP_529 ();
 b15ztpn00an1n08x5 TAP_530 ();
 b15ztpn00an1n08x5 TAP_531 ();
 b15ztpn00an1n08x5 TAP_532 ();
 b15ztpn00an1n08x5 TAP_533 ();
 b15ztpn00an1n08x5 TAP_534 ();
 b15ztpn00an1n08x5 TAP_535 ();
 b15ztpn00an1n08x5 TAP_536 ();
 b15ztpn00an1n08x5 TAP_537 ();
 b15ztpn00an1n08x5 TAP_538 ();
 b15ztpn00an1n08x5 TAP_539 ();
 b15ztpn00an1n08x5 TAP_540 ();
 b15ztpn00an1n08x5 TAP_541 ();
 b15ztpn00an1n08x5 TAP_542 ();
 b15ztpn00an1n08x5 TAP_543 ();
 b15ztpn00an1n08x5 TAP_544 ();
 b15ztpn00an1n08x5 TAP_545 ();
 b15ztpn00an1n08x5 TAP_546 ();
 b15ztpn00an1n08x5 TAP_547 ();
 b15ztpn00an1n08x5 TAP_548 ();
 b15ztpn00an1n08x5 TAP_549 ();
 b15ztpn00an1n08x5 TAP_550 ();
 b15ztpn00an1n08x5 TAP_551 ();
 b15ztpn00an1n08x5 TAP_552 ();
 b15ztpn00an1n08x5 TAP_553 ();
 b15ztpn00an1n08x5 TAP_554 ();
 b15ztpn00an1n08x5 TAP_555 ();
 b15ztpn00an1n08x5 TAP_556 ();
 b15ztpn00an1n08x5 TAP_557 ();
 b15ztpn00an1n08x5 TAP_558 ();
 b15ztpn00an1n08x5 TAP_559 ();
 b15ztpn00an1n08x5 TAP_560 ();
 b15ztpn00an1n08x5 TAP_561 ();
 b15ztpn00an1n08x5 TAP_562 ();
 b15ztpn00an1n08x5 TAP_563 ();
 b15ztpn00an1n08x5 TAP_564 ();
 b15ztpn00an1n08x5 TAP_565 ();
 b15ztpn00an1n08x5 TAP_566 ();
 b15ztpn00an1n08x5 TAP_567 ();
 b15ztpn00an1n08x5 TAP_568 ();
 b15ztpn00an1n08x5 TAP_569 ();
 b15ztpn00an1n08x5 TAP_570 ();
 b15ztpn00an1n08x5 TAP_571 ();
 b15ztpn00an1n08x5 TAP_572 ();
 b15ztpn00an1n08x5 TAP_573 ();
 b15ztpn00an1n08x5 TAP_574 ();
 b15ztpn00an1n08x5 TAP_575 ();
 b15ztpn00an1n08x5 TAP_576 ();
 b15ztpn00an1n08x5 TAP_577 ();
 b15ztpn00an1n08x5 TAP_578 ();
 b15ztpn00an1n08x5 TAP_579 ();
 b15ztpn00an1n08x5 TAP_580 ();
 b15ztpn00an1n08x5 TAP_581 ();
 b15ztpn00an1n08x5 TAP_582 ();
 b15ztpn00an1n08x5 TAP_583 ();
 b15ztpn00an1n08x5 TAP_584 ();
 b15ztpn00an1n08x5 TAP_585 ();
 b15ztpn00an1n08x5 TAP_586 ();
 b15ztpn00an1n08x5 TAP_587 ();
 b15ztpn00an1n08x5 TAP_588 ();
 b15ztpn00an1n08x5 TAP_589 ();
 b15ztpn00an1n08x5 TAP_590 ();
 b15ztpn00an1n08x5 TAP_591 ();
 b15ztpn00an1n08x5 TAP_592 ();
 b15ztpn00an1n08x5 TAP_593 ();
 b15ztpn00an1n08x5 TAP_594 ();
 b15ztpn00an1n08x5 TAP_595 ();
 b15ztpn00an1n08x5 TAP_596 ();
 b15ztpn00an1n08x5 TAP_597 ();
 b15ztpn00an1n08x5 TAP_598 ();
 b15ztpn00an1n08x5 TAP_599 ();
 b15ztpn00an1n08x5 TAP_600 ();
 b15ztpn00an1n08x5 TAP_601 ();
 b15ztpn00an1n08x5 TAP_602 ();
 b15ztpn00an1n08x5 TAP_603 ();
 b15ztpn00an1n08x5 TAP_604 ();
 b15ztpn00an1n08x5 TAP_605 ();
 b15ztpn00an1n08x5 TAP_606 ();
 b15ztpn00an1n08x5 TAP_607 ();
 b15ztpn00an1n08x5 TAP_608 ();
 b15ztpn00an1n08x5 TAP_609 ();
 b15ztpn00an1n08x5 TAP_610 ();
 b15ztpn00an1n08x5 TAP_611 ();
 b15ztpn00an1n08x5 TAP_612 ();
 b15ztpn00an1n08x5 TAP_613 ();
 b15ztpn00an1n08x5 TAP_614 ();
 b15ztpn00an1n08x5 TAP_615 ();
 b15ztpn00an1n08x5 TAP_616 ();
 b15ztpn00an1n08x5 TAP_617 ();
 b15ztpn00an1n08x5 TAP_618 ();
 b15ztpn00an1n08x5 TAP_619 ();
 b15ztpn00an1n08x5 TAP_620 ();
 b15ztpn00an1n08x5 TAP_621 ();
 b15ztpn00an1n08x5 TAP_622 ();
 b15ztpn00an1n08x5 TAP_623 ();
 b15ztpn00an1n08x5 TAP_624 ();
 b15ztpn00an1n08x5 TAP_625 ();
 b15ztpn00an1n08x5 TAP_626 ();
 b15ztpn00an1n08x5 TAP_627 ();
 b15ztpn00an1n08x5 TAP_628 ();
 b15ztpn00an1n08x5 TAP_629 ();
 b15ztpn00an1n08x5 TAP_630 ();
 b15ztpn00an1n08x5 TAP_631 ();
 b15ztpn00an1n08x5 TAP_632 ();
 b15ztpn00an1n08x5 TAP_633 ();
 b15ztpn00an1n08x5 TAP_634 ();
 b15ztpn00an1n08x5 TAP_635 ();
 b15ztpn00an1n08x5 TAP_636 ();
 b15ztpn00an1n08x5 TAP_637 ();
 b15ztpn00an1n08x5 TAP_638 ();
 b15ztpn00an1n08x5 TAP_639 ();
 b15ztpn00an1n08x5 TAP_640 ();
 b15ztpn00an1n08x5 TAP_641 ();
 b15ztpn00an1n08x5 TAP_642 ();
 b15ztpn00an1n08x5 TAP_643 ();
 b15ztpn00an1n08x5 TAP_644 ();
 b15ztpn00an1n08x5 TAP_645 ();
 b15ztpn00an1n08x5 TAP_646 ();
 b15ztpn00an1n08x5 TAP_647 ();
 b15ztpn00an1n08x5 TAP_648 ();
 b15ztpn00an1n08x5 TAP_649 ();
 b15ztpn00an1n08x5 TAP_650 ();
 b15ztpn00an1n08x5 TAP_651 ();
 b15ztpn00an1n08x5 TAP_652 ();
 b15ztpn00an1n08x5 TAP_653 ();
 b15ztpn00an1n08x5 TAP_654 ();
 b15ztpn00an1n08x5 TAP_655 ();
 b15ztpn00an1n08x5 TAP_656 ();
 b15ztpn00an1n08x5 TAP_657 ();
 b15ztpn00an1n08x5 TAP_658 ();
 b15ztpn00an1n08x5 TAP_659 ();
 b15ztpn00an1n08x5 TAP_660 ();
 b15ztpn00an1n08x5 TAP_661 ();
 b15ztpn00an1n08x5 TAP_662 ();
 b15ztpn00an1n08x5 TAP_663 ();
 b15ztpn00an1n08x5 TAP_664 ();
 b15ztpn00an1n08x5 TAP_665 ();
 b15ztpn00an1n08x5 TAP_666 ();
 b15ztpn00an1n08x5 TAP_667 ();
 b15ztpn00an1n08x5 TAP_668 ();
 b15ztpn00an1n08x5 TAP_669 ();
 b15ztpn00an1n08x5 TAP_670 ();
 b15ztpn00an1n08x5 TAP_671 ();
 b15ztpn00an1n08x5 TAP_672 ();
 b15ztpn00an1n08x5 TAP_673 ();
 b15ztpn00an1n08x5 TAP_674 ();
 b15ztpn00an1n08x5 TAP_675 ();
 b15ztpn00an1n08x5 TAP_676 ();
 b15ztpn00an1n08x5 TAP_677 ();
 b15ztpn00an1n08x5 TAP_678 ();
 b15ztpn00an1n08x5 TAP_679 ();
 b15ztpn00an1n08x5 TAP_680 ();
 b15ztpn00an1n08x5 TAP_681 ();
 b15ztpn00an1n08x5 TAP_682 ();
 b15ztpn00an1n08x5 TAP_683 ();
 b15ztpn00an1n08x5 TAP_684 ();
 b15ztpn00an1n08x5 TAP_685 ();
 b15ztpn00an1n08x5 TAP_686 ();
 b15ztpn00an1n08x5 TAP_687 ();
 b15ztpn00an1n08x5 TAP_688 ();
 b15ztpn00an1n08x5 TAP_689 ();
 b15ztpn00an1n08x5 TAP_690 ();
 b15ztpn00an1n08x5 TAP_691 ();
 b15ztpn00an1n08x5 TAP_692 ();
 b15ztpn00an1n08x5 TAP_693 ();
 b15ztpn00an1n08x5 TAP_694 ();
 b15ztpn00an1n08x5 TAP_695 ();
 b15ztpn00an1n08x5 TAP_696 ();
 b15ztpn00an1n08x5 TAP_697 ();
 b15ztpn00an1n08x5 TAP_698 ();
 b15ztpn00an1n08x5 TAP_699 ();
 b15ztpn00an1n08x5 TAP_700 ();
 b15ztpn00an1n08x5 TAP_701 ();
 b15ztpn00an1n08x5 TAP_702 ();
 b15ztpn00an1n08x5 TAP_703 ();
 b15ztpn00an1n08x5 TAP_704 ();
 b15ztpn00an1n08x5 TAP_705 ();
 b15ztpn00an1n08x5 TAP_706 ();
 b15ztpn00an1n08x5 TAP_707 ();
 b15ztpn00an1n08x5 TAP_708 ();
 b15ztpn00an1n08x5 TAP_709 ();
 b15ztpn00an1n08x5 TAP_710 ();
 b15ztpn00an1n08x5 TAP_711 ();
 b15ztpn00an1n08x5 TAP_712 ();
 b15ztpn00an1n08x5 TAP_713 ();
 b15ztpn00an1n08x5 TAP_714 ();
 b15ztpn00an1n08x5 TAP_715 ();
 b15ztpn00an1n08x5 TAP_716 ();
 b15ztpn00an1n08x5 TAP_717 ();
 b15ztpn00an1n08x5 TAP_718 ();
 b15ztpn00an1n08x5 TAP_719 ();
 b15ztpn00an1n08x5 TAP_720 ();
 b15ztpn00an1n08x5 TAP_721 ();
 b15ztpn00an1n08x5 TAP_722 ();
 b15ztpn00an1n08x5 TAP_723 ();
 b15ztpn00an1n08x5 TAP_724 ();
 b15ztpn00an1n08x5 TAP_725 ();
 b15ztpn00an1n08x5 TAP_726 ();
 b15ztpn00an1n08x5 TAP_727 ();
 b15ztpn00an1n08x5 TAP_728 ();
 b15ztpn00an1n08x5 TAP_729 ();
 b15ztpn00an1n08x5 TAP_730 ();
 b15ztpn00an1n08x5 TAP_731 ();
 b15ztpn00an1n08x5 TAP_732 ();
 b15ztpn00an1n08x5 TAP_733 ();
 b15ztpn00an1n08x5 TAP_734 ();
 b15ztpn00an1n08x5 TAP_735 ();
 b15ztpn00an1n08x5 TAP_736 ();
 b15ztpn00an1n08x5 TAP_737 ();
 b15ztpn00an1n08x5 TAP_738 ();
 b15ztpn00an1n08x5 TAP_739 ();
 b15ztpn00an1n08x5 TAP_740 ();
 b15ztpn00an1n08x5 TAP_741 ();
 b15ztpn00an1n08x5 TAP_742 ();
 b15ztpn00an1n08x5 TAP_743 ();
 b15ztpn00an1n08x5 TAP_744 ();
 b15ztpn00an1n08x5 TAP_745 ();
 b15ztpn00an1n08x5 TAP_746 ();
 b15ztpn00an1n08x5 TAP_747 ();
 b15ztpn00an1n08x5 TAP_748 ();
 b15ztpn00an1n08x5 TAP_749 ();
 b15ztpn00an1n08x5 TAP_750 ();
 b15ztpn00an1n08x5 TAP_751 ();
 b15ztpn00an1n08x5 TAP_752 ();
 b15ztpn00an1n08x5 TAP_753 ();
 b15ztpn00an1n08x5 TAP_754 ();
 b15ztpn00an1n08x5 TAP_755 ();
 b15ztpn00an1n08x5 TAP_756 ();
 b15ztpn00an1n08x5 TAP_757 ();
 b15ztpn00an1n08x5 TAP_758 ();
 b15ztpn00an1n08x5 TAP_759 ();
 b15ztpn00an1n08x5 TAP_760 ();
 b15ztpn00an1n08x5 TAP_761 ();
 b15ztpn00an1n08x5 TAP_762 ();
 b15ztpn00an1n08x5 TAP_763 ();
 b15ztpn00an1n08x5 TAP_764 ();
 b15ztpn00an1n08x5 TAP_765 ();
 b15ztpn00an1n08x5 TAP_766 ();
 b15ztpn00an1n08x5 TAP_767 ();
 b15ztpn00an1n08x5 TAP_768 ();
 b15ztpn00an1n08x5 TAP_769 ();
 b15ztpn00an1n08x5 TAP_770 ();
 b15ztpn00an1n08x5 TAP_771 ();
 b15ztpn00an1n08x5 TAP_772 ();
 b15ztpn00an1n08x5 TAP_773 ();
 b15ztpn00an1n08x5 TAP_774 ();
 b15ztpn00an1n08x5 TAP_775 ();
 b15ztpn00an1n08x5 TAP_776 ();
 b15ztpn00an1n08x5 TAP_777 ();
 b15ztpn00an1n08x5 TAP_778 ();
 b15ztpn00an1n08x5 TAP_779 ();
 b15ztpn00an1n08x5 TAP_780 ();
 b15bfn001as1n06x5 input1 (.a(alert_rx_i[0]),
    .o(net1));
 b15bfn001as1n06x5 input2 (.a(alert_rx_i[1]),
    .o(net2));
 b15bfn000ah1n06x5 input3 (.a(alert_rx_i[2]),
    .o(net3));
 b15bfn000ah1n06x5 input4 (.a(alert_rx_i[3]),
    .o(net4));
 b15bfn001aq1n06x5 input5 (.a(cio_gpio_i[0]),
    .o(net5));
 b15bfn000as1n06x5 input6 (.a(cio_gpio_i[10]),
    .o(net6));
 b15bfn000as1n04x5 input7 (.a(cio_gpio_i[11]),
    .o(net7));
 b15bfn000ah1n04x5 input8 (.a(cio_gpio_i[12]),
    .o(net8));
 b15bfn000an1n02x5 input9 (.a(cio_gpio_i[13]),
    .o(net9));
 b15bfn001as1n06x5 input10 (.a(cio_gpio_i[14]),
    .o(net10));
 b15bfn000ah1n06x5 input11 (.a(cio_gpio_i[15]),
    .o(net11));
 b15bfn000as1n06x5 input12 (.a(cio_gpio_i[16]),
    .o(net12));
 b15bfn000ah1n06x5 input13 (.a(cio_gpio_i[17]),
    .o(net13));
 b15bfn000ah1n02x5 input14 (.a(cio_gpio_i[18]),
    .o(net14));
 b15bfn000an1n02x5 input15 (.a(cio_gpio_i[19]),
    .o(net15));
 b15bfn000ah1n04x5 input16 (.a(cio_gpio_i[1]),
    .o(net16));
 b15bfn000al1n02x5 input17 (.a(cio_gpio_i[20]),
    .o(net17));
 b15bfn000as1n04x5 input18 (.a(cio_gpio_i[21]),
    .o(net18));
 b15bfn001ah1n08x5 input19 (.a(cio_gpio_i[22]),
    .o(net19));
 b15bfn000as1n02x5 input20 (.a(cio_gpio_i[23]),
    .o(net20));
 b15bfn001ah1n08x5 input21 (.a(cio_gpio_i[24]),
    .o(net21));
 b15bfm201as1n04x5 input22 (.a(cio_gpio_i[25]),
    .o(net22));
 b15bfn000as1n03x5 input23 (.a(cio_gpio_i[26]),
    .o(net23));
 b15bfn001as1n08x5 input24 (.a(cio_gpio_i[27]),
    .o(net24));
 b15bfn000as1n03x5 input25 (.a(cio_gpio_i[28]),
    .o(net25));
 b15bfn000ah1n03x5 input26 (.a(cio_gpio_i[29]),
    .o(net26));
 b15bfn001aq1n06x5 input27 (.a(cio_gpio_i[2]),
    .o(net27));
 b15bfn000ah1n02x5 input28 (.a(cio_gpio_i[30]),
    .o(net28));
 b15bfn001as1n06x5 input29 (.a(cio_gpio_i[31]),
    .o(net29));
 b15bfn000ah1n03x5 input30 (.a(cio_gpio_i[3]),
    .o(net30));
 b15bfn000ah1n03x5 input31 (.a(cio_gpio_i[4]),
    .o(net31));
 b15bfn000as1n04x5 input32 (.a(cio_gpio_i[5]),
    .o(net32));
 b15bfn000ah1n06x5 input33 (.a(cio_gpio_i[6]),
    .o(net33));
 b15bfn001ah1n12x5 input34 (.a(cio_gpio_i[7]),
    .o(net34));
 b15bfn001ah1n08x5 input35 (.a(cio_gpio_i[8]),
    .o(net35));
 b15bfn000as1n04x5 input36 (.a(cio_gpio_i[9]),
    .o(net36));
 b15bfn001as1n48x5 input37 (.a(net2444),
    .o(net37));
 b15bfn000aq1n02x5 input38 (.a(tl_i[0]),
    .o(net38));
 b15bfn001as1n12x5 input39 (.a(tl_i[100]),
    .o(net39));
 b15bfn001as1n12x5 input40 (.a(tl_i[101]),
    .o(net40));
 b15bfn001as1n12x5 input41 (.a(tl_i[105]),
    .o(net41));
 b15bfn001as1n08x5 input42 (.a(tl_i[106]),
    .o(net42));
 b15bfn001as1n16x5 input43 (.a(tl_i[107]),
    .o(net43));
 b15bfn001ah1n12x5 input44 (.a(tl_i[108]),
    .o(net44));
 b15bfn000ah1n04x5 input45 (.a(tl_i[10]),
    .o(net45));
 b15bfm201as1n04x5 input46 (.a(tl_i[11]),
    .o(net46));
 b15bfn000ah1n06x5 input47 (.a(tl_i[12]),
    .o(net47));
 b15bfn000ah1n04x5 input48 (.a(tl_i[13]),
    .o(net48));
 b15bfn000as1n04x5 input49 (.a(tl_i[14]),
    .o(net49));
 b15bfn001ah1n12x5 input50 (.a(tl_i[15]),
    .o(net50));
 b15bfn001as1n12x5 input51 (.a(tl_i[16]),
    .o(net51));
 b15bfn001as1n08x5 input52 (.a(tl_i[17]),
    .o(net52));
 b15bfn000as1n12x5 input53 (.a(tl_i[18]),
    .o(net53));
 b15bfn001as1n16x5 input54 (.a(tl_i[1]),
    .o(net54));
 b15bfn001as1n24x5 input55 (.a(tl_i[24]),
    .o(net55));
 b15bfn001as1n24x5 input56 (.a(tl_i[25]),
    .o(net56));
 b15bfn001as1n06x5 input57 (.a(tl_i[26]),
    .o(net57));
 b15bfn001as1n24x5 input58 (.a(tl_i[27]),
    .o(net58));
 b15bfn001as1n16x5 input59 (.a(tl_i[28]),
    .o(net59));
 b15bfn001as1n24x5 input60 (.a(tl_i[29]),
    .o(net60));
 b15bfn001as1n06x5 input61 (.a(tl_i[2]),
    .o(net61));
 b15bfn001as1n32x5 input62 (.a(tl_i[30]),
    .o(net62));
 b15bfn001ah1n48x5 input63 (.a(tl_i[31]),
    .o(net63));
 b15bfn001as1n24x5 input64 (.a(tl_i[32]),
    .o(net64));
 b15bfn001as1n32x5 input65 (.a(tl_i[33]),
    .o(net65));
 b15bfn001as1n32x5 input66 (.a(tl_i[34]),
    .o(net66));
 b15bfn001as1n32x5 input67 (.a(tl_i[35]),
    .o(net67));
 b15bfn001ah1n48x5 input68 (.a(tl_i[36]),
    .o(net68));
 b15bfn000as1n32x5 input69 (.a(tl_i[37]),
    .o(net69));
 b15bfn001as1n24x5 input70 (.a(tl_i[38]),
    .o(net70));
 b15bfn001as1n16x5 input71 (.a(tl_i[39]),
    .o(net71));
 b15bfn001as1n12x5 input72 (.a(tl_i[3]),
    .o(net72));
 b15bfn001ah1n64x5 input73 (.a(tl_i[40]),
    .o(net73));
 b15bfn001as1n48x5 input74 (.a(tl_i[41]),
    .o(net74));
 b15bfn001as1n48x5 input75 (.a(tl_i[42]),
    .o(net75));
 b15bfn001as1n48x5 input76 (.a(tl_i[43]),
    .o(net76));
 b15bfn001ah1n32x5 input77 (.a(tl_i[44]),
    .o(net77));
 b15bfn001as1n32x5 input78 (.a(tl_i[45]),
    .o(net78));
 b15bfn001ah1n48x5 input79 (.a(tl_i[46]),
    .o(net79));
 b15bfn001as1n48x5 input80 (.a(tl_i[47]),
    .o(net80));
 b15bfn001as1n24x5 input81 (.a(tl_i[48]),
    .o(net81));
 b15bfn001as1n24x5 input82 (.a(tl_i[49]),
    .o(net82));
 b15bfn000ah1n06x5 input83 (.a(tl_i[4]),
    .o(net83));
 b15bfn000ah1n48x5 input84 (.a(tl_i[50]),
    .o(net84));
 b15bfn001ah1n48x5 input85 (.a(tl_i[51]),
    .o(net85));
 b15bfn001as1n48x5 input86 (.a(tl_i[52]),
    .o(net86));
 b15bfn001as1n32x5 input87 (.a(tl_i[53]),
    .o(net87));
 b15bfn001ah1n48x5 input88 (.a(tl_i[54]),
    .o(net88));
 b15bfn001ah1n48x5 input89 (.a(tl_i[55]),
    .o(net89));
 b15bfn001ah1n16x5 input90 (.a(tl_i[56]),
    .o(net90));
 b15bfn001as1n12x5 input91 (.a(tl_i[57]),
    .o(net91));
 b15bfn001as1n12x5 input92 (.a(tl_i[58]),
    .o(net92));
 b15bfn001ah1n16x5 input93 (.a(tl_i[59]),
    .o(net93));
 b15bfn001ah1n16x5 input94 (.a(tl_i[5]),
    .o(net94));
 b15bfn001as1n16x5 input95 (.a(tl_i[60]),
    .o(net95));
 b15bfn001ah1n12x5 input96 (.a(tl_i[61]),
    .o(net96));
 b15bfn001as1n12x5 input97 (.a(tl_i[62]),
    .o(net97));
 b15bfn001as1n32x5 input98 (.a(tl_i[63]),
    .o(net98));
 b15bfn001as1n24x5 input99 (.a(tl_i[64]),
    .o(net99));
 b15bfn001ah1n48x5 input100 (.a(tl_i[65]),
    .o(net100));
 b15bfn001as1n08x5 input101 (.a(tl_i[66]),
    .o(net101));
 b15bfn001ah1n08x5 input102 (.a(tl_i[67]),
    .o(net102));
 b15bfn001ah1n08x5 input103 (.a(tl_i[68]),
    .o(net103));
 b15bfn001aq1n06x5 input104 (.a(tl_i[69]),
    .o(net104));
 b15bfn001as1n16x5 input105 (.a(tl_i[6]),
    .o(net105));
 b15bfn000ah1n06x5 input106 (.a(tl_i[70]),
    .o(net106));
 b15bfn001as1n06x5 input107 (.a(tl_i[71]),
    .o(net107));
 b15bfn001ah1n12x5 input108 (.a(tl_i[72]),
    .o(net108));
 b15bfn001ah1n08x5 input109 (.a(tl_i[73]),
    .o(net109));
 b15bfn001ah1n08x5 input110 (.a(tl_i[74]),
    .o(net110));
 b15bfn001as1n08x5 input111 (.a(tl_i[75]),
    .o(net111));
 b15bfn001ah1n08x5 input112 (.a(tl_i[76]),
    .o(net112));
 b15bfn001ah1n08x5 input113 (.a(tl_i[77]),
    .o(net113));
 b15bfn001ah1n12x5 input114 (.a(tl_i[78]),
    .o(net114));
 b15bfn001as1n06x5 input115 (.a(tl_i[79]),
    .o(net115));
 b15bfn001as1n12x5 input116 (.a(tl_i[7]),
    .o(net116));
 b15bfn001as1n08x5 input117 (.a(tl_i[80]),
    .o(net117));
 b15bfn001as1n08x5 input118 (.a(tl_i[81]),
    .o(net118));
 b15bfn001as1n08x5 input119 (.a(tl_i[82]),
    .o(net119));
 b15bfn001ah1n12x5 input120 (.a(tl_i[83]),
    .o(net120));
 b15bfn001ah1n08x5 input121 (.a(tl_i[84]),
    .o(net121));
 b15bfn001ah1n08x5 input122 (.a(tl_i[85]),
    .o(net122));
 b15bfn001as1n08x5 input123 (.a(tl_i[86]),
    .o(net123));
 b15bfn001as1n12x5 input124 (.a(tl_i[87]),
    .o(net124));
 b15bfn001ah1n12x5 input125 (.a(tl_i[88]),
    .o(net125));
 b15bfn001ah1n08x5 input126 (.a(tl_i[89]),
    .o(net126));
 b15bfn001aq1n06x5 input127 (.a(tl_i[8]),
    .o(net127));
 b15bfn001as1n08x5 input128 (.a(tl_i[90]),
    .o(net128));
 b15bfn001ah1n16x5 input129 (.a(tl_i[91]),
    .o(net129));
 b15bfn000as1n02x5 input130 (.a(tl_i[92]),
    .o(net130));
 b15bfn000as1n02x5 input131 (.a(tl_i[93]),
    .o(net131));
 b15bfn000as1n02x5 input132 (.a(tl_i[94]),
    .o(net132));
 b15bfn000as1n02x5 input133 (.a(tl_i[95]),
    .o(net133));
 b15bfn000ah1n02x5 input134 (.a(tl_i[96]),
    .o(net134));
 b15bfn000ah1n02x5 input135 (.a(tl_i[97]),
    .o(net135));
 b15bfn000as1n02x5 input136 (.a(tl_i[98]),
    .o(net136));
 b15bfn000as1n02x5 input137 (.a(tl_i[99]),
    .o(net137));
 b15bfn001aq1n06x5 input138 (.a(tl_i[9]),
    .o(net138));
 b15bfn000ah1n03x5 output139 (.a(net2517),
    .o(net1922));
 b15bfn000ah1n03x5 output140 (.a(net2515),
    .o(net1917));
 b15bfn000ah1n03x5 output141 (.a(net666),
    .o(cio_gpio_en_o[0]));
 b15bfn000ah1n03x5 output142 (.a(net142),
    .o(cio_gpio_en_o[10]));
 b15bfn000ah1n03x5 output143 (.a(net143),
    .o(cio_gpio_en_o[11]));
 b15bfn000ah1n03x5 output144 (.a(net660),
    .o(cio_gpio_en_o[12]));
 b15bfn000ah1n03x5 output145 (.a(net145),
    .o(cio_gpio_en_o[13]));
 b15bfn000ah1n03x5 output146 (.a(net146),
    .o(cio_gpio_en_o[14]));
 b15bfn000ah1n03x5 output147 (.a(net2477),
    .o(cio_gpio_en_o[15]));
 b15bfn000ah1n03x5 output148 (.a(net659),
    .o(cio_gpio_en_o[16]));
 b15bfn000ah1n03x5 output149 (.a(net2148),
    .o(cio_gpio_en_o[17]));
 b15bfn000ah1n03x5 output150 (.a(net2039),
    .o(net2040));
 b15bfn000ah1n03x5 output151 (.a(net2173),
    .o(cio_gpio_en_o[19]));
 b15bfn000ah1n03x5 output152 (.a(net663),
    .o(cio_gpio_en_o[1]));
 b15bfn000ah1n03x5 output153 (.a(net656),
    .o(cio_gpio_en_o[20]));
 b15bfn000ah1n03x5 output154 (.a(net2084),
    .o(cio_gpio_en_o[21]));
 b15bfn000ah1n03x5 output155 (.a(net653),
    .o(cio_gpio_en_o[22]));
 b15bfn000ah1n03x5 output156 (.a(net2051),
    .o(cio_gpio_en_o[23]));
 b15bfn000ah1n03x5 output157 (.a(net649),
    .o(cio_gpio_en_o[24]));
 b15bfn000ah1n03x5 output158 (.a(net648),
    .o(cio_gpio_en_o[25]));
 b15bfn000ah1n03x5 output159 (.a(net647),
    .o(cio_gpio_en_o[26]));
 b15bfn000ah1n03x5 output160 (.a(net2099),
    .o(cio_gpio_en_o[27]));
 b15bfn000ah1n03x5 output161 (.a(net2060),
    .o(net2061));
 b15bfn000ah1n03x5 output162 (.a(net2081),
    .o(net2082));
 b15bfn000ah1n03x5 output163 (.a(net2445),
    .o(cio_gpio_en_o[2]));
 b15bfn000ah1n03x5 output164 (.a(net2183),
    .o(cio_gpio_en_o[30]));
 b15bfn000ah1n03x5 output165 (.a(net2041),
    .o(net2042));
 b15bfn000ah1n03x5 output166 (.a(net2439),
    .o(cio_gpio_en_o[3]));
 b15bfn000ah1n03x5 output167 (.a(net642),
    .o(cio_gpio_en_o[4]));
 b15bfn000ah1n03x5 output168 (.a(net641),
    .o(cio_gpio_en_o[5]));
 b15bfn000ah1n03x5 output169 (.a(net169),
    .o(cio_gpio_en_o[6]));
 b15bfn000ah1n03x5 output170 (.a(net170),
    .o(cio_gpio_en_o[7]));
 b15bfn000ah1n03x5 output171 (.a(net171),
    .o(cio_gpio_en_o[8]));
 b15bfn000ah1n03x5 output172 (.a(net172),
    .o(cio_gpio_en_o[9]));
 b15bfn000ah1n03x5 output173 (.a(net2020),
    .o(net2021));
 b15bfn000ah1n03x5 output174 (.a(net2240),
    .o(cio_gpio_o[10]));
 b15bfn000ah1n03x5 output175 (.a(net2069),
    .o(cio_gpio_o[11]));
 b15bfn000ah1n03x5 output176 (.a(net2185),
    .o(cio_gpio_o[12]));
 b15bfn000ah1n03x5 output177 (.a(net635),
    .o(cio_gpio_o[13]));
 b15bfn000ah1n03x5 output178 (.a(net633),
    .o(cio_gpio_o[14]));
 b15bfn000ah1n03x5 output179 (.a(net2235),
    .o(cio_gpio_o[15]));
 b15bfn000ah1n03x5 output180 (.a(net180),
    .o(cio_gpio_o[16]));
 b15bfn000ah1n03x5 output181 (.a(net181),
    .o(cio_gpio_o[17]));
 b15bfn000ah1n03x5 output182 (.a(net632),
    .o(cio_gpio_o[18]));
 b15bfn000ah1n03x5 output183 (.a(net629),
    .o(cio_gpio_o[19]));
 b15bfn000ah1n03x5 output184 (.a(net2026),
    .o(net2027));
 b15bfn000ah1n03x5 output185 (.a(net628),
    .o(cio_gpio_o[20]));
 b15bfn000ah1n03x5 output186 (.a(net627),
    .o(cio_gpio_o[21]));
 b15bfn000ah1n03x5 output187 (.a(net625),
    .o(cio_gpio_o[22]));
 b15bfn000ah1n03x5 output188 (.a(net623),
    .o(cio_gpio_o[23]));
 b15bfn000ah1n03x5 output189 (.a(net622),
    .o(cio_gpio_o[24]));
 b15bfn000ah1n03x5 output190 (.a(net621),
    .o(cio_gpio_o[25]));
 b15bfn000ah1n03x5 output191 (.a(net619),
    .o(cio_gpio_o[26]));
 b15bfn000ah1n03x5 output192 (.a(net618),
    .o(cio_gpio_o[27]));
 b15bfn000ah1n03x5 output193 (.a(net2379),
    .o(cio_gpio_o[28]));
 b15bfn000ah1n03x5 output194 (.a(net616),
    .o(cio_gpio_o[29]));
 b15bfn000ah1n03x5 output195 (.a(net2077),
    .o(net2078));
 b15bfn000ah1n03x5 output196 (.a(net196),
    .o(cio_gpio_o[30]));
 b15bfn000ah1n03x5 output197 (.a(net197),
    .o(cio_gpio_o[31]));
 b15bfn000ah1n03x5 output198 (.a(net2096),
    .o(net2097));
 b15bfn000ah1n03x5 output199 (.a(net615),
    .o(cio_gpio_o[4]));
 b15bfn000ah1n03x5 output200 (.a(net2323),
    .o(cio_gpio_o[5]));
 b15bfn000ah1n03x5 output201 (.a(net2116),
    .o(cio_gpio_o[6]));
 b15bfn000ah1n03x5 output202 (.a(net612),
    .o(cio_gpio_o[7]));
 b15bfn000ah1n03x5 output203 (.a(net2036),
    .o(net2037));
 b15bfn000ah1n03x5 output204 (.a(net2111),
    .o(cio_gpio_o[9]));
 b15bfn000ah1n03x5 output205 (.a(net2521),
    .o(net1924));
 b15bfn000ah1n03x5 output206 (.a(net2529),
    .o(net1936));
 b15bfn000ah1n03x5 output207 (.a(net2533),
    .o(net1943));
 b15bfn000ah1n03x5 output208 (.a(net2505),
    .o(net1911));
 b15bfn000ah1n03x5 output209 (.a(net2501),
    .o(net1909));
 b15bfn000ah1n03x5 output210 (.a(net1937),
    .o(net1938));
 b15bfn000ah1n03x5 output211 (.a(net1939),
    .o(net1940));
 b15bfn000ah1n03x5 output212 (.a(net2486),
    .o(net1889));
 b15bfn000ah1n03x5 output213 (.a(net2483),
    .o(net1887));
 b15bfn000ah1n03x5 output214 (.a(net2503),
    .o(net1907));
 b15bfn000ah1n03x5 output215 (.a(net2527),
    .o(net1932));
 b15bfn000ah1n03x5 output216 (.a(net2499),
    .o(net1901));
 b15bfn000ah1n03x5 output217 (.a(net2531),
    .o(net1934));
 b15bfn000ah1n03x5 output218 (.a(net2513),
    .o(net1905));
 b15bfn000ah1n03x5 output219 (.a(net2491),
    .o(net1893));
 b15bfn000ah1n03x5 output220 (.a(net2489),
    .o(net1891));
 b15bfn000ah1n03x5 output221 (.a(net1966),
    .o(net1967));
 b15bfn000ah1n03x5 output222 (.a(net1968),
    .o(net1969));
 b15bfn000ah1n03x5 output223 (.a(net1972),
    .o(net1973));
 b15bfn000ah1n03x5 output224 (.a(net1974),
    .o(net1975));
 b15bfn000ah1n03x5 output225 (.a(net2495),
    .o(net1897));
 b15bfn000ah1n03x5 output226 (.a(net2493),
    .o(net1895));
 b15bfn000ah1n03x5 output227 (.a(net2497),
    .o(net1899));
 b15bfn000ah1n03x5 output228 (.a(net2511),
    .o(net1903));
 b15bfn000ah1n03x5 output229 (.a(net2535),
    .o(net1945));
 b15bfn000ah1n03x5 output230 (.a(net2509),
    .o(net1915));
 b15bfn000ah1n03x5 output231 (.a(net2519),
    .o(net1926));
 b15bfn000ah1n03x5 output232 (.a(net2523),
    .o(net1928));
 b15bfn000ah1n03x5 output233 (.a(net1979),
    .o(net1980));
 b15bfn000ah1n03x5 output234 (.a(net1987),
    .o(net1988));
 b15bfn000ah1n03x5 output235 (.a(net2507),
    .o(net1913));
 b15bfn000ah1n03x5 output236 (.a(net2525),
    .o(net1930));
 b15bfn000ah1n03x5 output237 (.a(net237),
    .o(tl_o[0]));
 b15bfn000ah1n03x5 output238 (.a(net1993),
    .o(tl_o[10]));
 b15bfn000ah1n03x5 output239 (.a(net1977),
    .o(net1978));
 b15bfn000ah1n03x5 output240 (.a(net1983),
    .o(net1984));
 b15bfn000ah1n03x5 output241 (.a(net241),
    .o(tl_o[13]));
 b15bfn000ah1n03x5 output242 (.a(net242),
    .o(tl_o[14]));
 b15bfn000ah1n03x5 output243 (.a(net243),
    .o(tl_o[15]));
 b15bfn000ah1n03x5 output244 (.a(net2024),
    .o(net2025));
 b15bfn000ah1n03x5 output245 (.a(net2093),
    .o(tl_o[17]));
 b15bfn000ah1n03x5 output246 (.a(net468),
    .o(tl_o[18]));
 b15bfn000ah1n03x5 output247 (.a(net2067),
    .o(tl_o[19]));
 b15bfn000ah1n03x5 output248 (.a(net1986),
    .o(tl_o[1]));
 b15bfn000ah1n03x5 output249 (.a(net464),
    .o(tl_o[20]));
 b15bfn000ah1n03x5 output250 (.a(net2055),
    .o(tl_o[21]));
 b15bfn000ah1n03x5 output251 (.a(net459),
    .o(tl_o[22]));
 b15bfn000ah1n03x5 output252 (.a(net2031),
    .o(tl_o[23]));
 b15bfn000ah1n03x5 output253 (.a(net2143),
    .o(tl_o[24]));
 b15bfn000ah1n03x5 output254 (.a(net2144),
    .o(tl_o[25]));
 b15bfn000ah1n03x5 output255 (.a(net2131),
    .o(tl_o[26]));
 b15bfn000ah1n03x5 output256 (.a(net2029),
    .o(tl_o[27]));
 b15bfn000ah1n03x5 output257 (.a(net2201),
    .o(tl_o[28]));
 b15bfn000ah1n03x5 output258 (.a(net493),
    .o(tl_o[29]));
 b15bfn000ah1n03x5 output259 (.a(net2114),
    .o(tl_o[2]));
 b15bfn000ah1n03x5 output260 (.a(net488),
    .o(tl_o[30]));
 b15bfn000ah1n03x5 output261 (.a(net484),
    .o(tl_o[31]));
 b15bfn000ah1n03x5 output262 (.a(net2146),
    .o(net2147));
 b15bfn000ah1n03x5 output263 (.a(net2018),
    .o(net2019));
 b15bfn000ah1n03x5 output264 (.a(net481),
    .o(tl_o[34]));
 b15bfn000ah1n03x5 output265 (.a(net2009),
    .o(tl_o[35]));
 b15bfn000ah1n03x5 output266 (.a(net2022),
    .o(net2023));
 b15bfn000ah1n03x5 output267 (.a(net1999),
    .o(net2000));
 b15bfn000ah1n03x5 output268 (.a(net2044),
    .o(tl_o[38]));
 b15bfn000ah1n03x5 output269 (.a(net2133),
    .o(tl_o[39]));
 b15bfn000ah1n03x5 output270 (.a(net2160),
    .o(tl_o[3]));
 b15bfn000ah1n03x5 output271 (.a(net2012),
    .o(net2013));
 b15bfn000ah1n03x5 output272 (.a(net2071),
    .o(net2072));
 b15bfn000ah1n03x5 output273 (.a(net2010),
    .o(net2011));
 b15bfn000ah1n03x5 output274 (.a(net2001),
    .o(net2002));
 b15bfn000ah1n03x5 output275 (.a(net2109),
    .o(net2110));
 b15bfn000ah1n03x5 output276 (.a(net2003),
    .o(net2004));
 b15bfn000ah1n03x5 output277 (.a(net2085),
    .o(net2086));
 b15bfn000ah1n03x5 output278 (.a(net2136),
    .o(net2137));
 b15bfn000ah1n03x5 output279 (.a(net1962),
    .o(net1963));
 b15bfn000ah1n03x5 output280 (.a(net2188),
    .o(tl_o[4]));
 b15bfn000ah1n03x5 output281 (.a(net1958),
    .o(net1959));
 b15bfn000ah1n03x5 output282 (.a(net1956),
    .o(net1957));
 b15bfn000ah1n03x5 output283 (.a(net1952),
    .o(net1953));
 b15bfn000ah1n03x5 output284 (.a(net1946),
    .o(net1947));
 b15bfn000ah1n03x5 output285 (.a(net1948),
    .o(net1949));
 b15bfn000ah1n03x5 output286 (.a(net1964),
    .o(net1965));
 b15bfn000ah1n03x5 output287 (.a(net1960),
    .o(net1961));
 b15bfn000ah1n03x5 output288 (.a(net1970),
    .o(net1971));
 b15bfn000ah1n03x5 output289 (.a(net1954),
    .o(net1955));
 b15bfn000ah1n03x5 output290 (.a(net290),
    .o(tl_o[5]));
 b15bfn000ah1n03x5 output291 (.a(net2035),
    .o(tl_o[62]));
 b15bfn000ah1n03x5 output292 (.a(net1919),
    .o(net1920));
 b15bfn000ah1n03x5 output293 (.a(net1982),
    .o(net1951));
 b15bfn000ah1n03x5 output294 (.a(net1997),
    .o(net1998));
 b15bfn000ah1n03x5 output295 (.a(net2219),
    .o(tl_o[6]));
 b15bfn000ah1n03x5 output296 (.a(net2120),
    .o(tl_o[7]));
 b15bfn000ah1n03x5 output297 (.a(net297),
    .o(tl_o[8]));
 b15bfn000ah1n03x5 output298 (.a(net298),
    .o(tl_o[9]));
 b15bfn001as1n24x5 wire299 (.a(N53),
    .o(net299));
 b15bfn001as1n32x5 wire300 (.a(N38),
    .o(net300));
 b15bfn001ah1n24x5 wire301 (.a(N65),
    .o(net301));
 b15bfn001as1n16x5 wire302 (.a(u_reg_u_reg_if_N30),
    .o(net302));
 b15bfn001ah1n24x5 wire303 (.a(N121),
    .o(net303));
 b15bfn001ah1n48x5 load_slew304 (.a(net305),
    .o(net304));
 b15bfn001ah1n48x5 max_length305 (.a(n3812),
    .o(net305));
 b15bfn001as1n24x5 wire306 (.a(n3488),
    .o(net306));
 b15bfn001ah1n64x5 fanout307 (.a(net310),
    .o(net307));
 b15bfn001ah1n48x5 load_slew308 (.a(net307),
    .o(net308));
 b15bfn001as1n64x5 fanout309 (.a(n3494),
    .o(net309));
 b15bfn001ah1n48x5 load_slew310 (.a(net311),
    .o(net310));
 b15bfn000as1n32x5 max_length311 (.a(net309),
    .o(net311));
 b15bfn001ah1n24x5 fanout312 (.a(n3448),
    .o(net312));
 b15bfn001ah1n24x5 fanout313 (.a(n3448),
    .o(net313));
 b15bfn001as1n16x5 wire314 (.a(net2432),
    .o(net314));
 b15bfn001as1n24x5 wire315 (.a(u_reg_u_reg_if_N28),
    .o(net315));
 b15bfn001as1n16x5 wire316 (.a(u_reg_u_reg_if_N17),
    .o(net316));
 b15bfn001as1n16x5 wire317 (.a(net2141),
    .o(net317));
 b15bfn001as1n24x5 wire318 (.a(n4188),
    .o(net318));
 b15bfn001as1n16x5 fanout319 (.a(n4187),
    .o(net319));
 b15bfn001ah1n24x5 fanout320 (.a(n4187),
    .o(net320));
 b15bfn001ah1n24x5 wire321 (.a(net322),
    .o(net321));
 b15bfn001as1n32x5 wire322 (.a(n4186),
    .o(net322));
 b15bfn001ah1n32x5 wire323 (.a(net324),
    .o(net323));
 b15bfn001as1n32x5 max_length324 (.a(n3861),
    .o(net324));
 b15bfn001as1n24x5 wire325 (.a(n3715),
    .o(net325));
 b15bfn001as1n48x5 fanout326 (.a(n3754),
    .o(net326));
 b15bfn001ah1n24x5 max_length327 (.a(net326),
    .o(net327));
 b15bfn001ah1n48x5 max_length328 (.a(net326),
    .o(net328));
 b15bfn001as1n24x5 wire329 (.a(n3754),
    .o(net329));
 b15bfn001ah1n32x5 max_length330 (.a(net331),
    .o(net330));
 b15bfn001as1n32x5 max_length331 (.a(n4181),
    .o(net331));
 b15bfn001ah1n32x5 wire332 (.a(net333),
    .o(net332));
 b15bfn001as1n24x5 max_length333 (.a(n3859),
    .o(net333));
 b15bfn001ah1n24x5 fanout334 (.a(net335),
    .o(net334));
 b15bfn001as1n32x5 fanout335 (.a(n3513),
    .o(net335));
 b15bfn001ah1n48x5 fanout336 (.a(n3343),
    .o(net336));
 b15bfn001ah1n16x5 fanout337 (.a(n3343),
    .o(net337));
 b15bfn001ah1n32x5 fanout338 (.a(net339),
    .o(net338));
 b15bfn001ah1n32x5 fanout339 (.a(n3344),
    .o(net339));
 b15bfn001as1n48x5 wire340 (.a(net341),
    .o(net340));
 b15bfn001ah1n32x5 max_length341 (.a(N113),
    .o(net341));
 b15bfn001as1n24x5 wire342 (.a(N113),
    .o(net342));
 b15bfn001as1n24x5 wire343 (.a(N113),
    .o(net343));
 b15bfn001ah1n24x5 fanout344 (.a(net345),
    .o(net344));
 b15bfn001as1n24x5 fanout345 (.a(n3307),
    .o(net345));
 b15bfn001as1n32x5 wire346 (.a(net345),
    .o(net346));
 b15bfn001as1n32x5 fanout347 (.a(n3305),
    .o(net347));
 b15bfn001as1n24x5 fanout348 (.a(n3305),
    .o(net348));
 b15bfn001ah1n64x5 fanout349 (.a(net350),
    .o(net349));
 b15bfn001as1n32x5 fanout350 (.a(n4179),
    .o(net350));
 b15bfn000as1n32x5 wire351 (.a(net350),
    .o(net351));
 b15bfn001as1n48x5 fanout352 (.a(n4178),
    .o(net352));
 b15bfn001ah1n32x5 wire353 (.a(net354),
    .o(net353));
 b15bfn001as1n32x5 wire354 (.a(net352),
    .o(net354));
 b15bfn001as1n24x5 max_length355 (.a(net356),
    .o(net355));
 b15bfn001as1n32x5 max_length356 (.a(net357),
    .o(net356));
 b15bfn001as1n32x5 load_slew357 (.a(n4024),
    .o(net357));
 b15bfn001ah1n48x5 load_slew358 (.a(net359),
    .o(net358));
 b15bfn001ah1n32x5 max_length359 (.a(n3821),
    .o(net359));
 b15bfn001as1n16x5 wire360 (.a(gen_filter_14__u_filter_diff_ctr_d[2]),
    .o(net360));
 b15bfn001ah1n24x5 wire361 (.a(n3947),
    .o(net361));
 b15bfn001ah1n24x5 wire362 (.a(n3869),
    .o(net362));
 b15bfn001ah1n24x5 wire363 (.a(n3009),
    .o(net363));
 b15bfn001as1n24x5 wire364 (.a(u_reg_u_data_in_wr_data[7]),
    .o(net364));
 b15bfn001as1n24x5 wire365 (.a(u_reg_u_data_in_wr_data[0]),
    .o(net365));
 b15bfn001ah1n48x5 max_length366 (.a(n3886),
    .o(net366));
 b15bfn001ah1n48x5 max_length367 (.a(n3886),
    .o(net367));
 b15bfn001as1n80x5 fanout368 (.a(net369),
    .o(net368));
 b15bfn001as1n64x5 fanout369 (.a(n3318),
    .o(net369));
 b15bfn001ah1n48x5 max_length370 (.a(net371),
    .o(net370));
 b15bfn001as1n48x5 wire371 (.a(net369),
    .o(net371));
 b15bfn001as1n32x5 max_length372 (.a(net369),
    .o(net372));
 b15bfn001as1n64x5 fanout373 (.a(net381),
    .o(net373));
 b15bfn001as1n24x5 wire374 (.a(net375),
    .o(net374));
 b15bfn001as1n24x5 max_length375 (.a(net376),
    .o(net375));
 b15bfn001as1n32x5 max_length376 (.a(net373),
    .o(net376));
 b15bfn001as1n64x5 fanout377 (.a(n3316),
    .o(net377));
 b15bfn001ah1n32x5 wire378 (.a(net380),
    .o(net378));
 b15bfn001ah1n48x5 wire379 (.a(net380),
    .o(net379));
 b15bfn001ah1n48x5 wire380 (.a(net377),
    .o(net380));
 b15bfn001ah1n32x5 max_length381 (.a(net377),
    .o(net381));
 b15bfn001as1n32x5 fanout382 (.a(net385),
    .o(net382));
 b15bfn001as1n32x5 wire383 (.a(net384),
    .o(net383));
 b15bfn001ah1n48x5 wire384 (.a(net382),
    .o(net384));
 b15bfn001as1n64x5 fanout385 (.a(n3314),
    .o(net385));
 b15bfn001ah1n48x5 wire386 (.a(net385),
    .o(net386));
 b15bfn001ah1n24x5 max_length387 (.a(net388),
    .o(net387));
 b15bfn001as1n24x5 max_length388 (.a(net385),
    .o(net388));
 b15bfn001ah1n24x5 wire389 (.a(n3314),
    .o(net389));
 b15bfn001as1n64x5 fanout390 (.a(n3909),
    .o(net390));
 b15bfn001ah1n32x5 max_length391 (.a(net393),
    .o(net391));
 b15bfn001ah1n48x5 load_slew392 (.a(net394),
    .o(net392));
 b15bfn001as1n32x5 max_length393 (.a(net394),
    .o(net393));
 b15bfn001ah1n48x5 max_length394 (.a(net390),
    .o(net394));
 b15bfn001as1n48x5 fanout395 (.a(net399),
    .o(net395));
 b15bfn001as1n32x5 wire396 (.a(net397),
    .o(net396));
 b15bfn001ah1n24x5 max_length397 (.a(net395),
    .o(net397));
 b15bfn000as1n32x5 fanout398 (.a(net399),
    .o(net398));
 b15bfn001as1n80x5 fanout399 (.a(n3304),
    .o(net399));
 b15bfn001as1n16x5 wire400 (.a(n3051),
    .o(net400));
 b15bfn001ah1n32x5 wire401 (.a(n3032),
    .o(net401));
 b15bfn001ah1n32x5 wire402 (.a(n3065),
    .o(net402));
 b15bfn001ah1n24x5 wire403 (.a(n3063),
    .o(net403));
 b15bfn001ah1n24x5 wire404 (.a(n3054),
    .o(net404));
 b15bfn001as1n48x5 fanout405 (.a(n4175),
    .o(net405));
 b15bfn001as1n32x5 wire406 (.a(net408),
    .o(net406));
 b15bfn001as1n48x5 max_length407 (.a(net405),
    .o(net407));
 b15bfn001as1n48x5 max_length408 (.a(net405),
    .o(net408));
 b15bfn001as1n24x5 wire409 (.a(net405),
    .o(net409));
 b15bfn001as1n48x5 wire410 (.a(net411),
    .o(net410));
 b15bfn001as1n32x5 max_length411 (.a(n4175),
    .o(net411));
 b15bfn001ah1n48x5 wire412 (.a(net413),
    .o(net412));
 b15bfn001ah1n48x5 wire413 (.a(net414),
    .o(net413));
 b15bfn001ah1n48x5 max_length414 (.a(n4026),
    .o(net414));
 b15bfn001ah1n24x5 wire415 (.a(n3934),
    .o(net415));
 b15bfn001as1n32x5 wire416 (.a(n3935),
    .o(net416));
 b15bfn001as1n64x5 fanout417 (.a(net421),
    .o(net417));
 b15bfn001ah1n32x5 max_length418 (.a(net419),
    .o(net418));
 b15bfn001ah1n32x5 max_length419 (.a(net420),
    .o(net419));
 b15bfn001as1n32x5 max_length420 (.a(net417),
    .o(net420));
 b15bfn001as1n64x5 fanout421 (.a(n3413),
    .o(net421));
 b15bfn001ah1n48x5 max_length422 (.a(net424),
    .o(net422));
 b15bfn001as1n32x5 max_length423 (.a(net424),
    .o(net423));
 b15bfn001as1n32x5 max_length424 (.a(net421),
    .o(net424));
 b15bfn001as1n64x5 fanout425 (.a(n3915),
    .o(net425));
 b15bfn000ah1n48x5 wire426 (.a(net427),
    .o(net426));
 b15bfn001ah1n64x5 wire427 (.a(net428),
    .o(net427));
 b15bfn001ah1n48x5 load_slew428 (.a(net425),
    .o(net428));
 b15bfn001as1n64x5 fanout429 (.a(n3908),
    .o(net429));
 b15bfn001as1n48x5 wire430 (.a(net431),
    .o(net430));
 b15bfn001as1n32x5 wire431 (.a(net432),
    .o(net431));
 b15bfn001as1n32x5 max_length432 (.a(net429),
    .o(net432));
 b15bfn001as1n80x5 fanout433 (.a(net436),
    .o(net433));
 b15bfn001as1n64x5 fanout434 (.a(n3309),
    .o(net434));
 b15bfn000ah1n48x5 wire435 (.a(net436),
    .o(net435));
 b15bfn001ah1n48x5 max_length436 (.a(net434),
    .o(net436));
 b15bfn001as1n80x5 fanout437 (.a(net438),
    .o(net437));
 b15bfn001as1n64x5 fanout438 (.a(net441),
    .o(net438));
 b15bfn001as1n32x5 wire439 (.a(net440),
    .o(net439));
 b15bfn001ah1n48x5 wire440 (.a(net438),
    .o(net440));
 b15bfn001ah1n32x5 wire441 (.a(n3415),
    .o(net441));
 b15bfn001as1n48x5 fanout442 (.a(net445),
    .o(net442));
 b15bfn001as1n32x5 max_length443 (.a(net444),
    .o(net443));
 b15bfn001ah1n48x5 max_length444 (.a(net442),
    .o(net444));
 b15bfn001as1n64x5 fanout445 (.a(n3306),
    .o(net445));
 b15bfn001ah1n32x5 wire446 (.a(net445),
    .o(net446));
 b15bfn001ah1n32x5 wire447 (.a(net448),
    .o(net447));
 b15bfn001ah1n32x5 wire448 (.a(net445),
    .o(net448));
 b15bfn000as1n24x5 wire449 (.a(n3306),
    .o(net449));
 b15bfn001ah1n24x5 wire450 (.a(n3042),
    .o(net450));
 b15bfn001as1n32x5 wire451 (.a(n3029),
    .o(net451));
 b15bfn001ah1n24x5 wire452 (.a(n3026),
    .o(net452));
 b15bfn001ah1n24x5 wire453 (.a(n3050),
    .o(net453));
 b15bfn001as1n24x5 wire454 (.a(n2992),
    .o(net454));
 b15bfn001ah1n12x5 wire455 (.a(net2142),
    .o(net455));
 b15bfn001ah1n12x5 load_slew456 (.a(net457),
    .o(net456));
 b15bfn001ah1n12x5 wire457 (.a(net2030),
    .o(net457));
 b15bfn001as1n16x5 wire458 (.a(net251),
    .o(net458));
 b15bfn001as1n12x5 wire459 (.a(net2175),
    .o(net459));
 b15bfn001ah1n16x5 wire460 (.a(net2054),
    .o(net460));
 b15bfn001as1n12x5 max_cap461 (.a(net462),
    .o(net461));
 b15bfn001ah1n24x5 wire462 (.a(net463),
    .o(net462));
 b15bfn001ah1n12x5 load_slew463 (.a(net2054),
    .o(net463));
 b15bfn001ah1n12x5 load_slew464 (.a(net2033),
    .o(net464));
 b15bfn001as1n08x5 wire465 (.a(net2032),
    .o(net465));
 b15bfn001ah1n12x5 wire466 (.a(net2066),
    .o(net466));
 b15bfn001as1n12x5 max_cap467 (.a(net246),
    .o(net467));
 b15bfn001ah1n16x5 max_cap468 (.a(net2124),
    .o(net468));
 b15bfn001ah1n12x5 wire469 (.a(net2003),
    .o(net469));
 b15bfn001as1n12x5 wire470 (.a(net471),
    .o(net470));
 b15bfn001ah1n06x5 load_slew471 (.a(net2001),
    .o(net471));
 b15bfn000as1n24x5 wire472 (.a(net473),
    .o(net472));
 b15bfn001ah1n12x5 wire473 (.a(net273),
    .o(net473));
 b15bfn001as1n08x5 wire474 (.a(net2010),
    .o(net474));
 b15bfn001ah1n12x5 wire475 (.a(net2043),
    .o(net475));
 b15bfn001ah1n12x5 wire476 (.a(net477),
    .o(net476));
 b15bfn001ah1n12x5 load_slew477 (.a(net478),
    .o(net477));
 b15bfn001ah1n12x5 wire478 (.a(net1999),
    .o(net478));
 b15bfn001ah1n16x5 wire479 (.a(net2008),
    .o(net479));
 b15bfn001ah1n16x5 wire480 (.a(net2052),
    .o(net480));
 b15bfn001ah1n12x5 wire481 (.a(net2053),
    .o(net481));
 b15bfn001as1n12x5 wire482 (.a(net2052),
    .o(net482));
 b15bfn001as1n16x5 wire483 (.a(net261),
    .o(net483));
 b15bfn001as1n12x5 max_cap484 (.a(net485),
    .o(net484));
 b15bfn001ah1n12x5 load_slew485 (.a(net486),
    .o(net485));
 b15bfn001ah1n12x5 wire486 (.a(net2211),
    .o(net486));
 b15bfn001ah1n24x5 wire487 (.a(net490),
    .o(net487));
 b15bfn001ah1n08x5 load_slew488 (.a(net2049),
    .o(net488));
 b15bfn001ah1n12x5 wire489 (.a(net2048),
    .o(net489));
 b15bfn001ah1n08x5 load_slew490 (.a(net2048),
    .o(net490));
 b15bfn001as1n24x5 wire491 (.a(net492),
    .o(net491));
 b15bfn001ah1n12x5 wire492 (.a(net258),
    .o(net492));
 b15bfn001as1n12x5 load_slew493 (.a(net2091),
    .o(net493));
 b15bfn001as1n12x5 wire494 (.a(net2090),
    .o(net494));
 b15bfn001ah1n24x5 wire495 (.a(net2200),
    .o(net495));
 b15bfn001as1n12x5 wire496 (.a(net2028),
    .o(net496));
 b15bfn001as1n08x5 load_slew497 (.a(net498),
    .o(net497));
 b15bfn001ah1n16x5 wire498 (.a(net2028),
    .o(net498));
 b15bfn000ah1n12x5 wire499 (.a(net2130),
    .o(net499));
 b15bfn001as1n12x5 max_cap500 (.a(net2130),
    .o(net500));
 b15bfn001as1n12x5 max_cap501 (.a(net2092),
    .o(net501));
 b15bfn001ah1n24x5 wire502 (.a(net503),
    .o(net502));
 b15bfn001ah1n12x5 wire503 (.a(net504),
    .o(net503));
 b15bfn001ah1n08x5 load_slew504 (.a(net2024),
    .o(net504));
 b15bfn001as1n12x5 wire505 (.a(reg2hw_intr_state__q__6_),
    .o(net505));
 b15bfn001as1n12x5 wire506 (.a(net507),
    .o(net506));
 b15bfn001ah1n16x5 wire507 (.a(reg2hw_intr_state__q__5_),
    .o(net507));
 b15bfn000as1n12x5 wire508 (.a(net2236),
    .o(net508));
 b15bfn001ah1n12x5 wire509 (.a(reg2hw_intr_state__q__3_),
    .o(net509));
 b15bfn001as1n12x5 wire510 (.a(reg2hw_intr_state__q__29_),
    .o(net510));
 b15bfn001as1n08x5 wire511 (.a(reg2hw_intr_state__q__15_),
    .o(net511));
 b15bfn001as1n12x5 wire512 (.a(reg2hw_intr_state__q__13_),
    .o(net512));
 b15bfn001ah1n12x5 wire513 (.a(reg2hw_intr_state__q__12_),
    .o(net513));
 b15bfn001ah1n24x5 wire514 (.a(net515),
    .o(net514));
 b15bfn001as1n16x5 wire515 (.a(reg2hw_intr_state__q__11_),
    .o(net515));
 b15bfn001as1n16x5 wire516 (.a(reg2hw_intr_state__q__10_),
    .o(net516));
 b15bfn001ah1n12x5 wire517 (.a(reg2hw_intr_state__q__1_),
    .o(net517));
 b15bfn001ah1n16x5 wire518 (.a(reg2hw_intr_enable__q__5_),
    .o(net518));
 b15bfn001ah1n16x5 wire519 (.a(net2227),
    .o(net519));
 b15bfn001as1n16x5 wire520 (.a(reg2hw_intr_enable__q__25_),
    .o(net520));
 b15bfn001as1n16x5 wire521 (.a(net2220),
    .o(net521));
 b15bfn001ah1n12x5 wire522 (.a(reg2hw_intr_enable__q__16_),
    .o(net522));
 b15bfn001as1n16x5 wire523 (.a(reg2hw_intr_enable__q__13_),
    .o(net523));
 b15bfn001as1n16x5 wire524 (.a(reg2hw_intr_enable__q__12_),
    .o(net524));
 b15bfn001ah1n16x5 wire525 (.a(reg2hw_intr_ctrl_en_rising__q__27_),
    .o(net525));
 b15bfn001ah1n12x5 wire526 (.a(reg2hw_intr_ctrl_en_rising__q__14_),
    .o(net526));
 b15bfn001ah1n12x5 wire527 (.a(net528),
    .o(net527));
 b15bfn000ah1n12x5 wire528 (.a(reg2hw_intr_ctrl_en_rising__q__13_),
    .o(net528));
 b15bfn001ah1n16x5 wire529 (.a(reg2hw_intr_ctrl_en_rising__q__1_),
    .o(net529));
 b15bfn001as1n24x5 wire530 (.a(net531),
    .o(net530));
 b15bfn001as1n12x5 wire531 (.a(reg2hw_intr_ctrl_en_lvllow__q__7_),
    .o(net531));
 b15bfn001as1n16x5 wire532 (.a(net533),
    .o(net532));
 b15bfn001ah1n12x5 wire533 (.a(reg2hw_intr_ctrl_en_lvllow__q__6_),
    .o(net533));
 b15bfn001as1n12x5 wire534 (.a(reg2hw_intr_ctrl_en_lvllow__q__25_),
    .o(net534));
 b15bfn001ah1n24x5 wire535 (.a(reg2hw_intr_ctrl_en_lvllow__q__15_),
    .o(net535));
 b15bfn001ah1n12x5 wire536 (.a(reg2hw_intr_ctrl_en_lvllow__q__15_),
    .o(net536));
 b15bfn001as1n16x5 wire537 (.a(reg2hw_intr_ctrl_en_lvllow__q__14_),
    .o(net537));
 b15bfn001ah1n16x5 wire538 (.a(net2350),
    .o(net538));
 b15bfn001as1n12x5 wire539 (.a(reg2hw_intr_ctrl_en_lvllow__q__10_),
    .o(net539));
 b15bfn001ah1n12x5 wire540 (.a(reg2hw_intr_ctrl_en_lvllow__q__0_),
    .o(net540));
 b15bfn001ah1n16x5 wire541 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__7_),
    .o(net541));
 b15bfn001as1n16x5 wire542 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__6_),
    .o(net542));
 b15bfn001as1n16x5 wire543 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__5_),
    .o(net543));
 b15bfn000ah1n24x5 wire544 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__4_),
    .o(net544));
 b15bfn001ah1n12x5 wire545 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__31_),
    .o(net545));
 b15bfn001ah1n16x5 wire546 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__21_),
    .o(net546));
 b15bfn001ah1n16x5 wire547 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__16_),
    .o(net547));
 b15bfn001ah1n12x5 wire548 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__13_),
    .o(net548));
 b15bfn001ah1n16x5 wire549 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__11_),
    .o(net549));
 b15bfn001ah1n16x5 wire550 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__10_),
    .o(net550));
 b15bfn001ah1n16x5 wire551 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__0_),
    .o(net551));
 b15bfn001as1n12x5 wire552 (.a(reg2hw_intr_ctrl_en_falling__q__4_),
    .o(net552));
 b15bfn001ah1n16x5 wire553 (.a(reg2hw_intr_ctrl_en_falling__q__3_),
    .o(net553));
 b15bfn001ah1n16x5 wire554 (.a(reg2hw_intr_ctrl_en_falling__q__2_),
    .o(net554));
 b15bfn001ah1n16x5 wire555 (.a(reg2hw_intr_ctrl_en_falling__q__27_),
    .o(net555));
 b15bfn001ah1n16x5 wire556 (.a(reg2hw_intr_ctrl_en_falling__q__18_),
    .o(net556));
 b15bfn001ah1n16x5 wire557 (.a(reg2hw_intr_ctrl_en_falling__q__15_),
    .o(net557));
 b15bfn001as1n16x5 wire558 (.a(reg2hw_intr_ctrl_en_falling__q__13_),
    .o(net558));
 b15bfn001ah1n16x5 wire559 (.a(reg2hw_intr_ctrl_en_falling__q__12_),
    .o(net559));
 b15bfn001as1n08x5 wire560 (.a(net561),
    .o(net560));
 b15bfn001as1n12x5 wire561 (.a(reg2hw_intr_ctrl_en_falling__q__1_),
    .o(net561));
 b15bfn001ah1n16x5 wire562 (.a(reg2hw_intr_ctrl_en_falling__q__0_),
    .o(net562));
 b15bfn001ah1n16x5 wire563 (.a(net564),
    .o(net563));
 b15bfn001ah1n16x5 wire564 (.a(reg2hw_ctrl_en_input_filter__q__8_),
    .o(net564));
 b15bfn001ah1n16x5 wire565 (.a(reg2hw_ctrl_en_input_filter__q__7_),
    .o(net565));
 b15bfn001as1n16x5 wire566 (.a(reg2hw_ctrl_en_input_filter__q__7_),
    .o(net566));
 b15bfn001ah1n24x5 wire567 (.a(reg2hw_ctrl_en_input_filter__q__6_),
    .o(net567));
 b15bfn001ah1n12x5 load_slew568 (.a(net569),
    .o(net568));
 b15bfn001ah1n12x5 wire569 (.a(reg2hw_ctrl_en_input_filter__q__5_),
    .o(net569));
 b15bfn001ah1n24x5 wire570 (.a(net571),
    .o(net570));
 b15bfn001ah1n16x5 max_cap571 (.a(reg2hw_ctrl_en_input_filter__q__4_),
    .o(net571));
 b15bfn001ah1n16x5 max_cap572 (.a(reg2hw_ctrl_en_input_filter__q__4_),
    .o(net572));
 b15bfn001ah1n12x5 wire573 (.a(reg2hw_ctrl_en_input_filter__q__31_),
    .o(net573));
 b15bfn001as1n12x5 max_cap574 (.a(net575),
    .o(net574));
 b15bfn001as1n16x5 wire575 (.a(reg2hw_ctrl_en_input_filter__q__30_),
    .o(net575));
 b15bfn001as1n08x5 wire576 (.a(reg2hw_ctrl_en_input_filter__q__3_),
    .o(net576));
 b15bfn001ah1n12x5 wire577 (.a(reg2hw_ctrl_en_input_filter__q__3_),
    .o(net577));
 b15bfn001ah1n24x5 wire578 (.a(reg2hw_ctrl_en_input_filter__q__29_),
    .o(net578));
 b15bfn001as1n16x5 wire579 (.a(reg2hw_ctrl_en_input_filter__q__28_),
    .o(net579));
 b15bfn001ah1n12x5 load_slew580 (.a(net581),
    .o(net580));
 b15bfn001ah1n08x5 load_slew581 (.a(reg2hw_ctrl_en_input_filter__q__26_),
    .o(net581));
 b15bfn001as1n16x5 wire582 (.a(net583),
    .o(net582));
 b15bfn001as1n06x5 load_slew583 (.a(reg2hw_ctrl_en_input_filter__q__24_),
    .o(net583));
 b15bfn001ah1n24x5 wire584 (.a(reg2hw_ctrl_en_input_filter__q__23_),
    .o(net584));
 b15bfn001as1n12x5 wire585 (.a(net586),
    .o(net585));
 b15bfn001as1n12x5 wire586 (.a(reg2hw_ctrl_en_input_filter__q__22_),
    .o(net586));
 b15bfn001ah1n16x5 wire587 (.a(reg2hw_ctrl_en_input_filter__q__21_),
    .o(net587));
 b15bfn001as1n24x5 wire588 (.a(net589),
    .o(net588));
 b15bfn001as1n12x5 wire589 (.a(reg2hw_ctrl_en_input_filter__q__19_),
    .o(net589));
 b15bfn001as1n24x5 wire590 (.a(net591),
    .o(net590));
 b15bfn001ah1n16x5 wire591 (.a(reg2hw_ctrl_en_input_filter__q__18_),
    .o(net591));
 b15bfn001as1n24x5 wire592 (.a(net593),
    .o(net592));
 b15bfn001as1n12x5 wire593 (.a(reg2hw_ctrl_en_input_filter__q__17_),
    .o(net593));
 b15bfn001as1n24x5 wire594 (.a(net595),
    .o(net594));
 b15bfn001as1n12x5 wire595 (.a(reg2hw_ctrl_en_input_filter__q__16_),
    .o(net595));
 b15bfn001as1n08x5 load_slew596 (.a(net597),
    .o(net596));
 b15bfn001as1n16x5 wire597 (.a(reg2hw_ctrl_en_input_filter__q__15_),
    .o(net597));
 b15bfn001ah1n12x5 load_slew598 (.a(net599),
    .o(net598));
 b15bfn001as1n12x5 wire599 (.a(reg2hw_ctrl_en_input_filter__q__14_),
    .o(net599));
 b15bfn001ah1n12x5 wire600 (.a(net601),
    .o(net600));
 b15bfn000as1n24x5 wire601 (.a(net602),
    .o(net601));
 b15bfn001ah1n12x5 wire602 (.a(reg2hw_ctrl_en_input_filter__q__13_),
    .o(net602));
 b15bfn001ah1n12x5 load_slew603 (.a(net604),
    .o(net603));
 b15bfn001ah1n24x5 wire604 (.a(net605),
    .o(net604));
 b15bfn001as1n08x5 wire605 (.a(reg2hw_ctrl_en_input_filter__q__12_),
    .o(net605));
 b15bfn001ah1n24x5 wire606 (.a(net607),
    .o(net606));
 b15bfn001ah1n12x5 load_slew607 (.a(reg2hw_ctrl_en_input_filter__q__11_),
    .o(net607));
 b15bfn001as1n12x5 max_cap608 (.a(reg2hw_ctrl_en_input_filter__q__10_),
    .o(net608));
 b15bfn001ah1n12x5 load_slew609 (.a(reg2hw_ctrl_en_input_filter__q__1_),
    .o(net609));
 b15bfn001as1n08x5 load_slew610 (.a(reg2hw_ctrl_en_input_filter__q__1_),
    .o(net610));
 b15bfn001ah1n12x5 wire611 (.a(reg2hw_ctrl_en_input_filter__q__0_),
    .o(net611));
 b15bfn001ah1n08x5 load_slew612 (.a(net2108),
    .o(net612));
 b15bfn001ah1n12x5 wire613 (.a(net2107),
    .o(net613));
 b15bfn001as1n16x5 wire614 (.a(net2115),
    .o(net614));
 b15bfn001ah1n12x5 wire615 (.a(net2245),
    .o(net615));
 b15bfn001ah1n16x5 max_cap616 (.a(net194),
    .o(net616));
 b15bfn001ah1n12x5 wire617 (.a(net193),
    .o(net617));
 b15bfn001as1n12x5 wire618 (.a(net192),
    .o(net618));
 b15bfn001ah1n12x5 load_slew619 (.a(net620),
    .o(net619));
 b15bfn001ah1n12x5 load_slew620 (.a(net191),
    .o(net620));
 b15bfn001as1n08x5 load_slew621 (.a(net190),
    .o(net621));
 b15bfn001as1n12x5 max_cap622 (.a(net2458),
    .o(net622));
 b15bfn001ah1n12x5 wire623 (.a(net2399),
    .o(net623));
 b15bfn001ah1n12x5 wire624 (.a(net188),
    .o(net624));
 b15bfn001as1n24x5 wire625 (.a(net626),
    .o(net625));
 b15bfn001as1n12x5 wire626 (.a(net2419),
    .o(net626));
 b15bfn001ah1n16x5 wire627 (.a(net2459),
    .o(net627));
 b15bfn001as1n16x5 wire628 (.a(net185),
    .o(net628));
 b15bfn001ah1n12x5 wire629 (.a(net630),
    .o(net629));
 b15bfn001ah1n24x5 wire630 (.a(net631),
    .o(net630));
 b15bfn001as1n08x5 wire631 (.a(net183),
    .o(net631));
 b15bfn001as1n12x5 wire632 (.a(net182),
    .o(net632));
 b15bfn000as1n32x5 wire633 (.a(net634),
    .o(net633));
 b15bfn001as1n16x5 wire634 (.a(net2251),
    .o(net634));
 b15bfn001ah1n12x5 load_slew635 (.a(net2151),
    .o(net635));
 b15bfn001as1n16x5 wire636 (.a(net2150),
    .o(net636));
 b15bfn001as1n16x5 wire637 (.a(net2184),
    .o(net637));
 b15bfn001ah1n16x5 wire638 (.a(net2068),
    .o(net638));
 b15bfn001as1n08x5 load_slew639 (.a(net170),
    .o(net639));
 b15bfn001ah1n12x5 load_slew640 (.a(net169),
    .o(net640));
 b15bfn001ah1n16x5 max_cap641 (.a(net168),
    .o(net641));
 b15bfn001ah1n16x5 max_cap642 (.a(net167),
    .o(net642));
 b15bfn001ah1n12x5 wire643 (.a(net165),
    .o(net643));
 b15bfn001as1n12x5 max_cap644 (.a(net162),
    .o(net644));
 b15bfn001as1n12x5 max_cap645 (.a(net161),
    .o(net645));
 b15bfn001as1n12x5 wire646 (.a(net2098),
    .o(net646));
 b15bfn001as1n16x5 wire647 (.a(net2174),
    .o(net647));
 b15bfn001as1n12x5 wire648 (.a(net2106),
    .o(net648));
 b15bfn001as1n12x5 max_cap649 (.a(net2080),
    .o(net649));
 b15bfn001as1n08x5 load_slew650 (.a(net2079),
    .o(net650));
 b15bfn001ah1n12x5 wire651 (.a(net156),
    .o(net651));
 b15bfn001ah1n12x5 wire652 (.a(net2050),
    .o(net652));
 b15bfn001as1n08x5 wire653 (.a(net2129),
    .o(net653));
 b15bfn001as1n12x5 wire654 (.a(net2128),
    .o(net654));
 b15bfn001ah1n12x5 load_slew655 (.a(net2083),
    .o(net655));
 b15bfn001as1n16x5 wire656 (.a(net2095),
    .o(net656));
 b15bfn001as1n12x5 wire657 (.a(net2094),
    .o(net657));
 b15bfn001as1n12x5 max_cap658 (.a(net150),
    .o(net658));
 b15bfn001as1n12x5 max_cap659 (.a(net2132),
    .o(net659));
 b15bfn001ah1n12x5 wire660 (.a(net144),
    .o(net660));
 b15bfn001ah1n12x5 load_slew661 (.a(net143),
    .o(net661));
 b15bfn001ah1n16x5 max_cap662 (.a(net142),
    .o(net662));
 b15bfn001ah1n12x5 load_slew663 (.a(net664),
    .o(net663));
 b15bfn001ah1n12x5 wire664 (.a(net2267),
    .o(net664));
 b15bfn001ah1n12x5 wire665 (.a(net666),
    .o(net665));
 b15bfn001as1n12x5 wire666 (.a(net2217),
    .o(net666));
 b15bfn001as1n32x5 wire667 (.a(n3732),
    .o(net667));
 b15bfn001ah1n24x5 wire668 (.a(n3716),
    .o(net668));
 b15bfn001as1n32x5 wire669 (.a(n3701),
    .o(net669));
 b15bfn001as1n32x5 wire670 (.a(n3822),
    .o(net670));
 b15bfn001ah1n24x5 max_length671 (.a(net672),
    .o(net671));
 b15bfn001as1n24x5 wire672 (.a(u_reg_u_reg_if_a_ack),
    .o(net672));
 b15bfn001as1n16x5 wire673 (.a(u_reg_data_in_qs[30]),
    .o(net673));
 b15bfn001ah1n24x5 wire674 (.a(net675),
    .o(net674));
 b15bfn001as1n08x5 wire675 (.a(net1919),
    .o(net675));
 b15bfn001ah1n12x5 wire676 (.a(net1918),
    .o(net676));
 b15bfn001ah1n16x5 wire677 (.a(net2138),
    .o(net677));
 b15bfn001ah1n16x5 wire678 (.a(net2274),
    .o(net678));
 b15bfn001ah1n16x5 wire679 (.a(net2208),
    .o(net679));
 b15bfn001ah1n16x5 wire680 (.a(net681),
    .o(net680));
 b15bfn001as1n16x5 wire681 (.a(net2409),
    .o(net681));
 b15bfn001as1n12x5 wire682 (.a(gen_filter_3__u_filter_filter_synced),
    .o(net682));
 b15bfn001as1n08x5 wire683 (.a(net684),
    .o(net683));
 b15bfn001ah1n24x5 wire684 (.a(gen_filter_26__u_filter_filter_synced),
    .o(net684));
 b15bfn001ah1n16x5 wire685 (.a(net2291),
    .o(net685));
 b15bfn001as1n16x5 wire686 (.a(gen_filter_19__u_filter_filter_synced),
    .o(net686));
 b15bfn001ah1n24x5 wire687 (.a(gen_filter_14__u_filter_diff_ctr_q[2]),
    .o(net687));
 b15bfn001as1n32x5 max_length688 (.a(net689),
    .o(net688));
 b15bfn001ah1n48x5 max_length689 (.a(n3814),
    .o(net689));
 b15bfn001ah1n24x5 wire690 (.a(net692),
    .o(net690));
 b15bfn001as1n48x5 max_length691 (.a(n4143),
    .o(net691));
 b15bfn001ah1n48x5 max_length692 (.a(n4143),
    .o(net692));
 b15bfn001ah1n32x5 wire693 (.a(n4140),
    .o(net693));
 b15bfn001as1n64x5 fanout694 (.a(n4139),
    .o(net694));
 b15bfn001as1n32x5 wire695 (.a(net696),
    .o(net695));
 b15bfn001as1n32x5 max_length696 (.a(net697),
    .o(net696));
 b15bfn001ah1n32x5 max_length697 (.a(net694),
    .o(net697));
 b15bfn001ah1n24x5 max_length698 (.a(net699),
    .o(net698));
 b15bfn001as1n24x5 wire699 (.a(n4134),
    .o(net699));
 b15bfn001as1n16x5 max_length700 (.a(net701),
    .o(net700));
 b15bfn001as1n32x5 max_length701 (.a(n4129),
    .o(net701));
 b15bfn001ah1n24x5 max_length702 (.a(net703),
    .o(net702));
 b15bfn001as1n24x5 max_length703 (.a(n4128),
    .o(net703));
 b15bfn001as1n24x5 wire704 (.a(n4117),
    .o(net704));
 b15bfn001as1n24x5 wire705 (.a(net706),
    .o(net705));
 b15bfn001as1n24x5 wire706 (.a(n4116),
    .o(net706));
 b15bfn001as1n48x5 fanout707 (.a(net710),
    .o(net707));
 b15bfn001as1n48x5 load_slew708 (.a(net709),
    .o(net708));
 b15bfn001as1n48x5 wire709 (.a(net707),
    .o(net709));
 b15bfn001ah1n32x5 wire710 (.a(net97),
    .o(net710));
 b15bfn001as1n32x5 wire711 (.a(net86),
    .o(net711));
 b15bfn001ah1n48x5 wire712 (.a(net81),
    .o(net712));
 b15bfn001ah1n48x5 max_length713 (.a(net78),
    .o(net713));
 b15bfn001ah1n48x5 wire714 (.a(net76),
    .o(net714));
 b15bfn001as1n48x5 wire715 (.a(net74),
    .o(net715));
 b15bfn001ah1n32x5 wire716 (.a(net73),
    .o(net716));
 b15bfn001ah1n48x5 wire717 (.a(net71),
    .o(net717));
 b15bfn000as1n32x5 wire718 (.a(net70),
    .o(net718));
 b15bfn001as1n32x5 wire719 (.a(net64),
    .o(net719));
 b15bfn001ah1n48x5 wire720 (.a(net60),
    .o(net720));
 b15bfn001as1n32x5 wire721 (.a(net58),
    .o(net721));
 b15bfn000ah1n48x5 wire722 (.a(net57),
    .o(net722));
 b15bfn001ah1n48x5 wire723 (.a(net56),
    .o(net723));
 b15bfn001as1n32x5 wire724 (.a(net55),
    .o(net724));
 b15bfn001ah1n64x5 fanout725 (.a(net732),
    .o(net725));
 b15bfn001as1n48x5 fanout726 (.a(net727),
    .o(net726));
 b15bfn001as1n48x5 fanout727 (.a(net731),
    .o(net727));
 b15bfn001as1n48x5 fanout728 (.a(net732),
    .o(net728));
 b15bfn001as1n32x5 fanout729 (.a(net732),
    .o(net729));
 b15bfn001as1n48x5 fanout730 (.a(net733),
    .o(net730));
 b15bfn001as1n64x5 fanout731 (.a(net759),
    .o(net731));
 b15bfn001ah1n48x5 wire732 (.a(net731),
    .o(net732));
 b15bfn001as1n32x5 max_length733 (.a(net731),
    .o(net733));
 b15bfn001as1n48x5 fanout734 (.a(net741),
    .o(net734));
 b15bfn001as1n48x5 fanout735 (.a(net740),
    .o(net735));
 b15bfn001as1n48x5 fanout736 (.a(net740),
    .o(net736));
 b15bfn001as1n48x5 fanout737 (.a(net738),
    .o(net737));
 b15bfn001as1n48x5 fanout738 (.a(net741),
    .o(net738));
 b15bfn001ah1n48x5 max_length739 (.a(net738),
    .o(net739));
 b15bfn001ah1n48x5 fanout740 (.a(net37),
    .o(net740));
 b15bfn001as1n32x5 max_length741 (.a(net740),
    .o(net741));
 b15bfn001ah1n64x5 fanout742 (.a(net745),
    .o(net742));
 b15bfn001as1n24x5 fanout743 (.a(net745),
    .o(net743));
 b15bfn001ah1n64x5 fanout744 (.a(net745),
    .o(net744));
 b15bfn001ah1n48x5 fanout745 (.a(net758),
    .o(net745));
 b15bfn001as1n48x5 fanout746 (.a(net748),
    .o(net746));
 b15bfn001as1n48x5 fanout747 (.a(net748),
    .o(net747));
 b15bfn001as1n48x5 fanout748 (.a(net758),
    .o(net748));
 b15bfn001as1n48x5 fanout749 (.a(net752),
    .o(net749));
 b15bfn001as1n32x5 fanout750 (.a(net752),
    .o(net750));
 b15bfn001as1n64x5 fanout751 (.a(net752),
    .o(net751));
 b15bfn001as1n48x5 fanout752 (.a(net760),
    .o(net752));
 b15bfn001ah1n64x5 fanout753 (.a(net757),
    .o(net753));
 b15bfn001as1n48x5 fanout754 (.a(net755),
    .o(net754));
 b15bfn001as1n48x5 fanout755 (.a(net756),
    .o(net755));
 b15bfn001as1n48x5 fanout756 (.a(net760),
    .o(net756));
 b15bfn001ah1n48x5 wire757 (.a(net756),
    .o(net757));
 b15bfn000ah1n48x5 wire758 (.a(net759),
    .o(net758));
 b15bfn001ah1n32x5 wire759 (.a(net37),
    .o(net759));
 b15bfn001as1n24x5 wire760 (.a(net37),
    .o(net760));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_0__cio_gpio_en_q_reg_1__761 (.o(net761));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_0__cio_gpio_en_q_reg_1__762 (.o(net762));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_10__cio_gpio_en_q_reg_11__763 (.o(net763));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_10__cio_gpio_en_q_reg_11__764 (.o(net764));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_12__cio_gpio_en_q_reg_13__765 (.o(net765));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_12__cio_gpio_en_q_reg_13__766 (.o(net766));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_14__cio_gpio_en_q_reg_15__767 (.o(net767));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_14__cio_gpio_en_q_reg_15__768 (.o(net768));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_16__cio_gpio_en_q_reg_17__769 (.o(net769));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_16__cio_gpio_en_q_reg_17__770 (.o(net770));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_18__cio_gpio_en_q_reg_19__771 (.o(net771));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_18__cio_gpio_en_q_reg_19__772 (.o(net772));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_20__cio_gpio_en_q_reg_21__773 (.o(net773));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_20__cio_gpio_en_q_reg_21__774 (.o(net774));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_22__cio_gpio_en_q_reg_23__775 (.o(net775));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_22__cio_gpio_en_q_reg_23__776 (.o(net776));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_24__cio_gpio_en_q_reg_25__777 (.o(net777));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_24__cio_gpio_en_q_reg_25__778 (.o(net778));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_26__cio_gpio_en_q_reg_27__779 (.o(net779));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_26__cio_gpio_en_q_reg_27__780 (.o(net780));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_28__cio_gpio_en_q_reg_29__781 (.o(net781));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_28__cio_gpio_en_q_reg_29__782 (.o(net782));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_2__cio_gpio_en_q_reg_3__783 (.o(net783));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_2__cio_gpio_en_q_reg_3__784 (.o(net784));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_30__cio_gpio_en_q_reg_31__785 (.o(net785));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_30__cio_gpio_en_q_reg_31__786 (.o(net786));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_4__cio_gpio_en_q_reg_5__787 (.o(net787));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_4__cio_gpio_en_q_reg_5__788 (.o(net788));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_6__cio_gpio_en_q_reg_7__789 (.o(net789));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_6__cio_gpio_en_q_reg_7__790 (.o(net790));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_8__cio_gpio_en_q_reg_9__791 (.o(net791));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_8__cio_gpio_en_q_reg_9__792 (.o(net792));
 b15tilo00an1n03x5 cio_gpio_q_reg_0__cio_gpio_q_reg_1__793 (.o(net793));
 b15tilo00an1n03x5 cio_gpio_q_reg_0__cio_gpio_q_reg_1__794 (.o(net794));
 b15tilo00an1n03x5 cio_gpio_q_reg_10__cio_gpio_q_reg_11__795 (.o(net795));
 b15tilo00an1n03x5 cio_gpio_q_reg_10__cio_gpio_q_reg_11__796 (.o(net796));
 b15tilo00an1n03x5 cio_gpio_q_reg_12__cio_gpio_q_reg_13__797 (.o(net797));
 b15tilo00an1n03x5 cio_gpio_q_reg_12__cio_gpio_q_reg_13__798 (.o(net798));
 b15tilo00an1n03x5 cio_gpio_q_reg_14__cio_gpio_q_reg_15__799 (.o(net799));
 b15tilo00an1n03x5 cio_gpio_q_reg_14__cio_gpio_q_reg_15__800 (.o(net800));
 b15tilo00an1n03x5 cio_gpio_q_reg_16__cio_gpio_q_reg_17__801 (.o(net801));
 b15tilo00an1n03x5 cio_gpio_q_reg_16__cio_gpio_q_reg_17__802 (.o(net802));
 b15tilo00an1n03x5 cio_gpio_q_reg_18__cio_gpio_q_reg_19__803 (.o(net803));
 b15tilo00an1n03x5 cio_gpio_q_reg_18__cio_gpio_q_reg_19__804 (.o(net804));
 b15tilo00an1n03x5 cio_gpio_q_reg_20__cio_gpio_q_reg_21__805 (.o(net805));
 b15tilo00an1n03x5 cio_gpio_q_reg_20__cio_gpio_q_reg_21__806 (.o(net806));
 b15tilo00an1n03x5 cio_gpio_q_reg_22__cio_gpio_q_reg_23__807 (.o(net807));
 b15tilo00an1n03x5 cio_gpio_q_reg_22__cio_gpio_q_reg_23__808 (.o(net808));
 b15tilo00an1n03x5 cio_gpio_q_reg_24__cio_gpio_q_reg_25__809 (.o(net809));
 b15tilo00an1n03x5 cio_gpio_q_reg_24__cio_gpio_q_reg_25__810 (.o(net810));
 b15tilo00an1n03x5 cio_gpio_q_reg_26__cio_gpio_q_reg_27__811 (.o(net811));
 b15tilo00an1n03x5 cio_gpio_q_reg_26__cio_gpio_q_reg_27__812 (.o(net812));
 b15tilo00an1n03x5 cio_gpio_q_reg_28__cio_gpio_q_reg_29__813 (.o(net813));
 b15tilo00an1n03x5 cio_gpio_q_reg_28__cio_gpio_q_reg_29__814 (.o(net814));
 b15tilo00an1n03x5 cio_gpio_q_reg_2__cio_gpio_q_reg_3__815 (.o(net815));
 b15tilo00an1n03x5 cio_gpio_q_reg_2__cio_gpio_q_reg_3__816 (.o(net816));
 b15tilo00an1n03x5 cio_gpio_q_reg_30__cio_gpio_q_reg_31__817 (.o(net817));
 b15tilo00an1n03x5 cio_gpio_q_reg_30__cio_gpio_q_reg_31__818 (.o(net818));
 b15tilo00an1n03x5 cio_gpio_q_reg_4__cio_gpio_q_reg_5__819 (.o(net819));
 b15tilo00an1n03x5 cio_gpio_q_reg_4__cio_gpio_q_reg_5__820 (.o(net820));
 b15tilo00an1n03x5 cio_gpio_q_reg_6__cio_gpio_q_reg_7__821 (.o(net821));
 b15tilo00an1n03x5 cio_gpio_q_reg_6__cio_gpio_q_reg_7__822 (.o(net822));
 b15tilo00an1n03x5 cio_gpio_q_reg_8__cio_gpio_q_reg_9__823 (.o(net823));
 b15tilo00an1n03x5 cio_gpio_q_reg_8__cio_gpio_q_reg_9__824 (.o(net824));
 b15tilo00an1n03x5 clk_gate_cio_gpio_en_q_reg_0_latch_825 (.o(net825));
 b15tilo00an1n03x5 clk_gate_cio_gpio_en_q_reg_latch_826 (.o(net826));
 b15tilo00an1n03x5 clk_gate_cio_gpio_q_reg_0_latch_827 (.o(net827));
 b15tilo00an1n03x5 clk_gate_cio_gpio_q_reg_latch_828 (.o(net828));
 b15tilo00an1n03x5 data_in_q_reg_0__data_in_q_reg_1__829 (.o(net829));
 b15tilo00an1n03x5 data_in_q_reg_0__data_in_q_reg_1__830 (.o(net830));
 b15tilo00an1n03x5 data_in_q_reg_10__data_in_q_reg_11__831 (.o(net831));
 b15tilo00an1n03x5 data_in_q_reg_10__data_in_q_reg_11__832 (.o(net832));
 b15tilo00an1n03x5 data_in_q_reg_12__data_in_q_reg_13__833 (.o(net833));
 b15tilo00an1n03x5 data_in_q_reg_12__data_in_q_reg_13__834 (.o(net834));
 b15tilo00an1n03x5 data_in_q_reg_14__data_in_q_reg_15__835 (.o(net835));
 b15tilo00an1n03x5 data_in_q_reg_14__data_in_q_reg_15__836 (.o(net836));
 b15tilo00an1n03x5 data_in_q_reg_16__data_in_q_reg_17__837 (.o(net837));
 b15tilo00an1n03x5 data_in_q_reg_16__data_in_q_reg_17__838 (.o(net838));
 b15tilo00an1n03x5 data_in_q_reg_18__data_in_q_reg_19__839 (.o(net839));
 b15tilo00an1n03x5 data_in_q_reg_18__data_in_q_reg_19__840 (.o(net840));
 b15tilo00an1n03x5 data_in_q_reg_20__data_in_q_reg_21__841 (.o(net841));
 b15tilo00an1n03x5 data_in_q_reg_20__data_in_q_reg_21__842 (.o(net842));
 b15tilo00an1n03x5 data_in_q_reg_22__data_in_q_reg_23__843 (.o(net843));
 b15tilo00an1n03x5 data_in_q_reg_22__data_in_q_reg_23__844 (.o(net844));
 b15tilo00an1n03x5 data_in_q_reg_24__data_in_q_reg_25__845 (.o(net845));
 b15tilo00an1n03x5 data_in_q_reg_24__data_in_q_reg_25__846 (.o(net846));
 b15tilo00an1n03x5 data_in_q_reg_26__data_in_q_reg_27__847 (.o(net847));
 b15tilo00an1n03x5 data_in_q_reg_26__data_in_q_reg_27__848 (.o(net848));
 b15tilo00an1n03x5 data_in_q_reg_28__data_in_q_reg_29__849 (.o(net849));
 b15tilo00an1n03x5 data_in_q_reg_28__data_in_q_reg_29__850 (.o(net850));
 b15tilo00an1n03x5 data_in_q_reg_2__data_in_q_reg_3__851 (.o(net851));
 b15tilo00an1n03x5 data_in_q_reg_2__data_in_q_reg_3__852 (.o(net852));
 b15tilo00an1n03x5 data_in_q_reg_30__data_in_q_reg_31__853 (.o(net853));
 b15tilo00an1n03x5 data_in_q_reg_30__data_in_q_reg_31__854 (.o(net854));
 b15tilo00an1n03x5 data_in_q_reg_4__data_in_q_reg_5__855 (.o(net855));
 b15tilo00an1n03x5 data_in_q_reg_4__data_in_q_reg_5__856 (.o(net856));
 b15tilo00an1n03x5 data_in_q_reg_6__data_in_q_reg_7__857 (.o(net857));
 b15tilo00an1n03x5 data_in_q_reg_6__data_in_q_reg_7__858 (.o(net858));
 b15tilo00an1n03x5 data_in_q_reg_8__data_in_q_reg_9__859 (.o(net859));
 b15tilo00an1n03x5 data_in_q_reg_8__data_in_q_reg_9__860 (.o(net860));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg_861 (.o(net861));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg_862 (.o(net862));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg_863 (.o(net863));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg_864 (.o(net864));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0__gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1__865 (.o(net865));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0__gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1__866 (.o(net866));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__867 (.o(net867));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__868 (.o(net868));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq_reg_869 (.o(net869));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__870 (.o(net870));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__871 (.o(net871));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg_872 (.o(net872));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg_873 (.o(net873));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_0__874 (.o(net874));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_1__875 (.o(net875));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq_reg_876 (.o(net876));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__877 (.o(net877));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__878 (.o(net878));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__879 (.o(net879));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__880 (.o(net880));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg_881 (.o(net881));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg_882 (.o(net882));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_0__883 (.o(net883));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_1__884 (.o(net884));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__885 (.o(net885));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__886 (.o(net886));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_1__887 (.o(net887));
 b15tilo00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_0__gen_filter_0__u_filter_diff_ctr_q_reg_1__888 (.o(net888));
 b15tilo00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_0__gen_filter_0__u_filter_diff_ctr_q_reg_1__889 (.o(net889));
 b15tilo00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_2__gen_filter_0__u_filter_diff_ctr_q_reg_3__890 (.o(net890));
 b15tilo00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_2__gen_filter_0__u_filter_diff_ctr_q_reg_3__891 (.o(net891));
 b15tilo00an1n03x5 gen_filter_0__u_filter_filter_q_reg_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__892 (.o(net892));
 b15tilo00an1n03x5 gen_filter_0__u_filter_filter_q_reg_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__893 (.o(net893));
 b15tilo00an1n03x5 gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_1__u_filter_diff_ctr_q_reg_0__894 (.o(net894));
 b15tilo00an1n03x5 gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_1__u_filter_diff_ctr_q_reg_0__895 (.o(net895));
 b15tilo00an1n03x5 gen_filter_0__u_filter_stored_value_q_reg_896 (.o(net896));
 b15tilo00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_1__gen_filter_10__u_filter_diff_ctr_q_reg_2__897 (.o(net897));
 b15tilo00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_1__gen_filter_10__u_filter_diff_ctr_q_reg_2__898 (.o(net898));
 b15tilo00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_filter_q_reg_899 (.o(net899));
 b15tilo00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_filter_q_reg_900 (.o(net900));
 b15tilo00an1n03x5 gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__901 (.o(net901));
 b15tilo00an1n03x5 gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__902 (.o(net902));
 b15tilo00an1n03x5 gen_filter_10__u_filter_stored_value_q_reg_903 (.o(net903));
 b15tilo00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_0__gen_filter_12__u_filter_diff_ctr_q_reg_0__904 (.o(net904));
 b15tilo00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_0__gen_filter_12__u_filter_diff_ctr_q_reg_0__905 (.o(net905));
 b15tilo00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_2__gen_filter_11__u_filter_diff_ctr_q_reg_3__906 (.o(net906));
 b15tilo00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_2__gen_filter_11__u_filter_diff_ctr_q_reg_3__907 (.o(net907));
 b15tilo00an1n03x5 gen_filter_11__u_filter_filter_q_reg_gen_filter_12__u_filter_filter_q_reg_908 (.o(net908));
 b15tilo00an1n03x5 gen_filter_11__u_filter_filter_q_reg_gen_filter_12__u_filter_filter_q_reg_909 (.o(net909));
 b15tilo00an1n03x5 gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_3__910 (.o(net910));
 b15tilo00an1n03x5 gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_3__911 (.o(net911));
 b15tilo00an1n03x5 gen_filter_11__u_filter_stored_value_q_reg_912 (.o(net912));
 b15tilo00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_1__gen_filter_12__u_filter_diff_ctr_q_reg_2__913 (.o(net913));
 b15tilo00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_1__gen_filter_12__u_filter_diff_ctr_q_reg_2__914 (.o(net914));
 b15tilo00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_diff_ctr_q_reg_0__915 (.o(net915));
 b15tilo00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_diff_ctr_q_reg_0__916 (.o(net916));
 b15tilo00an1n03x5 gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__917 (.o(net917));
 b15tilo00an1n03x5 gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__918 (.o(net918));
 b15tilo00an1n03x5 gen_filter_12__u_filter_stored_value_q_reg_919 (.o(net919));
 b15tilo00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_1__gen_filter_13__u_filter_diff_ctr_q_reg_2__920 (.o(net920));
 b15tilo00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_1__gen_filter_13__u_filter_diff_ctr_q_reg_2__921 (.o(net921));
 b15tilo00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_filter_q_reg_922 (.o(net922));
 b15tilo00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_filter_q_reg_923 (.o(net923));
 b15tilo00an1n03x5 gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__924 (.o(net924));
 b15tilo00an1n03x5 gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__925 (.o(net925));
 b15tilo00an1n03x5 gen_filter_13__u_filter_stored_value_q_reg_926 (.o(net926));
 b15tilo00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_1__927 (.o(net927));
 b15tilo00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_1__928 (.o(net928));
 b15tilo00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_2__gen_filter_26__u_filter_diff_ctr_q_reg_0__929 (.o(net929));
 b15tilo00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_2__gen_filter_26__u_filter_diff_ctr_q_reg_0__930 (.o(net930));
 b15tilo00an1n03x5 gen_filter_14__u_filter_filter_q_reg_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__931 (.o(net931));
 b15tilo00an1n03x5 gen_filter_14__u_filter_filter_q_reg_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__932 (.o(net932));
 b15tilo00an1n03x5 gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_diff_ctr_q_reg_0__933 (.o(net933));
 b15tilo00an1n03x5 gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_diff_ctr_q_reg_0__934 (.o(net934));
 b15tilo00an1n03x5 gen_filter_14__u_filter_stored_value_q_reg_935 (.o(net935));
 b15tilo00an1n03x5 gen_filter_15__u_filter_diff_ctr_q_reg_1__gen_filter_15__u_filter_diff_ctr_q_reg_2__936 (.o(net936));
 b15tilo00an1n03x5 gen_filter_15__u_filter_diff_ctr_q_reg_1__gen_filter_15__u_filter_diff_ctr_q_reg_2__937 (.o(net937));
 b15tilo00an1n03x5 gen_filter_15__u_filter_filter_q_reg_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__938 (.o(net938));
 b15tilo00an1n03x5 gen_filter_15__u_filter_filter_q_reg_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__939 (.o(net939));
 b15tilo00an1n03x5 gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_diff_ctr_q_reg_0__940 (.o(net940));
 b15tilo00an1n03x5 gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_diff_ctr_q_reg_0__941 (.o(net941));
 b15tilo00an1n03x5 gen_filter_15__u_filter_stored_value_q_reg_942 (.o(net942));
 b15tilo00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_0__gen_filter_16__u_filter_diff_ctr_q_reg_1__943 (.o(net943));
 b15tilo00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_0__gen_filter_16__u_filter_diff_ctr_q_reg_1__944 (.o(net944));
 b15tilo00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_2__gen_filter_16__u_filter_diff_ctr_q_reg_3__945 (.o(net945));
 b15tilo00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_2__gen_filter_16__u_filter_diff_ctr_q_reg_3__946 (.o(net946));
 b15tilo00an1n03x5 gen_filter_16__u_filter_filter_q_reg_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__947 (.o(net947));
 b15tilo00an1n03x5 gen_filter_16__u_filter_filter_q_reg_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__948 (.o(net948));
 b15tilo00an1n03x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__949 (.o(net949));
 b15tilo00an1n03x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__950 (.o(net950));
 b15tilo00an1n03x5 gen_filter_16__u_filter_stored_value_q_reg_951 (.o(net951));
 b15tilo00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_1__gen_filter_17__u_filter_diff_ctr_q_reg_2__952 (.o(net952));
 b15tilo00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_1__gen_filter_17__u_filter_diff_ctr_q_reg_2__953 (.o(net953));
 b15tilo00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_3__gen_filter_17__u_filter_filter_q_reg_954 (.o(net954));
 b15tilo00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_3__gen_filter_17__u_filter_filter_q_reg_955 (.o(net955));
 b15tilo00an1n03x5 gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_18__u_filter_diff_ctr_q_reg_0__956 (.o(net956));
 b15tilo00an1n03x5 gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_18__u_filter_diff_ctr_q_reg_0__957 (.o(net957));
 b15tilo00an1n03x5 gen_filter_17__u_filter_stored_value_q_reg_958 (.o(net958));
 b15tilo00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_1__gen_filter_18__u_filter_diff_ctr_q_reg_2__959 (.o(net959));
 b15tilo00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_1__gen_filter_18__u_filter_diff_ctr_q_reg_2__960 (.o(net960));
 b15tilo00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_3__gen_filter_18__u_filter_filter_q_reg_961 (.o(net961));
 b15tilo00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_3__gen_filter_18__u_filter_filter_q_reg_962 (.o(net962));
 b15tilo00an1n03x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__963 (.o(net963));
 b15tilo00an1n03x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__964 (.o(net964));
 b15tilo00an1n03x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__965 (.o(net965));
 b15tilo00an1n03x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__966 (.o(net966));
 b15tilo00an1n03x5 gen_filter_18__u_filter_stored_value_q_reg_967 (.o(net967));
 b15tilo00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_1__gen_filter_19__u_filter_diff_ctr_q_reg_2__968 (.o(net968));
 b15tilo00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_1__gen_filter_19__u_filter_diff_ctr_q_reg_2__969 (.o(net969));
 b15tilo00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_3__gen_filter_19__u_filter_filter_q_reg_970 (.o(net970));
 b15tilo00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_3__gen_filter_19__u_filter_filter_q_reg_971 (.o(net971));
 b15tilo00an1n03x5 gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__972 (.o(net972));
 b15tilo00an1n03x5 gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__973 (.o(net973));
 b15tilo00an1n03x5 gen_filter_19__u_filter_stored_value_q_reg_974 (.o(net974));
 b15tilo00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_1__gen_filter_1__u_filter_diff_ctr_q_reg_2__975 (.o(net975));
 b15tilo00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_1__gen_filter_1__u_filter_diff_ctr_q_reg_2__976 (.o(net976));
 b15tilo00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_3__gen_filter_1__u_filter_filter_q_reg_977 (.o(net977));
 b15tilo00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_3__gen_filter_1__u_filter_filter_q_reg_978 (.o(net978));
 b15tilo00an1n03x5 gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__979 (.o(net979));
 b15tilo00an1n03x5 gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__980 (.o(net980));
 b15tilo00an1n03x5 gen_filter_1__u_filter_stored_value_q_reg_981 (.o(net981));
 b15tilo00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_0__gen_filter_20__u_filter_diff_ctr_q_reg_1__982 (.o(net982));
 b15tilo00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_0__gen_filter_20__u_filter_diff_ctr_q_reg_1__983 (.o(net983));
 b15tilo00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_2__gen_filter_20__u_filter_diff_ctr_q_reg_3__984 (.o(net984));
 b15tilo00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_2__gen_filter_20__u_filter_diff_ctr_q_reg_3__985 (.o(net985));
 b15tilo00an1n03x5 gen_filter_20__u_filter_filter_q_reg_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__986 (.o(net986));
 b15tilo00an1n03x5 gen_filter_20__u_filter_filter_q_reg_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__987 (.o(net987));
 b15tilo00an1n03x5 gen_filter_20__u_filter_stored_value_q_reg_988 (.o(net988));
 b15tilo00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_0__gen_filter_21__u_filter_diff_ctr_q_reg_1__989 (.o(net989));
 b15tilo00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_0__gen_filter_21__u_filter_diff_ctr_q_reg_1__990 (.o(net990));
 b15tilo00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_2__gen_filter_21__u_filter_diff_ctr_q_reg_3__991 (.o(net991));
 b15tilo00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_2__gen_filter_21__u_filter_diff_ctr_q_reg_3__992 (.o(net992));
 b15tilo00an1n03x5 gen_filter_21__u_filter_filter_q_reg_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__993 (.o(net993));
 b15tilo00an1n03x5 gen_filter_21__u_filter_filter_q_reg_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__994 (.o(net994));
 b15tilo00an1n03x5 gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_diff_ctr_q_reg_0__995 (.o(net995));
 b15tilo00an1n03x5 gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_diff_ctr_q_reg_0__996 (.o(net996));
 b15tilo00an1n03x5 gen_filter_21__u_filter_stored_value_q_reg_997 (.o(net997));
 b15tilo00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_0__gen_filter_22__u_filter_diff_ctr_q_reg_1__998 (.o(net998));
 b15tilo00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_0__gen_filter_22__u_filter_diff_ctr_q_reg_1__999 (.o(net999));
 b15tilo00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_2__gen_filter_22__u_filter_diff_ctr_q_reg_3__1000 (.o(net1000));
 b15tilo00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_2__gen_filter_22__u_filter_diff_ctr_q_reg_3__1001 (.o(net1001));
 b15tilo00an1n03x5 gen_filter_22__u_filter_filter_q_reg_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1002 (.o(net1002));
 b15tilo00an1n03x5 gen_filter_22__u_filter_filter_q_reg_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1003 (.o(net1003));
 b15tilo00an1n03x5 gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_diff_ctr_q_reg_0__1004 (.o(net1004));
 b15tilo00an1n03x5 gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_diff_ctr_q_reg_0__1005 (.o(net1005));
 b15tilo00an1n03x5 gen_filter_22__u_filter_stored_value_q_reg_1006 (.o(net1006));
 b15tilo00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_1__gen_filter_23__u_filter_diff_ctr_q_reg_2__1007 (.o(net1007));
 b15tilo00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_1__gen_filter_23__u_filter_diff_ctr_q_reg_2__1008 (.o(net1008));
 b15tilo00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_3__gen_filter_23__u_filter_filter_q_reg_1009 (.o(net1009));
 b15tilo00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_3__gen_filter_23__u_filter_filter_q_reg_1010 (.o(net1010));
 b15tilo00an1n03x5 gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1011 (.o(net1011));
 b15tilo00an1n03x5 gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1012 (.o(net1012));
 b15tilo00an1n03x5 gen_filter_23__u_filter_stored_value_q_reg_1013 (.o(net1013));
 b15tilo00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_0__gen_filter_24__u_filter_diff_ctr_q_reg_1__1014 (.o(net1014));
 b15tilo00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_0__gen_filter_24__u_filter_diff_ctr_q_reg_1__1015 (.o(net1015));
 b15tilo00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_2__gen_filter_24__u_filter_diff_ctr_q_reg_3__1016 (.o(net1016));
 b15tilo00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_2__gen_filter_24__u_filter_diff_ctr_q_reg_3__1017 (.o(net1017));
 b15tilo00an1n03x5 gen_filter_24__u_filter_filter_q_reg_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1018 (.o(net1018));
 b15tilo00an1n03x5 gen_filter_24__u_filter_filter_q_reg_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1019 (.o(net1019));
 b15tilo00an1n03x5 gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_25__u_filter_diff_ctr_q_reg_0__1020 (.o(net1020));
 b15tilo00an1n03x5 gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_25__u_filter_diff_ctr_q_reg_0__1021 (.o(net1021));
 b15tilo00an1n03x5 gen_filter_24__u_filter_stored_value_q_reg_1022 (.o(net1022));
 b15tilo00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_1__gen_filter_25__u_filter_diff_ctr_q_reg_2__1023 (.o(net1023));
 b15tilo00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_1__gen_filter_25__u_filter_diff_ctr_q_reg_2__1024 (.o(net1024));
 b15tilo00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_3__gen_filter_25__u_filter_filter_q_reg_1025 (.o(net1025));
 b15tilo00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_3__gen_filter_25__u_filter_filter_q_reg_1026 (.o(net1026));
 b15tilo00an1n03x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_0__1027 (.o(net1027));
 b15tilo00an1n03x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_0__1028 (.o(net1028));
 b15tilo00an1n03x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_27__u_filter_diff_ctr_q_reg_0__1029 (.o(net1029));
 b15tilo00an1n03x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_27__u_filter_diff_ctr_q_reg_0__1030 (.o(net1030));
 b15tilo00an1n03x5 gen_filter_25__u_filter_stored_value_q_reg_1031 (.o(net1031));
 b15tilo00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_1__gen_filter_26__u_filter_diff_ctr_q_reg_2__1032 (.o(net1032));
 b15tilo00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_1__gen_filter_26__u_filter_diff_ctr_q_reg_2__1033 (.o(net1033));
 b15tilo00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_3__gen_filter_26__u_filter_filter_q_reg_1034 (.o(net1034));
 b15tilo00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_3__gen_filter_26__u_filter_filter_q_reg_1035 (.o(net1035));
 b15tilo00an1n03x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1036 (.o(net1036));
 b15tilo00an1n03x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1037 (.o(net1037));
 b15tilo00an1n03x5 gen_filter_26__u_filter_stored_value_q_reg_1038 (.o(net1038));
 b15tilo00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_1__gen_filter_27__u_filter_diff_ctr_q_reg_2__1039 (.o(net1039));
 b15tilo00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_1__gen_filter_27__u_filter_diff_ctr_q_reg_2__1040 (.o(net1040));
 b15tilo00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_3__gen_filter_27__u_filter_filter_q_reg_1041 (.o(net1041));
 b15tilo00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_3__gen_filter_27__u_filter_filter_q_reg_1042 (.o(net1042));
 b15tilo00an1n03x5 gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1043 (.o(net1043));
 b15tilo00an1n03x5 gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1044 (.o(net1044));
 b15tilo00an1n03x5 gen_filter_27__u_filter_stored_value_q_reg_1045 (.o(net1045));
 b15tilo00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_1__gen_filter_28__u_filter_diff_ctr_q_reg_2__1046 (.o(net1046));
 b15tilo00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_1__gen_filter_28__u_filter_diff_ctr_q_reg_2__1047 (.o(net1047));
 b15tilo00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_3__gen_filter_28__u_filter_filter_q_reg_1048 (.o(net1048));
 b15tilo00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_3__gen_filter_28__u_filter_filter_q_reg_1049 (.o(net1049));
 b15tilo00an1n03x5 gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1050 (.o(net1050));
 b15tilo00an1n03x5 gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1051 (.o(net1051));
 b15tilo00an1n03x5 gen_filter_28__u_filter_stored_value_q_reg_1052 (.o(net1052));
 b15tilo00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_0__gen_filter_29__u_filter_diff_ctr_q_reg_1__1053 (.o(net1053));
 b15tilo00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_0__gen_filter_29__u_filter_diff_ctr_q_reg_1__1054 (.o(net1054));
 b15tilo00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_2__gen_filter_29__u_filter_diff_ctr_q_reg_3__1055 (.o(net1055));
 b15tilo00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_2__gen_filter_29__u_filter_diff_ctr_q_reg_3__1056 (.o(net1056));
 b15tilo00an1n03x5 gen_filter_29__u_filter_filter_q_reg_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1057 (.o(net1057));
 b15tilo00an1n03x5 gen_filter_29__u_filter_filter_q_reg_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1058 (.o(net1058));
 b15tilo00an1n03x5 gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1059 (.o(net1059));
 b15tilo00an1n03x5 gen_filter_29__u_filter_stored_value_q_reg_1060 (.o(net1060));
 b15tilo00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_0__gen_filter_2__u_filter_diff_ctr_q_reg_1__1061 (.o(net1061));
 b15tilo00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_0__gen_filter_2__u_filter_diff_ctr_q_reg_1__1062 (.o(net1062));
 b15tilo00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_2__gen_filter_2__u_filter_diff_ctr_q_reg_3__1063 (.o(net1063));
 b15tilo00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_2__gen_filter_2__u_filter_diff_ctr_q_reg_3__1064 (.o(net1064));
 b15tilo00an1n03x5 gen_filter_2__u_filter_filter_q_reg_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1065 (.o(net1065));
 b15tilo00an1n03x5 gen_filter_2__u_filter_filter_q_reg_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1066 (.o(net1066));
 b15tilo00an1n03x5 gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1067 (.o(net1067));
 b15tilo00an1n03x5 gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1068 (.o(net1068));
 b15tilo00an1n03x5 gen_filter_2__u_filter_stored_value_q_reg_1069 (.o(net1069));
 b15tilo00an1n03x5 gen_filter_30__u_filter_diff_ctr_q_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_1__1070 (.o(net1070));
 b15tilo00an1n03x5 gen_filter_30__u_filter_diff_ctr_q_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_1__1071 (.o(net1071));
 b15tilo00an1n03x5 gen_filter_30__u_filter_diff_ctr_q_reg_2__gen_filter_30__u_filter_diff_ctr_q_reg_3__1072 (.o(net1072));
 b15tilo00an1n03x5 gen_filter_30__u_filter_diff_ctr_q_reg_2__gen_filter_30__u_filter_diff_ctr_q_reg_3__1073 (.o(net1073));
 b15tilo00an1n03x5 gen_filter_30__u_filter_filter_q_reg_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1074 (.o(net1074));
 b15tilo00an1n03x5 gen_filter_30__u_filter_filter_q_reg_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1075 (.o(net1075));
 b15tilo00an1n03x5 gen_filter_30__u_filter_stored_value_q_reg_1076 (.o(net1076));
 b15tilo00an1n03x5 gen_filter_31__u_filter_diff_ctr_q_reg_0__gen_filter_31__u_filter_diff_ctr_q_reg_1__1077 (.o(net1077));
 b15tilo00an1n03x5 gen_filter_31__u_filter_diff_ctr_q_reg_0__gen_filter_31__u_filter_diff_ctr_q_reg_1__1078 (.o(net1078));
 b15tilo00an1n03x5 gen_filter_31__u_filter_diff_ctr_q_reg_2__gen_filter_31__u_filter_diff_ctr_q_reg_3__1079 (.o(net1079));
 b15tilo00an1n03x5 gen_filter_31__u_filter_diff_ctr_q_reg_2__gen_filter_31__u_filter_diff_ctr_q_reg_3__1080 (.o(net1080));
 b15tilo00an1n03x5 gen_filter_31__u_filter_filter_q_reg_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1081 (.o(net1081));
 b15tilo00an1n03x5 gen_filter_31__u_filter_filter_q_reg_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1082 (.o(net1082));
 b15tilo00an1n03x5 gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_3__1083 (.o(net1083));
 b15tilo00an1n03x5 gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_3__1084 (.o(net1084));
 b15tilo00an1n03x5 gen_filter_31__u_filter_stored_value_q_reg_1085 (.o(net1085));
 b15tilo00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_0__gen_filter_3__u_filter_diff_ctr_q_reg_1__1086 (.o(net1086));
 b15tilo00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_0__gen_filter_3__u_filter_diff_ctr_q_reg_1__1087 (.o(net1087));
 b15tilo00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_2__gen_filter_3__u_filter_diff_ctr_q_reg_3__1088 (.o(net1088));
 b15tilo00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_2__gen_filter_3__u_filter_diff_ctr_q_reg_3__1089 (.o(net1089));
 b15tilo00an1n03x5 gen_filter_3__u_filter_filter_q_reg_gen_filter_4__u_filter_diff_ctr_q_reg_0__1090 (.o(net1090));
 b15tilo00an1n03x5 gen_filter_3__u_filter_filter_q_reg_gen_filter_4__u_filter_diff_ctr_q_reg_0__1091 (.o(net1091));
 b15tilo00an1n03x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1092 (.o(net1092));
 b15tilo00an1n03x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1093 (.o(net1093));
 b15tilo00an1n03x5 gen_filter_3__u_filter_stored_value_q_reg_1094 (.o(net1094));
 b15tilo00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_1__gen_filter_4__u_filter_diff_ctr_q_reg_2__1095 (.o(net1095));
 b15tilo00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_1__gen_filter_4__u_filter_diff_ctr_q_reg_2__1096 (.o(net1096));
 b15tilo00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_diff_ctr_q_reg_0__1097 (.o(net1097));
 b15tilo00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_diff_ctr_q_reg_0__1098 (.o(net1098));
 b15tilo00an1n03x5 gen_filter_4__u_filter_filter_q_reg_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1099 (.o(net1099));
 b15tilo00an1n03x5 gen_filter_4__u_filter_filter_q_reg_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1100 (.o(net1100));
 b15tilo00an1n03x5 gen_filter_4__u_filter_stored_value_q_reg_1101 (.o(net1101));
 b15tilo00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_0__gen_filter_5__u_filter_diff_ctr_q_reg_1__1102 (.o(net1102));
 b15tilo00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_0__gen_filter_5__u_filter_diff_ctr_q_reg_1__1103 (.o(net1103));
 b15tilo00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_2__gen_filter_5__u_filter_filter_q_reg_1104 (.o(net1104));
 b15tilo00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_2__gen_filter_5__u_filter_filter_q_reg_1105 (.o(net1105));
 b15tilo00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_3__gen_filter_6__u_filter_diff_ctr_q_reg_0__1106 (.o(net1106));
 b15tilo00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_3__gen_filter_6__u_filter_diff_ctr_q_reg_0__1107 (.o(net1107));
 b15tilo00an1n03x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_diff_ctr_q_reg_0__1108 (.o(net1108));
 b15tilo00an1n03x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_diff_ctr_q_reg_0__1109 (.o(net1109));
 b15tilo00an1n03x5 gen_filter_5__u_filter_stored_value_q_reg_1110 (.o(net1110));
 b15tilo00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_1__gen_filter_6__u_filter_diff_ctr_q_reg_2__1111 (.o(net1111));
 b15tilo00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_1__gen_filter_6__u_filter_diff_ctr_q_reg_2__1112 (.o(net1112));
 b15tilo00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_3__gen_filter_6__u_filter_filter_q_reg_1113 (.o(net1113));
 b15tilo00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_3__gen_filter_6__u_filter_filter_q_reg_1114 (.o(net1114));
 b15tilo00an1n03x5 gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1115 (.o(net1115));
 b15tilo00an1n03x5 gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1116 (.o(net1116));
 b15tilo00an1n03x5 gen_filter_6__u_filter_stored_value_q_reg_1117 (.o(net1117));
 b15tilo00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_0__gen_filter_7__u_filter_diff_ctr_q_reg_1__1118 (.o(net1118));
 b15tilo00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_0__gen_filter_7__u_filter_diff_ctr_q_reg_1__1119 (.o(net1119));
 b15tilo00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_2__gen_filter_7__u_filter_diff_ctr_q_reg_3__1120 (.o(net1120));
 b15tilo00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_2__gen_filter_7__u_filter_diff_ctr_q_reg_3__1121 (.o(net1121));
 b15tilo00an1n03x5 gen_filter_7__u_filter_filter_q_reg_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1122 (.o(net1122));
 b15tilo00an1n03x5 gen_filter_7__u_filter_filter_q_reg_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1123 (.o(net1123));
 b15tilo00an1n03x5 gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_diff_ctr_q_reg_3__1124 (.o(net1124));
 b15tilo00an1n03x5 gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_diff_ctr_q_reg_3__1125 (.o(net1125));
 b15tilo00an1n03x5 gen_filter_7__u_filter_stored_value_q_reg_1126 (.o(net1126));
 b15tilo00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_0__gen_filter_8__u_filter_diff_ctr_q_reg_1__1127 (.o(net1127));
 b15tilo00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_0__gen_filter_8__u_filter_diff_ctr_q_reg_1__1128 (.o(net1128));
 b15tilo00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_2__gen_filter_8__u_filter_diff_ctr_q_reg_3__1129 (.o(net1129));
 b15tilo00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_2__gen_filter_8__u_filter_diff_ctr_q_reg_3__1130 (.o(net1130));
 b15tilo00an1n03x5 gen_filter_8__u_filter_filter_q_reg_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1131 (.o(net1131));
 b15tilo00an1n03x5 gen_filter_8__u_filter_filter_q_reg_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1132 (.o(net1132));
 b15tilo00an1n03x5 gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_diff_ctr_q_reg_0__1133 (.o(net1133));
 b15tilo00an1n03x5 gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_diff_ctr_q_reg_0__1134 (.o(net1134));
 b15tilo00an1n03x5 gen_filter_8__u_filter_stored_value_q_reg_1135 (.o(net1135));
 b15tilo00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_1__gen_filter_9__u_filter_diff_ctr_q_reg_2__1136 (.o(net1136));
 b15tilo00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_1__gen_filter_9__u_filter_diff_ctr_q_reg_2__1137 (.o(net1137));
 b15tilo00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_3__gen_filter_9__u_filter_filter_q_reg_1138 (.o(net1138));
 b15tilo00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_3__gen_filter_9__u_filter_filter_q_reg_1139 (.o(net1139));
 b15tilo00an1n03x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_1__1140 (.o(net1140));
 b15tilo00an1n03x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_1__1141 (.o(net1141));
 b15tilo00an1n03x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1142 (.o(net1142));
 b15tilo00an1n03x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1143 (.o(net1143));
 b15tilo00an1n03x5 gen_filter_9__u_filter_stored_value_q_reg_1144 (.o(net1144));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_10__intr_hw_intr_o_reg_11__1145 (.o(net1145));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_10__intr_hw_intr_o_reg_11__1146 (.o(net1146));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_12__intr_hw_intr_o_reg_13__1147 (.o(net1147));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_12__intr_hw_intr_o_reg_13__1148 (.o(net1148));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_14__intr_hw_intr_o_reg_15__1149 (.o(net1149));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_14__intr_hw_intr_o_reg_15__1150 (.o(net1150));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_16__intr_hw_intr_o_reg_17__1151 (.o(net1151));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_16__intr_hw_intr_o_reg_17__1152 (.o(net1152));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_19__intr_hw_intr_o_reg_20__1153 (.o(net1153));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_19__intr_hw_intr_o_reg_20__1154 (.o(net1154));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_1__intr_hw_intr_o_reg_2__1155 (.o(net1155));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_1__intr_hw_intr_o_reg_2__1156 (.o(net1156));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_21__intr_hw_intr_o_reg_30__1157 (.o(net1157));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_21__intr_hw_intr_o_reg_30__1158 (.o(net1158));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_22__intr_hw_intr_o_reg_23__1159 (.o(net1159));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_22__intr_hw_intr_o_reg_23__1160 (.o(net1160));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_24__intr_hw_intr_o_reg_25__1161 (.o(net1161));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_24__intr_hw_intr_o_reg_25__1162 (.o(net1162));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_26__intr_hw_intr_o_reg_27__1163 (.o(net1163));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_26__intr_hw_intr_o_reg_27__1164 (.o(net1164));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_28__intr_hw_intr_o_reg_29__1165 (.o(net1165));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_28__intr_hw_intr_o_reg_29__1166 (.o(net1166));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_31__u_reg_u_data_in_q_reg_3__1167 (.o(net1167));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_31__u_reg_u_data_in_q_reg_3__1168 (.o(net1168));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_4__intr_hw_intr_o_reg_5__1169 (.o(net1169));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_4__intr_hw_intr_o_reg_5__1170 (.o(net1170));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_6__intr_hw_intr_o_reg_7__1171 (.o(net1171));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_6__intr_hw_intr_o_reg_7__1172 (.o(net1172));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_8__intr_hw_intr_o_reg_18__1173 (.o(net1173));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_8__intr_hw_intr_o_reg_18__1174 (.o(net1174));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_9__u_reg_u_data_in_q_reg_5__1175 (.o(net1175));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_9__u_reg_u_data_in_q_reg_5__1176 (.o(net1176));
 b15tilo00an1n03x5 u_reg_err_q_reg_u_reg_u_data_in_q_reg_6__1177 (.o(net1177));
 b15tilo00an1n03x5 u_reg_err_q_reg_u_reg_u_data_in_q_reg_6__1178 (.o(net1178));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_0_latch_1179 (.o(net1179));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_latch_1180 (.o(net1180));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_0__u_reg_u_ctrl_en_input_filter_q_reg_1__1181 (.o(net1181));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_0__u_reg_u_ctrl_en_input_filter_q_reg_1__1182 (.o(net1182));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_10__u_reg_u_ctrl_en_input_filter_q_reg_11__1183 (.o(net1183));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_10__u_reg_u_ctrl_en_input_filter_q_reg_11__1184 (.o(net1184));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_12__u_reg_u_ctrl_en_input_filter_q_reg_13__1185 (.o(net1185));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_12__u_reg_u_ctrl_en_input_filter_q_reg_13__1186 (.o(net1186));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_14__u_reg_u_ctrl_en_input_filter_q_reg_15__1187 (.o(net1187));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_14__u_reg_u_ctrl_en_input_filter_q_reg_15__1188 (.o(net1188));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_16__u_reg_u_ctrl_en_input_filter_q_reg_17__1189 (.o(net1189));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_16__u_reg_u_ctrl_en_input_filter_q_reg_17__1190 (.o(net1190));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_18__u_reg_u_ctrl_en_input_filter_q_reg_19__1191 (.o(net1191));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_18__u_reg_u_ctrl_en_input_filter_q_reg_19__1192 (.o(net1192));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_20__u_reg_u_ctrl_en_input_filter_q_reg_21__1193 (.o(net1193));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_20__u_reg_u_ctrl_en_input_filter_q_reg_21__1194 (.o(net1194));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_22__u_reg_u_ctrl_en_input_filter_q_reg_23__1195 (.o(net1195));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_22__u_reg_u_ctrl_en_input_filter_q_reg_23__1196 (.o(net1196));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_24__u_reg_u_ctrl_en_input_filter_q_reg_25__1197 (.o(net1197));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_24__u_reg_u_ctrl_en_input_filter_q_reg_25__1198 (.o(net1198));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_26__u_reg_u_ctrl_en_input_filter_q_reg_27__1199 (.o(net1199));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_26__u_reg_u_ctrl_en_input_filter_q_reg_27__1200 (.o(net1200));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_28__u_reg_u_ctrl_en_input_filter_q_reg_29__1201 (.o(net1201));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_28__u_reg_u_ctrl_en_input_filter_q_reg_29__1202 (.o(net1202));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_2__u_reg_u_ctrl_en_input_filter_q_reg_3__1203 (.o(net1203));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_2__u_reg_u_ctrl_en_input_filter_q_reg_3__1204 (.o(net1204));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_30__u_reg_u_ctrl_en_input_filter_q_reg_31__1205 (.o(net1205));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_30__u_reg_u_ctrl_en_input_filter_q_reg_31__1206 (.o(net1206));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_4__u_reg_u_ctrl_en_input_filter_q_reg_5__1207 (.o(net1207));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_4__u_reg_u_ctrl_en_input_filter_q_reg_5__1208 (.o(net1208));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_6__u_reg_u_ctrl_en_input_filter_q_reg_7__1209 (.o(net1209));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_6__u_reg_u_ctrl_en_input_filter_q_reg_7__1210 (.o(net1210));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_8__u_reg_u_ctrl_en_input_filter_q_reg_9__1211 (.o(net1211));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_8__u_reg_u_ctrl_en_input_filter_q_reg_9__1212 (.o(net1212));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_0__u_reg_u_data_in_q_reg_1__1213 (.o(net1213));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_0__u_reg_u_data_in_q_reg_1__1214 (.o(net1214));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_11__u_reg_u_data_in_q_reg_16__1215 (.o(net1215));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_11__u_reg_u_data_in_q_reg_16__1216 (.o(net1216));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_12__u_reg_u_data_in_q_reg_17__1217 (.o(net1217));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_12__u_reg_u_data_in_q_reg_17__1218 (.o(net1218));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_13__u_reg_u_data_in_q_reg_14__1219 (.o(net1219));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_13__u_reg_u_data_in_q_reg_14__1220 (.o(net1220));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_18__u_reg_u_data_in_q_reg_19__1221 (.o(net1221));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_18__u_reg_u_data_in_q_reg_19__1222 (.o(net1222));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_20__u_reg_u_data_in_q_reg_21__1223 (.o(net1223));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_20__u_reg_u_data_in_q_reg_21__1224 (.o(net1224));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_22__u_reg_u_data_in_q_reg_23__1225 (.o(net1225));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_22__u_reg_u_data_in_q_reg_23__1226 (.o(net1226));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_24__u_reg_u_data_in_q_reg_25__1227 (.o(net1227));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_24__u_reg_u_data_in_q_reg_25__1228 (.o(net1228));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_26__u_reg_u_reg_if_rspop_q_reg_1__1229 (.o(net1229));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_26__u_reg_u_reg_if_rspop_q_reg_1__1230 (.o(net1230));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_27__1231 (.o(net1231));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_28__u_reg_u_data_in_q_reg_29__1232 (.o(net1232));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_28__u_reg_u_data_in_q_reg_29__1233 (.o(net1233));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_2__u_reg_u_data_in_q_reg_8__1234 (.o(net1234));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_2__u_reg_u_data_in_q_reg_8__1235 (.o(net1235));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_30__u_reg_u_reg_if_rspop_q_reg_2__1236 (.o(net1236));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_30__u_reg_u_reg_if_rspop_q_reg_2__1237 (.o(net1237));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_4__u_reg_u_data_in_q_reg_10__1238 (.o(net1238));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_4__u_reg_u_data_in_q_reg_10__1239 (.o(net1239));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_7__u_reg_u_data_in_q_reg_31__1240 (.o(net1240));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_7__u_reg_u_data_in_q_reg_31__1241 (.o(net1241));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_9__u_reg_u_data_in_q_reg_15__1242 (.o(net1242));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_9__u_reg_u_data_in_q_reg_15__1243 (.o(net1243));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_0_latch_1244 (.o(net1244));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_latch_1245 (.o(net1245));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_0__u_reg_u_intr_ctrl_en_falling_q_reg_1__1246 (.o(net1246));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_0__u_reg_u_intr_ctrl_en_falling_q_reg_1__1247 (.o(net1247));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_10__u_reg_u_intr_ctrl_en_falling_q_reg_11__1248 (.o(net1248));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_10__u_reg_u_intr_ctrl_en_falling_q_reg_11__1249 (.o(net1249));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_12__u_reg_u_intr_ctrl_en_falling_q_reg_13__1250 (.o(net1250));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_12__u_reg_u_intr_ctrl_en_falling_q_reg_13__1251 (.o(net1251));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_14__u_reg_u_intr_ctrl_en_falling_q_reg_15__1252 (.o(net1252));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_14__u_reg_u_intr_ctrl_en_falling_q_reg_15__1253 (.o(net1253));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_16__u_reg_u_intr_ctrl_en_falling_q_reg_17__1254 (.o(net1254));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_16__u_reg_u_intr_ctrl_en_falling_q_reg_17__1255 (.o(net1255));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_18__u_reg_u_intr_ctrl_en_falling_q_reg_19__1256 (.o(net1256));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_18__u_reg_u_intr_ctrl_en_falling_q_reg_19__1257 (.o(net1257));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_20__u_reg_u_intr_ctrl_en_falling_q_reg_21__1258 (.o(net1258));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_20__u_reg_u_intr_ctrl_en_falling_q_reg_21__1259 (.o(net1259));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_22__u_reg_u_intr_ctrl_en_falling_q_reg_23__1260 (.o(net1260));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_22__u_reg_u_intr_ctrl_en_falling_q_reg_23__1261 (.o(net1261));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_24__u_reg_u_intr_ctrl_en_falling_q_reg_25__1262 (.o(net1262));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_24__u_reg_u_intr_ctrl_en_falling_q_reg_25__1263 (.o(net1263));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_26__u_reg_u_intr_ctrl_en_falling_q_reg_27__1264 (.o(net1264));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_26__u_reg_u_intr_ctrl_en_falling_q_reg_27__1265 (.o(net1265));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_28__u_reg_u_intr_ctrl_en_falling_q_reg_29__1266 (.o(net1266));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_28__u_reg_u_intr_ctrl_en_falling_q_reg_29__1267 (.o(net1267));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_2__u_reg_u_intr_ctrl_en_falling_q_reg_3__1268 (.o(net1268));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_2__u_reg_u_intr_ctrl_en_falling_q_reg_3__1269 (.o(net1269));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_30__u_reg_u_intr_ctrl_en_falling_q_reg_31__1270 (.o(net1270));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_30__u_reg_u_intr_ctrl_en_falling_q_reg_31__1271 (.o(net1271));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_4__u_reg_u_intr_ctrl_en_falling_q_reg_5__1272 (.o(net1272));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_4__u_reg_u_intr_ctrl_en_falling_q_reg_5__1273 (.o(net1273));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_6__u_reg_u_intr_ctrl_en_falling_q_reg_7__1274 (.o(net1274));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_6__u_reg_u_intr_ctrl_en_falling_q_reg_7__1275 (.o(net1275));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_8__u_reg_u_intr_ctrl_en_falling_q_reg_9__1276 (.o(net1276));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_8__u_reg_u_intr_ctrl_en_falling_q_reg_9__1277 (.o(net1277));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_0_latch_1278 (.o(net1278));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_latch_1279 (.o(net1279));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1__1280 (.o(net1280));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1__1281 (.o(net1281));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11__1282 (.o(net1282));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11__1283 (.o(net1283));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13__1284 (.o(net1284));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13__1285 (.o(net1285));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15__1286 (.o(net1286));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15__1287 (.o(net1287));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17__1288 (.o(net1288));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17__1289 (.o(net1289));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19__1290 (.o(net1290));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19__1291 (.o(net1291));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21__1292 (.o(net1292));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21__1293 (.o(net1293));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23__1294 (.o(net1294));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23__1295 (.o(net1295));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25__1296 (.o(net1296));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25__1297 (.o(net1297));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27__1298 (.o(net1298));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27__1299 (.o(net1299));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29__1300 (.o(net1300));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29__1301 (.o(net1301));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3__1302 (.o(net1302));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3__1303 (.o(net1303));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31__1304 (.o(net1304));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31__1305 (.o(net1305));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5__1306 (.o(net1306));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5__1307 (.o(net1307));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7__1308 (.o(net1308));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7__1309 (.o(net1309));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9__1310 (.o(net1310));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9__1311 (.o(net1311));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_0_latch_1312 (.o(net1312));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_latch_1313 (.o(net1313));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_reg_u_intr_ctrl_en_lvllow_q_reg_1__1314 (.o(net1314));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_reg_u_intr_ctrl_en_lvllow_q_reg_1__1315 (.o(net1315));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_reg_u_intr_ctrl_en_lvllow_q_reg_11__1316 (.o(net1316));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_reg_u_intr_ctrl_en_lvllow_q_reg_11__1317 (.o(net1317));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_reg_u_intr_ctrl_en_lvllow_q_reg_13__1318 (.o(net1318));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_reg_u_intr_ctrl_en_lvllow_q_reg_13__1319 (.o(net1319));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_reg_u_intr_ctrl_en_lvllow_q_reg_15__1320 (.o(net1320));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_reg_u_intr_ctrl_en_lvllow_q_reg_15__1321 (.o(net1321));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_reg_u_intr_ctrl_en_lvllow_q_reg_17__1322 (.o(net1322));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_reg_u_intr_ctrl_en_lvllow_q_reg_17__1323 (.o(net1323));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_reg_u_intr_ctrl_en_lvllow_q_reg_19__1324 (.o(net1324));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_reg_u_intr_ctrl_en_lvllow_q_reg_19__1325 (.o(net1325));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_reg_u_intr_ctrl_en_lvllow_q_reg_21__1326 (.o(net1326));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_reg_u_intr_ctrl_en_lvllow_q_reg_21__1327 (.o(net1327));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_reg_u_intr_ctrl_en_lvllow_q_reg_23__1328 (.o(net1328));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_reg_u_intr_ctrl_en_lvllow_q_reg_23__1329 (.o(net1329));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_reg_u_intr_ctrl_en_lvllow_q_reg_25__1330 (.o(net1330));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_reg_u_intr_ctrl_en_lvllow_q_reg_25__1331 (.o(net1331));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_reg_u_intr_ctrl_en_lvllow_q_reg_27__1332 (.o(net1332));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_reg_u_intr_ctrl_en_lvllow_q_reg_27__1333 (.o(net1333));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_reg_u_intr_ctrl_en_lvllow_q_reg_29__1334 (.o(net1334));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_reg_u_intr_ctrl_en_lvllow_q_reg_29__1335 (.o(net1335));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_reg_u_intr_ctrl_en_lvllow_q_reg_3__1336 (.o(net1336));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_reg_u_intr_ctrl_en_lvllow_q_reg_3__1337 (.o(net1337));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_reg_u_intr_ctrl_en_lvllow_q_reg_31__1338 (.o(net1338));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_reg_u_intr_ctrl_en_lvllow_q_reg_31__1339 (.o(net1339));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_reg_u_intr_ctrl_en_lvllow_q_reg_5__1340 (.o(net1340));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_reg_u_intr_ctrl_en_lvllow_q_reg_5__1341 (.o(net1341));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_reg_u_intr_ctrl_en_lvllow_q_reg_7__1342 (.o(net1342));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_reg_u_intr_ctrl_en_lvllow_q_reg_7__1343 (.o(net1343));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_reg_u_intr_ctrl_en_lvllow_q_reg_9__1344 (.o(net1344));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_reg_u_intr_ctrl_en_lvllow_q_reg_9__1345 (.o(net1345));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_0_latch_1346 (.o(net1346));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_latch_1347 (.o(net1347));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_0__u_reg_u_intr_ctrl_en_rising_q_reg_1__1348 (.o(net1348));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_0__u_reg_u_intr_ctrl_en_rising_q_reg_1__1349 (.o(net1349));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_10__u_reg_u_intr_ctrl_en_rising_q_reg_11__1350 (.o(net1350));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_10__u_reg_u_intr_ctrl_en_rising_q_reg_11__1351 (.o(net1351));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_12__u_reg_u_intr_ctrl_en_rising_q_reg_13__1352 (.o(net1352));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_12__u_reg_u_intr_ctrl_en_rising_q_reg_13__1353 (.o(net1353));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_14__u_reg_u_intr_ctrl_en_rising_q_reg_15__1354 (.o(net1354));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_14__u_reg_u_intr_ctrl_en_rising_q_reg_15__1355 (.o(net1355));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_16__u_reg_u_intr_ctrl_en_rising_q_reg_17__1356 (.o(net1356));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_16__u_reg_u_intr_ctrl_en_rising_q_reg_17__1357 (.o(net1357));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_18__u_reg_u_intr_ctrl_en_rising_q_reg_19__1358 (.o(net1358));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_18__u_reg_u_intr_ctrl_en_rising_q_reg_19__1359 (.o(net1359));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_20__u_reg_u_intr_ctrl_en_rising_q_reg_21__1360 (.o(net1360));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_20__u_reg_u_intr_ctrl_en_rising_q_reg_21__1361 (.o(net1361));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_22__u_reg_u_intr_ctrl_en_rising_q_reg_23__1362 (.o(net1362));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_22__u_reg_u_intr_ctrl_en_rising_q_reg_23__1363 (.o(net1363));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_24__u_reg_u_intr_ctrl_en_rising_q_reg_25__1364 (.o(net1364));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_24__u_reg_u_intr_ctrl_en_rising_q_reg_25__1365 (.o(net1365));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_26__u_reg_u_intr_ctrl_en_rising_q_reg_27__1366 (.o(net1366));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_26__u_reg_u_intr_ctrl_en_rising_q_reg_27__1367 (.o(net1367));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_28__u_reg_u_intr_ctrl_en_rising_q_reg_29__1368 (.o(net1368));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_28__u_reg_u_intr_ctrl_en_rising_q_reg_29__1369 (.o(net1369));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_2__u_reg_u_intr_ctrl_en_rising_q_reg_3__1370 (.o(net1370));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_2__u_reg_u_intr_ctrl_en_rising_q_reg_3__1371 (.o(net1371));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_30__u_reg_u_intr_ctrl_en_rising_q_reg_31__1372 (.o(net1372));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_30__u_reg_u_intr_ctrl_en_rising_q_reg_31__1373 (.o(net1373));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_4__u_reg_u_intr_ctrl_en_rising_q_reg_5__1374 (.o(net1374));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_4__u_reg_u_intr_ctrl_en_rising_q_reg_5__1375 (.o(net1375));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_6__u_reg_u_intr_ctrl_en_rising_q_reg_7__1376 (.o(net1376));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_6__u_reg_u_intr_ctrl_en_rising_q_reg_7__1377 (.o(net1377));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_8__u_reg_u_intr_ctrl_en_rising_q_reg_9__1378 (.o(net1378));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_8__u_reg_u_intr_ctrl_en_rising_q_reg_9__1379 (.o(net1379));
 b15tilo00an1n03x5 u_reg_u_intr_enable_clk_gate_q_reg_0_latch_1380 (.o(net1380));
 b15tilo00an1n03x5 u_reg_u_intr_enable_clk_gate_q_reg_latch_1381 (.o(net1381));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_0__u_reg_u_intr_enable_q_reg_1__1382 (.o(net1382));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_0__u_reg_u_intr_enable_q_reg_1__1383 (.o(net1383));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_10__u_reg_u_intr_enable_q_reg_11__1384 (.o(net1384));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_10__u_reg_u_intr_enable_q_reg_11__1385 (.o(net1385));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_12__u_reg_u_intr_enable_q_reg_13__1386 (.o(net1386));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_12__u_reg_u_intr_enable_q_reg_13__1387 (.o(net1387));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_14__u_reg_u_intr_enable_q_reg_15__1388 (.o(net1388));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_14__u_reg_u_intr_enable_q_reg_15__1389 (.o(net1389));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_16__u_reg_u_intr_enable_q_reg_17__1390 (.o(net1390));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_16__u_reg_u_intr_enable_q_reg_17__1391 (.o(net1391));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_18__u_reg_u_intr_enable_q_reg_19__1392 (.o(net1392));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_18__u_reg_u_intr_enable_q_reg_19__1393 (.o(net1393));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_20__u_reg_u_intr_enable_q_reg_21__1394 (.o(net1394));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_20__u_reg_u_intr_enable_q_reg_21__1395 (.o(net1395));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_22__u_reg_u_intr_enable_q_reg_23__1396 (.o(net1396));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_22__u_reg_u_intr_enable_q_reg_23__1397 (.o(net1397));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_24__u_reg_u_intr_enable_q_reg_25__1398 (.o(net1398));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_24__u_reg_u_intr_enable_q_reg_25__1399 (.o(net1399));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_26__u_reg_u_intr_enable_q_reg_27__1400 (.o(net1400));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_26__u_reg_u_intr_enable_q_reg_27__1401 (.o(net1401));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_28__u_reg_u_intr_enable_q_reg_29__1402 (.o(net1402));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_28__u_reg_u_intr_enable_q_reg_29__1403 (.o(net1403));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_2__u_reg_u_intr_enable_q_reg_3__1404 (.o(net1404));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_2__u_reg_u_intr_enable_q_reg_3__1405 (.o(net1405));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_30__u_reg_u_intr_enable_q_reg_31__1406 (.o(net1406));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_30__u_reg_u_intr_enable_q_reg_31__1407 (.o(net1407));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_4__u_reg_u_intr_enable_q_reg_5__1408 (.o(net1408));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_4__u_reg_u_intr_enable_q_reg_5__1409 (.o(net1409));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_6__u_reg_u_intr_enable_q_reg_7__1410 (.o(net1410));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_6__u_reg_u_intr_enable_q_reg_7__1411 (.o(net1411));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_8__u_reg_u_intr_enable_q_reg_9__1412 (.o(net1412));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_8__u_reg_u_intr_enable_q_reg_9__1413 (.o(net1413));
 b15tilo00an1n03x5 u_reg_u_intr_state_clk_gate_q_reg_0_latch_1414 (.o(net1414));
 b15tilo00an1n03x5 u_reg_u_intr_state_clk_gate_q_reg_latch_1415 (.o(net1415));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_0__u_reg_u_intr_state_q_reg_1__1416 (.o(net1416));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_0__u_reg_u_intr_state_q_reg_1__1417 (.o(net1417));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_10__u_reg_u_intr_state_q_reg_11__1418 (.o(net1418));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_10__u_reg_u_intr_state_q_reg_11__1419 (.o(net1419));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_12__u_reg_u_intr_state_q_reg_13__1420 (.o(net1420));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_12__u_reg_u_intr_state_q_reg_13__1421 (.o(net1421));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_14__u_reg_u_intr_state_q_reg_15__1422 (.o(net1422));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_14__u_reg_u_intr_state_q_reg_15__1423 (.o(net1423));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_16__u_reg_u_intr_state_q_reg_17__1424 (.o(net1424));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_16__u_reg_u_intr_state_q_reg_17__1425 (.o(net1425));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_18__u_reg_u_intr_state_q_reg_19__1426 (.o(net1426));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_18__u_reg_u_intr_state_q_reg_19__1427 (.o(net1427));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_20__u_reg_u_intr_state_q_reg_21__1428 (.o(net1428));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_20__u_reg_u_intr_state_q_reg_21__1429 (.o(net1429));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_22__u_reg_u_intr_state_q_reg_23__1430 (.o(net1430));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_22__u_reg_u_intr_state_q_reg_23__1431 (.o(net1431));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_24__u_reg_u_intr_state_q_reg_25__1432 (.o(net1432));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_24__u_reg_u_intr_state_q_reg_25__1433 (.o(net1433));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_26__u_reg_u_intr_state_q_reg_27__1434 (.o(net1434));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_26__u_reg_u_intr_state_q_reg_27__1435 (.o(net1435));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_28__u_reg_u_intr_state_q_reg_29__1436 (.o(net1436));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_28__u_reg_u_intr_state_q_reg_29__1437 (.o(net1437));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_2__u_reg_u_intr_state_q_reg_3__1438 (.o(net1438));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_2__u_reg_u_intr_state_q_reg_3__1439 (.o(net1439));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_30__u_reg_u_intr_state_q_reg_31__1440 (.o(net1440));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_30__u_reg_u_intr_state_q_reg_31__1441 (.o(net1441));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_4__u_reg_u_intr_state_q_reg_5__1442 (.o(net1442));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_4__u_reg_u_intr_state_q_reg_5__1443 (.o(net1443));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_6__u_reg_u_intr_state_q_reg_7__1444 (.o(net1444));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_6__u_reg_u_intr_state_q_reg_7__1445 (.o(net1445));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_8__u_reg_u_intr_state_q_reg_9__1446 (.o(net1446));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_8__u_reg_u_intr_state_q_reg_9__1447 (.o(net1447));
 b15tilo00an1n03x5 u_reg_u_reg_if_clk_gate_rdata_q_reg_0_latch_1448 (.o(net1448));
 b15tilo00an1n03x5 u_reg_u_reg_if_clk_gate_rdata_q_reg_latch_1449 (.o(net1449));
 b15tilo00an1n03x5 u_reg_u_reg_if_clk_gate_reqid_q_reg_latch_1450 (.o(net1450));
 b15tilo00an1n03x5 u_reg_u_reg_if_error_q_reg_1451 (.o(net1451));
 b15tilo00an1n03x5 u_reg_u_reg_if_outstanding_q_reg_1452 (.o(net1452));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_0__u_reg_u_reg_if_rdata_q_reg_1__1453 (.o(net1453));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_0__u_reg_u_reg_if_rdata_q_reg_1__1454 (.o(net1454));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_10__u_reg_u_reg_if_rdata_q_reg_11__1455 (.o(net1455));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_10__u_reg_u_reg_if_rdata_q_reg_11__1456 (.o(net1456));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_12__u_reg_u_reg_if_rdata_q_reg_13__1457 (.o(net1457));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_12__u_reg_u_reg_if_rdata_q_reg_13__1458 (.o(net1458));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_14__u_reg_u_reg_if_rdata_q_reg_15__1459 (.o(net1459));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_14__u_reg_u_reg_if_rdata_q_reg_15__1460 (.o(net1460));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_16__u_reg_u_reg_if_rdata_q_reg_17__1461 (.o(net1461));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_16__u_reg_u_reg_if_rdata_q_reg_17__1462 (.o(net1462));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_18__u_reg_u_reg_if_rdata_q_reg_19__1463 (.o(net1463));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_18__u_reg_u_reg_if_rdata_q_reg_19__1464 (.o(net1464));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_20__u_reg_u_reg_if_rdata_q_reg_21__1465 (.o(net1465));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_20__u_reg_u_reg_if_rdata_q_reg_21__1466 (.o(net1466));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_22__u_reg_u_reg_if_rdata_q_reg_23__1467 (.o(net1467));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_22__u_reg_u_reg_if_rdata_q_reg_23__1468 (.o(net1468));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_24__u_reg_u_reg_if_rdata_q_reg_25__1469 (.o(net1469));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_24__u_reg_u_reg_if_rdata_q_reg_25__1470 (.o(net1470));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_26__u_reg_u_reg_if_rdata_q_reg_27__1471 (.o(net1471));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_26__u_reg_u_reg_if_rdata_q_reg_27__1472 (.o(net1472));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_28__u_reg_u_reg_if_rdata_q_reg_29__1473 (.o(net1473));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_28__u_reg_u_reg_if_rdata_q_reg_29__1474 (.o(net1474));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_2__u_reg_u_reg_if_rdata_q_reg_3__1475 (.o(net1475));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_2__u_reg_u_reg_if_rdata_q_reg_3__1476 (.o(net1476));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_30__u_reg_u_reg_if_rdata_q_reg_31__1477 (.o(net1477));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_30__u_reg_u_reg_if_rdata_q_reg_31__1478 (.o(net1478));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_4__u_reg_u_reg_if_rdata_q_reg_5__1479 (.o(net1479));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_4__u_reg_u_reg_if_rdata_q_reg_5__1480 (.o(net1480));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_6__u_reg_u_reg_if_rdata_q_reg_7__1481 (.o(net1481));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_6__u_reg_u_reg_if_rdata_q_reg_7__1482 (.o(net1482));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_8__u_reg_u_reg_if_rdata_q_reg_9__1483 (.o(net1483));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_q_reg_8__u_reg_u_reg_if_rdata_q_reg_9__1484 (.o(net1484));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_q_reg_0__u_reg_u_reg_if_reqid_q_reg_1__1485 (.o(net1485));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_q_reg_0__u_reg_u_reg_if_reqid_q_reg_1__1486 (.o(net1486));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_q_reg_2__u_reg_u_reg_if_reqid_q_reg_3__1487 (.o(net1487));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_q_reg_2__u_reg_u_reg_if_reqid_q_reg_3__1488 (.o(net1488));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_q_reg_4__u_reg_u_reg_if_reqid_q_reg_5__1489 (.o(net1489));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_q_reg_4__u_reg_u_reg_if_reqid_q_reg_5__1490 (.o(net1490));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_q_reg_6__u_reg_u_reg_if_reqid_q_reg_7__1491 (.o(net1491));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_q_reg_6__u_reg_u_reg_if_reqid_q_reg_7__1492 (.o(net1492));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqsz_q_reg_0__1493 (.o(net1493));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqsz_q_reg_1__1494 (.o(net1494));
 b15tilo00an1n03x5 u_reg_u_reg_if_rspop_q_reg_0__1495 (.o(net1495));
 b15tihi00an1n03x5 U3362_1497 (.o(net1497));
 b15tihi00an1n03x5 U3364_1498 (.o(net1498));
 b15tihi00an1n03x5 U3366_1499 (.o(net1499));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_0__cio_gpio_en_q_reg_1__1500 (.o(net1500));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_10__cio_gpio_en_q_reg_11__1501 (.o(net1501));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_12__cio_gpio_en_q_reg_13__1502 (.o(net1502));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_14__cio_gpio_en_q_reg_15__1503 (.o(net1503));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_16__cio_gpio_en_q_reg_17__1504 (.o(net1504));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_18__cio_gpio_en_q_reg_19__1505 (.o(net1505));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_20__cio_gpio_en_q_reg_21__1506 (.o(net1506));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_22__cio_gpio_en_q_reg_23__1507 (.o(net1507));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_24__cio_gpio_en_q_reg_25__1508 (.o(net1508));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_26__cio_gpio_en_q_reg_27__1509 (.o(net1509));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_28__cio_gpio_en_q_reg_29__1510 (.o(net1510));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_2__cio_gpio_en_q_reg_3__1511 (.o(net1511));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_30__cio_gpio_en_q_reg_31__1512 (.o(net1512));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_4__cio_gpio_en_q_reg_5__1513 (.o(net1513));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_6__cio_gpio_en_q_reg_7__1514 (.o(net1514));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_8__cio_gpio_en_q_reg_9__1515 (.o(net1515));
 b15tihi00an1n03x5 cio_gpio_q_reg_0__cio_gpio_q_reg_1__1516 (.o(net1516));
 b15tihi00an1n03x5 cio_gpio_q_reg_10__cio_gpio_q_reg_11__1517 (.o(net1517));
 b15tihi00an1n03x5 cio_gpio_q_reg_12__cio_gpio_q_reg_13__1518 (.o(net1518));
 b15tihi00an1n03x5 cio_gpio_q_reg_14__cio_gpio_q_reg_15__1519 (.o(net1519));
 b15tihi00an1n03x5 cio_gpio_q_reg_16__cio_gpio_q_reg_17__1520 (.o(net1520));
 b15tihi00an1n03x5 cio_gpio_q_reg_18__cio_gpio_q_reg_19__1521 (.o(net1521));
 b15tihi00an1n03x5 cio_gpio_q_reg_20__cio_gpio_q_reg_21__1522 (.o(net1522));
 b15tihi00an1n03x5 cio_gpio_q_reg_22__cio_gpio_q_reg_23__1523 (.o(net1523));
 b15tihi00an1n03x5 cio_gpio_q_reg_24__cio_gpio_q_reg_25__1524 (.o(net1524));
 b15tihi00an1n03x5 cio_gpio_q_reg_26__cio_gpio_q_reg_27__1525 (.o(net1525));
 b15tihi00an1n03x5 cio_gpio_q_reg_28__cio_gpio_q_reg_29__1526 (.o(net1526));
 b15tihi00an1n03x5 cio_gpio_q_reg_2__cio_gpio_q_reg_3__1527 (.o(net1527));
 b15tihi00an1n03x5 cio_gpio_q_reg_30__cio_gpio_q_reg_31__1528 (.o(net1528));
 b15tihi00an1n03x5 cio_gpio_q_reg_4__cio_gpio_q_reg_5__1529 (.o(net1529));
 b15tihi00an1n03x5 cio_gpio_q_reg_6__cio_gpio_q_reg_7__1530 (.o(net1530));
 b15tihi00an1n03x5 cio_gpio_q_reg_8__cio_gpio_q_reg_9__1531 (.o(net1531));
 b15tihi00an1n03x5 data_in_q_reg_0__data_in_q_reg_1__1532 (.o(net1532));
 b15tihi00an1n03x5 data_in_q_reg_10__data_in_q_reg_11__1533 (.o(net1533));
 b15tihi00an1n03x5 data_in_q_reg_12__data_in_q_reg_13__1534 (.o(net1534));
 b15tihi00an1n03x5 data_in_q_reg_14__data_in_q_reg_15__1535 (.o(net1535));
 b15tihi00an1n03x5 data_in_q_reg_16__data_in_q_reg_17__1536 (.o(net1536));
 b15tihi00an1n03x5 data_in_q_reg_18__data_in_q_reg_19__1537 (.o(net1537));
 b15tihi00an1n03x5 data_in_q_reg_20__data_in_q_reg_21__1538 (.o(net1538));
 b15tihi00an1n03x5 data_in_q_reg_22__data_in_q_reg_23__1539 (.o(net1539));
 b15tihi00an1n03x5 data_in_q_reg_24__data_in_q_reg_25__1540 (.o(net1540));
 b15tihi00an1n03x5 data_in_q_reg_26__data_in_q_reg_27__1541 (.o(net1541));
 b15tihi00an1n03x5 data_in_q_reg_28__data_in_q_reg_29__1542 (.o(net1542));
 b15tihi00an1n03x5 data_in_q_reg_2__data_in_q_reg_3__1543 (.o(net1543));
 b15tihi00an1n03x5 data_in_q_reg_30__data_in_q_reg_31__1544 (.o(net1544));
 b15tihi00an1n03x5 data_in_q_reg_4__data_in_q_reg_5__1545 (.o(net1545));
 b15tihi00an1n03x5 data_in_q_reg_6__data_in_q_reg_7__1546 (.o(net1546));
 b15tihi00an1n03x5 data_in_q_reg_8__data_in_q_reg_9__1547 (.o(net1547));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg_1548 (.o(net1548));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg_1549 (.o(net1549));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0__gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1__1550 (.o(net1550));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1551 (.o(net1551));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq_reg_1552 (.o(net1552));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1553 (.o(net1553));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1554 (.o(net1554));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg_1555 (.o(net1555));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_0__1556 (.o(net1556));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_1__1557 (.o(net1557));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq_reg_1558 (.o(net1558));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1559 (.o(net1559));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1560 (.o(net1560));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1561 (.o(net1561));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg_1562 (.o(net1562));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_0__1563 (.o(net1563));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_1__1564 (.o(net1564));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1565 (.o(net1565));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_1__1566 (.o(net1566));
 b15tihi00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_0__gen_filter_0__u_filter_diff_ctr_q_reg_1__1567 (.o(net1567));
 b15tihi00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_2__gen_filter_0__u_filter_diff_ctr_q_reg_3__1568 (.o(net1568));
 b15tihi00an1n03x5 gen_filter_0__u_filter_filter_q_reg_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1569 (.o(net1569));
 b15tihi00an1n03x5 gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_1__u_filter_diff_ctr_q_reg_0__1570 (.o(net1570));
 b15tihi00an1n03x5 gen_filter_0__u_filter_stored_value_q_reg_1571 (.o(net1571));
 b15tihi00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_1__gen_filter_10__u_filter_diff_ctr_q_reg_2__1572 (.o(net1572));
 b15tihi00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_filter_q_reg_1573 (.o(net1573));
 b15tihi00an1n03x5 gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1574 (.o(net1574));
 b15tihi00an1n03x5 gen_filter_10__u_filter_stored_value_q_reg_1575 (.o(net1575));
 b15tihi00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_0__gen_filter_12__u_filter_diff_ctr_q_reg_0__1576 (.o(net1576));
 b15tihi00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_2__gen_filter_11__u_filter_diff_ctr_q_reg_3__1577 (.o(net1577));
 b15tihi00an1n03x5 gen_filter_11__u_filter_filter_q_reg_gen_filter_12__u_filter_filter_q_reg_1578 (.o(net1578));
 b15tihi00an1n03x5 gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_3__1579 (.o(net1579));
 b15tihi00an1n03x5 gen_filter_11__u_filter_stored_value_q_reg_1580 (.o(net1580));
 b15tihi00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_1__gen_filter_12__u_filter_diff_ctr_q_reg_2__1581 (.o(net1581));
 b15tihi00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_diff_ctr_q_reg_0__1582 (.o(net1582));
 b15tihi00an1n03x5 gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1583 (.o(net1583));
 b15tihi00an1n03x5 gen_filter_12__u_filter_stored_value_q_reg_1584 (.o(net1584));
 b15tihi00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_1__gen_filter_13__u_filter_diff_ctr_q_reg_2__1585 (.o(net1585));
 b15tihi00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_filter_q_reg_1586 (.o(net1586));
 b15tihi00an1n03x5 gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1587 (.o(net1587));
 b15tihi00an1n03x5 gen_filter_13__u_filter_stored_value_q_reg_1588 (.o(net1588));
 b15tihi00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_1__1589 (.o(net1589));
 b15tihi00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_2__gen_filter_26__u_filter_diff_ctr_q_reg_0__1590 (.o(net1590));
 b15tihi00an1n03x5 gen_filter_14__u_filter_filter_q_reg_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1591 (.o(net1591));
 b15tihi00an1n03x5 gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_diff_ctr_q_reg_0__1592 (.o(net1592));
 b15tihi00an1n03x5 gen_filter_14__u_filter_stored_value_q_reg_1593 (.o(net1593));
 b15tihi00an1n03x5 gen_filter_15__u_filter_diff_ctr_q_reg_1__gen_filter_15__u_filter_diff_ctr_q_reg_2__1594 (.o(net1594));
 b15tihi00an1n03x5 gen_filter_15__u_filter_filter_q_reg_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1595 (.o(net1595));
 b15tihi00an1n03x5 gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_diff_ctr_q_reg_0__1596 (.o(net1596));
 b15tihi00an1n03x5 gen_filter_15__u_filter_stored_value_q_reg_1597 (.o(net1597));
 b15tihi00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_0__gen_filter_16__u_filter_diff_ctr_q_reg_1__1598 (.o(net1598));
 b15tihi00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_2__gen_filter_16__u_filter_diff_ctr_q_reg_3__1599 (.o(net1599));
 b15tihi00an1n03x5 gen_filter_16__u_filter_filter_q_reg_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1600 (.o(net1600));
 b15tihi00an1n03x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1601 (.o(net1601));
 b15tihi00an1n03x5 gen_filter_16__u_filter_stored_value_q_reg_1602 (.o(net1602));
 b15tihi00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_1__gen_filter_17__u_filter_diff_ctr_q_reg_2__1603 (.o(net1603));
 b15tihi00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_3__gen_filter_17__u_filter_filter_q_reg_1604 (.o(net1604));
 b15tihi00an1n03x5 gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_18__u_filter_diff_ctr_q_reg_0__1605 (.o(net1605));
 b15tihi00an1n03x5 gen_filter_17__u_filter_stored_value_q_reg_1606 (.o(net1606));
 b15tihi00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_1__gen_filter_18__u_filter_diff_ctr_q_reg_2__1607 (.o(net1607));
 b15tihi00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_3__gen_filter_18__u_filter_filter_q_reg_1608 (.o(net1608));
 b15tihi00an1n03x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1609 (.o(net1609));
 b15tihi00an1n03x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1610 (.o(net1610));
 b15tihi00an1n03x5 gen_filter_18__u_filter_stored_value_q_reg_1611 (.o(net1611));
 b15tihi00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_1__gen_filter_19__u_filter_diff_ctr_q_reg_2__1612 (.o(net1612));
 b15tihi00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_3__gen_filter_19__u_filter_filter_q_reg_1613 (.o(net1613));
 b15tihi00an1n03x5 gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1614 (.o(net1614));
 b15tihi00an1n03x5 gen_filter_19__u_filter_stored_value_q_reg_1615 (.o(net1615));
 b15tihi00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_1__gen_filter_1__u_filter_diff_ctr_q_reg_2__1616 (.o(net1616));
 b15tihi00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_3__gen_filter_1__u_filter_filter_q_reg_1617 (.o(net1617));
 b15tihi00an1n03x5 gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1618 (.o(net1618));
 b15tihi00an1n03x5 gen_filter_1__u_filter_stored_value_q_reg_1619 (.o(net1619));
 b15tihi00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_0__gen_filter_20__u_filter_diff_ctr_q_reg_1__1620 (.o(net1620));
 b15tihi00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_2__gen_filter_20__u_filter_diff_ctr_q_reg_3__1621 (.o(net1621));
 b15tihi00an1n03x5 gen_filter_20__u_filter_filter_q_reg_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1622 (.o(net1622));
 b15tihi00an1n03x5 gen_filter_20__u_filter_stored_value_q_reg_1623 (.o(net1623));
 b15tihi00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_0__gen_filter_21__u_filter_diff_ctr_q_reg_1__1624 (.o(net1624));
 b15tihi00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_2__gen_filter_21__u_filter_diff_ctr_q_reg_3__1625 (.o(net1625));
 b15tihi00an1n03x5 gen_filter_21__u_filter_filter_q_reg_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1626 (.o(net1626));
 b15tihi00an1n03x5 gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_diff_ctr_q_reg_0__1627 (.o(net1627));
 b15tihi00an1n03x5 gen_filter_21__u_filter_stored_value_q_reg_1628 (.o(net1628));
 b15tihi00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_0__gen_filter_22__u_filter_diff_ctr_q_reg_1__1629 (.o(net1629));
 b15tihi00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_2__gen_filter_22__u_filter_diff_ctr_q_reg_3__1630 (.o(net1630));
 b15tihi00an1n03x5 gen_filter_22__u_filter_filter_q_reg_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1631 (.o(net1631));
 b15tihi00an1n03x5 gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_diff_ctr_q_reg_0__1632 (.o(net1632));
 b15tihi00an1n03x5 gen_filter_22__u_filter_stored_value_q_reg_1633 (.o(net1633));
 b15tihi00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_1__gen_filter_23__u_filter_diff_ctr_q_reg_2__1634 (.o(net1634));
 b15tihi00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_3__gen_filter_23__u_filter_filter_q_reg_1635 (.o(net1635));
 b15tihi00an1n03x5 gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1636 (.o(net1636));
 b15tihi00an1n03x5 gen_filter_23__u_filter_stored_value_q_reg_1637 (.o(net1637));
 b15tihi00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_0__gen_filter_24__u_filter_diff_ctr_q_reg_1__1638 (.o(net1638));
 b15tihi00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_2__gen_filter_24__u_filter_diff_ctr_q_reg_3__1639 (.o(net1639));
 b15tihi00an1n03x5 gen_filter_24__u_filter_filter_q_reg_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1640 (.o(net1640));
 b15tihi00an1n03x5 gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_25__u_filter_diff_ctr_q_reg_0__1641 (.o(net1641));
 b15tihi00an1n03x5 gen_filter_24__u_filter_stored_value_q_reg_1642 (.o(net1642));
 b15tihi00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_1__gen_filter_25__u_filter_diff_ctr_q_reg_2__1643 (.o(net1643));
 b15tihi00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_3__gen_filter_25__u_filter_filter_q_reg_1644 (.o(net1644));
 b15tihi00an1n03x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_0__1645 (.o(net1645));
 b15tihi00an1n03x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_27__u_filter_diff_ctr_q_reg_0__1646 (.o(net1646));
 b15tihi00an1n03x5 gen_filter_25__u_filter_stored_value_q_reg_1647 (.o(net1647));
 b15tihi00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_1__gen_filter_26__u_filter_diff_ctr_q_reg_2__1648 (.o(net1648));
 b15tihi00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_3__gen_filter_26__u_filter_filter_q_reg_1649 (.o(net1649));
 b15tihi00an1n03x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1650 (.o(net1650));
 b15tihi00an1n03x5 gen_filter_26__u_filter_stored_value_q_reg_1651 (.o(net1651));
 b15tihi00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_1__gen_filter_27__u_filter_diff_ctr_q_reg_2__1652 (.o(net1652));
 b15tihi00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_3__gen_filter_27__u_filter_filter_q_reg_1653 (.o(net1653));
 b15tihi00an1n03x5 gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1654 (.o(net1654));
 b15tihi00an1n03x5 gen_filter_27__u_filter_stored_value_q_reg_1655 (.o(net1655));
 b15tihi00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_1__gen_filter_28__u_filter_diff_ctr_q_reg_2__1656 (.o(net1656));
 b15tihi00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_3__gen_filter_28__u_filter_filter_q_reg_1657 (.o(net1657));
 b15tihi00an1n03x5 gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1658 (.o(net1658));
 b15tihi00an1n03x5 gen_filter_28__u_filter_stored_value_q_reg_1659 (.o(net1659));
 b15tihi00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_0__gen_filter_29__u_filter_diff_ctr_q_reg_1__1660 (.o(net1660));
 b15tihi00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_2__gen_filter_29__u_filter_diff_ctr_q_reg_3__1661 (.o(net1661));
 b15tihi00an1n03x5 gen_filter_29__u_filter_filter_q_reg_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1662 (.o(net1662));
 b15tihi00an1n03x5 gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1663 (.o(net1663));
 b15tihi00an1n03x5 gen_filter_29__u_filter_stored_value_q_reg_1664 (.o(net1664));
 b15tihi00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_0__gen_filter_2__u_filter_diff_ctr_q_reg_1__1665 (.o(net1665));
 b15tihi00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_2__gen_filter_2__u_filter_diff_ctr_q_reg_3__1666 (.o(net1666));
 b15tihi00an1n03x5 gen_filter_2__u_filter_filter_q_reg_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1667 (.o(net1667));
 b15tihi00an1n03x5 gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1668 (.o(net1668));
 b15tihi00an1n03x5 gen_filter_2__u_filter_stored_value_q_reg_1669 (.o(net1669));
 b15tihi00an1n03x5 gen_filter_30__u_filter_diff_ctr_q_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_1__1670 (.o(net1670));
 b15tihi00an1n03x5 gen_filter_30__u_filter_diff_ctr_q_reg_2__gen_filter_30__u_filter_diff_ctr_q_reg_3__1671 (.o(net1671));
 b15tihi00an1n03x5 gen_filter_30__u_filter_filter_q_reg_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1672 (.o(net1672));
 b15tihi00an1n03x5 gen_filter_30__u_filter_stored_value_q_reg_1673 (.o(net1673));
 b15tihi00an1n03x5 gen_filter_31__u_filter_diff_ctr_q_reg_0__gen_filter_31__u_filter_diff_ctr_q_reg_1__1674 (.o(net1674));
 b15tihi00an1n03x5 gen_filter_31__u_filter_diff_ctr_q_reg_2__gen_filter_31__u_filter_diff_ctr_q_reg_3__1675 (.o(net1675));
 b15tihi00an1n03x5 gen_filter_31__u_filter_filter_q_reg_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1676 (.o(net1676));
 b15tihi00an1n03x5 gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_3__1677 (.o(net1677));
 b15tihi00an1n03x5 gen_filter_31__u_filter_stored_value_q_reg_1678 (.o(net1678));
 b15tihi00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_0__gen_filter_3__u_filter_diff_ctr_q_reg_1__1679 (.o(net1679));
 b15tihi00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_2__gen_filter_3__u_filter_diff_ctr_q_reg_3__1680 (.o(net1680));
 b15tihi00an1n03x5 gen_filter_3__u_filter_filter_q_reg_gen_filter_4__u_filter_diff_ctr_q_reg_0__1681 (.o(net1681));
 b15tihi00an1n03x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1682 (.o(net1682));
 b15tihi00an1n03x5 gen_filter_3__u_filter_stored_value_q_reg_1683 (.o(net1683));
 b15tihi00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_1__gen_filter_4__u_filter_diff_ctr_q_reg_2__1684 (.o(net1684));
 b15tihi00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_diff_ctr_q_reg_0__1685 (.o(net1685));
 b15tihi00an1n03x5 gen_filter_4__u_filter_filter_q_reg_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1686 (.o(net1686));
 b15tihi00an1n03x5 gen_filter_4__u_filter_stored_value_q_reg_1687 (.o(net1687));
 b15tihi00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_0__gen_filter_5__u_filter_diff_ctr_q_reg_1__1688 (.o(net1688));
 b15tihi00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_2__gen_filter_5__u_filter_filter_q_reg_1689 (.o(net1689));
 b15tihi00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_3__gen_filter_6__u_filter_diff_ctr_q_reg_0__1690 (.o(net1690));
 b15tihi00an1n03x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_diff_ctr_q_reg_0__1691 (.o(net1691));
 b15tihi00an1n03x5 gen_filter_5__u_filter_stored_value_q_reg_1692 (.o(net1692));
 b15tihi00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_1__gen_filter_6__u_filter_diff_ctr_q_reg_2__1693 (.o(net1693));
 b15tihi00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_3__gen_filter_6__u_filter_filter_q_reg_1694 (.o(net1694));
 b15tihi00an1n03x5 gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1695 (.o(net1695));
 b15tihi00an1n03x5 gen_filter_6__u_filter_stored_value_q_reg_1696 (.o(net1696));
 b15tihi00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_0__gen_filter_7__u_filter_diff_ctr_q_reg_1__1697 (.o(net1697));
 b15tihi00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_2__gen_filter_7__u_filter_diff_ctr_q_reg_3__1698 (.o(net1698));
 b15tihi00an1n03x5 gen_filter_7__u_filter_filter_q_reg_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1699 (.o(net1699));
 b15tihi00an1n03x5 gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_diff_ctr_q_reg_3__1700 (.o(net1700));
 b15tihi00an1n03x5 gen_filter_7__u_filter_stored_value_q_reg_1701 (.o(net1701));
 b15tihi00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_0__gen_filter_8__u_filter_diff_ctr_q_reg_1__1702 (.o(net1702));
 b15tihi00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_2__gen_filter_8__u_filter_diff_ctr_q_reg_3__1703 (.o(net1703));
 b15tihi00an1n03x5 gen_filter_8__u_filter_filter_q_reg_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1704 (.o(net1704));
 b15tihi00an1n03x5 gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_diff_ctr_q_reg_0__1705 (.o(net1705));
 b15tihi00an1n03x5 gen_filter_8__u_filter_stored_value_q_reg_1706 (.o(net1706));
 b15tihi00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_1__gen_filter_9__u_filter_diff_ctr_q_reg_2__1707 (.o(net1707));
 b15tihi00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_3__gen_filter_9__u_filter_filter_q_reg_1708 (.o(net1708));
 b15tihi00an1n03x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_1__1709 (.o(net1709));
 b15tihi00an1n03x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1710 (.o(net1710));
 b15tihi00an1n03x5 gen_filter_9__u_filter_stored_value_q_reg_1711 (.o(net1711));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_10__intr_hw_intr_o_reg_11__1712 (.o(net1712));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_12__intr_hw_intr_o_reg_13__1713 (.o(net1713));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_14__intr_hw_intr_o_reg_15__1714 (.o(net1714));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_16__intr_hw_intr_o_reg_17__1715 (.o(net1715));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_19__intr_hw_intr_o_reg_20__1716 (.o(net1716));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_1__intr_hw_intr_o_reg_2__1717 (.o(net1717));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_21__intr_hw_intr_o_reg_30__1718 (.o(net1718));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_22__intr_hw_intr_o_reg_23__1719 (.o(net1719));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_24__intr_hw_intr_o_reg_25__1720 (.o(net1720));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_26__intr_hw_intr_o_reg_27__1721 (.o(net1721));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_28__intr_hw_intr_o_reg_29__1722 (.o(net1722));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_31__u_reg_u_data_in_q_reg_3__1723 (.o(net1723));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_4__intr_hw_intr_o_reg_5__1724 (.o(net1724));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_6__intr_hw_intr_o_reg_7__1725 (.o(net1725));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_8__intr_hw_intr_o_reg_18__1726 (.o(net1726));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_9__u_reg_u_data_in_q_reg_5__1727 (.o(net1727));
 b15tihi00an1n03x5 u_reg_err_q_reg_u_reg_u_data_in_q_reg_6__1728 (.o(net1728));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_0__u_reg_u_ctrl_en_input_filter_q_reg_1__1729 (.o(net1729));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_10__u_reg_u_ctrl_en_input_filter_q_reg_11__1730 (.o(net1730));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_12__u_reg_u_ctrl_en_input_filter_q_reg_13__1731 (.o(net1731));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_14__u_reg_u_ctrl_en_input_filter_q_reg_15__1732 (.o(net1732));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_16__u_reg_u_ctrl_en_input_filter_q_reg_17__1733 (.o(net1733));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_18__u_reg_u_ctrl_en_input_filter_q_reg_19__1734 (.o(net1734));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_20__u_reg_u_ctrl_en_input_filter_q_reg_21__1735 (.o(net1735));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_22__u_reg_u_ctrl_en_input_filter_q_reg_23__1736 (.o(net1736));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_24__u_reg_u_ctrl_en_input_filter_q_reg_25__1737 (.o(net1737));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_26__u_reg_u_ctrl_en_input_filter_q_reg_27__1738 (.o(net1738));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_28__u_reg_u_ctrl_en_input_filter_q_reg_29__1739 (.o(net1739));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_2__u_reg_u_ctrl_en_input_filter_q_reg_3__1740 (.o(net1740));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_30__u_reg_u_ctrl_en_input_filter_q_reg_31__1741 (.o(net1741));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_4__u_reg_u_ctrl_en_input_filter_q_reg_5__1742 (.o(net1742));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_6__u_reg_u_ctrl_en_input_filter_q_reg_7__1743 (.o(net1743));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_8__u_reg_u_ctrl_en_input_filter_q_reg_9__1744 (.o(net1744));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_0__u_reg_u_data_in_q_reg_1__1745 (.o(net1745));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_11__u_reg_u_data_in_q_reg_16__1746 (.o(net1746));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_12__u_reg_u_data_in_q_reg_17__1747 (.o(net1747));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_13__u_reg_u_data_in_q_reg_14__1748 (.o(net1748));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_18__u_reg_u_data_in_q_reg_19__1749 (.o(net1749));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_20__u_reg_u_data_in_q_reg_21__1750 (.o(net1750));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_22__u_reg_u_data_in_q_reg_23__1751 (.o(net1751));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_24__u_reg_u_data_in_q_reg_25__1752 (.o(net1752));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_26__u_reg_u_reg_if_rspop_q_reg_1__1753 (.o(net1753));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_27__1754 (.o(net1754));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_28__u_reg_u_data_in_q_reg_29__1755 (.o(net1755));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_2__u_reg_u_data_in_q_reg_8__1756 (.o(net1756));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_30__u_reg_u_reg_if_rspop_q_reg_2__1757 (.o(net1757));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_4__u_reg_u_data_in_q_reg_10__1758 (.o(net1758));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_7__u_reg_u_data_in_q_reg_31__1759 (.o(net1759));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_9__u_reg_u_data_in_q_reg_15__1760 (.o(net1760));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_0__u_reg_u_intr_ctrl_en_falling_q_reg_1__1761 (.o(net1761));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_10__u_reg_u_intr_ctrl_en_falling_q_reg_11__1762 (.o(net1762));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_12__u_reg_u_intr_ctrl_en_falling_q_reg_13__1763 (.o(net1763));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_14__u_reg_u_intr_ctrl_en_falling_q_reg_15__1764 (.o(net1764));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_16__u_reg_u_intr_ctrl_en_falling_q_reg_17__1765 (.o(net1765));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_18__u_reg_u_intr_ctrl_en_falling_q_reg_19__1766 (.o(net1766));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_20__u_reg_u_intr_ctrl_en_falling_q_reg_21__1767 (.o(net1767));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_22__u_reg_u_intr_ctrl_en_falling_q_reg_23__1768 (.o(net1768));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_24__u_reg_u_intr_ctrl_en_falling_q_reg_25__1769 (.o(net1769));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_26__u_reg_u_intr_ctrl_en_falling_q_reg_27__1770 (.o(net1770));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_28__u_reg_u_intr_ctrl_en_falling_q_reg_29__1771 (.o(net1771));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_2__u_reg_u_intr_ctrl_en_falling_q_reg_3__1772 (.o(net1772));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_30__u_reg_u_intr_ctrl_en_falling_q_reg_31__1773 (.o(net1773));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_4__u_reg_u_intr_ctrl_en_falling_q_reg_5__1774 (.o(net1774));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_6__u_reg_u_intr_ctrl_en_falling_q_reg_7__1775 (.o(net1775));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_8__u_reg_u_intr_ctrl_en_falling_q_reg_9__1776 (.o(net1776));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1__1777 (.o(net1777));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11__1778 (.o(net1778));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13__1779 (.o(net1779));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15__1780 (.o(net1780));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17__1781 (.o(net1781));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19__1782 (.o(net1782));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21__1783 (.o(net1783));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23__1784 (.o(net1784));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25__1785 (.o(net1785));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27__1786 (.o(net1786));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29__1787 (.o(net1787));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3__1788 (.o(net1788));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31__1789 (.o(net1789));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5__1790 (.o(net1790));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7__1791 (.o(net1791));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9__1792 (.o(net1792));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_reg_u_intr_ctrl_en_lvllow_q_reg_1__1793 (.o(net1793));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_reg_u_intr_ctrl_en_lvllow_q_reg_11__1794 (.o(net1794));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_reg_u_intr_ctrl_en_lvllow_q_reg_13__1795 (.o(net1795));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_reg_u_intr_ctrl_en_lvllow_q_reg_15__1796 (.o(net1796));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_reg_u_intr_ctrl_en_lvllow_q_reg_17__1797 (.o(net1797));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_reg_u_intr_ctrl_en_lvllow_q_reg_19__1798 (.o(net1798));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_reg_u_intr_ctrl_en_lvllow_q_reg_21__1799 (.o(net1799));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_reg_u_intr_ctrl_en_lvllow_q_reg_23__1800 (.o(net1800));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_reg_u_intr_ctrl_en_lvllow_q_reg_25__1801 (.o(net1801));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_reg_u_intr_ctrl_en_lvllow_q_reg_27__1802 (.o(net1802));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_reg_u_intr_ctrl_en_lvllow_q_reg_29__1803 (.o(net1803));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_reg_u_intr_ctrl_en_lvllow_q_reg_3__1804 (.o(net1804));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_reg_u_intr_ctrl_en_lvllow_q_reg_31__1805 (.o(net1805));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_reg_u_intr_ctrl_en_lvllow_q_reg_5__1806 (.o(net1806));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_reg_u_intr_ctrl_en_lvllow_q_reg_7__1807 (.o(net1807));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_reg_u_intr_ctrl_en_lvllow_q_reg_9__1808 (.o(net1808));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_0__u_reg_u_intr_ctrl_en_rising_q_reg_1__1809 (.o(net1809));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_10__u_reg_u_intr_ctrl_en_rising_q_reg_11__1810 (.o(net1810));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_12__u_reg_u_intr_ctrl_en_rising_q_reg_13__1811 (.o(net1811));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_14__u_reg_u_intr_ctrl_en_rising_q_reg_15__1812 (.o(net1812));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_16__u_reg_u_intr_ctrl_en_rising_q_reg_17__1813 (.o(net1813));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_18__u_reg_u_intr_ctrl_en_rising_q_reg_19__1814 (.o(net1814));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_20__u_reg_u_intr_ctrl_en_rising_q_reg_21__1815 (.o(net1815));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_22__u_reg_u_intr_ctrl_en_rising_q_reg_23__1816 (.o(net1816));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_24__u_reg_u_intr_ctrl_en_rising_q_reg_25__1817 (.o(net1817));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_26__u_reg_u_intr_ctrl_en_rising_q_reg_27__1818 (.o(net1818));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_28__u_reg_u_intr_ctrl_en_rising_q_reg_29__1819 (.o(net1819));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_2__u_reg_u_intr_ctrl_en_rising_q_reg_3__1820 (.o(net1820));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_30__u_reg_u_intr_ctrl_en_rising_q_reg_31__1821 (.o(net1821));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_4__u_reg_u_intr_ctrl_en_rising_q_reg_5__1822 (.o(net1822));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_6__u_reg_u_intr_ctrl_en_rising_q_reg_7__1823 (.o(net1823));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_8__u_reg_u_intr_ctrl_en_rising_q_reg_9__1824 (.o(net1824));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_0__u_reg_u_intr_enable_q_reg_1__1825 (.o(net1825));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_10__u_reg_u_intr_enable_q_reg_11__1826 (.o(net1826));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_12__u_reg_u_intr_enable_q_reg_13__1827 (.o(net1827));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_14__u_reg_u_intr_enable_q_reg_15__1828 (.o(net1828));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_16__u_reg_u_intr_enable_q_reg_17__1829 (.o(net1829));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_18__u_reg_u_intr_enable_q_reg_19__1830 (.o(net1830));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_20__u_reg_u_intr_enable_q_reg_21__1831 (.o(net1831));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_22__u_reg_u_intr_enable_q_reg_23__1832 (.o(net1832));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_24__u_reg_u_intr_enable_q_reg_25__1833 (.o(net1833));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_26__u_reg_u_intr_enable_q_reg_27__1834 (.o(net1834));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_28__u_reg_u_intr_enable_q_reg_29__1835 (.o(net1835));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_2__u_reg_u_intr_enable_q_reg_3__1836 (.o(net1836));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_30__u_reg_u_intr_enable_q_reg_31__1837 (.o(net1837));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_4__u_reg_u_intr_enable_q_reg_5__1838 (.o(net1838));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_6__u_reg_u_intr_enable_q_reg_7__1839 (.o(net1839));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_8__u_reg_u_intr_enable_q_reg_9__1840 (.o(net1840));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_0__u_reg_u_intr_state_q_reg_1__1841 (.o(net1841));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_10__u_reg_u_intr_state_q_reg_11__1842 (.o(net1842));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_12__u_reg_u_intr_state_q_reg_13__1843 (.o(net1843));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_14__u_reg_u_intr_state_q_reg_15__1844 (.o(net1844));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_16__u_reg_u_intr_state_q_reg_17__1845 (.o(net1845));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_18__u_reg_u_intr_state_q_reg_19__1846 (.o(net1846));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_20__u_reg_u_intr_state_q_reg_21__1847 (.o(net1847));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_22__u_reg_u_intr_state_q_reg_23__1848 (.o(net1848));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_24__u_reg_u_intr_state_q_reg_25__1849 (.o(net1849));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_26__u_reg_u_intr_state_q_reg_27__1850 (.o(net1850));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_28__u_reg_u_intr_state_q_reg_29__1851 (.o(net1851));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_2__u_reg_u_intr_state_q_reg_3__1852 (.o(net1852));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_30__u_reg_u_intr_state_q_reg_31__1853 (.o(net1853));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_4__u_reg_u_intr_state_q_reg_5__1854 (.o(net1854));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_6__u_reg_u_intr_state_q_reg_7__1855 (.o(net1855));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_8__u_reg_u_intr_state_q_reg_9__1856 (.o(net1856));
 b15tihi00an1n03x5 u_reg_u_reg_if_error_q_reg_1857 (.o(net1857));
 b15tihi00an1n03x5 u_reg_u_reg_if_outstanding_q_reg_1858 (.o(net1858));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_0__u_reg_u_reg_if_rdata_q_reg_1__1859 (.o(net1859));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_10__u_reg_u_reg_if_rdata_q_reg_11__1860 (.o(net1860));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_12__u_reg_u_reg_if_rdata_q_reg_13__1861 (.o(net1861));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_14__u_reg_u_reg_if_rdata_q_reg_15__1862 (.o(net1862));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_16__u_reg_u_reg_if_rdata_q_reg_17__1863 (.o(net1863));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_18__u_reg_u_reg_if_rdata_q_reg_19__1864 (.o(net1864));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_20__u_reg_u_reg_if_rdata_q_reg_21__1865 (.o(net1865));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_22__u_reg_u_reg_if_rdata_q_reg_23__1866 (.o(net1866));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_24__u_reg_u_reg_if_rdata_q_reg_25__1867 (.o(net1867));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_26__u_reg_u_reg_if_rdata_q_reg_27__1868 (.o(net1868));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_28__u_reg_u_reg_if_rdata_q_reg_29__1869 (.o(net1869));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_2__u_reg_u_reg_if_rdata_q_reg_3__1870 (.o(net1870));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_30__u_reg_u_reg_if_rdata_q_reg_31__1871 (.o(net1871));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_4__u_reg_u_reg_if_rdata_q_reg_5__1872 (.o(net1872));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_6__u_reg_u_reg_if_rdata_q_reg_7__1873 (.o(net1873));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_q_reg_8__u_reg_u_reg_if_rdata_q_reg_9__1874 (.o(net1874));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqid_q_reg_0__u_reg_u_reg_if_reqid_q_reg_1__1875 (.o(net1875));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqid_q_reg_2__u_reg_u_reg_if_reqid_q_reg_3__1876 (.o(net1876));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqid_q_reg_4__u_reg_u_reg_if_reqid_q_reg_5__1877 (.o(net1877));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqid_q_reg_6__u_reg_u_reg_if_reqid_q_reg_7__1878 (.o(net1878));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqsz_q_reg_0__1879 (.o(net1879));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqsz_q_reg_1__1880 (.o(net1880));
 b15tihi00an1n03x5 u_reg_u_reg_if_rspop_q_reg_0__1881 (.o(net1881));
 b15cbf000an1n16x5 clkbuf_leaf_1_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_1_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_2_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_2_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_3_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_3_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_4_clk_i (.clk(net1885),
    .clkout(clknet_leaf_4_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_5_clk_i (.clk(net1883),
    .clkout(clknet_leaf_5_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_6_clk_i (.clk(net1883),
    .clkout(clknet_leaf_6_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_7_clk_i (.clk(clknet_1_1__leaf_clk_i),
    .clkout(clknet_leaf_7_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_8_clk_i (.clk(net1884),
    .clkout(clknet_leaf_8_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_9_clk_i (.clk(clknet_1_1__leaf_clk_i),
    .clkout(clknet_leaf_9_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_10_clk_i (.clk(net1884),
    .clkout(clknet_leaf_10_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_11_clk_i (.clk(net1884),
    .clkout(clknet_leaf_11_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_12_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_12_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_13_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_13_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_14_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_14_clk_i));
 b15cbf000an1n16x5 clkbuf_0_clk_i (.clk(net1882),
    .clkout(clknet_0_clk_i));
 b15cbf000an1n16x5 clkbuf_1_0__f_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_1_0__leaf_clk_i));
 b15cbf000an1n16x5 clkbuf_1_1__f_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_1_1__leaf_clk_i));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_reg_if_net2138 (.clk(u_reg_u_reg_if_net2138),
    .clkout(clknet_0_u_reg_u_reg_if_net2138));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_reg_if_net2138 (.clk(clknet_0_u_reg_u_reg_if_net2138),
    .clkout(clknet_1_0__leaf_u_reg_u_reg_if_net2138));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_reg_if_net2138 (.clk(clknet_0_u_reg_u_reg_if_net2138),
    .clkout(clknet_1_1__leaf_u_reg_u_reg_if_net2138));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_reg_if_net2144 (.clk(u_reg_u_reg_if_net2144),
    .clkout(clknet_0_u_reg_u_reg_if_net2144));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_reg_if_net2144 (.clk(clknet_0_u_reg_u_reg_if_net2144),
    .clkout(clknet_1_0__leaf_u_reg_u_reg_if_net2144));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_reg_if_net2144 (.clk(clknet_0_u_reg_u_reg_if_net2144),
    .clkout(clknet_1_1__leaf_u_reg_u_reg_if_net2144));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_reg_if_net2149 (.clk(u_reg_u_reg_if_net2149),
    .clkout(clknet_0_u_reg_u_reg_if_net2149));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_reg_if_net2149 (.clk(clknet_0_u_reg_u_reg_if_net2149),
    .clkout(clknet_1_0__leaf_u_reg_u_reg_if_net2149));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_reg_if_net2149 (.clk(clknet_0_u_reg_u_reg_if_net2149),
    .clkout(clknet_1_1__leaf_u_reg_u_reg_if_net2149));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_state_net2115 (.clk(u_reg_u_intr_state_net2115),
    .clkout(clknet_0_u_reg_u_intr_state_net2115));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_state_net2115 (.clk(clknet_0_u_reg_u_intr_state_net2115),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_state_net2115));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_state_net2115 (.clk(clknet_0_u_reg_u_intr_state_net2115),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_state_net2115));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_state_net2121 (.clk(u_reg_u_intr_state_net2121),
    .clkout(clknet_0_u_reg_u_intr_state_net2121));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_state_net2121 (.clk(clknet_0_u_reg_u_intr_state_net2121),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_state_net2121));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_state_net2121 (.clk(clknet_0_u_reg_u_intr_state_net2121),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_state_net2121));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_enable_net2092 (.clk(u_reg_u_intr_enable_net2092),
    .clkout(clknet_0_u_reg_u_intr_enable_net2092));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_enable_net2092 (.clk(clknet_0_u_reg_u_intr_enable_net2092),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_enable_net2092));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_enable_net2092 (.clk(clknet_0_u_reg_u_intr_enable_net2092),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_enable_net2092));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_enable_net2098 (.clk(u_reg_u_intr_enable_net2098),
    .clkout(clknet_0_u_reg_u_intr_enable_net2098));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_enable_net2098 (.clk(clknet_0_u_reg_u_intr_enable_net2098),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_enable_net2098));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_enable_net2098 (.clk(clknet_0_u_reg_u_intr_enable_net2098),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_enable_net2098));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_rising_net2092 (.clk(u_reg_u_intr_ctrl_en_rising_net2092),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_rising_net2092));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_rising_net2092 (.clk(clknet_0_u_reg_u_intr_ctrl_en_rising_net2092),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2092));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_rising_net2092 (.clk(clknet_0_u_reg_u_intr_ctrl_en_rising_net2092),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2092));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_rising_net2098 (.clk(u_reg_u_intr_ctrl_en_rising_net2098),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_rising_net2098));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_rising_net2098 (.clk(clknet_0_u_reg_u_intr_ctrl_en_rising_net2098),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2098));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_rising_net2098 (.clk(clknet_0_u_reg_u_intr_ctrl_en_rising_net2098),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2098));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_lvllow_net2092 (.clk(u_reg_u_intr_ctrl_en_lvllow_net2092),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2092));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_lvllow_net2092 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2092),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_lvllow_net2092 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2092),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2092));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_lvllow_net2098 (.clk(u_reg_u_intr_ctrl_en_lvllow_net2098),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2098));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_lvllow_net2098 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2098),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_lvllow_net2098 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2098),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2098));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_lvlhigh_net2092 (.clk(u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2092));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_lvlhigh_net2092 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_lvlhigh_net2092 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2092),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2092));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_lvlhigh_net2098 (.clk(u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2098));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_lvlhigh_net2098 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_lvlhigh_net2098 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2098),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2098));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_falling_net2092 (.clk(u_reg_u_intr_ctrl_en_falling_net2092),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_falling_net2092));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_falling_net2092 (.clk(clknet_0_u_reg_u_intr_ctrl_en_falling_net2092),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2092));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_falling_net2092 (.clk(clknet_0_u_reg_u_intr_ctrl_en_falling_net2092),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2092));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_falling_net2098 (.clk(u_reg_u_intr_ctrl_en_falling_net2098),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_falling_net2098));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_falling_net2098 (.clk(clknet_0_u_reg_u_intr_ctrl_en_falling_net2098),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2098));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_falling_net2098 (.clk(clknet_0_u_reg_u_intr_ctrl_en_falling_net2098),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2098));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_ctrl_en_input_filter_net2092 (.clk(u_reg_u_ctrl_en_input_filter_net2092),
    .clkout(clknet_0_u_reg_u_ctrl_en_input_filter_net2092));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_ctrl_en_input_filter_net2092 (.clk(clknet_0_u_reg_u_ctrl_en_input_filter_net2092),
    .clkout(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2092));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_ctrl_en_input_filter_net2092 (.clk(clknet_0_u_reg_u_ctrl_en_input_filter_net2092),
    .clkout(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2092));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_ctrl_en_input_filter_net2098 (.clk(u_reg_u_ctrl_en_input_filter_net2098),
    .clkout(clknet_0_u_reg_u_ctrl_en_input_filter_net2098));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_ctrl_en_input_filter_net2098 (.clk(clknet_0_u_reg_u_ctrl_en_input_filter_net2098),
    .clkout(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2098));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_ctrl_en_input_filter_net2098 (.clk(clknet_0_u_reg_u_ctrl_en_input_filter_net2098),
    .clkout(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2098));
 b15cbf000an1n16x5 clkbuf_0_net2059 (.clk(net2059),
    .clkout(clknet_0_net2059));
 b15cbf000an1n16x5 clkbuf_1_0__f_net2059 (.clk(clknet_0_net2059),
    .clkout(clknet_1_0__leaf_net2059));
 b15cbf000an1n16x5 clkbuf_1_1__f_net2059 (.clk(clknet_0_net2059),
    .clkout(clknet_1_1__leaf_net2059));
 b15cbf000an1n16x5 clkbuf_0_net2065 (.clk(net2065),
    .clkout(clknet_0_net2065));
 b15cbf000an1n16x5 clkbuf_1_0__f_net2065 (.clk(clknet_0_net2065),
    .clkout(clknet_1_0__leaf_net2065));
 b15cbf000an1n16x5 clkbuf_1_1__f_net2065 (.clk(clknet_0_net2065),
    .clkout(clknet_1_1__leaf_net2065));
 b15cbf000an1n16x5 clkbuf_0_net2070 (.clk(net2070),
    .clkout(clknet_0_net2070));
 b15cbf000an1n16x5 clkbuf_1_0__f_net2070 (.clk(clknet_0_net2070),
    .clkout(clknet_1_0__leaf_net2070));
 b15cbf000an1n16x5 clkbuf_1_1__f_net2070 (.clk(clknet_0_net2070),
    .clkout(clknet_1_1__leaf_net2070));
 b15cbf000an1n16x5 clkbuf_0_net2075 (.clk(net2075),
    .clkout(clknet_0_net2075));
 b15cbf000an1n16x5 clkbuf_1_0__f_net2075 (.clk(clknet_0_net2075),
    .clkout(clknet_1_0__leaf_net2075));
 b15cbf000an1n16x5 clkbuf_1_1__f_net2075 (.clk(clknet_0_net2075),
    .clkout(clknet_1_1__leaf_net2075));
 b15bfn001ah1n32x5 wire1 (.a(clk_i),
    .o(net1882));
 b15bfn001ah1n16x5 max_length2 (.a(clknet_1_1__leaf_clk_i),
    .o(net1883));
 b15bfn001ah1n24x5 wire3 (.a(net1885),
    .o(net1884));
 b15bfn001as1n16x5 max_length4 (.a(clknet_1_1__leaf_clk_i),
    .o(net1885));
 b15cbf034ar1n64x5 hold5 (.clk(net2482),
    .clkout(net1886));
 b15cbf034ar1n64x5 hold6 (.clk(net2484),
    .clkout(intr_gpio_o[17]));
 b15cbf034ar1n64x5 hold7 (.clk(net2485),
    .clkout(net1888));
 b15cbf034ar1n64x5 hold8 (.clk(net2487),
    .clkout(intr_gpio_o[16]));
 b15cbf034ar1n64x5 hold9 (.clk(net2488),
    .clkout(net1890));
 b15cbf034ar1n64x5 hold10 (.clk(net1891),
    .clkout(intr_gpio_o[23]));
 b15cbf034ar1n64x5 hold11 (.clk(net2490),
    .clkout(net1892));
 b15cbf034ar1n64x5 hold12 (.clk(net1893),
    .clkout(intr_gpio_o[22]));
 b15cbf034ar1n64x5 hold13 (.clk(net2492),
    .clkout(net1894));
 b15cbf034ar1n64x5 hold14 (.clk(net1895),
    .clkout(intr_gpio_o[29]));
 b15cbf034ar1n64x5 hold15 (.clk(net2494),
    .clkout(net1896));
 b15cbf034ar1n64x5 hold16 (.clk(net1897),
    .clkout(intr_gpio_o[28]));
 b15cbf034ar1n64x5 hold17 (.clk(net2496),
    .clkout(net1898));
 b15cbf034ar1n64x5 hold18 (.clk(net1899),
    .clkout(intr_gpio_o[2]));
 b15cbf034ar1n64x5 hold19 (.clk(net2498),
    .clkout(net1900));
 b15cbf034ar1n64x5 hold20 (.clk(net1901),
    .clkout(intr_gpio_o[1]));
 b15cbf034ar1n64x5 hold21 (.clk(net2510),
    .clkout(net1902));
 b15cbf034ar1n64x5 hold22 (.clk(net1903),
    .clkout(intr_gpio_o[30]));
 b15cbf034ar1n64x5 hold23 (.clk(net2512),
    .clkout(net1904));
 b15cbf034ar1n64x5 hold24 (.clk(net1905),
    .clkout(intr_gpio_o[21]));
 b15cbf034ar1n64x5 hold25 (.clk(net2502),
    .clkout(net1906));
 b15cbf034ar1n64x5 hold26 (.clk(net1907),
    .clkout(intr_gpio_o[18]));
 b15cbf034ar1n64x5 hold27 (.clk(net2500),
    .clkout(net1908));
 b15cbf034ar1n64x5 hold28 (.clk(net1909),
    .clkout(intr_gpio_o[13]));
 b15cbf034ar1n64x5 hold29 (.clk(net2504),
    .clkout(net1910));
 b15cbf034ar1n64x5 hold30 (.clk(net1911),
    .clkout(intr_gpio_o[12]));
 b15cbf034ar1n64x5 hold31 (.clk(net2506),
    .clkout(net1912));
 b15cbf034ar1n64x5 hold32 (.clk(net1913),
    .clkout(intr_gpio_o[8]));
 b15cbf034ar1n64x5 hold33 (.clk(net2508),
    .clkout(net1914));
 b15cbf034ar1n64x5 hold34 (.clk(net1915),
    .clkout(intr_gpio_o[3]));
 b15cbf034ar1n64x5 hold35 (.clk(net2514),
    .clkout(net1916));
 b15cbf034ar1n64x5 hold36 (.clk(net1917),
    .clkout(alert_tx_o[1]));
 b15cbf034ar1n64x5 hold37 (.clk(net1941),
    .clkout(net1918));
 b15cbf034ar1n64x5 hold38 (.clk(net676),
    .clkout(net1919));
 b15cbf034ar1n64x5 hold39 (.clk(net1920),
    .clkout(tl_o[63]));
 b15cbf034ar1n64x5 hold40 (.clk(net2516),
    .clkout(net1921));
 b15cbf034ar1n64x5 hold41 (.clk(net1922),
    .clkout(alert_tx_o[0]));
 b15cbf034ar1n64x5 hold42 (.clk(net2520),
    .clkout(net1923));
 b15cbf034ar1n64x5 hold43 (.clk(net1924),
    .clkout(intr_gpio_o[0]));
 b15cbf034ar1n64x5 hold44 (.clk(net2518),
    .clkout(net1925));
 b15cbf034ar1n64x5 hold45 (.clk(net1926),
    .clkout(intr_gpio_o[4]));
 b15cbf034ar1n64x5 hold46 (.clk(net2522),
    .clkout(net1927));
 b15cbf034ar1n64x5 hold47 (.clk(net1928),
    .clkout(intr_gpio_o[5]));
 b15cbf034ar1n64x5 hold48 (.clk(net2524),
    .clkout(net1929));
 b15cbf034ar1n64x5 hold49 (.clk(net1930),
    .clkout(intr_gpio_o[9]));
 b15cbf034ar1n64x5 hold50 (.clk(net2526),
    .clkout(net1931));
 b15cbf034ar1n64x5 hold51 (.clk(net1932),
    .clkout(intr_gpio_o[19]));
 b15cbf034ar1n64x5 hold52 (.clk(net2530),
    .clkout(net1933));
 b15cbf034ar1n64x5 hold53 (.clk(net1934),
    .clkout(intr_gpio_o[20]));
 b15cbf034ar1n64x5 hold54 (.clk(net2528),
    .clkout(net1935));
 b15cbf034ar1n64x5 hold55 (.clk(net1936),
    .clkout(intr_gpio_o[10]));
 b15cbf034ar1n64x5 hold56 (.clk(net2537),
    .clkout(net1937));
 b15cbf034ar1n64x5 hold57 (.clk(net1938),
    .clkout(intr_gpio_o[14]));
 b15cbf034ar1n64x5 hold58 (.clk(net2536),
    .clkout(net1939));
 b15cbf034ar1n64x5 hold59 (.clk(net1940),
    .clkout(intr_gpio_o[15]));
 b15cbf034ar1n64x5 hold60 (.clk(net292),
    .clkout(net1941));
 b15cbf034ar1n64x5 hold61 (.clk(net2532),
    .clkout(net1942));
 b15cbf034ar1n64x5 hold62 (.clk(net1943),
    .clkout(intr_gpio_o[11]));
 b15cbf034ar1n64x5 hold63 (.clk(net2534),
    .clkout(net1944));
 b15cbf034ar1n64x5 hold64 (.clk(net1945),
    .clkout(intr_gpio_o[31]));
 b15cbf034ar1n64x5 hold65 (.clk(net2543),
    .clkout(net1946));
 b15cbf034ar1n64x5 hold66 (.clk(net1947),
    .clkout(tl_o[53]));
 b15cbf034ar1n64x5 hold67 (.clk(net2542),
    .clkout(net1948));
 b15cbf034ar1n64x5 hold68 (.clk(net1949),
    .clkout(tl_o[54]));
 b15cbf034ar1n64x5 hold69 (.clk(net1981),
    .clkout(net1950));
 b15cbf034ar1n64x5 hold70 (.clk(net1951),
    .clkout(tl_o[64]));
 b15cbf034ar1n64x5 hold71 (.clk(net2544),
    .clkout(net1952));
 b15cbf034ar1n64x5 hold72 (.clk(net1953),
    .clkout(tl_o[52]));
 b15cbf034ar1n64x5 hold73 (.clk(net1989),
    .clkout(net1954));
 b15cbf034ar1n64x5 hold74 (.clk(net1955),
    .clkout(tl_o[58]));
 b15cbf034ar1n64x5 hold75 (.clk(net2545),
    .clkout(net1956));
 b15cbf034ar1n64x5 hold76 (.clk(net1957),
    .clkout(tl_o[51]));
 b15cbf034ar1n64x5 hold77 (.clk(net2546),
    .clkout(net1958));
 b15cbf034ar1n64x5 hold78 (.clk(net1959),
    .clkout(tl_o[50]));
 b15cbf034ar1n64x5 hold79 (.clk(net2548),
    .clkout(net1960));
 b15cbf034ar1n64x5 hold80 (.clk(net1961),
    .clkout(tl_o[56]));
 b15cbf034ar1n64x5 hold81 (.clk(net2547),
    .clkout(net1962));
 b15cbf034ar1n64x5 hold82 (.clk(net1963),
    .clkout(tl_o[49]));
 b15cbf034ar1n64x5 hold83 (.clk(net2549),
    .clkout(net1964));
 b15cbf034ar1n64x5 hold84 (.clk(net1965),
    .clkout(tl_o[55]));
 b15cbf034ar1n64x5 hold85 (.clk(net2538),
    .clkout(net1966));
 b15cbf034ar1n64x5 hold86 (.clk(net1967),
    .clkout(intr_gpio_o[24]));
 b15cbf034ar1n64x5 hold87 (.clk(net2539),
    .clkout(net1968));
 b15cbf034ar1n64x5 hold88 (.clk(net1969),
    .clkout(intr_gpio_o[25]));
 b15cbf034ar1n64x5 hold89 (.clk(net1991),
    .clkout(net1970));
 b15cbf034ar1n64x5 hold90 (.clk(net1971),
    .clkout(tl_o[57]));
 b15cbf034ar1n64x5 hold91 (.clk(net2540),
    .clkout(net1972));
 b15cbf034ar1n64x5 hold92 (.clk(net1973),
    .clkout(intr_gpio_o[26]));
 b15cbf034ar1n64x5 hold93 (.clk(net2541),
    .clkout(net1974));
 b15cbf034ar1n64x5 hold94 (.clk(net1975),
    .clkout(intr_gpio_o[27]));
 b15cbf034ar1n64x5 hold95 (.clk(net1985),
    .clkout(net1976));
 b15cbf034ar1n64x5 hold96 (.clk(net239),
    .clkout(net1977));
 b15cbf034ar1n64x5 hold97 (.clk(net1978),
    .clkout(tl_o[11]));
 b15cbf034ar1n64x5 hold98 (.clk(net2550),
    .clkout(net1979));
 b15cbf034ar1n64x5 hold99 (.clk(net1980),
    .clkout(intr_gpio_o[6]));
 b15cbf034ar1n64x5 hold100 (.clk(net293),
    .clkout(net1981));
 b15cbf034ar1n64x5 hold101 (.clk(net1950),
    .clkout(net1982));
 b15cbf034ar1n64x5 hold102 (.clk(net240),
    .clkout(net1983));
 b15cbf034ar1n64x5 hold103 (.clk(net1984),
    .clkout(tl_o[12]));
 b15cbf034ar1n64x5 hold104 (.clk(net248),
    .clkout(net1985));
 b15cbf034ar1n64x5 hold105 (.clk(net1976),
    .clkout(net1986));
 b15cbf034ar1n64x5 hold106 (.clk(net2551),
    .clkout(net1987));
 b15cbf034ar1n64x5 hold107 (.clk(net1988),
    .clkout(intr_gpio_o[7]));
 b15cbf034ar1n64x5 hold108 (.clk(net289),
    .clkout(net1989));
 b15cbf034ar1n64x5 hold109 (.clk(net1954),
    .clkout(net1990));
 b15cbf034ar1n64x5 hold110 (.clk(net288),
    .clkout(net1991));
 b15cbf034ar1n64x5 hold111 (.clk(net1970),
    .clkout(net1992));
 b15cbf034ar1n64x5 hold112 (.clk(net238),
    .clkout(net1993));
 b15cbf034ar1n64x5 hold113 (.clk(net2034),
    .clkout(net1994));
 b15cbf034ar1n64x5 hold114 (.clk(n2954),
    .clkout(net1995));
 b15cbf034ar1n64x5 hold115 (.clk(n2956),
    .clkout(net1996));
 b15cbf034ar1n64x5 hold116 (.clk(net2038),
    .clkout(net1997));
 b15cbf034ar1n64x5 hold117 (.clk(net1998),
    .clkout(tl_o[65]));
 b15cbf034ar1n64x5 hold118 (.clk(net2555),
    .clkout(net1999));
 b15cbf034ar1n64x5 hold119 (.clk(net2000),
    .clkout(tl_o[37]));
 b15cbf034ar1n64x5 hold120 (.clk(net2564),
    .clkout(net2001));
 b15cbf034ar1n64x5 hold121 (.clk(net2002),
    .clkout(tl_o[43]));
 b15cbf034ar1n64x5 hold122 (.clk(net2557),
    .clkout(net2003));
 b15cbf034ar1n64x5 hold123 (.clk(net2004),
    .clkout(tl_o[45]));
 b15cbf034ar1n64x5 hold124 (.clk(u_reg_data_in_qs[19]),
    .clkout(net2005));
 b15cbf034ar1n64x5 hold125 (.clk(n3941),
    .clkout(net2006));
 b15cbf034ar1n64x5 hold126 (.clk(u_reg_u_reg_if_N33),
    .clkout(net2007));
 b15cbf034ar1n64x5 hold127 (.clk(net265),
    .clkout(net2008));
 b15cbf034ar1n64x5 hold128 (.clk(net479),
    .clkout(net2009));
 b15cbf034ar1n64x5 hold129 (.clk(net273),
    .clkout(net2010));
 b15cbf034ar1n64x5 hold130 (.clk(net2011),
    .clkout(tl_o[42]));
 b15cbf034ar1n64x5 hold131 (.clk(net2117),
    .clkout(net2012));
 b15cbf034ar1n64x5 hold132 (.clk(net2013),
    .clkout(tl_o[40]));
 b15cbf034ar1n64x5 hold133 (.clk(u_reg_data_in_qs[18]),
    .clkout(net2014));
 b15cbf034ar1n64x5 hold134 (.clk(n3933),
    .clkout(net2015));
 b15cbf034ar1n64x5 hold135 (.clk(n3937),
    .clkout(net2016));
 b15cbf034ar1n64x5 hold136 (.clk(u_reg_u_reg_if_N32),
    .clkout(net2017));
 b15cbf034ar1n64x5 hold137 (.clk(net2112),
    .clkout(net2018));
 b15cbf034ar1n64x5 hold138 (.clk(net2019),
    .clkout(tl_o[33]));
 b15cbf034ar1n64x5 hold139 (.clk(net173),
    .clkout(net2020));
 b15cbf034ar1n64x5 hold140 (.clk(net2021),
    .clkout(cio_gpio_o[0]));
 b15cbf034ar1n64x5 hold141 (.clk(net2556),
    .clkout(net2022));
 b15cbf034ar1n64x5 hold142 (.clk(net2023),
    .clkout(tl_o[36]));
 b15cbf034ar1n64x5 hold143 (.clk(net244),
    .clkout(net2024));
 b15cbf034ar1n64x5 hold144 (.clk(net2025),
    .clkout(tl_o[16]));
 b15cbf034ar1n64x5 hold145 (.clk(net184),
    .clkout(net2026));
 b15cbf034ar1n64x5 hold146 (.clk(net2027),
    .clkout(cio_gpio_o[1]));
 b15cbf034ar1n64x5 hold147 (.clk(net256),
    .clkout(net2028));
 b15cbf034ar1n64x5 hold148 (.clk(net496),
    .clkout(net2029));
 b15cbf034ar1n64x5 hold149 (.clk(net252),
    .clkout(net2030));
 b15cbf034ar1n64x5 hold150 (.clk(net457),
    .clkout(net2031));
 b15cbf034ar1n64x5 hold151 (.clk(net249),
    .clkout(net2032));
 b15cbf034ar1n64x5 hold152 (.clk(net465),
    .clkout(net2033));
 b15cbf034ar1n64x5 hold153 (.clk(net291),
    .clkout(net2034));
 b15cbf034ar1n64x5 hold154 (.clk(net1994),
    .clkout(net2035));
 b15cbf034ar1n64x5 hold155 (.clk(net203),
    .clkout(net2036));
 b15cbf034ar1n64x5 hold156 (.clk(net2037),
    .clkout(cio_gpio_o[8]));
 b15cbf034ar1n64x5 hold157 (.clk(net294),
    .clkout(net2038));
 b15cbf034ar1n64x5 hold158 (.clk(net150),
    .clkout(net2039));
 b15cbf034ar1n64x5 hold159 (.clk(net2040),
    .clkout(cio_gpio_en_o[18]));
 b15cbf034ar1n64x5 hold160 (.clk(net165),
    .clkout(net2041));
 b15cbf034ar1n64x5 hold161 (.clk(net2042),
    .clkout(cio_gpio_en_o[31]));
 b15cbf034ar1n64x5 hold162 (.clk(net268),
    .clkout(net2043));
 b15cbf034ar1n64x5 hold163 (.clk(net475),
    .clkout(net2044));
 b15cbf034ar1n64x5 hold164 (.clk(u_reg_data_in_qs[25]),
    .clkout(net2045));
 b15cbf034ar1n64x5 hold165 (.clk(n3985),
    .clkout(net2046));
 b15cbf034ar1n64x5 hold166 (.clk(u_reg_u_reg_if_N39),
    .clkout(net2047));
 b15cbf034ar1n64x5 hold167 (.clk(net260),
    .clkout(net2048));
 b15cbf034ar1n64x5 hold168 (.clk(net489),
    .clkout(net2049));
 b15cbf034ar1n64x5 hold169 (.clk(net156),
    .clkout(net2050));
 b15cbf034ar1n64x5 hold170 (.clk(net652),
    .clkout(net2051));
 b15cbf034ar1n64x5 hold171 (.clk(net264),
    .clkout(net2052));
 b15cbf034ar1n64x5 hold172 (.clk(net482),
    .clkout(net2053));
 b15cbf034ar1n64x5 hold173 (.clk(net250),
    .clkout(net2054));
 b15cbf034ar1n64x5 hold174 (.clk(net460),
    .clkout(net2055));
 b15cbf034ar1n64x5 hold175 (.clk(u_reg_data_in_qs[20]),
    .clkout(net2056));
 b15cbf034ar1n64x5 hold176 (.clk(n3950),
    .clkout(net2057));
 b15cbf034ar1n64x5 hold177 (.clk(u_reg_u_reg_if_N34),
    .clkout(net2058));
 b15cbf034ar1n64x5 hold178 (.clk(net161),
    .clkout(net2060));
 b15cbf034ar1n64x5 hold179 (.clk(net2061),
    .clkout(cio_gpio_en_o[28]));
 b15cbf034ar1n64x5 hold180 (.clk(u_reg_data_in_qs[28]),
    .clkout(net2062));
 b15cbf034ar1n64x5 hold181 (.clk(n4004),
    .clkout(net2063));
 b15cbf034ar1n64x5 hold182 (.clk(u_reg_u_reg_if_N42),
    .clkout(net2064));
 b15cbf034ar1n64x5 hold183 (.clk(net247),
    .clkout(net2066));
 b15cbf034ar1n64x5 hold184 (.clk(net466),
    .clkout(net2067));
 b15cbf034ar1n64x5 hold185 (.clk(net175),
    .clkout(net2068));
 b15cbf034ar1n64x5 hold186 (.clk(net638),
    .clkout(net2069));
 b15cbf034ar1n64x5 hold187 (.clk(net2218),
    .clkout(net2071));
 b15cbf034ar1n64x5 hold188 (.clk(net2072),
    .clkout(tl_o[41]));
 b15cbf034ar1n64x5 hold189 (.clk(u_reg_data_in_qs[7]),
    .clkout(net2073));
 b15cbf034ar1n64x5 hold190 (.clk(n3412),
    .clkout(net2074));
 b15cbf034ar1n64x5 hold191 (.clk(u_reg_u_reg_if_N21),
    .clkout(net2076));
 b15cbf034ar1n64x5 hold192 (.clk(net195),
    .clkout(net2077));
 b15cbf034ar1n64x5 hold193 (.clk(net2078),
    .clkout(cio_gpio_o[2]));
 b15cbf034ar1n64x5 hold194 (.clk(net157),
    .clkout(net2079));
 b15cbf034ar1n64x5 hold195 (.clk(net650),
    .clkout(net2080));
 b15cbf034ar1n64x5 hold196 (.clk(net162),
    .clkout(net2081));
 b15cbf034ar1n64x5 hold197 (.clk(net2082),
    .clkout(cio_gpio_en_o[29]));
 b15cbf034ar1n64x5 hold198 (.clk(net154),
    .clkout(net2083));
 b15cbf034ar1n64x5 hold199 (.clk(net655),
    .clkout(net2084));
 b15cbf034ar1n64x5 hold200 (.clk(net277),
    .clkout(net2085));
 b15cbf034ar1n64x5 hold201 (.clk(net2086),
    .clkout(tl_o[46]));
 b15cbf034ar1n64x5 hold202 (.clk(u_reg_data_in_qs[21]),
    .clkout(net2087));
 b15cbf034ar1n64x5 hold203 (.clk(n3957),
    .clkout(net2088));
 b15cbf034ar1n64x5 hold204 (.clk(u_reg_u_reg_if_N35),
    .clkout(net2089));
 b15cbf034ar1n64x5 hold205 (.clk(net258),
    .clkout(net2090));
 b15cbf034ar1n64x5 hold206 (.clk(net494),
    .clkout(net2091));
 b15cbf034ar1n64x5 hold207 (.clk(net245),
    .clkout(net2092));
 b15cbf034ar1n64x5 hold208 (.clk(net501),
    .clkout(net2093));
 b15cbf034ar1n64x5 hold209 (.clk(net153),
    .clkout(net2094));
 b15cbf034ar1n64x5 hold210 (.clk(net657),
    .clkout(net2095));
 b15cbf034ar1n64x5 hold211 (.clk(net198),
    .clkout(net2096));
 b15cbf034ar1n64x5 hold212 (.clk(net2097),
    .clkout(cio_gpio_o[3]));
 b15cbf034ar1n64x5 hold213 (.clk(net160),
    .clkout(net2098));
 b15cbf034ar1n64x5 hold214 (.clk(net646),
    .clkout(net2099));
 b15cbf034ar1n64x5 hold215 (.clk(u_reg_data_in_qs[12]),
    .clkout(net2100));
 b15cbf034ar1n64x5 hold216 (.clk(n3400),
    .clkout(net2101));
 b15cbf034ar1n64x5 hold217 (.clk(u_reg_u_reg_if_N26),
    .clkout(net2102));
 b15cbf034ar1n64x5 hold218 (.clk(u_reg_data_in_qs[6]),
    .clkout(net2103));
 b15cbf034ar1n64x5 hold219 (.clk(n3377),
    .clkout(net2104));
 b15cbf034ar1n64x5 hold220 (.clk(u_reg_u_reg_if_N20),
    .clkout(net2105));
 b15cbf034ar1n64x5 hold221 (.clk(net158),
    .clkout(net2106));
 b15cbf034ar1n64x5 hold222 (.clk(net202),
    .clkout(net2107));
 b15cbf034ar1n64x5 hold223 (.clk(net613),
    .clkout(net2108));
 b15cbf034ar1n64x5 hold224 (.clk(net2214),
    .clkout(net2109));
 b15cbf034ar1n64x5 hold225 (.clk(net2110),
    .clkout(tl_o[44]));
 b15cbf034ar1n64x5 hold226 (.clk(net204),
    .clkout(net2111));
 b15cbf034ar1n64x5 hold227 (.clk(net263),
    .clkout(net2112));
 b15cbf034ar1n64x5 hold228 (.clk(n3044),
    .clkout(net2113));
 b15cbf034ar1n64x5 hold229 (.clk(net259),
    .clkout(net2114));
 b15cbf034ar1n64x5 hold230 (.clk(net201),
    .clkout(net2115));
 b15cbf034ar1n64x5 hold231 (.clk(net614),
    .clkout(net2116));
 b15cbf034ar1n64x5 hold232 (.clk(net271),
    .clkout(net2117));
 b15cbf034ar1n64x5 hold233 (.clk(n2989),
    .clkout(net2118));
 b15cbf034ar1n64x5 hold234 (.clk(n3019),
    .clkout(net2119));
 b15cbf034ar1n64x5 hold235 (.clk(net296),
    .clkout(net2120));
 b15cbf034ar1n64x5 hold236 (.clk(gen_filter_17__u_filter_filter_q),
    .clkout(net2121));
 b15cbf034ar1n64x5 hold237 (.clk(n2879),
    .clkout(net2122));
 b15cbf034ar1n64x5 hold238 (.clk(gen_filter_17__u_filter_diff_ctr_d[1]),
    .clkout(net2123));
 b15cbf034ar1n64x5 hold239 (.clk(net246),
    .clkout(net2124));
 b15cbf034ar1n64x5 hold240 (.clk(net2561),
    .clkout(net2125));
 b15cbf034ar1n64x5 hold241 (.clk(u_reg_data_in_qs[16]),
    .clkout(net2126));
 b15cbf034ar1n64x5 hold242 (.clk(n3925),
    .clkout(net2127));
 b15cbf034ar1n64x5 hold243 (.clk(net155),
    .clkout(net2128));
 b15cbf034ar1n64x5 hold244 (.clk(net654),
    .clkout(net2129));
 b15cbf034ar1n64x5 hold245 (.clk(net255),
    .clkout(net2130));
 b15cbf034ar1n64x5 hold246 (.clk(net499),
    .clkout(net2131));
 b15cbf034ar1n64x5 hold247 (.clk(net148),
    .clkout(net2132));
 b15cbf034ar1n64x5 hold248 (.clk(net269),
    .clkout(net2133));
 b15cbf034ar1n64x5 hold249 (.clk(reg2hw_intr_enable__q__29_),
    .clkout(net2134));
 b15cbf034ar1n64x5 hold250 (.clk(u_reg_u_reg_if_N43),
    .clkout(net2135));
 b15cbf034ar1n64x5 hold251 (.clk(net2158),
    .clkout(net2136));
 b15cbf034ar1n64x5 hold252 (.clk(net2137),
    .clkout(tl_o[47]));
 b15cbf034ar1n64x5 hold253 (.clk(u_reg_data_in_qs[11]),
    .clkout(net2138));
 b15cbf034ar1n64x5 hold254 (.clk(net677),
    .clkout(net2139));
 b15cbf034ar1n64x5 hold255 (.clk(n3368),
    .clkout(net2140));
 b15cbf034ar1n64x5 hold256 (.clk(u_reg_u_reg_if_N25),
    .clkout(net2141));
 b15cbf034ar1n64x5 hold257 (.clk(net2186),
    .clkout(net2142));
 b15cbf034ar1n64x5 hold258 (.clk(net455),
    .clkout(net2143));
 b15cbf034ar1n64x5 hold259 (.clk(net254),
    .clkout(net2144));
 b15cbf034ar1n64x5 hold260 (.clk(gen_filter_14__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2145));
 b15cbf034ar1n64x5 hold261 (.clk(net2209),
    .clkout(net2146));
 b15cbf034ar1n64x5 hold262 (.clk(net2147),
    .clkout(tl_o[32]));
 b15cbf034ar1n64x5 hold263 (.clk(net149),
    .clkout(net2148));
 b15cbf034ar1n64x5 hold264 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_intq_0_),
    .clkout(net2149));
 b15cbf034ar1n64x5 hold265 (.clk(net177),
    .clkout(net2150));
 b15cbf034ar1n64x5 hold266 (.clk(net636),
    .clkout(net2151));
 b15cbf034ar1n64x5 hold267 (.clk(gen_filter_15__u_filter_diff_ctr_q[3]),
    .clkout(net2152));
 b15cbf034ar1n64x5 hold268 (.clk(n2918),
    .clkout(net2153));
 b15cbf034ar1n64x5 hold269 (.clk(gen_filter_15__u_filter_diff_ctr_d[0]),
    .clkout(net2154));
 b15cbf034ar1n64x5 hold270 (.clk(gen_filter_17__u_filter_diff_ctr_q[3]),
    .clkout(net2155));
 b15cbf034ar1n64x5 hold271 (.clk(gen_filter_17__u_filter_diff_ctr_d[2]),
    .clkout(net2156));
 b15cbf034ar1n64x5 hold272 (.clk(gen_filter_29__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2157));
 b15cbf034ar1n64x5 hold273 (.clk(net278),
    .clkout(net2158));
 b15cbf034ar1n64x5 hold274 (.clk(n3062),
    .clkout(net2159));
 b15cbf034ar1n64x5 hold275 (.clk(net270),
    .clkout(net2160));
 b15cbf034ar1n64x5 hold276 (.clk(gen_filter_23__u_filter_filter_q),
    .clkout(net2161));
 b15cbf034ar1n64x5 hold277 (.clk(n2885),
    .clkout(net2162));
 b15cbf034ar1n64x5 hold278 (.clk(gen_filter_23__u_filter_diff_ctr_d[1]),
    .clkout(net2163));
 b15cbf034ar1n64x5 hold279 (.clk(gen_filter_23__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2164));
 b15cbf034ar1n64x5 hold280 (.clk(gen_filter_25__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2165));
 b15cbf034ar1n64x5 hold281 (.clk(gen_filter_10__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2166));
 b15cbf034ar1n64x5 hold282 (.clk(gen_filter_12__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2167));
 b15cbf034ar1n64x5 hold283 (.clk(gen_filter_1__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2168));
 b15cbf034ar1n64x5 hold284 (.clk(gen_filter_13__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2169));
 b15cbf034ar1n64x5 hold285 (.clk(gen_filter_27__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2170));
 b15cbf034ar1n64x5 hold286 (.clk(gen_filter_6__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2171));
 b15cbf034ar1n64x5 hold287 (.clk(gen_filter_26__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2172));
 b15cbf034ar1n64x5 hold288 (.clk(net151),
    .clkout(net2173));
 b15cbf034ar1n64x5 hold289 (.clk(net159),
    .clkout(net2174));
 b15cbf034ar1n64x5 hold290 (.clk(net251),
    .clkout(net2175));
 b15cbf034ar1n64x5 hold291 (.clk(gen_filter_28__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2176));
 b15cbf034ar1n64x5 hold292 (.clk(gen_filter_23__u_filter_diff_ctr_q[3]),
    .clkout(net2177));
 b15cbf034ar1n64x5 hold293 (.clk(gen_filter_23__u_filter_diff_ctr_d[0]),
    .clkout(net2178));
 b15cbf034ar1n64x5 hold294 (.clk(gen_filter_8__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2179));
 b15cbf034ar1n64x5 hold295 (.clk(gen_filter_15__u_filter_filter_q),
    .clkout(net2180));
 b15cbf034ar1n64x5 hold296 (.clk(n2915),
    .clkout(net2181));
 b15cbf034ar1n64x5 hold297 (.clk(gen_filter_15__u_filter_diff_ctr_d[2]),
    .clkout(net2182));
 b15cbf034ar1n64x5 hold298 (.clk(net164),
    .clkout(net2183));
 b15cbf034ar1n64x5 hold299 (.clk(net176),
    .clkout(net2184));
 b15cbf034ar1n64x5 hold300 (.clk(net637),
    .clkout(net2185));
 b15cbf034ar1n64x5 hold301 (.clk(net253),
    .clkout(net2186));
 b15cbf034ar1n64x5 hold302 (.clk(n3036),
    .clkout(net2187));
 b15cbf034ar1n64x5 hold303 (.clk(net280),
    .clkout(net2188));
 b15cbf034ar1n64x5 hold304 (.clk(gen_filter_24__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2189));
 b15cbf034ar1n64x5 hold305 (.clk(gen_filter_16__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2190));
 b15cbf034ar1n64x5 hold306 (.clk(u_reg_data_in_qs[5]),
    .clkout(net2191));
 b15cbf034ar1n64x5 hold307 (.clk(n3432),
    .clkout(net2192));
 b15cbf034ar1n64x5 hold308 (.clk(n3437),
    .clkout(net2193));
 b15cbf034ar1n64x5 hold309 (.clk(u_reg_u_reg_if_N19),
    .clkout(net2194));
 b15cbf034ar1n64x5 hold310 (.clk(u_reg_data_in_qs[23]),
    .clkout(net2195));
 b15cbf034ar1n64x5 hold311 (.clk(n3969),
    .clkout(net2196));
 b15cbf034ar1n64x5 hold312 (.clk(u_reg_u_reg_if_N37),
    .clkout(net2197));
 b15cbf034ar1n64x5 hold313 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_intq_0_),
    .clkout(net2198));
 b15cbf034ar1n64x5 hold314 (.clk(gen_filter_22__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2199));
 b15cbf034ar1n64x5 hold315 (.clk(net257),
    .clkout(net2200));
 b15cbf034ar1n64x5 hold316 (.clk(net495),
    .clkout(net2201));
 b15cbf034ar1n64x5 hold317 (.clk(gen_filter_15__u_filter_diff_ctr_q[1]),
    .clkout(net2202));
 b15cbf034ar1n64x5 hold318 (.clk(n2916),
    .clkout(net2203));
 b15cbf034ar1n64x5 hold319 (.clk(gen_filter_15__u_filter_diff_ctr_d[1]),
    .clkout(net2204));
 b15cbf034ar1n64x5 hold320 (.clk(u_reg_data_in_qs[22]),
    .clkout(net2205));
 b15cbf034ar1n64x5 hold321 (.clk(n3963),
    .clkout(net2206));
 b15cbf034ar1n64x5 hold322 (.clk(u_reg_u_reg_if_N36),
    .clkout(net2207));
 b15cbf034ar1n64x5 hold323 (.clk(gen_filter_6__u_filter_filter_synced),
    .clkout(net2208));
 b15cbf034ar1n64x5 hold324 (.clk(net262),
    .clkout(net2209));
 b15cbf034ar1n64x5 hold325 (.clk(gen_filter_0__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2210));
 b15cbf034ar1n64x5 hold326 (.clk(net261),
    .clkout(net2211));
 b15cbf034ar1n64x5 hold327 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_intq_0_),
    .clkout(net2212));
 b15cbf034ar1n64x5 hold328 (.clk(gen_filter_9__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2213));
 b15cbf034ar1n64x5 hold329 (.clk(net275),
    .clkout(net2214));
 b15cbf034ar1n64x5 hold330 (.clk(n2988),
    .clkout(net2215));
 b15cbf034ar1n64x5 hold331 (.clk(gen_filter_8__u_filter_filter_synced),
    .clkout(net2216));
 b15cbf034ar1n64x5 hold332 (.clk(net141),
    .clkout(net2217));
 b15cbf034ar1n64x5 hold333 (.clk(net272),
    .clkout(net2218));
 b15cbf034ar1n64x5 hold334 (.clk(net295),
    .clkout(net2219));
 b15cbf034ar1n64x5 hold335 (.clk(reg2hw_intr_enable__q__24_),
    .clkout(net2220));
 b15cbf034ar1n64x5 hold336 (.clk(n3978),
    .clkout(net2221));
 b15cbf034ar1n64x5 hold337 (.clk(u_reg_u_reg_if_N38),
    .clkout(net2222));
 b15cbf034ar1n64x5 hold338 (.clk(data_in_q[15]),
    .clkout(net2223));
 b15cbf034ar1n64x5 hold339 (.clk(gen_filter_7__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2224));
 b15cbf034ar1n64x5 hold340 (.clk(gen_filter_3__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2225));
 b15cbf034ar1n64x5 hold341 (.clk(gen_filter_19__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2226));
 b15cbf034ar1n64x5 hold342 (.clk(reg2hw_intr_enable__q__27_),
    .clkout(net2227));
 b15cbf034ar1n64x5 hold343 (.clk(u_reg_u_reg_if_N41),
    .clkout(net2228));
 b15cbf034ar1n64x5 hold344 (.clk(u_reg_data_in_qs[3]),
    .clkout(net2229));
 b15cbf034ar1n64x5 hold345 (.clk(gen_filter_23__u_filter_stored_value_q),
    .clkout(net2230));
 b15cbf034ar1n64x5 hold346 (.clk(gen_filter_10__u_filter_diff_ctr_q[3]),
    .clkout(net2231));
 b15cbf034ar1n64x5 hold347 (.clk(n2845),
    .clkout(net2232));
 b15cbf034ar1n64x5 hold348 (.clk(gen_filter_10__u_filter_diff_ctr_d[2]),
    .clkout(net2233));
 b15cbf034ar1n64x5 hold349 (.clk(gen_filter_21__u_filter_stored_value_q),
    .clkout(net2234));
 b15cbf034ar1n64x5 hold350 (.clk(net179),
    .clkout(net2235));
 b15cbf034ar1n64x5 hold351 (.clk(reg2hw_intr_state__q__4_),
    .clkout(net2236));
 b15cbf034ar1n64x5 hold352 (.clk(u_reg_u_reg_if_N18),
    .clkout(net2237));
 b15cbf034ar1n64x5 hold353 (.clk(gen_alert_tx_0__u_prim_alert_sender_n1),
    .clkout(net2238));
 b15cbf034ar1n64x5 hold354 (.clk(gen_filter_21__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2239));
 b15cbf034ar1n64x5 hold355 (.clk(net174),
    .clkout(net2240));
 b15cbf034ar1n64x5 hold356 (.clk(gen_filter_24__u_filter_filter_q),
    .clkout(net2241));
 b15cbf034ar1n64x5 hold357 (.clk(gen_filter_24__u_filter_diff_ctr_d[0]),
    .clkout(net2242));
 b15cbf034ar1n64x5 hold358 (.clk(data_in_q[13]),
    .clkout(net2243));
 b15cbf034ar1n64x5 hold359 (.clk(n3785),
    .clkout(net2244));
 b15cbf034ar1n64x5 hold360 (.clk(net199),
    .clkout(net2245));
 b15cbf034ar1n64x5 hold361 (.clk(gen_filter_18__u_filter_stored_value_q),
    .clkout(net2246));
 b15cbf034ar1n64x5 hold362 (.clk(gen_filter_10__u_filter_filter_q),
    .clkout(net2247));
 b15cbf034ar1n64x5 hold363 (.clk(n2840),
    .clkout(net2248));
 b15cbf034ar1n64x5 hold364 (.clk(n2843),
    .clkout(net2249));
 b15cbf034ar1n64x5 hold365 (.clk(gen_filter_10__u_filter_diff_ctr_d[1]),
    .clkout(net2250));
 b15cbf034ar1n64x5 hold366 (.clk(net178),
    .clkout(net2251));
 b15cbf034ar1n64x5 hold367 (.clk(u_reg_data_in_qs[31]),
    .clkout(net2252));
 b15cbf034ar1n64x5 hold368 (.clk(u_reg_u_reg_if_N45),
    .clkout(net2253));
 b15cbf034ar1n64x5 hold369 (.clk(data_in_q[19]),
    .clkout(net2254));
 b15cbf034ar1n64x5 hold370 (.clk(n3771),
    .clkout(net2255));
 b15cbf034ar1n64x5 hold371 (.clk(u_reg_data_in_qs[9]),
    .clkout(net2256));
 b15cbf034ar1n64x5 hold372 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q),
    .clkout(net2257));
 b15cbf034ar1n64x5 hold373 (.clk(gen_filter_10__u_filter_diff_ctr_q[0]),
    .clkout(net2258));
 b15cbf034ar1n64x5 hold374 (.clk(gen_filter_29__u_filter_filter_synced),
    .clkout(net2259));
 b15cbf034ar1n64x5 hold375 (.clk(gen_filter_24__u_filter_diff_ctr_q[2]),
    .clkout(net2260));
 b15cbf034ar1n64x5 hold376 (.clk(n2741),
    .clkout(net2261));
 b15cbf034ar1n64x5 hold377 (.clk(gen_filter_24__u_filter_diff_ctr_d[2]),
    .clkout(net2262));
 b15cbf034ar1n64x5 hold378 (.clk(data_in_q[12]),
    .clkout(net2263));
 b15cbf034ar1n64x5 hold379 (.clk(gen_filter_16__u_filter_stored_value_q),
    .clkout(net2264));
 b15cbf034ar1n64x5 hold380 (.clk(gen_filter_6__u_filter_filter_q),
    .clkout(net2265));
 b15cbf034ar1n64x5 hold381 (.clk(gen_filter_6__u_filter_diff_ctr_d[0]),
    .clkout(net2266));
 b15cbf034ar1n64x5 hold382 (.clk(net152),
    .clkout(net2267));
 b15cbf034ar1n64x5 hold383 (.clk(gen_filter_27__u_filter_stored_value_q),
    .clkout(net2268));
 b15cbf034ar1n64x5 hold384 (.clk(reg2hw_intr_ctrl_en_falling__q__30_),
    .clkout(net2269));
 b15cbf034ar1n64x5 hold385 (.clk(u_reg_u_reg_if_N44),
    .clkout(net2270));
 b15cbf034ar1n64x5 hold386 (.clk(gen_filter_4__u_filter_diff_ctr_q[0]),
    .clkout(net2271));
 b15cbf034ar1n64x5 hold387 (.clk(gen_filter_4__u_filter_diff_ctr_d[1]),
    .clkout(net2272));
 b15cbf034ar1n64x5 hold388 (.clk(gen_filter_10__u_filter_filter_synced),
    .clkout(net2273));
 b15cbf034ar1n64x5 hold389 (.clk(u_reg_data_in_qs[0]),
    .clkout(net2274));
 b15cbf034ar1n64x5 hold390 (.clk(u_reg_data_in_qs[8]),
    .clkout(net2275));
 b15cbf034ar1n64x5 hold391 (.clk(gen_filter_19__u_filter_filter_q),
    .clkout(net2276));
 b15cbf034ar1n64x5 hold392 (.clk(gen_filter_19__u_filter_diff_ctr_d[0]),
    .clkout(net2277));
 b15cbf034ar1n64x5 hold393 (.clk(gen_filter_15__u_filter_filter_synced),
    .clkout(net2278));
 b15cbf034ar1n64x5 hold394 (.clk(gen_filter_9__u_filter_diff_ctr_q[3]),
    .clkout(net2279));
 b15cbf034ar1n64x5 hold395 (.clk(eq_x_136_n25),
    .clkout(net2280));
 b15cbf034ar1n64x5 hold396 (.clk(gen_filter_24__u_filter_diff_ctr_q[3]),
    .clkout(net2281));
 b15cbf034ar1n64x5 hold397 (.clk(gen_filter_22__u_filter_diff_ctr_q[3]),
    .clkout(net2282));
 b15cbf034ar1n64x5 hold398 (.clk(n2835),
    .clkout(net2283));
 b15cbf034ar1n64x5 hold399 (.clk(data_in_q[18]),
    .clkout(net2284));
 b15cbf034ar1n64x5 hold400 (.clk(n3786),
    .clkout(net2285));
 b15cbf034ar1n64x5 hold401 (.clk(gen_filter_31__u_filter_filter_q),
    .clkout(net2286));
 b15cbf034ar1n64x5 hold402 (.clk(gen_filter_31__u_filter_diff_ctr_d[3]),
    .clkout(net2287));
 b15cbf034ar1n64x5 hold403 (.clk(gen_filter_31__u_filter_diff_ctr_q[3]),
    .clkout(net2288));
 b15cbf034ar1n64x5 hold404 (.clk(gen_filter_31__u_filter_diff_ctr_d[2]),
    .clkout(net2289));
 b15cbf034ar1n64x5 hold405 (.clk(gen_filter_4__u_filter_filter_synced),
    .clkout(net2290));
 b15cbf034ar1n64x5 hold406 (.clk(gen_filter_20__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2291));
 b15cbf034ar1n64x5 hold407 (.clk(gen_filter_17__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2292));
 b15cbf034ar1n64x5 hold408 (.clk(gen_filter_17__u_filter_diff_ctr_q[0]),
    .clkout(net2293));
 b15cbf034ar1n64x5 hold409 (.clk(gen_filter_19__u_filter_diff_ctr_q[2]),
    .clkout(net2294));
 b15cbf034ar1n64x5 hold410 (.clk(n2786),
    .clkout(net2295));
 b15cbf034ar1n64x5 hold411 (.clk(gen_filter_19__u_filter_diff_ctr_d[3]),
    .clkout(net2296));
 b15cbf034ar1n64x5 hold412 (.clk(gen_filter_11__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2297));
 b15cbf034ar1n64x5 hold413 (.clk(gen_filter_8__u_filter_filter_q),
    .clkout(net2298));
 b15cbf034ar1n64x5 hold414 (.clk(n2869),
    .clkout(net2299));
 b15cbf034ar1n64x5 hold415 (.clk(gen_filter_8__u_filter_diff_ctr_d[2]),
    .clkout(net2300));
 b15cbf034ar1n64x5 hold416 (.clk(gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q),
    .clkout(net2301));
 b15cbf034ar1n64x5 hold417 (.clk(gen_filter_0__u_filter_filter_q),
    .clkout(net2302));
 b15cbf034ar1n64x5 hold418 (.clk(gen_filter_0__u_filter_diff_ctr_d[3]),
    .clkout(net2303));
 b15cbf034ar1n64x5 hold419 (.clk(gen_filter_0__u_filter_diff_ctr_q[0]),
    .clkout(net2304));
 b15cbf034ar1n64x5 hold420 (.clk(gen_filter_0__u_filter_diff_ctr_d[0]),
    .clkout(net2305));
 b15cbf034ar1n64x5 hold421 (.clk(gen_filter_19__u_filter_diff_ctr_q[2]),
    .clkout(net2306));
 b15cbf034ar1n64x5 hold422 (.clk(gen_filter_22__u_filter_diff_ctr_q[0]),
    .clkout(net2307));
 b15cbf034ar1n64x5 hold423 (.clk(gen_filter_18__u_filter_diff_ctr_q[2]),
    .clkout(net2308));
 b15cbf034ar1n64x5 hold424 (.clk(gen_filter_18__u_filter_diff_ctr_d[2]),
    .clkout(net2309));
 b15cbf034ar1n64x5 hold425 (.clk(gen_filter_4__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2310));
 b15cbf034ar1n64x5 hold426 (.clk(gen_filter_2__u_filter_diff_ctr_q[3]),
    .clkout(net2311));
 b15cbf034ar1n64x5 hold427 (.clk(gen_filter_2__u_filter_diff_ctr_d[0]),
    .clkout(net2312));
 b15cbf034ar1n64x5 hold428 (.clk(gen_filter_26__u_filter_stored_value_q),
    .clkout(net2313));
 b15cbf034ar1n64x5 hold429 (.clk(gen_filter_19__u_filter_diff_ctr_q[3]),
    .clkout(net2314));
 b15cbf034ar1n64x5 hold430 (.clk(u_reg_data_in_qs[10]),
    .clkout(net2315));
 b15cbf034ar1n64x5 hold431 (.clk(n3428),
    .clkout(net2316));
 b15cbf034ar1n64x5 hold432 (.clk(u_reg_u_reg_if_N24),
    .clkout(net2317));
 b15cbf034ar1n64x5 hold433 (.clk(gen_filter_25__u_filter_diff_ctr_q[2]),
    .clkout(net2318));
 b15cbf034ar1n64x5 hold434 (.clk(n2766),
    .clkout(net2319));
 b15cbf034ar1n64x5 hold435 (.clk(gen_filter_25__u_filter_diff_ctr_d[2]),
    .clkout(net2320));
 b15cbf034ar1n64x5 hold436 (.clk(gen_filter_16__u_filter_filter_q),
    .clkout(net2321));
 b15cbf034ar1n64x5 hold437 (.clk(gen_filter_16__u_filter_diff_ctr_d[0]),
    .clkout(net2322));
 b15cbf034ar1n64x5 hold438 (.clk(net200),
    .clkout(net2323));
 b15cbf034ar1n64x5 hold439 (.clk(gen_filter_13__u_filter_filter_q),
    .clkout(net2324));
 b15cbf034ar1n64x5 hold440 (.clk(gen_filter_13__u_filter_diff_ctr_d[1]),
    .clkout(net2325));
 b15cbf034ar1n64x5 hold441 (.clk(gen_filter_8__u_filter_diff_ctr_q[3]),
    .clkout(net2326));
 b15cbf034ar1n64x5 hold442 (.clk(gen_filter_6__u_filter_diff_ctr_q[1]),
    .clkout(net2327));
 b15cbf034ar1n64x5 hold443 (.clk(gen_filter_8__u_filter_diff_ctr_q[1]),
    .clkout(net2328));
 b15cbf034ar1n64x5 hold444 (.clk(gen_filter_2__u_filter_filter_q),
    .clkout(net2329));
 b15cbf034ar1n64x5 hold445 (.clk(gen_filter_27__u_filter_filter_synced),
    .clkout(net2330));
 b15cbf034ar1n64x5 hold446 (.clk(data_in_q[14]),
    .clkout(net2331));
 b15cbf034ar1n64x5 hold447 (.clk(gen_filter_9__u_filter_filter_q),
    .clkout(net2332));
 b15cbf034ar1n64x5 hold448 (.clk(gen_filter_16__u_filter_diff_ctr_q[3]),
    .clkout(net2333));
 b15cbf034ar1n64x5 hold449 (.clk(gen_filter_16__u_filter_diff_ctr_d[3]),
    .clkout(net2334));
 b15cbf034ar1n64x5 hold450 (.clk(gen_filter_8__u_filter_diff_ctr_q[0]),
    .clkout(net2335));
 b15cbf034ar1n64x5 hold451 (.clk(gen_filter_29__u_filter_diff_ctr_q[0]),
    .clkout(net2336));
 b15cbf034ar1n64x5 hold452 (.clk(gen_filter_29__u_filter_diff_ctr_d[0]),
    .clkout(net2337));
 b15cbf034ar1n64x5 hold453 (.clk(gen_filter_3__u_filter_diff_ctr_q[3]),
    .clkout(net2338));
 b15cbf034ar1n64x5 hold454 (.clk(gen_filter_28__u_filter_diff_ctr_q[0]),
    .clkout(net2339));
 b15cbf034ar1n64x5 hold455 (.clk(gen_filter_28__u_filter_diff_ctr_d[0]),
    .clkout(net2340));
 b15cbf034ar1n64x5 hold456 (.clk(gen_filter_7__u_filter_filter_synced),
    .clkout(net2341));
 b15cbf034ar1n64x5 hold457 (.clk(gen_filter_29__u_filter_diff_ctr_q[2]),
    .clkout(net2342));
 b15cbf034ar1n64x5 hold458 (.clk(n2824),
    .clkout(net2343));
 b15cbf034ar1n64x5 hold459 (.clk(gen_filter_29__u_filter_diff_ctr_d[2]),
    .clkout(net2344));
 b15cbf034ar1n64x5 hold460 (.clk(gen_filter_0__u_filter_diff_ctr_q[1]),
    .clkout(net2345));
 b15cbf034ar1n64x5 hold461 (.clk(gen_filter_16__u_filter_diff_ctr_q[1]),
    .clkout(net2346));
 b15cbf034ar1n64x5 hold462 (.clk(gen_filter_16__u_filter_diff_ctr_d[1]),
    .clkout(net2347));
 b15cbf034ar1n64x5 hold463 (.clk(gen_filter_11__u_filter_diff_ctr_q[3]),
    .clkout(net2348));
 b15cbf034ar1n64x5 hold464 (.clk(gen_filter_11__u_filter_diff_ctr_d[3]),
    .clkout(net2349));
 b15cbf034ar1n64x5 hold465 (.clk(reg2hw_intr_ctrl_en_lvllow__q__13_),
    .clkout(net2350));
 b15cbf034ar1n64x5 hold466 (.clk(u_reg_u_reg_if_N27),
    .clkout(net2351));
 b15cbf034ar1n64x5 hold467 (.clk(gen_filter_5__u_filter_diff_ctr_q[0]),
    .clkout(net2352));
 b15cbf034ar1n64x5 hold468 (.clk(gen_filter_5__u_filter_diff_ctr_d[0]),
    .clkout(net2353));
 b15cbf034ar1n64x5 hold469 (.clk(gen_filter_6__u_filter_diff_ctr_q[2]),
    .clkout(net2354));
 b15cbf034ar1n64x5 hold470 (.clk(n2708),
    .clkout(net2355));
 b15cbf034ar1n64x5 hold471 (.clk(gen_filter_18__u_filter_diff_ctr_q[1]),
    .clkout(net2356));
 b15cbf034ar1n64x5 hold472 (.clk(gen_filter_18__u_filter_diff_ctr_d[1]),
    .clkout(net2357));
 b15cbf034ar1n64x5 hold473 (.clk(gen_filter_9__u_filter_diff_ctr_q[2]),
    .clkout(net2358));
 b15cbf034ar1n64x5 hold474 (.clk(gen_filter_20__u_filter_filter_q),
    .clkout(net2359));
 b15cbf034ar1n64x5 hold475 (.clk(gen_filter_12__u_filter_filter_q),
    .clkout(net2360));
 b15cbf034ar1n64x5 hold476 (.clk(gen_filter_12__u_filter_diff_ctr_d[1]),
    .clkout(net2361));
 b15cbf034ar1n64x5 hold477 (.clk(gen_filter_29__u_filter_diff_ctr_q[1]),
    .clkout(net2362));
 b15cbf034ar1n64x5 hold478 (.clk(gen_filter_29__u_filter_diff_ctr_d[1]),
    .clkout(net2363));
 b15cbf034ar1n64x5 hold479 (.clk(gen_filter_13__u_filter_diff_ctr_q[0]),
    .clkout(net2364));
 b15cbf034ar1n64x5 hold480 (.clk(gen_filter_13__u_filter_diff_ctr_d[0]),
    .clkout(net2365));
 b15cbf034ar1n64x5 hold481 (.clk(gen_filter_3__u_filter_diff_ctr_q[0]),
    .clkout(net2366));
 b15cbf034ar1n64x5 hold482 (.clk(gen_filter_8__u_filter_stored_value_q),
    .clkout(net2367));
 b15cbf034ar1n64x5 hold483 (.clk(gen_filter_2__u_filter_diff_ctr_q[2]),
    .clkout(net2368));
 b15cbf034ar1n64x5 hold484 (.clk(gen_filter_1__u_filter_diff_ctr_q[2]),
    .clkout(net2369));
 b15cbf034ar1n64x5 hold485 (.clk(n2859),
    .clkout(net2370));
 b15cbf034ar1n64x5 hold486 (.clk(gen_filter_1__u_filter_diff_ctr_d[2]),
    .clkout(net2371));
 b15cbf034ar1n64x5 hold487 (.clk(gen_filter_25__u_filter_filter_q),
    .clkout(net2372));
 b15cbf034ar1n64x5 hold488 (.clk(gen_filter_25__u_filter_diff_ctr_d[1]),
    .clkout(net2373));
 b15cbf034ar1n64x5 hold489 (.clk(gen_filter_27__u_filter_diff_ctr_q[3]),
    .clkout(net2374));
 b15cbf034ar1n64x5 hold490 (.clk(gen_filter_27__u_filter_diff_ctr_d[3]),
    .clkout(net2375));
 b15cbf034ar1n64x5 hold491 (.clk(reg2hw_intr_ctrl_en_lvlhigh__q__17_),
    .clkout(net2376));
 b15cbf034ar1n64x5 hold492 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd),
    .clkout(net2377));
 b15cbf034ar1n64x5 hold493 (.clk(gen_filter_27__u_filter_filter_q),
    .clkout(net2378));
 b15cbf034ar1n64x5 hold494 (.clk(net193),
    .clkout(net2379));
 b15cbf034ar1n64x5 hold495 (.clk(gen_filter_14__u_filter_filter_synced),
    .clkout(net2380));
 b15cbf034ar1n64x5 hold496 (.clk(gen_filter_26__u_filter_diff_ctr_q[0]),
    .clkout(net2381));
 b15cbf034ar1n64x5 hold497 (.clk(gen_filter_27__u_filter_diff_ctr_q[2]),
    .clkout(net2382));
 b15cbf034ar1n64x5 hold498 (.clk(gen_filter_2__u_filter_diff_ctr_q[2]),
    .clkout(net2383));
 b15cbf034ar1n64x5 hold499 (.clk(gen_filter_27__u_filter_diff_ctr_q[2]),
    .clkout(net2384));
 b15cbf034ar1n64x5 hold500 (.clk(gen_filter_12__u_filter_diff_ctr_q[2]),
    .clkout(net2385));
 b15cbf034ar1n64x5 hold501 (.clk(n2774),
    .clkout(net2386));
 b15cbf034ar1n64x5 hold502 (.clk(gen_filter_1__u_filter_diff_ctr_q[0]),
    .clkout(net2387));
 b15cbf034ar1n64x5 hold503 (.clk(gen_filter_1__u_filter_diff_ctr_d[0]),
    .clkout(net2388));
 b15cbf034ar1n64x5 hold504 (.clk(gen_filter_30__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2389));
 b15cbf034ar1n64x5 hold505 (.clk(gen_filter_21__u_filter_diff_ctr_q[0]),
    .clkout(net2390));
 b15cbf034ar1n64x5 hold506 (.clk(reg2hw_intr_state__q__1_),
    .clkout(net2391));
 b15cbf034ar1n64x5 hold507 (.clk(gen_filter_4__u_filter_filter_q),
    .clkout(net2392));
 b15cbf034ar1n64x5 hold508 (.clk(n2866),
    .clkout(net2393));
 b15cbf034ar1n64x5 hold509 (.clk(gen_filter_4__u_filter_diff_ctr_d[2]),
    .clkout(net2394));
 b15cbf034ar1n64x5 hold510 (.clk(gen_filter_13__u_filter_diff_ctr_q[2]),
    .clkout(net2395));
 b15cbf034ar1n64x5 hold511 (.clk(n2762),
    .clkout(net2396));
 b15cbf034ar1n64x5 hold512 (.clk(gen_filter_30__u_filter_diff_ctr_q[0]),
    .clkout(net2397));
 b15cbf034ar1n64x5 hold513 (.clk(gen_filter_30__u_filter_diff_ctr_d[0]),
    .clkout(net2398));
 b15cbf034ar1n64x5 hold514 (.clk(net188),
    .clkout(net2399));
 b15cbf034ar1n64x5 hold515 (.clk(reg2hw_intr_ctrl_en_lvlhigh__q__26_),
    .clkout(net2400));
 b15cbf034ar1n64x5 hold516 (.clk(u_reg_u_reg_if_N40),
    .clkout(net2401));
 b15cbf034ar1n64x5 hold517 (.clk(gen_filter_0__u_filter_diff_ctr_q[0]),
    .clkout(net2402));
 b15cbf034ar1n64x5 hold518 (.clk(n2772),
    .clkout(net2403));
 b15cbf034ar1n64x5 hold519 (.clk(gen_filter_0__u_filter_diff_ctr_d[2]),
    .clkout(net2404));
 b15cbf034ar1n64x5 hold520 (.clk(gen_filter_11__u_filter_diff_ctr_q[2]),
    .clkout(net2405));
 b15cbf034ar1n64x5 hold521 (.clk(gen_filter_11__u_filter_diff_ctr_d[2]),
    .clkout(net2406));
 b15cbf034ar1n64x5 hold522 (.clk(gen_filter_12__u_filter_diff_ctr_q[3]),
    .clkout(net2407));
 b15cbf034ar1n64x5 hold523 (.clk(gen_filter_12__u_filter_diff_ctr_d[2]),
    .clkout(net2408));
 b15cbf034ar1n64x5 hold524 (.clk(gen_filter_5__u_filter_filter_synced),
    .clkout(net2409));
 b15cbf034ar1n64x5 hold525 (.clk(gen_filter_5__u_filter_diff_ctr_q[3]),
    .clkout(net2410));
 b15cbf034ar1n64x5 hold526 (.clk(gen_filter_5__u_filter_diff_ctr_d[2]),
    .clkout(net2411));
 b15cbf034ar1n64x5 hold527 (.clk(gen_filter_1__u_filter_diff_ctr_q[3]),
    .clkout(net2412));
 b15cbf034ar1n64x5 hold528 (.clk(gen_filter_1__u_filter_diff_ctr_d[1]),
    .clkout(net2413));
 b15cbf034ar1n64x5 hold529 (.clk(gen_filter_30__u_filter_diff_ctr_q[2]),
    .clkout(net2414));
 b15cbf034ar1n64x5 hold530 (.clk(n2828),
    .clkout(net2415));
 b15cbf034ar1n64x5 hold531 (.clk(gen_filter_30__u_filter_diff_ctr_d[1]),
    .clkout(net2416));
 b15cbf034ar1n64x5 hold532 (.clk(gen_filter_18__u_filter_diff_ctr_q[3]),
    .clkout(net2417));
 b15cbf034ar1n64x5 hold533 (.clk(gen_filter_18__u_filter_diff_ctr_d[3]),
    .clkout(net2418));
 b15cbf034ar1n64x5 hold534 (.clk(net187),
    .clkout(net2419));
 b15cbf034ar1n64x5 hold535 (.clk(gen_filter_28__u_filter_diff_ctr_q[2]),
    .clkout(net2420));
 b15cbf034ar1n64x5 hold536 (.clk(gen_filter_28__u_filter_diff_ctr_d[2]),
    .clkout(net2421));
 b15cbf034ar1n64x5 hold537 (.clk(gen_filter_18__u_filter_diff_ctr_q[0]),
    .clkout(net2422));
 b15cbf034ar1n64x5 hold538 (.clk(gen_filter_18__u_filter_diff_ctr_d[0]),
    .clkout(net2423));
 b15cbf034ar1n64x5 hold539 (.clk(gen_filter_10__u_filter_filter_synced),
    .clkout(net2424));
 b15cbf034ar1n64x5 hold540 (.clk(gen_filter_26__u_filter_filter_q),
    .clkout(net2425));
 b15cbf034ar1n64x5 hold541 (.clk(gen_filter_26__u_filter_diff_ctr_d[3]),
    .clkout(net2426));
 b15cbf034ar1n64x5 hold542 (.clk(gen_filter_12__u_filter_diff_ctr_q[0]),
    .clkout(net2427));
 b15cbf034ar1n64x5 hold543 (.clk(gen_filter_12__u_filter_diff_ctr_d[0]),
    .clkout(net2428));
 b15cbf034ar1n64x5 hold544 (.clk(gen_filter_22__u_filter_filter_synced),
    .clkout(net2429));
 b15cbf034ar1n64x5 hold545 (.clk(gen_filter_6__u_filter_stored_value_q),
    .clkout(net2430));
 b15cbf034ar1n64x5 hold546 (.clk(u_reg_data_in_qs[1]),
    .clkout(net2431));
 b15cbf034ar1n64x5 hold547 (.clk(u_reg_u_reg_if_N15),
    .clkout(net2432));
 b15cbf034ar1n64x5 hold548 (.clk(gen_filter_5__u_filter_filter_q),
    .clkout(net2433));
 b15cbf034ar1n64x5 hold549 (.clk(reg2hw_intr_state__q__6_),
    .clkout(net2434));
 b15cbf034ar1n64x5 hold550 (.clk(gen_filter_31__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2435));
 b15cbf034ar1n64x5 hold551 (.clk(gen_filter_25__u_filter_diff_ctr_q[3]),
    .clkout(net2436));
 b15cbf034ar1n64x5 hold552 (.clk(gen_filter_0__u_filter_diff_ctr_q[3]),
    .clkout(net2437));
 b15cbf034ar1n64x5 hold553 (.clk(reg2hw_intr_state__q__10_),
    .clkout(net2438));
 b15cbf034ar1n64x5 hold554 (.clk(net166),
    .clkout(net2439));
 b15cbf034ar1n64x5 hold555 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .clkout(net2440));
 b15cbf034ar1n64x5 hold556 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .clkout(net2441));
 b15cbf034ar1n64x5 hold557 (.clk(gen_filter_14__u_filter_diff_ctr_q[3]),
    .clkout(net2442));
 b15cbf034ar1n64x5 hold558 (.clk(gen_filter_14__u_filter_diff_ctr_d[3]),
    .clkout(net2443));
 b15cbf034ar1n64x5 hold559 (.clk(rst_ni),
    .clkout(net2444));
 b15cbf034ar1n64x5 hold560 (.clk(net163),
    .clkout(net2445));
 b15cbf034ar1n64x5 hold561 (.clk(gen_filter_29__u_filter_stored_value_q),
    .clkout(net2446));
 b15cbf034ar1n64x5 hold562 (.clk(gen_filter_2__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2447));
 b15cbf034ar1n64x5 hold563 (.clk(gen_filter_2__u_filter_diff_ctr_q[2]),
    .clkout(net2448));
 b15cbf034ar1n64x5 hold564 (.clk(gen_filter_15__u_filter_stored_value_q),
    .clkout(net2449));
 b15cbf034ar1n64x5 hold565 (.clk(gen_filter_30__u_filter_diff_ctr_q[3]),
    .clkout(net2450));
 b15cbf034ar1n64x5 hold566 (.clk(gen_filter_22__u_filter_stored_value_q),
    .clkout(net2451));
 b15cbf034ar1n64x5 hold567 (.clk(gen_filter_29__u_filter_diff_ctr_q[3]),
    .clkout(net2452));
 b15cbf034ar1n64x5 hold568 (.clk(reg2hw_intr_state__q__29_),
    .clkout(net2453));
 b15cbf034ar1n64x5 hold569 (.clk(gen_filter_25__u_filter_diff_ctr_q[3]),
    .clkout(net2454));
 b15cbf034ar1n64x5 hold570 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q),
    .clkout(net2455));
 b15cbf034ar1n64x5 hold571 (.clk(gen_filter_6__u_filter_diff_ctr_q[1]),
    .clkout(net2456));
 b15cbf034ar1n64x5 hold572 (.clk(gen_filter_15__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2457));
 b15cbf034ar1n64x5 hold573 (.clk(net189),
    .clkout(net2458));
 b15cbf034ar1n64x5 hold574 (.clk(net186),
    .clkout(net2459));
 b15cbf034ar1n64x5 hold575 (.clk(gen_filter_20__u_filter_stored_value_q),
    .clkout(net2460));
 b15cbf034ar1n64x5 hold576 (.clk(gen_filter_28__u_filter_diff_ctr_q[3]),
    .clkout(net2461));
 b15cbf034ar1n64x5 hold577 (.clk(gen_filter_28__u_filter_diff_ctr_d[1]),
    .clkout(net2462));
 b15cbf034ar1n64x5 hold578 (.clk(gen_filter_26__u_filter_diff_ctr_q[2]),
    .clkout(net2463));
 b15cbf034ar1n64x5 hold579 (.clk(reg2hw_intr_state__q__5_),
    .clkout(net2464));
 b15cbf034ar1n64x5 hold580 (.clk(gen_filter_28__u_filter_stored_value_q),
    .clkout(net2465));
 b15cbf034ar1n64x5 hold581 (.clk(gen_filter_25__u_filter_stored_value_q),
    .clkout(net2466));
 b15cbf034ar1n64x5 hold582 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[0]),
    .clkout(net2467));
 b15cbf034ar1n64x5 hold583 (.clk(gen_filter_1__u_filter_filter_synced),
    .clkout(net2468));
 b15cbf034ar1n64x5 hold584 (.clk(gen_filter_26__u_filter_diff_ctr_q[0]),
    .clkout(net2469));
 b15cbf034ar1n64x5 hold585 (.clk(gen_filter_1__u_filter_diff_ctr_q[3]),
    .clkout(net2470));
 b15cbf034ar1n64x5 hold586 (.clk(gen_filter_13__u_filter_filter_synced),
    .clkout(net2471));
 b15cbf034ar1n64x5 hold587 (.clk(u_reg_err_q),
    .clkout(net2472));
 b15cbf034ar1n64x5 hold588 (.clk(gen_filter_21__u_filter_diff_ctr_q[3]),
    .clkout(net2473));
 b15cbf034ar1n64x5 hold589 (.clk(reg2hw_intr_enable__q__30_),
    .clkout(net2474));
 b15cbf034ar1n64x5 hold590 (.clk(data_in_q[16]),
    .clkout(net2475));
 b15cbf034ar1n64x5 hold591 (.clk(gen_filter_30__u_filter_filter_synced),
    .clkout(net2476));
 b15cbf034ar1n64x5 hold592 (.clk(net147),
    .clkout(net2477));
 b15cbf034ar1n64x5 hold593 (.clk(gen_filter_7__u_filter_diff_ctr_q[3]),
    .clkout(net2478));
 b15cbf034ar1n64x5 hold594 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .clkout(net2479));
 b15cbf034ar1n64x5 hold595 (.clk(gen_filter_9__u_filter_stored_value_q),
    .clkout(net2480));
 b15cbf034ar1n64x5 hold596 (.clk(gen_filter_2__u_filter_stored_value_q),
    .clkout(net2481));
 b15cbf034ar1n64x5 hold597 (.clk(net213),
    .clkout(net2482));
 b15cbf034ar1n64x5 hold598 (.clk(net1886),
    .clkout(net2483));
 b15cbf034ar1n64x5 hold599 (.clk(net1887),
    .clkout(net2484));
 b15cbf034ar1n64x5 hold600 (.clk(net212),
    .clkout(net2485));
 b15cbf034ar1n64x5 hold601 (.clk(net1888),
    .clkout(net2486));
 b15cbf034ar1n64x5 hold602 (.clk(net1889),
    .clkout(net2487));
 b15cbf034ar1n64x5 hold603 (.clk(net220),
    .clkout(net2488));
 b15cbf034ar1n64x5 hold604 (.clk(net1890),
    .clkout(net2489));
 b15cbf034ar1n64x5 hold605 (.clk(net219),
    .clkout(net2490));
 b15cbf034ar1n64x5 hold606 (.clk(net1892),
    .clkout(net2491));
 b15cbf034ar1n64x5 hold607 (.clk(net226),
    .clkout(net2492));
 b15cbf034ar1n64x5 hold608 (.clk(net1894),
    .clkout(net2493));
 b15cbf034ar1n64x5 hold609 (.clk(net225),
    .clkout(net2494));
 b15cbf034ar1n64x5 hold610 (.clk(net1896),
    .clkout(net2495));
 b15cbf034ar1n64x5 hold611 (.clk(net227),
    .clkout(net2496));
 b15cbf034ar1n64x5 hold612 (.clk(net1898),
    .clkout(net2497));
 b15cbf034ar1n64x5 hold613 (.clk(net216),
    .clkout(net2498));
 b15cbf034ar1n64x5 hold614 (.clk(net1900),
    .clkout(net2499));
 b15cbf034ar1n64x5 hold615 (.clk(net209),
    .clkout(net2500));
 b15cbf034ar1n64x5 hold616 (.clk(net1908),
    .clkout(net2501));
 b15cbf034ar1n64x5 hold617 (.clk(net214),
    .clkout(net2502));
 b15cbf034ar1n64x5 hold618 (.clk(net1906),
    .clkout(net2503));
 b15cbf034ar1n64x5 hold619 (.clk(net208),
    .clkout(net2504));
 b15cbf034ar1n64x5 hold620 (.clk(net1910),
    .clkout(net2505));
 b15cbf034ar1n64x5 hold621 (.clk(net235),
    .clkout(net2506));
 b15cbf034ar1n64x5 hold622 (.clk(net1912),
    .clkout(net2507));
 b15cbf034ar1n64x5 hold623 (.clk(net230),
    .clkout(net2508));
 b15cbf034ar1n64x5 hold624 (.clk(net1914),
    .clkout(net2509));
 b15cbf034ar1n64x5 hold625 (.clk(net228),
    .clkout(net2510));
 b15cbf034ar1n64x5 hold626 (.clk(net1902),
    .clkout(net2511));
 b15cbf034ar1n64x5 hold627 (.clk(net218),
    .clkout(net2512));
 b15cbf034ar1n64x5 hold628 (.clk(net1904),
    .clkout(net2513));
 b15cbf034ar1n64x5 hold629 (.clk(net140),
    .clkout(net2514));
 b15cbf034ar1n64x5 hold630 (.clk(net1916),
    .clkout(net2515));
 b15cbf034ar1n64x5 hold631 (.clk(net139),
    .clkout(net2516));
 b15cbf034ar1n64x5 hold632 (.clk(net1921),
    .clkout(net2517));
 b15cbf034ar1n64x5 hold633 (.clk(net231),
    .clkout(net2518));
 b15cbf034ar1n64x5 hold634 (.clk(net1925),
    .clkout(net2519));
 b15cbf034ar1n64x5 hold635 (.clk(net205),
    .clkout(net2520));
 b15cbf034ar1n64x5 hold636 (.clk(net1923),
    .clkout(net2521));
 b15cbf034ar1n64x5 hold637 (.clk(net232),
    .clkout(net2522));
 b15cbf034ar1n64x5 hold638 (.clk(net1927),
    .clkout(net2523));
 b15cbf034ar1n64x5 hold639 (.clk(net236),
    .clkout(net2524));
 b15cbf034ar1n64x5 hold640 (.clk(net1929),
    .clkout(net2525));
 b15cbf034ar1n64x5 hold641 (.clk(net215),
    .clkout(net2526));
 b15cbf034ar1n64x5 hold642 (.clk(net1931),
    .clkout(net2527));
 b15cbf034ar1n64x5 hold643 (.clk(net206),
    .clkout(net2528));
 b15cbf034ar1n64x5 hold644 (.clk(net1935),
    .clkout(net2529));
 b15cbf034ar1n64x5 hold645 (.clk(net217),
    .clkout(net2530));
 b15cbf034ar1n64x5 hold646 (.clk(net1933),
    .clkout(net2531));
 b15cbf034ar1n64x5 hold647 (.clk(net207),
    .clkout(net2532));
 b15cbf034ar1n64x5 hold648 (.clk(net1942),
    .clkout(net2533));
 b15cbf034ar1n64x5 hold649 (.clk(net229),
    .clkout(net2534));
 b15cbf034ar1n64x5 hold650 (.clk(net1944),
    .clkout(net2535));
 b15cbf034ar1n64x5 hold651 (.clk(net211),
    .clkout(net2536));
 b15cbf034ar1n64x5 hold652 (.clk(net210),
    .clkout(net2537));
 b15cbf034ar1n64x5 hold653 (.clk(net221),
    .clkout(net2538));
 b15cbf034ar1n64x5 hold654 (.clk(net222),
    .clkout(net2539));
 b15cbf034ar1n64x5 hold655 (.clk(net223),
    .clkout(net2540));
 b15cbf034ar1n64x5 hold656 (.clk(net224),
    .clkout(net2541));
 b15cbf034ar1n64x5 hold657 (.clk(net285),
    .clkout(net2542));
 b15cbf034ar1n64x5 hold658 (.clk(net284),
    .clkout(net2543));
 b15cbf034ar1n64x5 hold659 (.clk(net283),
    .clkout(net2544));
 b15cbf034ar1n64x5 hold660 (.clk(net282),
    .clkout(net2545));
 b15cbf034ar1n64x5 hold661 (.clk(net281),
    .clkout(net2546));
 b15cbf034ar1n64x5 hold662 (.clk(net279),
    .clkout(net2547));
 b15cbf034ar1n64x5 hold663 (.clk(net287),
    .clkout(net2548));
 b15cbf034ar1n64x5 hold664 (.clk(net286),
    .clkout(net2549));
 b15cbf034ar1n64x5 hold665 (.clk(net233),
    .clkout(net2550));
 b15cbf034ar1n64x5 hold666 (.clk(net234),
    .clkout(net2551));
 b15cbf034ar1n64x5 hold667 (.clk(reg2hw_intr_ctrl_en_lvlhigh__q__19_),
    .clkout(net2552));
 b15cbf034ar1n64x5 hold668 (.clk(gen_filter_22__u_filter_diff_ctr_q[3]),
    .clkout(net2553));
 b15cbf034ar1n64x5 hold669 (.clk(net186),
    .clkout(net2554));
 b15cbf034ar1n64x5 hold670 (.clk(net267),
    .clkout(net2555));
 b15cbf034ar1n64x5 hold671 (.clk(net266),
    .clkout(net2556));
 b15cbf034ar1n64x5 hold672 (.clk(net276),
    .clkout(net2557));
 b15cbf034ar1n64x5 hold673 (.clk(net155),
    .clkout(net2558));
 b15cbf034ar1n64x5 hold674 (.clk(net188),
    .clkout(net2559));
 b15cbf034ar1n64x5 hold675 (.clk(gen_filter_7__u_filter_diff_ctr_q[3]),
    .clkout(net2560));
 b15cbf034ar1n64x5 hold676 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_intq_0_),
    .clkout(net2561));
 b15cbf034ar1n64x5 hold677 (.clk(gen_filter_28__u_filter_diff_ctr_q[2]),
    .clkout(net2562));
 b15cbf034ar1n64x5 hold678 (.clk(u_reg_data_in_qs[29]),
    .clkout(net2563));
 b15cbf034ar1n64x5 hold679 (.clk(net274),
    .clkout(net2564));
 b15cbf034ar1n64x5 hold680 (.clk(gen_filter_22__u_filter_diff_ctr_q[0]),
    .clkout(net2565));
 b15cbf034ar1n64x5 hold681 (.clk(gen_filter_6__u_filter_diff_ctr_q[1]),
    .clkout(net2566));
 b15cbf034ar1n64x5 hold682 (.clk(gen_filter_0__u_filter_diff_ctr_q[0]),
    .clkout(net2567));
 b15cbf034ar1n64x5 hold683 (.clk(gen_filter_24__u_filter_diff_ctr_q[2]),
    .clkout(net2568));
 b15cbf034ar1n64x5 hold684 (.clk(gen_filter_7__u_filter_diff_ctr_q[3]),
    .clkout(net2569));
 b15cbf034ar1n64x5 hold685 (.clk(gen_filter_6__u_filter_diff_ctr_q[1]),
    .clkout(net2570));
 b15zdnd11an1n64x5 FILLER_0_8 ();
 b15zdnd11an1n64x5 FILLER_0_72 ();
 b15zdnd11an1n64x5 FILLER_0_136 ();
 b15zdnd11an1n64x5 FILLER_0_200 ();
 b15zdnd11an1n64x5 FILLER_0_264 ();
 b15zdnd11an1n64x5 FILLER_0_328 ();
 b15zdnd11an1n64x5 FILLER_0_392 ();
 b15zdnd11an1n64x5 FILLER_0_456 ();
 b15zdnd11an1n64x5 FILLER_0_520 ();
 b15zdnd11an1n08x5 FILLER_0_584 ();
 b15zdnd00an1n02x5 FILLER_0_592 ();
 b15zdnd11an1n08x5 FILLER_0_598 ();
 b15zdnd00an1n01x5 FILLER_0_606 ();
 b15zdnd11an1n08x5 FILLER_0_611 ();
 b15zdnd11an1n04x5 FILLER_0_619 ();
 b15zdnd00an1n01x5 FILLER_0_623 ();
 b15zdnd11an1n32x5 FILLER_0_629 ();
 b15zdnd11an1n04x5 FILLER_0_661 ();
 b15zdnd00an1n02x5 FILLER_0_665 ();
 b15zdnd00an1n01x5 FILLER_0_667 ();
 b15zdnd11an1n32x5 FILLER_0_673 ();
 b15zdnd11an1n08x5 FILLER_0_705 ();
 b15zdnd11an1n04x5 FILLER_0_713 ();
 b15zdnd00an1n01x5 FILLER_0_717 ();
 b15zdnd11an1n64x5 FILLER_0_726 ();
 b15zdnd11an1n32x5 FILLER_0_790 ();
 b15zdnd11an1n16x5 FILLER_0_822 ();
 b15zdnd11an1n08x5 FILLER_0_838 ();
 b15zdnd11an1n08x5 FILLER_0_888 ();
 b15zdnd00an1n02x5 FILLER_0_896 ();
 b15zdnd11an1n08x5 FILLER_0_940 ();
 b15zdnd00an1n02x5 FILLER_0_948 ();
 b15zdnd11an1n08x5 FILLER_0_992 ();
 b15zdnd00an1n01x5 FILLER_0_1000 ();
 b15zdnd11an1n64x5 FILLER_0_1043 ();
 b15zdnd00an1n01x5 FILLER_0_1107 ();
 b15zdnd11an1n04x5 FILLER_0_1112 ();
 b15zdnd00an1n01x5 FILLER_0_1116 ();
 b15zdnd11an1n04x5 FILLER_0_1128 ();
 b15zdnd11an1n32x5 FILLER_0_1174 ();
 b15zdnd11an1n08x5 FILLER_0_1206 ();
 b15zdnd00an1n01x5 FILLER_0_1214 ();
 b15zdnd11an1n16x5 FILLER_0_1220 ();
 b15zdnd11an1n08x5 FILLER_0_1236 ();
 b15zdnd11an1n04x5 FILLER_0_1248 ();
 b15zdnd00an1n02x5 FILLER_0_1252 ();
 b15zdnd00an1n01x5 FILLER_0_1254 ();
 b15zdnd11an1n04x5 FILLER_0_1259 ();
 b15zdnd11an1n04x5 FILLER_0_1305 ();
 b15zdnd11an1n16x5 FILLER_0_1351 ();
 b15zdnd11an1n08x5 FILLER_0_1367 ();
 b15zdnd00an1n02x5 FILLER_0_1375 ();
 b15zdnd00an1n01x5 FILLER_0_1377 ();
 b15zdnd11an1n16x5 FILLER_0_1383 ();
 b15zdnd11an1n04x5 FILLER_0_1399 ();
 b15zdnd00an1n02x5 FILLER_0_1403 ();
 b15zdnd00an1n01x5 FILLER_0_1405 ();
 b15zdnd11an1n16x5 FILLER_0_1410 ();
 b15zdnd11an1n04x5 FILLER_0_1426 ();
 b15zdnd00an1n02x5 FILLER_0_1434 ();
 b15zdnd00an1n02x5 FILLER_0_1444 ();
 b15zdnd00an1n01x5 FILLER_0_1446 ();
 b15zdnd11an1n16x5 FILLER_0_1451 ();
 b15zdnd11an1n08x5 FILLER_0_1467 ();
 b15zdnd00an1n01x5 FILLER_0_1475 ();
 b15zdnd11an1n16x5 FILLER_0_1518 ();
 b15zdnd00an1n01x5 FILLER_0_1534 ();
 b15zdnd11an1n64x5 FILLER_0_1540 ();
 b15zdnd11an1n08x5 FILLER_0_1604 ();
 b15zdnd00an1n01x5 FILLER_0_1612 ();
 b15zdnd11an1n64x5 FILLER_0_1617 ();
 b15zdnd11an1n64x5 FILLER_0_1681 ();
 b15zdnd11an1n64x5 FILLER_0_1745 ();
 b15zdnd11an1n16x5 FILLER_0_1809 ();
 b15zdnd00an1n01x5 FILLER_0_1825 ();
 b15zdnd11an1n04x5 FILLER_0_1831 ();
 b15zdnd00an1n02x5 FILLER_0_1835 ();
 b15zdnd11an1n64x5 FILLER_0_1844 ();
 b15zdnd11an1n64x5 FILLER_0_1908 ();
 b15zdnd11an1n64x5 FILLER_0_1972 ();
 b15zdnd11an1n64x5 FILLER_0_2036 ();
 b15zdnd11an1n32x5 FILLER_0_2100 ();
 b15zdnd11an1n16x5 FILLER_0_2132 ();
 b15zdnd11an1n04x5 FILLER_0_2148 ();
 b15zdnd00an1n02x5 FILLER_0_2152 ();
 b15zdnd11an1n64x5 FILLER_0_2162 ();
 b15zdnd11an1n32x5 FILLER_0_2226 ();
 b15zdnd11an1n16x5 FILLER_0_2258 ();
 b15zdnd00an1n02x5 FILLER_0_2274 ();
 b15zdnd11an1n64x5 FILLER_1_0 ();
 b15zdnd11an1n64x5 FILLER_1_64 ();
 b15zdnd11an1n64x5 FILLER_1_128 ();
 b15zdnd11an1n64x5 FILLER_1_192 ();
 b15zdnd11an1n64x5 FILLER_1_256 ();
 b15zdnd11an1n64x5 FILLER_1_320 ();
 b15zdnd11an1n64x5 FILLER_1_384 ();
 b15zdnd11an1n64x5 FILLER_1_448 ();
 b15zdnd11an1n64x5 FILLER_1_512 ();
 b15zdnd11an1n64x5 FILLER_1_576 ();
 b15zdnd11an1n64x5 FILLER_1_640 ();
 b15zdnd11an1n64x5 FILLER_1_704 ();
 b15zdnd11an1n64x5 FILLER_1_768 ();
 b15zdnd11an1n08x5 FILLER_1_832 ();
 b15zdnd11an1n04x5 FILLER_1_840 ();
 b15zdnd00an1n02x5 FILLER_1_844 ();
 b15zdnd00an1n01x5 FILLER_1_846 ();
 b15zdnd11an1n16x5 FILLER_1_851 ();
 b15zdnd00an1n02x5 FILLER_1_867 ();
 b15zdnd11an1n04x5 FILLER_1_895 ();
 b15zdnd11an1n04x5 FILLER_1_903 ();
 b15zdnd00an1n02x5 FILLER_1_907 ();
 b15zdnd11an1n16x5 FILLER_1_913 ();
 b15zdnd11an1n08x5 FILLER_1_929 ();
 b15zdnd00an1n02x5 FILLER_1_937 ();
 b15zdnd00an1n01x5 FILLER_1_939 ();
 b15zdnd11an1n04x5 FILLER_1_944 ();
 b15zdnd11an1n04x5 FILLER_1_952 ();
 b15zdnd11an1n32x5 FILLER_1_961 ();
 b15zdnd11an1n08x5 FILLER_1_993 ();
 b15zdnd11an1n04x5 FILLER_1_1005 ();
 b15zdnd00an1n02x5 FILLER_1_1009 ();
 b15zdnd11an1n04x5 FILLER_1_1031 ();
 b15zdnd11an1n64x5 FILLER_1_1039 ();
 b15zdnd11an1n08x5 FILLER_1_1103 ();
 b15zdnd11an1n04x5 FILLER_1_1125 ();
 b15zdnd11an1n16x5 FILLER_1_1133 ();
 b15zdnd00an1n01x5 FILLER_1_1149 ();
 b15zdnd11an1n04x5 FILLER_1_1154 ();
 b15zdnd11an1n64x5 FILLER_1_1163 ();
 b15zdnd11an1n32x5 FILLER_1_1227 ();
 b15zdnd00an1n01x5 FILLER_1_1259 ();
 b15zdnd11an1n32x5 FILLER_1_1264 ();
 b15zdnd11an1n08x5 FILLER_1_1296 ();
 b15zdnd11an1n04x5 FILLER_1_1308 ();
 b15zdnd11an1n16x5 FILLER_1_1316 ();
 b15zdnd00an1n01x5 FILLER_1_1332 ();
 b15zdnd11an1n32x5 FILLER_1_1375 ();
 b15zdnd11an1n16x5 FILLER_1_1407 ();
 b15zdnd11an1n04x5 FILLER_1_1423 ();
 b15zdnd00an1n01x5 FILLER_1_1427 ();
 b15zdnd11an1n08x5 FILLER_1_1470 ();
 b15zdnd11an1n64x5 FILLER_1_1482 ();
 b15zdnd11an1n64x5 FILLER_1_1546 ();
 b15zdnd11an1n64x5 FILLER_1_1610 ();
 b15zdnd11an1n64x5 FILLER_1_1674 ();
 b15zdnd11an1n64x5 FILLER_1_1738 ();
 b15zdnd11an1n64x5 FILLER_1_1802 ();
 b15zdnd11an1n64x5 FILLER_1_1866 ();
 b15zdnd11an1n64x5 FILLER_1_1930 ();
 b15zdnd11an1n64x5 FILLER_1_1994 ();
 b15zdnd11an1n64x5 FILLER_1_2058 ();
 b15zdnd11an1n64x5 FILLER_1_2122 ();
 b15zdnd11an1n64x5 FILLER_1_2186 ();
 b15zdnd11an1n32x5 FILLER_1_2250 ();
 b15zdnd00an1n02x5 FILLER_1_2282 ();
 b15zdnd11an1n64x5 FILLER_2_8 ();
 b15zdnd11an1n64x5 FILLER_2_72 ();
 b15zdnd11an1n64x5 FILLER_2_136 ();
 b15zdnd11an1n64x5 FILLER_2_200 ();
 b15zdnd11an1n64x5 FILLER_2_264 ();
 b15zdnd11an1n64x5 FILLER_2_328 ();
 b15zdnd11an1n64x5 FILLER_2_392 ();
 b15zdnd11an1n64x5 FILLER_2_456 ();
 b15zdnd11an1n64x5 FILLER_2_520 ();
 b15zdnd11an1n64x5 FILLER_2_584 ();
 b15zdnd11an1n64x5 FILLER_2_648 ();
 b15zdnd11an1n04x5 FILLER_2_712 ();
 b15zdnd00an1n02x5 FILLER_2_716 ();
 b15zdnd11an1n64x5 FILLER_2_726 ();
 b15zdnd11an1n64x5 FILLER_2_790 ();
 b15zdnd11an1n64x5 FILLER_2_854 ();
 b15zdnd11an1n64x5 FILLER_2_918 ();
 b15zdnd11an1n64x5 FILLER_2_982 ();
 b15zdnd11an1n64x5 FILLER_2_1046 ();
 b15zdnd11an1n32x5 FILLER_2_1110 ();
 b15zdnd11an1n04x5 FILLER_2_1142 ();
 b15zdnd00an1n02x5 FILLER_2_1146 ();
 b15zdnd11an1n64x5 FILLER_2_1152 ();
 b15zdnd11an1n64x5 FILLER_2_1216 ();
 b15zdnd11an1n32x5 FILLER_2_1280 ();
 b15zdnd11an1n16x5 FILLER_2_1312 ();
 b15zdnd00an1n02x5 FILLER_2_1328 ();
 b15zdnd00an1n01x5 FILLER_2_1330 ();
 b15zdnd11an1n64x5 FILLER_2_1335 ();
 b15zdnd11an1n32x5 FILLER_2_1399 ();
 b15zdnd11an1n64x5 FILLER_2_1435 ();
 b15zdnd11an1n64x5 FILLER_2_1499 ();
 b15zdnd11an1n64x5 FILLER_2_1563 ();
 b15zdnd11an1n64x5 FILLER_2_1627 ();
 b15zdnd11an1n64x5 FILLER_2_1691 ();
 b15zdnd11an1n64x5 FILLER_2_1755 ();
 b15zdnd11an1n64x5 FILLER_2_1819 ();
 b15zdnd11an1n64x5 FILLER_2_1883 ();
 b15zdnd11an1n64x5 FILLER_2_1947 ();
 b15zdnd11an1n64x5 FILLER_2_2011 ();
 b15zdnd11an1n64x5 FILLER_2_2075 ();
 b15zdnd11an1n08x5 FILLER_2_2139 ();
 b15zdnd11an1n04x5 FILLER_2_2147 ();
 b15zdnd00an1n02x5 FILLER_2_2151 ();
 b15zdnd00an1n01x5 FILLER_2_2153 ();
 b15zdnd11an1n64x5 FILLER_2_2162 ();
 b15zdnd11an1n32x5 FILLER_2_2226 ();
 b15zdnd11an1n16x5 FILLER_2_2258 ();
 b15zdnd00an1n02x5 FILLER_2_2274 ();
 b15zdnd11an1n64x5 FILLER_3_0 ();
 b15zdnd11an1n64x5 FILLER_3_64 ();
 b15zdnd11an1n64x5 FILLER_3_128 ();
 b15zdnd11an1n64x5 FILLER_3_192 ();
 b15zdnd11an1n64x5 FILLER_3_256 ();
 b15zdnd11an1n64x5 FILLER_3_320 ();
 b15zdnd11an1n64x5 FILLER_3_384 ();
 b15zdnd11an1n64x5 FILLER_3_448 ();
 b15zdnd11an1n64x5 FILLER_3_512 ();
 b15zdnd11an1n64x5 FILLER_3_576 ();
 b15zdnd11an1n64x5 FILLER_3_640 ();
 b15zdnd11an1n64x5 FILLER_3_704 ();
 b15zdnd11an1n64x5 FILLER_3_768 ();
 b15zdnd11an1n64x5 FILLER_3_832 ();
 b15zdnd11an1n64x5 FILLER_3_896 ();
 b15zdnd11an1n64x5 FILLER_3_960 ();
 b15zdnd11an1n64x5 FILLER_3_1024 ();
 b15zdnd11an1n64x5 FILLER_3_1088 ();
 b15zdnd11an1n64x5 FILLER_3_1152 ();
 b15zdnd11an1n64x5 FILLER_3_1216 ();
 b15zdnd11an1n64x5 FILLER_3_1280 ();
 b15zdnd11an1n64x5 FILLER_3_1344 ();
 b15zdnd11an1n64x5 FILLER_3_1408 ();
 b15zdnd11an1n64x5 FILLER_3_1472 ();
 b15zdnd11an1n64x5 FILLER_3_1536 ();
 b15zdnd11an1n64x5 FILLER_3_1600 ();
 b15zdnd11an1n64x5 FILLER_3_1664 ();
 b15zdnd11an1n64x5 FILLER_3_1728 ();
 b15zdnd11an1n64x5 FILLER_3_1792 ();
 b15zdnd11an1n64x5 FILLER_3_1856 ();
 b15zdnd11an1n64x5 FILLER_3_1920 ();
 b15zdnd11an1n64x5 FILLER_3_1984 ();
 b15zdnd11an1n64x5 FILLER_3_2048 ();
 b15zdnd11an1n64x5 FILLER_3_2112 ();
 b15zdnd11an1n64x5 FILLER_3_2176 ();
 b15zdnd11an1n32x5 FILLER_3_2240 ();
 b15zdnd11an1n08x5 FILLER_3_2272 ();
 b15zdnd11an1n04x5 FILLER_3_2280 ();
 b15zdnd11an1n64x5 FILLER_4_8 ();
 b15zdnd11an1n64x5 FILLER_4_72 ();
 b15zdnd11an1n64x5 FILLER_4_136 ();
 b15zdnd11an1n64x5 FILLER_4_200 ();
 b15zdnd11an1n64x5 FILLER_4_264 ();
 b15zdnd11an1n64x5 FILLER_4_328 ();
 b15zdnd11an1n64x5 FILLER_4_392 ();
 b15zdnd11an1n64x5 FILLER_4_456 ();
 b15zdnd11an1n64x5 FILLER_4_520 ();
 b15zdnd11an1n64x5 FILLER_4_584 ();
 b15zdnd11an1n64x5 FILLER_4_648 ();
 b15zdnd11an1n04x5 FILLER_4_712 ();
 b15zdnd00an1n02x5 FILLER_4_716 ();
 b15zdnd11an1n64x5 FILLER_4_726 ();
 b15zdnd11an1n64x5 FILLER_4_790 ();
 b15zdnd11an1n64x5 FILLER_4_854 ();
 b15zdnd11an1n64x5 FILLER_4_918 ();
 b15zdnd11an1n64x5 FILLER_4_982 ();
 b15zdnd11an1n64x5 FILLER_4_1046 ();
 b15zdnd11an1n16x5 FILLER_4_1110 ();
 b15zdnd11an1n08x5 FILLER_4_1126 ();
 b15zdnd11an1n64x5 FILLER_4_1176 ();
 b15zdnd11an1n64x5 FILLER_4_1240 ();
 b15zdnd11an1n64x5 FILLER_4_1304 ();
 b15zdnd11an1n64x5 FILLER_4_1368 ();
 b15zdnd11an1n64x5 FILLER_4_1432 ();
 b15zdnd11an1n64x5 FILLER_4_1496 ();
 b15zdnd11an1n64x5 FILLER_4_1560 ();
 b15zdnd11an1n64x5 FILLER_4_1624 ();
 b15zdnd11an1n64x5 FILLER_4_1688 ();
 b15zdnd11an1n64x5 FILLER_4_1752 ();
 b15zdnd11an1n64x5 FILLER_4_1816 ();
 b15zdnd11an1n64x5 FILLER_4_1880 ();
 b15zdnd11an1n64x5 FILLER_4_1944 ();
 b15zdnd11an1n64x5 FILLER_4_2008 ();
 b15zdnd11an1n64x5 FILLER_4_2072 ();
 b15zdnd11an1n16x5 FILLER_4_2136 ();
 b15zdnd00an1n02x5 FILLER_4_2152 ();
 b15zdnd11an1n64x5 FILLER_4_2162 ();
 b15zdnd11an1n32x5 FILLER_4_2226 ();
 b15zdnd11an1n16x5 FILLER_4_2258 ();
 b15zdnd00an1n02x5 FILLER_4_2274 ();
 b15zdnd11an1n64x5 FILLER_5_0 ();
 b15zdnd11an1n64x5 FILLER_5_64 ();
 b15zdnd11an1n64x5 FILLER_5_128 ();
 b15zdnd11an1n64x5 FILLER_5_192 ();
 b15zdnd11an1n64x5 FILLER_5_256 ();
 b15zdnd11an1n64x5 FILLER_5_320 ();
 b15zdnd11an1n64x5 FILLER_5_384 ();
 b15zdnd11an1n64x5 FILLER_5_448 ();
 b15zdnd11an1n64x5 FILLER_5_512 ();
 b15zdnd11an1n64x5 FILLER_5_576 ();
 b15zdnd11an1n64x5 FILLER_5_640 ();
 b15zdnd11an1n64x5 FILLER_5_704 ();
 b15zdnd11an1n64x5 FILLER_5_768 ();
 b15zdnd11an1n16x5 FILLER_5_832 ();
 b15zdnd11an1n08x5 FILLER_5_848 ();
 b15zdnd11an1n04x5 FILLER_5_856 ();
 b15zdnd00an1n01x5 FILLER_5_860 ();
 b15zdnd11an1n08x5 FILLER_5_903 ();
 b15zdnd11an1n64x5 FILLER_5_953 ();
 b15zdnd11an1n64x5 FILLER_5_1017 ();
 b15zdnd11an1n64x5 FILLER_5_1081 ();
 b15zdnd11an1n16x5 FILLER_5_1145 ();
 b15zdnd11an1n04x5 FILLER_5_1161 ();
 b15zdnd00an1n02x5 FILLER_5_1165 ();
 b15zdnd11an1n32x5 FILLER_5_1209 ();
 b15zdnd11an1n16x5 FILLER_5_1241 ();
 b15zdnd11an1n04x5 FILLER_5_1257 ();
 b15zdnd00an1n02x5 FILLER_5_1261 ();
 b15zdnd00an1n01x5 FILLER_5_1263 ();
 b15zdnd11an1n04x5 FILLER_5_1306 ();
 b15zdnd11an1n08x5 FILLER_5_1352 ();
 b15zdnd11an1n04x5 FILLER_5_1360 ();
 b15zdnd00an1n02x5 FILLER_5_1364 ();
 b15zdnd11an1n64x5 FILLER_5_1408 ();
 b15zdnd11an1n64x5 FILLER_5_1472 ();
 b15zdnd11an1n64x5 FILLER_5_1536 ();
 b15zdnd11an1n64x5 FILLER_5_1600 ();
 b15zdnd11an1n64x5 FILLER_5_1664 ();
 b15zdnd11an1n64x5 FILLER_5_1728 ();
 b15zdnd11an1n64x5 FILLER_5_1792 ();
 b15zdnd11an1n64x5 FILLER_5_1856 ();
 b15zdnd11an1n64x5 FILLER_5_1920 ();
 b15zdnd11an1n64x5 FILLER_5_1984 ();
 b15zdnd11an1n64x5 FILLER_5_2048 ();
 b15zdnd11an1n64x5 FILLER_5_2112 ();
 b15zdnd11an1n64x5 FILLER_5_2176 ();
 b15zdnd11an1n32x5 FILLER_5_2240 ();
 b15zdnd11an1n08x5 FILLER_5_2272 ();
 b15zdnd11an1n04x5 FILLER_5_2280 ();
 b15zdnd11an1n64x5 FILLER_6_8 ();
 b15zdnd11an1n64x5 FILLER_6_72 ();
 b15zdnd11an1n64x5 FILLER_6_136 ();
 b15zdnd11an1n64x5 FILLER_6_200 ();
 b15zdnd11an1n64x5 FILLER_6_264 ();
 b15zdnd11an1n64x5 FILLER_6_328 ();
 b15zdnd11an1n64x5 FILLER_6_392 ();
 b15zdnd11an1n64x5 FILLER_6_456 ();
 b15zdnd11an1n64x5 FILLER_6_520 ();
 b15zdnd11an1n64x5 FILLER_6_584 ();
 b15zdnd11an1n64x5 FILLER_6_648 ();
 b15zdnd11an1n04x5 FILLER_6_712 ();
 b15zdnd00an1n02x5 FILLER_6_716 ();
 b15zdnd11an1n64x5 FILLER_6_726 ();
 b15zdnd11an1n64x5 FILLER_6_790 ();
 b15zdnd11an1n64x5 FILLER_6_854 ();
 b15zdnd11an1n64x5 FILLER_6_918 ();
 b15zdnd11an1n64x5 FILLER_6_982 ();
 b15zdnd11an1n64x5 FILLER_6_1046 ();
 b15zdnd11an1n64x5 FILLER_6_1110 ();
 b15zdnd11an1n64x5 FILLER_6_1174 ();
 b15zdnd11an1n64x5 FILLER_6_1238 ();
 b15zdnd11an1n64x5 FILLER_6_1302 ();
 b15zdnd11an1n64x5 FILLER_6_1366 ();
 b15zdnd11an1n64x5 FILLER_6_1430 ();
 b15zdnd11an1n64x5 FILLER_6_1494 ();
 b15zdnd11an1n64x5 FILLER_6_1558 ();
 b15zdnd11an1n64x5 FILLER_6_1622 ();
 b15zdnd11an1n64x5 FILLER_6_1686 ();
 b15zdnd11an1n64x5 FILLER_6_1750 ();
 b15zdnd11an1n64x5 FILLER_6_1814 ();
 b15zdnd11an1n64x5 FILLER_6_1878 ();
 b15zdnd11an1n64x5 FILLER_6_1942 ();
 b15zdnd11an1n64x5 FILLER_6_2006 ();
 b15zdnd11an1n64x5 FILLER_6_2070 ();
 b15zdnd11an1n16x5 FILLER_6_2134 ();
 b15zdnd11an1n04x5 FILLER_6_2150 ();
 b15zdnd11an1n64x5 FILLER_6_2162 ();
 b15zdnd11an1n32x5 FILLER_6_2226 ();
 b15zdnd11an1n16x5 FILLER_6_2258 ();
 b15zdnd00an1n02x5 FILLER_6_2274 ();
 b15zdnd11an1n64x5 FILLER_7_0 ();
 b15zdnd11an1n64x5 FILLER_7_64 ();
 b15zdnd11an1n64x5 FILLER_7_128 ();
 b15zdnd11an1n64x5 FILLER_7_192 ();
 b15zdnd11an1n64x5 FILLER_7_256 ();
 b15zdnd11an1n64x5 FILLER_7_320 ();
 b15zdnd11an1n64x5 FILLER_7_384 ();
 b15zdnd11an1n64x5 FILLER_7_448 ();
 b15zdnd11an1n64x5 FILLER_7_512 ();
 b15zdnd11an1n64x5 FILLER_7_576 ();
 b15zdnd11an1n64x5 FILLER_7_640 ();
 b15zdnd11an1n64x5 FILLER_7_704 ();
 b15zdnd11an1n64x5 FILLER_7_768 ();
 b15zdnd11an1n32x5 FILLER_7_832 ();
 b15zdnd11an1n16x5 FILLER_7_864 ();
 b15zdnd11an1n08x5 FILLER_7_880 ();
 b15zdnd11an1n04x5 FILLER_7_888 ();
 b15zdnd00an1n01x5 FILLER_7_892 ();
 b15zdnd11an1n16x5 FILLER_7_896 ();
 b15zdnd11an1n04x5 FILLER_7_912 ();
 b15zdnd00an1n02x5 FILLER_7_916 ();
 b15zdnd00an1n01x5 FILLER_7_918 ();
 b15zdnd11an1n64x5 FILLER_7_926 ();
 b15zdnd11an1n64x5 FILLER_7_990 ();
 b15zdnd11an1n64x5 FILLER_7_1054 ();
 b15zdnd11an1n32x5 FILLER_7_1118 ();
 b15zdnd11an1n08x5 FILLER_7_1150 ();
 b15zdnd11an1n04x5 FILLER_7_1158 ();
 b15zdnd11an1n16x5 FILLER_7_1165 ();
 b15zdnd11an1n08x5 FILLER_7_1181 ();
 b15zdnd11an1n04x5 FILLER_7_1189 ();
 b15zdnd00an1n01x5 FILLER_7_1193 ();
 b15zdnd11an1n32x5 FILLER_7_1202 ();
 b15zdnd11an1n16x5 FILLER_7_1234 ();
 b15zdnd00an1n02x5 FILLER_7_1250 ();
 b15zdnd00an1n01x5 FILLER_7_1252 ();
 b15zdnd11an1n16x5 FILLER_7_1256 ();
 b15zdnd11an1n08x5 FILLER_7_1272 ();
 b15zdnd00an1n02x5 FILLER_7_1280 ();
 b15zdnd11an1n04x5 FILLER_7_1285 ();
 b15zdnd11an1n64x5 FILLER_7_1292 ();
 b15zdnd11an1n64x5 FILLER_7_1356 ();
 b15zdnd11an1n64x5 FILLER_7_1420 ();
 b15zdnd11an1n64x5 FILLER_7_1484 ();
 b15zdnd11an1n64x5 FILLER_7_1548 ();
 b15zdnd11an1n64x5 FILLER_7_1612 ();
 b15zdnd11an1n64x5 FILLER_7_1676 ();
 b15zdnd11an1n64x5 FILLER_7_1740 ();
 b15zdnd11an1n64x5 FILLER_7_1804 ();
 b15zdnd11an1n32x5 FILLER_7_1868 ();
 b15zdnd11an1n16x5 FILLER_7_1900 ();
 b15zdnd11an1n08x5 FILLER_7_1916 ();
 b15zdnd11an1n04x5 FILLER_7_1924 ();
 b15zdnd11an1n64x5 FILLER_7_1931 ();
 b15zdnd11an1n64x5 FILLER_7_1995 ();
 b15zdnd11an1n64x5 FILLER_7_2059 ();
 b15zdnd11an1n64x5 FILLER_7_2123 ();
 b15zdnd11an1n08x5 FILLER_7_2187 ();
 b15zdnd00an1n02x5 FILLER_7_2195 ();
 b15zdnd00an1n01x5 FILLER_7_2197 ();
 b15zdnd11an1n04x5 FILLER_7_2201 ();
 b15zdnd11an1n64x5 FILLER_7_2208 ();
 b15zdnd11an1n08x5 FILLER_7_2272 ();
 b15zdnd11an1n04x5 FILLER_7_2280 ();
 b15zdnd11an1n64x5 FILLER_8_8 ();
 b15zdnd11an1n64x5 FILLER_8_72 ();
 b15zdnd11an1n64x5 FILLER_8_136 ();
 b15zdnd11an1n64x5 FILLER_8_200 ();
 b15zdnd11an1n64x5 FILLER_8_264 ();
 b15zdnd11an1n64x5 FILLER_8_328 ();
 b15zdnd11an1n64x5 FILLER_8_392 ();
 b15zdnd11an1n64x5 FILLER_8_456 ();
 b15zdnd11an1n64x5 FILLER_8_520 ();
 b15zdnd11an1n64x5 FILLER_8_584 ();
 b15zdnd11an1n64x5 FILLER_8_648 ();
 b15zdnd11an1n04x5 FILLER_8_712 ();
 b15zdnd00an1n02x5 FILLER_8_716 ();
 b15zdnd11an1n64x5 FILLER_8_726 ();
 b15zdnd11an1n32x5 FILLER_8_790 ();
 b15zdnd11an1n16x5 FILLER_8_822 ();
 b15zdnd11an1n08x5 FILLER_8_838 ();
 b15zdnd11an1n04x5 FILLER_8_846 ();
 b15zdnd00an1n02x5 FILLER_8_850 ();
 b15zdnd11an1n08x5 FILLER_8_858 ();
 b15zdnd11an1n04x5 FILLER_8_866 ();
 b15zdnd11an1n64x5 FILLER_8_922 ();
 b15zdnd11an1n64x5 FILLER_8_986 ();
 b15zdnd11an1n64x5 FILLER_8_1050 ();
 b15zdnd11an1n08x5 FILLER_8_1114 ();
 b15zdnd00an1n01x5 FILLER_8_1122 ();
 b15zdnd11an1n04x5 FILLER_8_1130 ();
 b15zdnd11an1n16x5 FILLER_8_1186 ();
 b15zdnd11an1n04x5 FILLER_8_1202 ();
 b15zdnd00an1n02x5 FILLER_8_1206 ();
 b15zdnd11an1n32x5 FILLER_8_1217 ();
 b15zdnd11an1n04x5 FILLER_8_1249 ();
 b15zdnd00an1n01x5 FILLER_8_1253 ();
 b15zdnd11an1n04x5 FILLER_8_1257 ();
 b15zdnd00an1n02x5 FILLER_8_1261 ();
 b15zdnd00an1n01x5 FILLER_8_1263 ();
 b15zdnd11an1n64x5 FILLER_8_1316 ();
 b15zdnd11an1n64x5 FILLER_8_1380 ();
 b15zdnd11an1n64x5 FILLER_8_1444 ();
 b15zdnd11an1n64x5 FILLER_8_1508 ();
 b15zdnd11an1n64x5 FILLER_8_1572 ();
 b15zdnd11an1n64x5 FILLER_8_1636 ();
 b15zdnd11an1n64x5 FILLER_8_1700 ();
 b15zdnd11an1n64x5 FILLER_8_1764 ();
 b15zdnd11an1n64x5 FILLER_8_1828 ();
 b15zdnd11an1n32x5 FILLER_8_1892 ();
 b15zdnd11an1n64x5 FILLER_8_1927 ();
 b15zdnd11an1n16x5 FILLER_8_1991 ();
 b15zdnd11an1n04x5 FILLER_8_2007 ();
 b15zdnd00an1n01x5 FILLER_8_2011 ();
 b15zdnd11an1n04x5 FILLER_8_2015 ();
 b15zdnd11an1n64x5 FILLER_8_2022 ();
 b15zdnd11an1n64x5 FILLER_8_2086 ();
 b15zdnd11an1n04x5 FILLER_8_2150 ();
 b15zdnd11an1n32x5 FILLER_8_2162 ();
 b15zdnd11an1n08x5 FILLER_8_2194 ();
 b15zdnd00an1n02x5 FILLER_8_2202 ();
 b15zdnd11an1n64x5 FILLER_8_2207 ();
 b15zdnd11an1n04x5 FILLER_8_2271 ();
 b15zdnd00an1n01x5 FILLER_8_2275 ();
 b15zdnd11an1n64x5 FILLER_9_0 ();
 b15zdnd11an1n64x5 FILLER_9_64 ();
 b15zdnd11an1n64x5 FILLER_9_128 ();
 b15zdnd11an1n64x5 FILLER_9_192 ();
 b15zdnd11an1n64x5 FILLER_9_256 ();
 b15zdnd11an1n64x5 FILLER_9_320 ();
 b15zdnd11an1n64x5 FILLER_9_384 ();
 b15zdnd11an1n64x5 FILLER_9_448 ();
 b15zdnd11an1n64x5 FILLER_9_512 ();
 b15zdnd11an1n64x5 FILLER_9_576 ();
 b15zdnd11an1n64x5 FILLER_9_640 ();
 b15zdnd11an1n64x5 FILLER_9_704 ();
 b15zdnd11an1n64x5 FILLER_9_768 ();
 b15zdnd11an1n32x5 FILLER_9_832 ();
 b15zdnd11an1n16x5 FILLER_9_864 ();
 b15zdnd11an1n08x5 FILLER_9_880 ();
 b15zdnd00an1n02x5 FILLER_9_888 ();
 b15zdnd11an1n04x5 FILLER_9_893 ();
 b15zdnd11an1n64x5 FILLER_9_900 ();
 b15zdnd11an1n64x5 FILLER_9_964 ();
 b15zdnd11an1n32x5 FILLER_9_1028 ();
 b15zdnd11an1n08x5 FILLER_9_1060 ();
 b15zdnd00an1n01x5 FILLER_9_1068 ();
 b15zdnd11an1n16x5 FILLER_9_1076 ();
 b15zdnd11an1n16x5 FILLER_9_1098 ();
 b15zdnd11an1n08x5 FILLER_9_1114 ();
 b15zdnd11an1n04x5 FILLER_9_1122 ();
 b15zdnd00an1n02x5 FILLER_9_1126 ();
 b15zdnd11an1n04x5 FILLER_9_1159 ();
 b15zdnd11an1n08x5 FILLER_9_1166 ();
 b15zdnd11an1n04x5 FILLER_9_1174 ();
 b15zdnd00an1n02x5 FILLER_9_1178 ();
 b15zdnd11an1n32x5 FILLER_9_1185 ();
 b15zdnd11an1n16x5 FILLER_9_1217 ();
 b15zdnd11an1n04x5 FILLER_9_1285 ();
 b15zdnd11an1n32x5 FILLER_9_1292 ();
 b15zdnd11an1n16x5 FILLER_9_1324 ();
 b15zdnd00an1n02x5 FILLER_9_1340 ();
 b15zdnd11an1n32x5 FILLER_9_1387 ();
 b15zdnd11an1n16x5 FILLER_9_1419 ();
 b15zdnd11an1n08x5 FILLER_9_1435 ();
 b15zdnd00an1n02x5 FILLER_9_1443 ();
 b15zdnd00an1n01x5 FILLER_9_1445 ();
 b15zdnd11an1n64x5 FILLER_9_1453 ();
 b15zdnd11an1n64x5 FILLER_9_1517 ();
 b15zdnd11an1n64x5 FILLER_9_1581 ();
 b15zdnd11an1n64x5 FILLER_9_1645 ();
 b15zdnd11an1n64x5 FILLER_9_1709 ();
 b15zdnd11an1n64x5 FILLER_9_1773 ();
 b15zdnd11an1n64x5 FILLER_9_1837 ();
 b15zdnd11an1n64x5 FILLER_9_1901 ();
 b15zdnd11an1n64x5 FILLER_9_1965 ();
 b15zdnd11an1n64x5 FILLER_9_2029 ();
 b15zdnd11an1n64x5 FILLER_9_2093 ();
 b15zdnd11an1n32x5 FILLER_9_2157 ();
 b15zdnd11an1n08x5 FILLER_9_2189 ();
 b15zdnd11an1n04x5 FILLER_9_2197 ();
 b15zdnd00an1n01x5 FILLER_9_2201 ();
 b15zdnd11an1n64x5 FILLER_9_2205 ();
 b15zdnd11an1n08x5 FILLER_9_2269 ();
 b15zdnd11an1n04x5 FILLER_9_2277 ();
 b15zdnd00an1n02x5 FILLER_9_2281 ();
 b15zdnd00an1n01x5 FILLER_9_2283 ();
 b15zdnd11an1n64x5 FILLER_10_8 ();
 b15zdnd11an1n64x5 FILLER_10_72 ();
 b15zdnd11an1n64x5 FILLER_10_136 ();
 b15zdnd11an1n64x5 FILLER_10_200 ();
 b15zdnd11an1n64x5 FILLER_10_264 ();
 b15zdnd11an1n64x5 FILLER_10_328 ();
 b15zdnd11an1n64x5 FILLER_10_392 ();
 b15zdnd11an1n64x5 FILLER_10_456 ();
 b15zdnd11an1n64x5 FILLER_10_520 ();
 b15zdnd11an1n64x5 FILLER_10_584 ();
 b15zdnd11an1n64x5 FILLER_10_648 ();
 b15zdnd11an1n04x5 FILLER_10_712 ();
 b15zdnd00an1n02x5 FILLER_10_716 ();
 b15zdnd11an1n64x5 FILLER_10_726 ();
 b15zdnd11an1n64x5 FILLER_10_790 ();
 b15zdnd11an1n64x5 FILLER_10_854 ();
 b15zdnd11an1n64x5 FILLER_10_918 ();
 b15zdnd11an1n64x5 FILLER_10_982 ();
 b15zdnd11an1n64x5 FILLER_10_1046 ();
 b15zdnd11an1n32x5 FILLER_10_1110 ();
 b15zdnd11an1n16x5 FILLER_10_1142 ();
 b15zdnd11an1n64x5 FILLER_10_1161 ();
 b15zdnd11an1n32x5 FILLER_10_1225 ();
 b15zdnd00an1n01x5 FILLER_10_1257 ();
 b15zdnd11an1n64x5 FILLER_10_1261 ();
 b15zdnd11an1n64x5 FILLER_10_1325 ();
 b15zdnd11an1n64x5 FILLER_10_1389 ();
 b15zdnd11an1n64x5 FILLER_10_1453 ();
 b15zdnd11an1n64x5 FILLER_10_1517 ();
 b15zdnd11an1n64x5 FILLER_10_1581 ();
 b15zdnd11an1n64x5 FILLER_10_1645 ();
 b15zdnd11an1n64x5 FILLER_10_1709 ();
 b15zdnd11an1n64x5 FILLER_10_1773 ();
 b15zdnd11an1n64x5 FILLER_10_1837 ();
 b15zdnd11an1n64x5 FILLER_10_1901 ();
 b15zdnd11an1n64x5 FILLER_10_1965 ();
 b15zdnd11an1n64x5 FILLER_10_2029 ();
 b15zdnd11an1n32x5 FILLER_10_2093 ();
 b15zdnd11an1n16x5 FILLER_10_2125 ();
 b15zdnd11an1n08x5 FILLER_10_2141 ();
 b15zdnd11an1n04x5 FILLER_10_2149 ();
 b15zdnd00an1n01x5 FILLER_10_2153 ();
 b15zdnd11an1n64x5 FILLER_10_2162 ();
 b15zdnd11an1n32x5 FILLER_10_2226 ();
 b15zdnd11an1n16x5 FILLER_10_2258 ();
 b15zdnd00an1n02x5 FILLER_10_2274 ();
 b15zdnd11an1n64x5 FILLER_11_0 ();
 b15zdnd11an1n64x5 FILLER_11_64 ();
 b15zdnd11an1n64x5 FILLER_11_128 ();
 b15zdnd11an1n64x5 FILLER_11_192 ();
 b15zdnd11an1n64x5 FILLER_11_256 ();
 b15zdnd11an1n64x5 FILLER_11_320 ();
 b15zdnd11an1n64x5 FILLER_11_384 ();
 b15zdnd11an1n64x5 FILLER_11_448 ();
 b15zdnd11an1n64x5 FILLER_11_512 ();
 b15zdnd11an1n64x5 FILLER_11_576 ();
 b15zdnd11an1n64x5 FILLER_11_640 ();
 b15zdnd11an1n64x5 FILLER_11_704 ();
 b15zdnd11an1n64x5 FILLER_11_768 ();
 b15zdnd11an1n64x5 FILLER_11_832 ();
 b15zdnd11an1n64x5 FILLER_11_896 ();
 b15zdnd11an1n64x5 FILLER_11_960 ();
 b15zdnd11an1n64x5 FILLER_11_1024 ();
 b15zdnd11an1n64x5 FILLER_11_1088 ();
 b15zdnd11an1n64x5 FILLER_11_1152 ();
 b15zdnd11an1n32x5 FILLER_11_1216 ();
 b15zdnd11an1n16x5 FILLER_11_1248 ();
 b15zdnd11an1n04x5 FILLER_11_1264 ();
 b15zdnd00an1n01x5 FILLER_11_1268 ();
 b15zdnd11an1n64x5 FILLER_11_1285 ();
 b15zdnd11an1n64x5 FILLER_11_1349 ();
 b15zdnd11an1n64x5 FILLER_11_1413 ();
 b15zdnd11an1n64x5 FILLER_11_1477 ();
 b15zdnd11an1n64x5 FILLER_11_1541 ();
 b15zdnd11an1n64x5 FILLER_11_1605 ();
 b15zdnd11an1n64x5 FILLER_11_1669 ();
 b15zdnd11an1n64x5 FILLER_11_1733 ();
 b15zdnd11an1n64x5 FILLER_11_1797 ();
 b15zdnd11an1n64x5 FILLER_11_1861 ();
 b15zdnd11an1n64x5 FILLER_11_1925 ();
 b15zdnd11an1n64x5 FILLER_11_1989 ();
 b15zdnd11an1n64x5 FILLER_11_2053 ();
 b15zdnd11an1n64x5 FILLER_11_2117 ();
 b15zdnd11an1n64x5 FILLER_11_2181 ();
 b15zdnd11an1n32x5 FILLER_11_2245 ();
 b15zdnd11an1n04x5 FILLER_11_2277 ();
 b15zdnd00an1n02x5 FILLER_11_2281 ();
 b15zdnd00an1n01x5 FILLER_11_2283 ();
 b15zdnd11an1n64x5 FILLER_12_8 ();
 b15zdnd11an1n64x5 FILLER_12_72 ();
 b15zdnd11an1n64x5 FILLER_12_136 ();
 b15zdnd11an1n64x5 FILLER_12_200 ();
 b15zdnd11an1n64x5 FILLER_12_264 ();
 b15zdnd11an1n64x5 FILLER_12_328 ();
 b15zdnd11an1n64x5 FILLER_12_392 ();
 b15zdnd11an1n64x5 FILLER_12_456 ();
 b15zdnd11an1n64x5 FILLER_12_520 ();
 b15zdnd11an1n64x5 FILLER_12_584 ();
 b15zdnd11an1n64x5 FILLER_12_648 ();
 b15zdnd11an1n04x5 FILLER_12_712 ();
 b15zdnd00an1n02x5 FILLER_12_716 ();
 b15zdnd11an1n64x5 FILLER_12_726 ();
 b15zdnd11an1n64x5 FILLER_12_790 ();
 b15zdnd11an1n64x5 FILLER_12_854 ();
 b15zdnd11an1n64x5 FILLER_12_918 ();
 b15zdnd11an1n64x5 FILLER_12_982 ();
 b15zdnd11an1n64x5 FILLER_12_1046 ();
 b15zdnd11an1n64x5 FILLER_12_1110 ();
 b15zdnd11an1n64x5 FILLER_12_1174 ();
 b15zdnd11an1n64x5 FILLER_12_1238 ();
 b15zdnd11an1n64x5 FILLER_12_1302 ();
 b15zdnd11an1n64x5 FILLER_12_1366 ();
 b15zdnd11an1n64x5 FILLER_12_1430 ();
 b15zdnd00an1n01x5 FILLER_12_1494 ();
 b15zdnd11an1n04x5 FILLER_12_1537 ();
 b15zdnd00an1n02x5 FILLER_12_1541 ();
 b15zdnd11an1n32x5 FILLER_12_1585 ();
 b15zdnd11an1n16x5 FILLER_12_1617 ();
 b15zdnd11an1n04x5 FILLER_12_1633 ();
 b15zdnd00an1n01x5 FILLER_12_1637 ();
 b15zdnd11an1n64x5 FILLER_12_1641 ();
 b15zdnd11an1n64x5 FILLER_12_1705 ();
 b15zdnd11an1n64x5 FILLER_12_1769 ();
 b15zdnd11an1n64x5 FILLER_12_1833 ();
 b15zdnd11an1n64x5 FILLER_12_1897 ();
 b15zdnd11an1n64x5 FILLER_12_1961 ();
 b15zdnd11an1n64x5 FILLER_12_2025 ();
 b15zdnd11an1n64x5 FILLER_12_2089 ();
 b15zdnd00an1n01x5 FILLER_12_2153 ();
 b15zdnd11an1n64x5 FILLER_12_2162 ();
 b15zdnd11an1n32x5 FILLER_12_2226 ();
 b15zdnd11an1n16x5 FILLER_12_2258 ();
 b15zdnd00an1n02x5 FILLER_12_2274 ();
 b15zdnd11an1n64x5 FILLER_13_0 ();
 b15zdnd11an1n64x5 FILLER_13_64 ();
 b15zdnd11an1n64x5 FILLER_13_128 ();
 b15zdnd11an1n64x5 FILLER_13_192 ();
 b15zdnd11an1n64x5 FILLER_13_256 ();
 b15zdnd11an1n64x5 FILLER_13_320 ();
 b15zdnd11an1n64x5 FILLER_13_384 ();
 b15zdnd11an1n64x5 FILLER_13_448 ();
 b15zdnd11an1n64x5 FILLER_13_512 ();
 b15zdnd11an1n64x5 FILLER_13_576 ();
 b15zdnd11an1n64x5 FILLER_13_640 ();
 b15zdnd11an1n64x5 FILLER_13_704 ();
 b15zdnd11an1n64x5 FILLER_13_768 ();
 b15zdnd11an1n64x5 FILLER_13_832 ();
 b15zdnd11an1n64x5 FILLER_13_896 ();
 b15zdnd11an1n08x5 FILLER_13_960 ();
 b15zdnd11an1n08x5 FILLER_13_1010 ();
 b15zdnd00an1n02x5 FILLER_13_1018 ();
 b15zdnd11an1n64x5 FILLER_13_1062 ();
 b15zdnd11an1n64x5 FILLER_13_1126 ();
 b15zdnd11an1n64x5 FILLER_13_1190 ();
 b15zdnd11an1n64x5 FILLER_13_1254 ();
 b15zdnd11an1n64x5 FILLER_13_1318 ();
 b15zdnd11an1n64x5 FILLER_13_1382 ();
 b15zdnd11an1n64x5 FILLER_13_1446 ();
 b15zdnd11an1n64x5 FILLER_13_1510 ();
 b15zdnd11an1n32x5 FILLER_13_1574 ();
 b15zdnd11an1n04x5 FILLER_13_1606 ();
 b15zdnd00an1n02x5 FILLER_13_1610 ();
 b15zdnd11an1n64x5 FILLER_13_1664 ();
 b15zdnd11an1n64x5 FILLER_13_1728 ();
 b15zdnd11an1n64x5 FILLER_13_1792 ();
 b15zdnd11an1n64x5 FILLER_13_1856 ();
 b15zdnd11an1n64x5 FILLER_13_1920 ();
 b15zdnd11an1n64x5 FILLER_13_1984 ();
 b15zdnd11an1n64x5 FILLER_13_2048 ();
 b15zdnd11an1n64x5 FILLER_13_2112 ();
 b15zdnd11an1n64x5 FILLER_13_2176 ();
 b15zdnd11an1n32x5 FILLER_13_2240 ();
 b15zdnd11an1n08x5 FILLER_13_2272 ();
 b15zdnd11an1n04x5 FILLER_13_2280 ();
 b15zdnd11an1n64x5 FILLER_14_8 ();
 b15zdnd11an1n64x5 FILLER_14_72 ();
 b15zdnd11an1n64x5 FILLER_14_136 ();
 b15zdnd11an1n64x5 FILLER_14_200 ();
 b15zdnd11an1n64x5 FILLER_14_264 ();
 b15zdnd11an1n64x5 FILLER_14_328 ();
 b15zdnd11an1n64x5 FILLER_14_392 ();
 b15zdnd11an1n64x5 FILLER_14_456 ();
 b15zdnd11an1n64x5 FILLER_14_520 ();
 b15zdnd11an1n64x5 FILLER_14_584 ();
 b15zdnd11an1n64x5 FILLER_14_648 ();
 b15zdnd11an1n04x5 FILLER_14_712 ();
 b15zdnd00an1n02x5 FILLER_14_716 ();
 b15zdnd11an1n64x5 FILLER_14_726 ();
 b15zdnd11an1n64x5 FILLER_14_790 ();
 b15zdnd11an1n64x5 FILLER_14_854 ();
 b15zdnd11an1n64x5 FILLER_14_918 ();
 b15zdnd11an1n64x5 FILLER_14_982 ();
 b15zdnd11an1n64x5 FILLER_14_1046 ();
 b15zdnd11an1n64x5 FILLER_14_1110 ();
 b15zdnd11an1n64x5 FILLER_14_1174 ();
 b15zdnd11an1n64x5 FILLER_14_1238 ();
 b15zdnd11an1n64x5 FILLER_14_1302 ();
 b15zdnd11an1n64x5 FILLER_14_1366 ();
 b15zdnd11an1n64x5 FILLER_14_1430 ();
 b15zdnd11an1n32x5 FILLER_14_1494 ();
 b15zdnd11an1n08x5 FILLER_14_1526 ();
 b15zdnd11an1n04x5 FILLER_14_1534 ();
 b15zdnd11an1n04x5 FILLER_14_1541 ();
 b15zdnd11an1n64x5 FILLER_14_1548 ();
 b15zdnd11an1n16x5 FILLER_14_1612 ();
 b15zdnd11an1n64x5 FILLER_14_1670 ();
 b15zdnd11an1n64x5 FILLER_14_1734 ();
 b15zdnd11an1n64x5 FILLER_14_1798 ();
 b15zdnd11an1n64x5 FILLER_14_1862 ();
 b15zdnd11an1n64x5 FILLER_14_1926 ();
 b15zdnd11an1n64x5 FILLER_14_1990 ();
 b15zdnd11an1n64x5 FILLER_14_2054 ();
 b15zdnd11an1n32x5 FILLER_14_2118 ();
 b15zdnd11an1n04x5 FILLER_14_2150 ();
 b15zdnd11an1n64x5 FILLER_14_2162 ();
 b15zdnd11an1n32x5 FILLER_14_2226 ();
 b15zdnd11an1n16x5 FILLER_14_2258 ();
 b15zdnd00an1n02x5 FILLER_14_2274 ();
 b15zdnd11an1n64x5 FILLER_15_0 ();
 b15zdnd11an1n64x5 FILLER_15_64 ();
 b15zdnd11an1n64x5 FILLER_15_128 ();
 b15zdnd11an1n64x5 FILLER_15_192 ();
 b15zdnd11an1n64x5 FILLER_15_256 ();
 b15zdnd11an1n64x5 FILLER_15_320 ();
 b15zdnd11an1n64x5 FILLER_15_384 ();
 b15zdnd11an1n64x5 FILLER_15_448 ();
 b15zdnd11an1n64x5 FILLER_15_512 ();
 b15zdnd11an1n64x5 FILLER_15_576 ();
 b15zdnd11an1n64x5 FILLER_15_640 ();
 b15zdnd11an1n64x5 FILLER_15_704 ();
 b15zdnd11an1n64x5 FILLER_15_768 ();
 b15zdnd11an1n64x5 FILLER_15_832 ();
 b15zdnd11an1n64x5 FILLER_15_896 ();
 b15zdnd11an1n64x5 FILLER_15_960 ();
 b15zdnd11an1n64x5 FILLER_15_1024 ();
 b15zdnd11an1n64x5 FILLER_15_1088 ();
 b15zdnd11an1n64x5 FILLER_15_1152 ();
 b15zdnd11an1n64x5 FILLER_15_1216 ();
 b15zdnd11an1n64x5 FILLER_15_1280 ();
 b15zdnd11an1n64x5 FILLER_15_1344 ();
 b15zdnd11an1n64x5 FILLER_15_1408 ();
 b15zdnd11an1n32x5 FILLER_15_1472 ();
 b15zdnd11an1n16x5 FILLER_15_1504 ();
 b15zdnd11an1n08x5 FILLER_15_1520 ();
 b15zdnd00an1n01x5 FILLER_15_1528 ();
 b15zdnd11an1n32x5 FILLER_15_1571 ();
 b15zdnd11an1n16x5 FILLER_15_1603 ();
 b15zdnd11an1n08x5 FILLER_15_1619 ();
 b15zdnd00an1n02x5 FILLER_15_1627 ();
 b15zdnd00an1n01x5 FILLER_15_1629 ();
 b15zdnd11an1n04x5 FILLER_15_1633 ();
 b15zdnd11an1n64x5 FILLER_15_1640 ();
 b15zdnd11an1n64x5 FILLER_15_1704 ();
 b15zdnd11an1n64x5 FILLER_15_1768 ();
 b15zdnd11an1n64x5 FILLER_15_1832 ();
 b15zdnd11an1n64x5 FILLER_15_1896 ();
 b15zdnd11an1n64x5 FILLER_15_1960 ();
 b15zdnd11an1n64x5 FILLER_15_2024 ();
 b15zdnd11an1n64x5 FILLER_15_2088 ();
 b15zdnd11an1n64x5 FILLER_15_2152 ();
 b15zdnd11an1n64x5 FILLER_15_2216 ();
 b15zdnd11an1n04x5 FILLER_15_2280 ();
 b15zdnd11an1n64x5 FILLER_16_8 ();
 b15zdnd11an1n64x5 FILLER_16_72 ();
 b15zdnd11an1n64x5 FILLER_16_136 ();
 b15zdnd11an1n64x5 FILLER_16_200 ();
 b15zdnd11an1n64x5 FILLER_16_264 ();
 b15zdnd11an1n64x5 FILLER_16_328 ();
 b15zdnd11an1n64x5 FILLER_16_392 ();
 b15zdnd11an1n64x5 FILLER_16_456 ();
 b15zdnd11an1n16x5 FILLER_16_520 ();
 b15zdnd11an1n08x5 FILLER_16_536 ();
 b15zdnd11an1n64x5 FILLER_16_547 ();
 b15zdnd11an1n64x5 FILLER_16_611 ();
 b15zdnd11an1n32x5 FILLER_16_675 ();
 b15zdnd11an1n08x5 FILLER_16_707 ();
 b15zdnd00an1n02x5 FILLER_16_715 ();
 b15zdnd00an1n01x5 FILLER_16_717 ();
 b15zdnd11an1n64x5 FILLER_16_726 ();
 b15zdnd11an1n16x5 FILLER_16_790 ();
 b15zdnd11an1n08x5 FILLER_16_806 ();
 b15zdnd11an1n04x5 FILLER_16_814 ();
 b15zdnd11an1n64x5 FILLER_16_821 ();
 b15zdnd11an1n16x5 FILLER_16_885 ();
 b15zdnd11an1n08x5 FILLER_16_901 ();
 b15zdnd11an1n04x5 FILLER_16_909 ();
 b15zdnd00an1n02x5 FILLER_16_913 ();
 b15zdnd11an1n64x5 FILLER_16_918 ();
 b15zdnd11an1n64x5 FILLER_16_982 ();
 b15zdnd11an1n64x5 FILLER_16_1046 ();
 b15zdnd11an1n64x5 FILLER_16_1110 ();
 b15zdnd11an1n64x5 FILLER_16_1174 ();
 b15zdnd11an1n64x5 FILLER_16_1238 ();
 b15zdnd11an1n64x5 FILLER_16_1302 ();
 b15zdnd11an1n64x5 FILLER_16_1366 ();
 b15zdnd11an1n32x5 FILLER_16_1430 ();
 b15zdnd11an1n16x5 FILLER_16_1462 ();
 b15zdnd11an1n08x5 FILLER_16_1478 ();
 b15zdnd11an1n04x5 FILLER_16_1486 ();
 b15zdnd00an1n02x5 FILLER_16_1490 ();
 b15zdnd11an1n16x5 FILLER_16_1495 ();
 b15zdnd00an1n02x5 FILLER_16_1511 ();
 b15zdnd11an1n64x5 FILLER_16_1565 ();
 b15zdnd11an1n64x5 FILLER_16_1629 ();
 b15zdnd11an1n64x5 FILLER_16_1693 ();
 b15zdnd11an1n64x5 FILLER_16_1757 ();
 b15zdnd11an1n64x5 FILLER_16_1821 ();
 b15zdnd11an1n64x5 FILLER_16_1885 ();
 b15zdnd11an1n64x5 FILLER_16_1949 ();
 b15zdnd11an1n64x5 FILLER_16_2013 ();
 b15zdnd11an1n64x5 FILLER_16_2077 ();
 b15zdnd11an1n08x5 FILLER_16_2141 ();
 b15zdnd11an1n04x5 FILLER_16_2149 ();
 b15zdnd00an1n01x5 FILLER_16_2153 ();
 b15zdnd11an1n64x5 FILLER_16_2162 ();
 b15zdnd11an1n32x5 FILLER_16_2226 ();
 b15zdnd11an1n16x5 FILLER_16_2258 ();
 b15zdnd00an1n02x5 FILLER_16_2274 ();
 b15zdnd11an1n64x5 FILLER_17_0 ();
 b15zdnd11an1n64x5 FILLER_17_64 ();
 b15zdnd11an1n64x5 FILLER_17_128 ();
 b15zdnd11an1n64x5 FILLER_17_192 ();
 b15zdnd11an1n64x5 FILLER_17_256 ();
 b15zdnd11an1n64x5 FILLER_17_320 ();
 b15zdnd11an1n64x5 FILLER_17_384 ();
 b15zdnd11an1n64x5 FILLER_17_448 ();
 b15zdnd11an1n04x5 FILLER_17_512 ();
 b15zdnd00an1n01x5 FILLER_17_516 ();
 b15zdnd11an1n64x5 FILLER_17_569 ();
 b15zdnd11an1n64x5 FILLER_17_633 ();
 b15zdnd11an1n64x5 FILLER_17_697 ();
 b15zdnd11an1n32x5 FILLER_17_761 ();
 b15zdnd11an1n08x5 FILLER_17_793 ();
 b15zdnd11an1n04x5 FILLER_17_801 ();
 b15zdnd00an1n02x5 FILLER_17_805 ();
 b15zdnd11an1n32x5 FILLER_17_849 ();
 b15zdnd11an1n04x5 FILLER_17_881 ();
 b15zdnd00an1n02x5 FILLER_17_885 ();
 b15zdnd00an1n01x5 FILLER_17_887 ();
 b15zdnd11an1n16x5 FILLER_17_940 ();
 b15zdnd11an1n08x5 FILLER_17_956 ();
 b15zdnd11an1n04x5 FILLER_17_964 ();
 b15zdnd00an1n01x5 FILLER_17_968 ();
 b15zdnd11an1n64x5 FILLER_17_972 ();
 b15zdnd11an1n64x5 FILLER_17_1036 ();
 b15zdnd11an1n64x5 FILLER_17_1100 ();
 b15zdnd11an1n64x5 FILLER_17_1164 ();
 b15zdnd11an1n64x5 FILLER_17_1228 ();
 b15zdnd11an1n64x5 FILLER_17_1292 ();
 b15zdnd11an1n64x5 FILLER_17_1356 ();
 b15zdnd11an1n64x5 FILLER_17_1420 ();
 b15zdnd11an1n08x5 FILLER_17_1484 ();
 b15zdnd11an1n04x5 FILLER_17_1495 ();
 b15zdnd11an1n32x5 FILLER_17_1502 ();
 b15zdnd11an1n04x5 FILLER_17_1534 ();
 b15zdnd11an1n64x5 FILLER_17_1541 ();
 b15zdnd11an1n64x5 FILLER_17_1605 ();
 b15zdnd11an1n64x5 FILLER_17_1669 ();
 b15zdnd11an1n64x5 FILLER_17_1733 ();
 b15zdnd11an1n64x5 FILLER_17_1797 ();
 b15zdnd11an1n64x5 FILLER_17_1861 ();
 b15zdnd11an1n64x5 FILLER_17_1925 ();
 b15zdnd11an1n64x5 FILLER_17_1989 ();
 b15zdnd11an1n64x5 FILLER_17_2053 ();
 b15zdnd11an1n64x5 FILLER_17_2117 ();
 b15zdnd11an1n64x5 FILLER_17_2181 ();
 b15zdnd11an1n32x5 FILLER_17_2245 ();
 b15zdnd11an1n04x5 FILLER_17_2277 ();
 b15zdnd00an1n02x5 FILLER_17_2281 ();
 b15zdnd00an1n01x5 FILLER_17_2283 ();
 b15zdnd11an1n64x5 FILLER_18_8 ();
 b15zdnd11an1n64x5 FILLER_18_72 ();
 b15zdnd11an1n64x5 FILLER_18_136 ();
 b15zdnd11an1n64x5 FILLER_18_200 ();
 b15zdnd11an1n64x5 FILLER_18_264 ();
 b15zdnd11an1n64x5 FILLER_18_328 ();
 b15zdnd11an1n64x5 FILLER_18_392 ();
 b15zdnd11an1n64x5 FILLER_18_456 ();
 b15zdnd11an1n16x5 FILLER_18_520 ();
 b15zdnd11an1n04x5 FILLER_18_539 ();
 b15zdnd11an1n64x5 FILLER_18_546 ();
 b15zdnd11an1n64x5 FILLER_18_610 ();
 b15zdnd11an1n32x5 FILLER_18_674 ();
 b15zdnd11an1n08x5 FILLER_18_706 ();
 b15zdnd11an1n04x5 FILLER_18_714 ();
 b15zdnd11an1n64x5 FILLER_18_726 ();
 b15zdnd00an1n01x5 FILLER_18_790 ();
 b15zdnd11an1n64x5 FILLER_18_843 ();
 b15zdnd11an1n04x5 FILLER_18_910 ();
 b15zdnd11an1n16x5 FILLER_18_917 ();
 b15zdnd11an1n08x5 FILLER_18_933 ();
 b15zdnd00an1n01x5 FILLER_18_941 ();
 b15zdnd11an1n64x5 FILLER_18_994 ();
 b15zdnd11an1n64x5 FILLER_18_1058 ();
 b15zdnd11an1n64x5 FILLER_18_1122 ();
 b15zdnd11an1n64x5 FILLER_18_1186 ();
 b15zdnd11an1n64x5 FILLER_18_1250 ();
 b15zdnd11an1n64x5 FILLER_18_1314 ();
 b15zdnd11an1n64x5 FILLER_18_1378 ();
 b15zdnd11an1n16x5 FILLER_18_1442 ();
 b15zdnd11an1n08x5 FILLER_18_1458 ();
 b15zdnd00an1n02x5 FILLER_18_1466 ();
 b15zdnd00an1n01x5 FILLER_18_1468 ();
 b15zdnd11an1n04x5 FILLER_18_1521 ();
 b15zdnd00an1n02x5 FILLER_18_1525 ();
 b15zdnd11an1n04x5 FILLER_18_1569 ();
 b15zdnd00an1n02x5 FILLER_18_1573 ();
 b15zdnd11an1n64x5 FILLER_18_1617 ();
 b15zdnd11an1n64x5 FILLER_18_1681 ();
 b15zdnd11an1n64x5 FILLER_18_1745 ();
 b15zdnd11an1n64x5 FILLER_18_1809 ();
 b15zdnd11an1n64x5 FILLER_18_1873 ();
 b15zdnd11an1n64x5 FILLER_18_1937 ();
 b15zdnd11an1n64x5 FILLER_18_2001 ();
 b15zdnd11an1n64x5 FILLER_18_2065 ();
 b15zdnd11an1n16x5 FILLER_18_2129 ();
 b15zdnd11an1n08x5 FILLER_18_2145 ();
 b15zdnd00an1n01x5 FILLER_18_2153 ();
 b15zdnd11an1n64x5 FILLER_18_2162 ();
 b15zdnd11an1n32x5 FILLER_18_2226 ();
 b15zdnd11an1n16x5 FILLER_18_2258 ();
 b15zdnd00an1n02x5 FILLER_18_2274 ();
 b15zdnd11an1n64x5 FILLER_19_0 ();
 b15zdnd11an1n64x5 FILLER_19_64 ();
 b15zdnd11an1n64x5 FILLER_19_128 ();
 b15zdnd11an1n64x5 FILLER_19_192 ();
 b15zdnd11an1n64x5 FILLER_19_256 ();
 b15zdnd11an1n64x5 FILLER_19_320 ();
 b15zdnd11an1n64x5 FILLER_19_384 ();
 b15zdnd11an1n64x5 FILLER_19_448 ();
 b15zdnd11an1n64x5 FILLER_19_512 ();
 b15zdnd11an1n64x5 FILLER_19_576 ();
 b15zdnd11an1n64x5 FILLER_19_640 ();
 b15zdnd11an1n64x5 FILLER_19_704 ();
 b15zdnd11an1n32x5 FILLER_19_768 ();
 b15zdnd11an1n08x5 FILLER_19_800 ();
 b15zdnd00an1n02x5 FILLER_19_808 ();
 b15zdnd11an1n04x5 FILLER_19_813 ();
 b15zdnd11an1n64x5 FILLER_19_820 ();
 b15zdnd11an1n16x5 FILLER_19_884 ();
 b15zdnd11an1n04x5 FILLER_19_900 ();
 b15zdnd11an1n08x5 FILLER_19_946 ();
 b15zdnd11an1n04x5 FILLER_19_954 ();
 b15zdnd00an1n02x5 FILLER_19_958 ();
 b15zdnd00an1n01x5 FILLER_19_960 ();
 b15zdnd11an1n04x5 FILLER_19_964 ();
 b15zdnd11an1n64x5 FILLER_19_971 ();
 b15zdnd11an1n64x5 FILLER_19_1035 ();
 b15zdnd11an1n64x5 FILLER_19_1099 ();
 b15zdnd11an1n64x5 FILLER_19_1163 ();
 b15zdnd11an1n64x5 FILLER_19_1227 ();
 b15zdnd11an1n64x5 FILLER_19_1291 ();
 b15zdnd11an1n64x5 FILLER_19_1355 ();
 b15zdnd11an1n64x5 FILLER_19_1419 ();
 b15zdnd11an1n64x5 FILLER_19_1483 ();
 b15zdnd11an1n64x5 FILLER_19_1547 ();
 b15zdnd11an1n64x5 FILLER_19_1611 ();
 b15zdnd11an1n64x5 FILLER_19_1675 ();
 b15zdnd11an1n64x5 FILLER_19_1739 ();
 b15zdnd11an1n64x5 FILLER_19_1803 ();
 b15zdnd11an1n64x5 FILLER_19_1867 ();
 b15zdnd11an1n64x5 FILLER_19_1931 ();
 b15zdnd11an1n64x5 FILLER_19_1995 ();
 b15zdnd11an1n64x5 FILLER_19_2059 ();
 b15zdnd11an1n64x5 FILLER_19_2123 ();
 b15zdnd11an1n64x5 FILLER_19_2187 ();
 b15zdnd11an1n32x5 FILLER_19_2251 ();
 b15zdnd00an1n01x5 FILLER_19_2283 ();
 b15zdnd11an1n64x5 FILLER_20_8 ();
 b15zdnd11an1n64x5 FILLER_20_72 ();
 b15zdnd11an1n64x5 FILLER_20_136 ();
 b15zdnd11an1n64x5 FILLER_20_200 ();
 b15zdnd11an1n64x5 FILLER_20_264 ();
 b15zdnd11an1n64x5 FILLER_20_328 ();
 b15zdnd11an1n64x5 FILLER_20_392 ();
 b15zdnd11an1n64x5 FILLER_20_456 ();
 b15zdnd11an1n64x5 FILLER_20_520 ();
 b15zdnd11an1n64x5 FILLER_20_584 ();
 b15zdnd11an1n64x5 FILLER_20_648 ();
 b15zdnd11an1n04x5 FILLER_20_712 ();
 b15zdnd00an1n02x5 FILLER_20_716 ();
 b15zdnd11an1n64x5 FILLER_20_726 ();
 b15zdnd11an1n08x5 FILLER_20_790 ();
 b15zdnd11an1n04x5 FILLER_20_798 ();
 b15zdnd00an1n02x5 FILLER_20_802 ();
 b15zdnd11an1n64x5 FILLER_20_846 ();
 b15zdnd11an1n64x5 FILLER_20_910 ();
 b15zdnd11an1n64x5 FILLER_20_974 ();
 b15zdnd11an1n64x5 FILLER_20_1038 ();
 b15zdnd11an1n64x5 FILLER_20_1102 ();
 b15zdnd11an1n64x5 FILLER_20_1166 ();
 b15zdnd11an1n64x5 FILLER_20_1230 ();
 b15zdnd11an1n32x5 FILLER_20_1294 ();
 b15zdnd11an1n16x5 FILLER_20_1326 ();
 b15zdnd11an1n08x5 FILLER_20_1342 ();
 b15zdnd00an1n02x5 FILLER_20_1350 ();
 b15zdnd11an1n04x5 FILLER_20_1394 ();
 b15zdnd11an1n64x5 FILLER_20_1401 ();
 b15zdnd11an1n64x5 FILLER_20_1465 ();
 b15zdnd11an1n64x5 FILLER_20_1529 ();
 b15zdnd11an1n64x5 FILLER_20_1593 ();
 b15zdnd11an1n64x5 FILLER_20_1657 ();
 b15zdnd11an1n64x5 FILLER_20_1721 ();
 b15zdnd11an1n64x5 FILLER_20_1785 ();
 b15zdnd11an1n64x5 FILLER_20_1849 ();
 b15zdnd11an1n64x5 FILLER_20_1913 ();
 b15zdnd11an1n64x5 FILLER_20_1977 ();
 b15zdnd11an1n64x5 FILLER_20_2041 ();
 b15zdnd11an1n32x5 FILLER_20_2105 ();
 b15zdnd11an1n16x5 FILLER_20_2137 ();
 b15zdnd00an1n01x5 FILLER_20_2153 ();
 b15zdnd11an1n64x5 FILLER_20_2162 ();
 b15zdnd11an1n32x5 FILLER_20_2226 ();
 b15zdnd11an1n16x5 FILLER_20_2258 ();
 b15zdnd00an1n02x5 FILLER_20_2274 ();
 b15zdnd11an1n64x5 FILLER_21_0 ();
 b15zdnd11an1n64x5 FILLER_21_64 ();
 b15zdnd11an1n64x5 FILLER_21_128 ();
 b15zdnd11an1n64x5 FILLER_21_192 ();
 b15zdnd11an1n32x5 FILLER_21_256 ();
 b15zdnd00an1n02x5 FILLER_21_288 ();
 b15zdnd00an1n01x5 FILLER_21_290 ();
 b15zdnd11an1n08x5 FILLER_21_294 ();
 b15zdnd11an1n04x5 FILLER_21_302 ();
 b15zdnd00an1n02x5 FILLER_21_306 ();
 b15zdnd00an1n01x5 FILLER_21_308 ();
 b15zdnd11an1n64x5 FILLER_21_312 ();
 b15zdnd11an1n64x5 FILLER_21_376 ();
 b15zdnd11an1n08x5 FILLER_21_440 ();
 b15zdnd11an1n04x5 FILLER_21_448 ();
 b15zdnd00an1n01x5 FILLER_21_452 ();
 b15zdnd11an1n64x5 FILLER_21_456 ();
 b15zdnd11an1n64x5 FILLER_21_520 ();
 b15zdnd11an1n64x5 FILLER_21_584 ();
 b15zdnd11an1n64x5 FILLER_21_648 ();
 b15zdnd11an1n16x5 FILLER_21_712 ();
 b15zdnd11an1n08x5 FILLER_21_728 ();
 b15zdnd00an1n01x5 FILLER_21_736 ();
 b15zdnd11an1n64x5 FILLER_21_789 ();
 b15zdnd11an1n64x5 FILLER_21_853 ();
 b15zdnd11an1n64x5 FILLER_21_917 ();
 b15zdnd11an1n64x5 FILLER_21_981 ();
 b15zdnd11an1n64x5 FILLER_21_1045 ();
 b15zdnd11an1n64x5 FILLER_21_1109 ();
 b15zdnd11an1n64x5 FILLER_21_1173 ();
 b15zdnd11an1n64x5 FILLER_21_1237 ();
 b15zdnd11an1n64x5 FILLER_21_1301 ();
 b15zdnd11an1n04x5 FILLER_21_1365 ();
 b15zdnd00an1n02x5 FILLER_21_1369 ();
 b15zdnd11an1n64x5 FILLER_21_1423 ();
 b15zdnd11an1n64x5 FILLER_21_1487 ();
 b15zdnd11an1n64x5 FILLER_21_1551 ();
 b15zdnd11an1n64x5 FILLER_21_1615 ();
 b15zdnd11an1n64x5 FILLER_21_1679 ();
 b15zdnd11an1n64x5 FILLER_21_1743 ();
 b15zdnd11an1n64x5 FILLER_21_1807 ();
 b15zdnd11an1n64x5 FILLER_21_1871 ();
 b15zdnd11an1n64x5 FILLER_21_1935 ();
 b15zdnd11an1n64x5 FILLER_21_1999 ();
 b15zdnd11an1n64x5 FILLER_21_2063 ();
 b15zdnd11an1n64x5 FILLER_21_2127 ();
 b15zdnd11an1n64x5 FILLER_21_2191 ();
 b15zdnd11an1n16x5 FILLER_21_2255 ();
 b15zdnd11an1n08x5 FILLER_21_2271 ();
 b15zdnd11an1n04x5 FILLER_21_2279 ();
 b15zdnd00an1n01x5 FILLER_21_2283 ();
 b15zdnd11an1n64x5 FILLER_22_8 ();
 b15zdnd11an1n64x5 FILLER_22_72 ();
 b15zdnd11an1n64x5 FILLER_22_136 ();
 b15zdnd11an1n64x5 FILLER_22_200 ();
 b15zdnd11an1n04x5 FILLER_22_264 ();
 b15zdnd00an1n02x5 FILLER_22_268 ();
 b15zdnd00an1n01x5 FILLER_22_270 ();
 b15zdnd11an1n64x5 FILLER_22_311 ();
 b15zdnd11an1n32x5 FILLER_22_375 ();
 b15zdnd11an1n16x5 FILLER_22_407 ();
 b15zdnd00an1n02x5 FILLER_22_423 ();
 b15zdnd00an1n01x5 FILLER_22_425 ();
 b15zdnd11an1n64x5 FILLER_22_478 ();
 b15zdnd11an1n64x5 FILLER_22_542 ();
 b15zdnd11an1n64x5 FILLER_22_606 ();
 b15zdnd11an1n32x5 FILLER_22_670 ();
 b15zdnd11an1n16x5 FILLER_22_702 ();
 b15zdnd11an1n16x5 FILLER_22_726 ();
 b15zdnd11an1n08x5 FILLER_22_742 ();
 b15zdnd11an1n04x5 FILLER_22_750 ();
 b15zdnd00an1n02x5 FILLER_22_754 ();
 b15zdnd00an1n01x5 FILLER_22_756 ();
 b15zdnd11an1n04x5 FILLER_22_760 ();
 b15zdnd11an1n64x5 FILLER_22_767 ();
 b15zdnd11an1n64x5 FILLER_22_831 ();
 b15zdnd11an1n64x5 FILLER_22_895 ();
 b15zdnd11an1n64x5 FILLER_22_959 ();
 b15zdnd11an1n04x5 FILLER_22_1023 ();
 b15zdnd00an1n02x5 FILLER_22_1027 ();
 b15zdnd00an1n01x5 FILLER_22_1029 ();
 b15zdnd11an1n64x5 FILLER_22_1033 ();
 b15zdnd11an1n64x5 FILLER_22_1097 ();
 b15zdnd11an1n64x5 FILLER_22_1161 ();
 b15zdnd11an1n64x5 FILLER_22_1225 ();
 b15zdnd11an1n32x5 FILLER_22_1289 ();
 b15zdnd11an1n08x5 FILLER_22_1321 ();
 b15zdnd11an1n16x5 FILLER_22_1371 ();
 b15zdnd11an1n08x5 FILLER_22_1387 ();
 b15zdnd00an1n01x5 FILLER_22_1395 ();
 b15zdnd11an1n04x5 FILLER_22_1399 ();
 b15zdnd11an1n64x5 FILLER_22_1406 ();
 b15zdnd11an1n64x5 FILLER_22_1470 ();
 b15zdnd11an1n64x5 FILLER_22_1534 ();
 b15zdnd11an1n64x5 FILLER_22_1598 ();
 b15zdnd11an1n64x5 FILLER_22_1662 ();
 b15zdnd11an1n64x5 FILLER_22_1726 ();
 b15zdnd11an1n32x5 FILLER_22_1790 ();
 b15zdnd11an1n16x5 FILLER_22_1822 ();
 b15zdnd11an1n08x5 FILLER_22_1838 ();
 b15zdnd00an1n02x5 FILLER_22_1846 ();
 b15zdnd11an1n04x5 FILLER_22_1851 ();
 b15zdnd11an1n64x5 FILLER_22_1858 ();
 b15zdnd11an1n64x5 FILLER_22_1922 ();
 b15zdnd11an1n64x5 FILLER_22_1986 ();
 b15zdnd11an1n64x5 FILLER_22_2050 ();
 b15zdnd11an1n32x5 FILLER_22_2114 ();
 b15zdnd11an1n08x5 FILLER_22_2146 ();
 b15zdnd11an1n64x5 FILLER_22_2162 ();
 b15zdnd11an1n32x5 FILLER_22_2226 ();
 b15zdnd11an1n16x5 FILLER_22_2258 ();
 b15zdnd00an1n02x5 FILLER_22_2274 ();
 b15zdnd11an1n64x5 FILLER_23_0 ();
 b15zdnd11an1n64x5 FILLER_23_64 ();
 b15zdnd11an1n64x5 FILLER_23_128 ();
 b15zdnd11an1n64x5 FILLER_23_192 ();
 b15zdnd11an1n64x5 FILLER_23_256 ();
 b15zdnd11an1n64x5 FILLER_23_320 ();
 b15zdnd11an1n32x5 FILLER_23_384 ();
 b15zdnd11an1n16x5 FILLER_23_416 ();
 b15zdnd11an1n08x5 FILLER_23_432 ();
 b15zdnd11an1n04x5 FILLER_23_440 ();
 b15zdnd11an1n04x5 FILLER_23_447 ();
 b15zdnd11an1n64x5 FILLER_23_454 ();
 b15zdnd11an1n64x5 FILLER_23_518 ();
 b15zdnd11an1n64x5 FILLER_23_582 ();
 b15zdnd11an1n64x5 FILLER_23_646 ();
 b15zdnd11an1n32x5 FILLER_23_710 ();
 b15zdnd11an1n08x5 FILLER_23_742 ();
 b15zdnd11an1n04x5 FILLER_23_750 ();
 b15zdnd00an1n02x5 FILLER_23_754 ();
 b15zdnd00an1n01x5 FILLER_23_756 ();
 b15zdnd11an1n64x5 FILLER_23_760 ();
 b15zdnd11an1n64x5 FILLER_23_824 ();
 b15zdnd11an1n64x5 FILLER_23_888 ();
 b15zdnd11an1n32x5 FILLER_23_952 ();
 b15zdnd00an1n02x5 FILLER_23_984 ();
 b15zdnd00an1n01x5 FILLER_23_986 ();
 b15zdnd11an1n08x5 FILLER_23_1029 ();
 b15zdnd11an1n64x5 FILLER_23_1040 ();
 b15zdnd11an1n64x5 FILLER_23_1104 ();
 b15zdnd11an1n64x5 FILLER_23_1168 ();
 b15zdnd11an1n32x5 FILLER_23_1232 ();
 b15zdnd11an1n16x5 FILLER_23_1264 ();
 b15zdnd00an1n02x5 FILLER_23_1280 ();
 b15zdnd11an1n04x5 FILLER_23_1285 ();
 b15zdnd11an1n04x5 FILLER_23_1292 ();
 b15zdnd00an1n02x5 FILLER_23_1296 ();
 b15zdnd00an1n01x5 FILLER_23_1298 ();
 b15zdnd11an1n64x5 FILLER_23_1341 ();
 b15zdnd11an1n64x5 FILLER_23_1405 ();
 b15zdnd11an1n32x5 FILLER_23_1469 ();
 b15zdnd11an1n08x5 FILLER_23_1501 ();
 b15zdnd11an1n04x5 FILLER_23_1551 ();
 b15zdnd11an1n64x5 FILLER_23_1607 ();
 b15zdnd11an1n16x5 FILLER_23_1671 ();
 b15zdnd11an1n08x5 FILLER_23_1729 ();
 b15zdnd00an1n01x5 FILLER_23_1737 ();
 b15zdnd11an1n04x5 FILLER_23_1741 ();
 b15zdnd11an1n64x5 FILLER_23_1748 ();
 b15zdnd11an1n16x5 FILLER_23_1812 ();
 b15zdnd00an1n02x5 FILLER_23_1828 ();
 b15zdnd11an1n64x5 FILLER_23_1882 ();
 b15zdnd11an1n64x5 FILLER_23_1946 ();
 b15zdnd11an1n64x5 FILLER_23_2010 ();
 b15zdnd11an1n64x5 FILLER_23_2074 ();
 b15zdnd11an1n64x5 FILLER_23_2138 ();
 b15zdnd11an1n64x5 FILLER_23_2202 ();
 b15zdnd11an1n16x5 FILLER_23_2266 ();
 b15zdnd00an1n02x5 FILLER_23_2282 ();
 b15zdnd11an1n64x5 FILLER_24_8 ();
 b15zdnd11an1n64x5 FILLER_24_72 ();
 b15zdnd11an1n64x5 FILLER_24_136 ();
 b15zdnd11an1n64x5 FILLER_24_200 ();
 b15zdnd11an1n64x5 FILLER_24_264 ();
 b15zdnd11an1n64x5 FILLER_24_328 ();
 b15zdnd11an1n64x5 FILLER_24_392 ();
 b15zdnd11an1n64x5 FILLER_24_456 ();
 b15zdnd11an1n64x5 FILLER_24_520 ();
 b15zdnd11an1n64x5 FILLER_24_584 ();
 b15zdnd11an1n64x5 FILLER_24_648 ();
 b15zdnd11an1n04x5 FILLER_24_712 ();
 b15zdnd00an1n02x5 FILLER_24_716 ();
 b15zdnd11an1n64x5 FILLER_24_726 ();
 b15zdnd11an1n64x5 FILLER_24_790 ();
 b15zdnd11an1n64x5 FILLER_24_854 ();
 b15zdnd11an1n64x5 FILLER_24_918 ();
 b15zdnd11an1n16x5 FILLER_24_982 ();
 b15zdnd11an1n04x5 FILLER_24_998 ();
 b15zdnd00an1n02x5 FILLER_24_1002 ();
 b15zdnd11an1n04x5 FILLER_24_1046 ();
 b15zdnd11an1n64x5 FILLER_24_1053 ();
 b15zdnd11an1n64x5 FILLER_24_1117 ();
 b15zdnd11an1n64x5 FILLER_24_1181 ();
 b15zdnd11an1n16x5 FILLER_24_1245 ();
 b15zdnd00an1n02x5 FILLER_24_1261 ();
 b15zdnd00an1n01x5 FILLER_24_1263 ();
 b15zdnd11an1n64x5 FILLER_24_1316 ();
 b15zdnd11an1n64x5 FILLER_24_1380 ();
 b15zdnd11an1n32x5 FILLER_24_1444 ();
 b15zdnd11an1n16x5 FILLER_24_1476 ();
 b15zdnd11an1n08x5 FILLER_24_1492 ();
 b15zdnd00an1n02x5 FILLER_24_1500 ();
 b15zdnd00an1n01x5 FILLER_24_1502 ();
 b15zdnd11an1n16x5 FILLER_24_1545 ();
 b15zdnd11an1n08x5 FILLER_24_1561 ();
 b15zdnd11an1n04x5 FILLER_24_1569 ();
 b15zdnd11an1n04x5 FILLER_24_1576 ();
 b15zdnd11an1n64x5 FILLER_24_1583 ();
 b15zdnd11an1n32x5 FILLER_24_1647 ();
 b15zdnd11an1n16x5 FILLER_24_1679 ();
 b15zdnd11an1n08x5 FILLER_24_1695 ();
 b15zdnd11an1n04x5 FILLER_24_1703 ();
 b15zdnd00an1n01x5 FILLER_24_1707 ();
 b15zdnd11an1n64x5 FILLER_24_1748 ();
 b15zdnd11an1n32x5 FILLER_24_1812 ();
 b15zdnd11an1n08x5 FILLER_24_1844 ();
 b15zdnd00an1n02x5 FILLER_24_1852 ();
 b15zdnd00an1n01x5 FILLER_24_1854 ();
 b15zdnd11an1n64x5 FILLER_24_1858 ();
 b15zdnd11an1n64x5 FILLER_24_1922 ();
 b15zdnd11an1n64x5 FILLER_24_1986 ();
 b15zdnd11an1n64x5 FILLER_24_2050 ();
 b15zdnd11an1n32x5 FILLER_24_2114 ();
 b15zdnd11an1n08x5 FILLER_24_2146 ();
 b15zdnd11an1n64x5 FILLER_24_2162 ();
 b15zdnd11an1n32x5 FILLER_24_2226 ();
 b15zdnd11an1n16x5 FILLER_24_2258 ();
 b15zdnd00an1n02x5 FILLER_24_2274 ();
 b15zdnd11an1n64x5 FILLER_25_0 ();
 b15zdnd11an1n64x5 FILLER_25_64 ();
 b15zdnd11an1n64x5 FILLER_25_128 ();
 b15zdnd11an1n64x5 FILLER_25_192 ();
 b15zdnd11an1n64x5 FILLER_25_256 ();
 b15zdnd11an1n64x5 FILLER_25_320 ();
 b15zdnd11an1n64x5 FILLER_25_384 ();
 b15zdnd11an1n64x5 FILLER_25_448 ();
 b15zdnd11an1n64x5 FILLER_25_512 ();
 b15zdnd11an1n64x5 FILLER_25_576 ();
 b15zdnd11an1n32x5 FILLER_25_640 ();
 b15zdnd11an1n16x5 FILLER_25_672 ();
 b15zdnd11an1n08x5 FILLER_25_688 ();
 b15zdnd11an1n04x5 FILLER_25_696 ();
 b15zdnd00an1n02x5 FILLER_25_700 ();
 b15zdnd00an1n01x5 FILLER_25_702 ();
 b15zdnd11an1n64x5 FILLER_25_745 ();
 b15zdnd11an1n64x5 FILLER_25_809 ();
 b15zdnd11an1n64x5 FILLER_25_873 ();
 b15zdnd11an1n16x5 FILLER_25_937 ();
 b15zdnd11an1n08x5 FILLER_25_995 ();
 b15zdnd11an1n04x5 FILLER_25_1003 ();
 b15zdnd00an1n01x5 FILLER_25_1007 ();
 b15zdnd11an1n64x5 FILLER_25_1060 ();
 b15zdnd11an1n64x5 FILLER_25_1124 ();
 b15zdnd11an1n64x5 FILLER_25_1188 ();
 b15zdnd11an1n32x5 FILLER_25_1252 ();
 b15zdnd00an1n02x5 FILLER_25_1284 ();
 b15zdnd11an1n04x5 FILLER_25_1328 ();
 b15zdnd00an1n02x5 FILLER_25_1332 ();
 b15zdnd00an1n01x5 FILLER_25_1334 ();
 b15zdnd11an1n64x5 FILLER_25_1377 ();
 b15zdnd11an1n32x5 FILLER_25_1441 ();
 b15zdnd11an1n16x5 FILLER_25_1473 ();
 b15zdnd00an1n02x5 FILLER_25_1489 ();
 b15zdnd11an1n32x5 FILLER_25_1533 ();
 b15zdnd11an1n16x5 FILLER_25_1565 ();
 b15zdnd11an1n64x5 FILLER_25_1584 ();
 b15zdnd11an1n64x5 FILLER_25_1648 ();
 b15zdnd11an1n64x5 FILLER_25_1712 ();
 b15zdnd11an1n64x5 FILLER_25_1776 ();
 b15zdnd11an1n64x5 FILLER_25_1840 ();
 b15zdnd11an1n64x5 FILLER_25_1904 ();
 b15zdnd11an1n64x5 FILLER_25_1968 ();
 b15zdnd11an1n64x5 FILLER_25_2032 ();
 b15zdnd11an1n64x5 FILLER_25_2096 ();
 b15zdnd11an1n64x5 FILLER_25_2160 ();
 b15zdnd11an1n32x5 FILLER_25_2224 ();
 b15zdnd11an1n16x5 FILLER_25_2256 ();
 b15zdnd11an1n08x5 FILLER_25_2272 ();
 b15zdnd11an1n04x5 FILLER_25_2280 ();
 b15zdnd11an1n64x5 FILLER_26_8 ();
 b15zdnd11an1n64x5 FILLER_26_72 ();
 b15zdnd11an1n64x5 FILLER_26_136 ();
 b15zdnd11an1n64x5 FILLER_26_200 ();
 b15zdnd11an1n64x5 FILLER_26_264 ();
 b15zdnd11an1n64x5 FILLER_26_328 ();
 b15zdnd11an1n32x5 FILLER_26_392 ();
 b15zdnd11an1n04x5 FILLER_26_424 ();
 b15zdnd11an1n32x5 FILLER_26_470 ();
 b15zdnd11an1n08x5 FILLER_26_502 ();
 b15zdnd11an1n04x5 FILLER_26_510 ();
 b15zdnd00an1n02x5 FILLER_26_514 ();
 b15zdnd00an1n01x5 FILLER_26_516 ();
 b15zdnd11an1n64x5 FILLER_26_559 ();
 b15zdnd11an1n64x5 FILLER_26_623 ();
 b15zdnd11an1n16x5 FILLER_26_687 ();
 b15zdnd11an1n08x5 FILLER_26_703 ();
 b15zdnd11an1n04x5 FILLER_26_711 ();
 b15zdnd00an1n02x5 FILLER_26_715 ();
 b15zdnd00an1n01x5 FILLER_26_717 ();
 b15zdnd11an1n64x5 FILLER_26_726 ();
 b15zdnd11an1n64x5 FILLER_26_790 ();
 b15zdnd11an1n64x5 FILLER_26_854 ();
 b15zdnd11an1n64x5 FILLER_26_918 ();
 b15zdnd11an1n64x5 FILLER_26_982 ();
 b15zdnd11an1n08x5 FILLER_26_1046 ();
 b15zdnd11an1n64x5 FILLER_26_1072 ();
 b15zdnd11an1n64x5 FILLER_26_1136 ();
 b15zdnd11an1n64x5 FILLER_26_1200 ();
 b15zdnd11an1n16x5 FILLER_26_1264 ();
 b15zdnd11an1n08x5 FILLER_26_1280 ();
 b15zdnd00an1n01x5 FILLER_26_1288 ();
 b15zdnd11an1n64x5 FILLER_26_1292 ();
 b15zdnd11an1n64x5 FILLER_26_1356 ();
 b15zdnd11an1n64x5 FILLER_26_1420 ();
 b15zdnd11an1n08x5 FILLER_26_1484 ();
 b15zdnd00an1n02x5 FILLER_26_1492 ();
 b15zdnd00an1n01x5 FILLER_26_1494 ();
 b15zdnd11an1n64x5 FILLER_26_1537 ();
 b15zdnd11an1n64x5 FILLER_26_1601 ();
 b15zdnd11an1n64x5 FILLER_26_1665 ();
 b15zdnd11an1n64x5 FILLER_26_1729 ();
 b15zdnd11an1n64x5 FILLER_26_1793 ();
 b15zdnd11an1n64x5 FILLER_26_1857 ();
 b15zdnd11an1n64x5 FILLER_26_1921 ();
 b15zdnd11an1n64x5 FILLER_26_1985 ();
 b15zdnd11an1n64x5 FILLER_26_2049 ();
 b15zdnd11an1n32x5 FILLER_26_2113 ();
 b15zdnd11an1n08x5 FILLER_26_2145 ();
 b15zdnd00an1n01x5 FILLER_26_2153 ();
 b15zdnd11an1n64x5 FILLER_26_2162 ();
 b15zdnd11an1n32x5 FILLER_26_2226 ();
 b15zdnd11an1n16x5 FILLER_26_2258 ();
 b15zdnd00an1n02x5 FILLER_26_2274 ();
 b15zdnd11an1n64x5 FILLER_27_0 ();
 b15zdnd11an1n64x5 FILLER_27_64 ();
 b15zdnd11an1n64x5 FILLER_27_128 ();
 b15zdnd11an1n64x5 FILLER_27_192 ();
 b15zdnd11an1n64x5 FILLER_27_256 ();
 b15zdnd11an1n64x5 FILLER_27_320 ();
 b15zdnd11an1n64x5 FILLER_27_384 ();
 b15zdnd11an1n64x5 FILLER_27_448 ();
 b15zdnd11an1n32x5 FILLER_27_512 ();
 b15zdnd11an1n16x5 FILLER_27_544 ();
 b15zdnd11an1n04x5 FILLER_27_560 ();
 b15zdnd00an1n01x5 FILLER_27_564 ();
 b15zdnd11an1n64x5 FILLER_27_568 ();
 b15zdnd11an1n64x5 FILLER_27_632 ();
 b15zdnd11an1n16x5 FILLER_27_696 ();
 b15zdnd11an1n08x5 FILLER_27_712 ();
 b15zdnd00an1n02x5 FILLER_27_720 ();
 b15zdnd00an1n01x5 FILLER_27_722 ();
 b15zdnd11an1n64x5 FILLER_27_765 ();
 b15zdnd11an1n64x5 FILLER_27_829 ();
 b15zdnd11an1n64x5 FILLER_27_893 ();
 b15zdnd11an1n64x5 FILLER_27_957 ();
 b15zdnd11an1n32x5 FILLER_27_1021 ();
 b15zdnd11an1n04x5 FILLER_27_1053 ();
 b15zdnd11an1n64x5 FILLER_27_1099 ();
 b15zdnd11an1n64x5 FILLER_27_1163 ();
 b15zdnd11an1n64x5 FILLER_27_1227 ();
 b15zdnd11an1n64x5 FILLER_27_1291 ();
 b15zdnd11an1n64x5 FILLER_27_1355 ();
 b15zdnd11an1n64x5 FILLER_27_1419 ();
 b15zdnd11an1n04x5 FILLER_27_1483 ();
 b15zdnd00an1n02x5 FILLER_27_1487 ();
 b15zdnd11an1n64x5 FILLER_27_1531 ();
 b15zdnd11an1n64x5 FILLER_27_1595 ();
 b15zdnd11an1n64x5 FILLER_27_1659 ();
 b15zdnd11an1n64x5 FILLER_27_1723 ();
 b15zdnd11an1n32x5 FILLER_27_1787 ();
 b15zdnd11an1n04x5 FILLER_27_1822 ();
 b15zdnd11an1n16x5 FILLER_27_1831 ();
 b15zdnd11an1n08x5 FILLER_27_1847 ();
 b15zdnd00an1n01x5 FILLER_27_1855 ();
 b15zdnd11an1n64x5 FILLER_27_1898 ();
 b15zdnd11an1n64x5 FILLER_27_1962 ();
 b15zdnd11an1n64x5 FILLER_27_2026 ();
 b15zdnd11an1n64x5 FILLER_27_2090 ();
 b15zdnd11an1n64x5 FILLER_27_2154 ();
 b15zdnd11an1n64x5 FILLER_27_2218 ();
 b15zdnd00an1n02x5 FILLER_27_2282 ();
 b15zdnd11an1n64x5 FILLER_28_8 ();
 b15zdnd11an1n64x5 FILLER_28_72 ();
 b15zdnd11an1n64x5 FILLER_28_136 ();
 b15zdnd11an1n64x5 FILLER_28_200 ();
 b15zdnd11an1n64x5 FILLER_28_264 ();
 b15zdnd11an1n64x5 FILLER_28_328 ();
 b15zdnd11an1n64x5 FILLER_28_392 ();
 b15zdnd11an1n64x5 FILLER_28_456 ();
 b15zdnd11an1n16x5 FILLER_28_520 ();
 b15zdnd00an1n02x5 FILLER_28_536 ();
 b15zdnd11an1n64x5 FILLER_28_590 ();
 b15zdnd11an1n16x5 FILLER_28_654 ();
 b15zdnd00an1n02x5 FILLER_28_670 ();
 b15zdnd00an1n01x5 FILLER_28_672 ();
 b15zdnd11an1n32x5 FILLER_28_676 ();
 b15zdnd11an1n08x5 FILLER_28_708 ();
 b15zdnd00an1n02x5 FILLER_28_716 ();
 b15zdnd11an1n64x5 FILLER_28_726 ();
 b15zdnd11an1n64x5 FILLER_28_790 ();
 b15zdnd11an1n64x5 FILLER_28_854 ();
 b15zdnd11an1n64x5 FILLER_28_918 ();
 b15zdnd11an1n08x5 FILLER_28_982 ();
 b15zdnd11an1n04x5 FILLER_28_990 ();
 b15zdnd00an1n02x5 FILLER_28_994 ();
 b15zdnd11an1n04x5 FILLER_28_999 ();
 b15zdnd00an1n01x5 FILLER_28_1003 ();
 b15zdnd11an1n64x5 FILLER_28_1010 ();
 b15zdnd11an1n64x5 FILLER_28_1074 ();
 b15zdnd11an1n16x5 FILLER_28_1138 ();
 b15zdnd11an1n04x5 FILLER_28_1154 ();
 b15zdnd11an1n04x5 FILLER_28_1198 ();
 b15zdnd11an1n32x5 FILLER_28_1205 ();
 b15zdnd11an1n04x5 FILLER_28_1237 ();
 b15zdnd11an1n64x5 FILLER_28_1252 ();
 b15zdnd11an1n64x5 FILLER_28_1316 ();
 b15zdnd11an1n64x5 FILLER_28_1380 ();
 b15zdnd11an1n64x5 FILLER_28_1444 ();
 b15zdnd00an1n02x5 FILLER_28_1508 ();
 b15zdnd11an1n64x5 FILLER_28_1515 ();
 b15zdnd11an1n64x5 FILLER_28_1579 ();
 b15zdnd11an1n32x5 FILLER_28_1643 ();
 b15zdnd11an1n16x5 FILLER_28_1675 ();
 b15zdnd00an1n02x5 FILLER_28_1691 ();
 b15zdnd11an1n64x5 FILLER_28_1701 ();
 b15zdnd11an1n32x5 FILLER_28_1765 ();
 b15zdnd11an1n16x5 FILLER_28_1797 ();
 b15zdnd00an1n02x5 FILLER_28_1813 ();
 b15zdnd00an1n01x5 FILLER_28_1815 ();
 b15zdnd11an1n08x5 FILLER_28_1819 ();
 b15zdnd00an1n02x5 FILLER_28_1827 ();
 b15zdnd11an1n04x5 FILLER_28_1832 ();
 b15zdnd11an1n64x5 FILLER_28_1878 ();
 b15zdnd11an1n64x5 FILLER_28_1942 ();
 b15zdnd11an1n64x5 FILLER_28_2006 ();
 b15zdnd11an1n64x5 FILLER_28_2070 ();
 b15zdnd11an1n16x5 FILLER_28_2134 ();
 b15zdnd11an1n04x5 FILLER_28_2150 ();
 b15zdnd11an1n64x5 FILLER_28_2162 ();
 b15zdnd11an1n32x5 FILLER_28_2226 ();
 b15zdnd11an1n16x5 FILLER_28_2258 ();
 b15zdnd00an1n02x5 FILLER_28_2274 ();
 b15zdnd11an1n64x5 FILLER_29_0 ();
 b15zdnd11an1n64x5 FILLER_29_64 ();
 b15zdnd11an1n64x5 FILLER_29_128 ();
 b15zdnd11an1n64x5 FILLER_29_192 ();
 b15zdnd11an1n64x5 FILLER_29_256 ();
 b15zdnd11an1n64x5 FILLER_29_320 ();
 b15zdnd11an1n32x5 FILLER_29_384 ();
 b15zdnd11an1n08x5 FILLER_29_416 ();
 b15zdnd00an1n02x5 FILLER_29_424 ();
 b15zdnd11an1n64x5 FILLER_29_441 ();
 b15zdnd11an1n08x5 FILLER_29_505 ();
 b15zdnd00an1n01x5 FILLER_29_513 ();
 b15zdnd11an1n08x5 FILLER_29_556 ();
 b15zdnd11an1n64x5 FILLER_29_567 ();
 b15zdnd11an1n32x5 FILLER_29_631 ();
 b15zdnd00an1n02x5 FILLER_29_663 ();
 b15zdnd11an1n04x5 FILLER_29_668 ();
 b15zdnd11an1n04x5 FILLER_29_675 ();
 b15zdnd00an1n01x5 FILLER_29_679 ();
 b15zdnd11an1n64x5 FILLER_29_722 ();
 b15zdnd11an1n64x5 FILLER_29_786 ();
 b15zdnd11an1n64x5 FILLER_29_850 ();
 b15zdnd11an1n64x5 FILLER_29_914 ();
 b15zdnd00an1n02x5 FILLER_29_978 ();
 b15zdnd11an1n04x5 FILLER_29_985 ();
 b15zdnd00an1n02x5 FILLER_29_989 ();
 b15zdnd00an1n01x5 FILLER_29_991 ();
 b15zdnd11an1n64x5 FILLER_29_1034 ();
 b15zdnd11an1n64x5 FILLER_29_1098 ();
 b15zdnd11an1n32x5 FILLER_29_1162 ();
 b15zdnd11an1n64x5 FILLER_29_1197 ();
 b15zdnd11an1n64x5 FILLER_29_1261 ();
 b15zdnd11an1n64x5 FILLER_29_1325 ();
 b15zdnd11an1n32x5 FILLER_29_1389 ();
 b15zdnd11an1n04x5 FILLER_29_1421 ();
 b15zdnd00an1n02x5 FILLER_29_1425 ();
 b15zdnd00an1n01x5 FILLER_29_1427 ();
 b15zdnd11an1n64x5 FILLER_29_1433 ();
 b15zdnd11an1n64x5 FILLER_29_1497 ();
 b15zdnd11an1n64x5 FILLER_29_1561 ();
 b15zdnd11an1n32x5 FILLER_29_1625 ();
 b15zdnd11an1n16x5 FILLER_29_1657 ();
 b15zdnd00an1n01x5 FILLER_29_1673 ();
 b15zdnd11an1n64x5 FILLER_29_1678 ();
 b15zdnd11an1n32x5 FILLER_29_1742 ();
 b15zdnd11an1n16x5 FILLER_29_1774 ();
 b15zdnd11an1n08x5 FILLER_29_1790 ();
 b15zdnd11an1n04x5 FILLER_29_1798 ();
 b15zdnd00an1n02x5 FILLER_29_1802 ();
 b15zdnd11an1n04x5 FILLER_29_1822 ();
 b15zdnd00an1n01x5 FILLER_29_1826 ();
 b15zdnd11an1n64x5 FILLER_29_1869 ();
 b15zdnd11an1n64x5 FILLER_29_1933 ();
 b15zdnd11an1n64x5 FILLER_29_1997 ();
 b15zdnd11an1n64x5 FILLER_29_2061 ();
 b15zdnd11an1n64x5 FILLER_29_2125 ();
 b15zdnd11an1n64x5 FILLER_29_2189 ();
 b15zdnd11an1n16x5 FILLER_29_2253 ();
 b15zdnd11an1n08x5 FILLER_29_2269 ();
 b15zdnd11an1n04x5 FILLER_29_2277 ();
 b15zdnd00an1n02x5 FILLER_29_2281 ();
 b15zdnd00an1n01x5 FILLER_29_2283 ();
 b15zdnd11an1n64x5 FILLER_30_8 ();
 b15zdnd11an1n64x5 FILLER_30_72 ();
 b15zdnd11an1n64x5 FILLER_30_136 ();
 b15zdnd11an1n64x5 FILLER_30_200 ();
 b15zdnd11an1n16x5 FILLER_30_264 ();
 b15zdnd11an1n08x5 FILLER_30_280 ();
 b15zdnd11an1n04x5 FILLER_30_288 ();
 b15zdnd00an1n01x5 FILLER_30_292 ();
 b15zdnd11an1n32x5 FILLER_30_296 ();
 b15zdnd11an1n16x5 FILLER_30_328 ();
 b15zdnd11an1n64x5 FILLER_30_386 ();
 b15zdnd11an1n64x5 FILLER_30_450 ();
 b15zdnd11an1n16x5 FILLER_30_514 ();
 b15zdnd00an1n02x5 FILLER_30_530 ();
 b15zdnd11an1n16x5 FILLER_30_536 ();
 b15zdnd11an1n04x5 FILLER_30_552 ();
 b15zdnd00an1n01x5 FILLER_30_556 ();
 b15zdnd11an1n64x5 FILLER_30_560 ();
 b15zdnd11an1n16x5 FILLER_30_624 ();
 b15zdnd11an1n04x5 FILLER_30_640 ();
 b15zdnd00an1n02x5 FILLER_30_644 ();
 b15zdnd11an1n04x5 FILLER_30_698 ();
 b15zdnd11an1n04x5 FILLER_30_711 ();
 b15zdnd00an1n02x5 FILLER_30_715 ();
 b15zdnd00an1n01x5 FILLER_30_717 ();
 b15zdnd11an1n64x5 FILLER_30_726 ();
 b15zdnd11an1n64x5 FILLER_30_790 ();
 b15zdnd11an1n64x5 FILLER_30_854 ();
 b15zdnd11an1n32x5 FILLER_30_918 ();
 b15zdnd11an1n08x5 FILLER_30_950 ();
 b15zdnd11an1n04x5 FILLER_30_958 ();
 b15zdnd00an1n01x5 FILLER_30_962 ();
 b15zdnd11an1n08x5 FILLER_30_967 ();
 b15zdnd00an1n02x5 FILLER_30_975 ();
 b15zdnd00an1n01x5 FILLER_30_977 ();
 b15zdnd11an1n64x5 FILLER_30_985 ();
 b15zdnd11an1n32x5 FILLER_30_1049 ();
 b15zdnd00an1n02x5 FILLER_30_1081 ();
 b15zdnd11an1n64x5 FILLER_30_1125 ();
 b15zdnd11an1n64x5 FILLER_30_1189 ();
 b15zdnd11an1n64x5 FILLER_30_1253 ();
 b15zdnd11an1n32x5 FILLER_30_1317 ();
 b15zdnd11an1n04x5 FILLER_30_1349 ();
 b15zdnd00an1n01x5 FILLER_30_1353 ();
 b15zdnd11an1n64x5 FILLER_30_1359 ();
 b15zdnd11an1n64x5 FILLER_30_1423 ();
 b15zdnd11an1n16x5 FILLER_30_1487 ();
 b15zdnd11an1n64x5 FILLER_30_1509 ();
 b15zdnd11an1n64x5 FILLER_30_1573 ();
 b15zdnd11an1n16x5 FILLER_30_1637 ();
 b15zdnd11an1n08x5 FILLER_30_1653 ();
 b15zdnd00an1n02x5 FILLER_30_1661 ();
 b15zdnd11an1n04x5 FILLER_30_1670 ();
 b15zdnd11an1n64x5 FILLER_30_1701 ();
 b15zdnd11an1n32x5 FILLER_30_1765 ();
 b15zdnd11an1n16x5 FILLER_30_1797 ();
 b15zdnd00an1n01x5 FILLER_30_1813 ();
 b15zdnd11an1n04x5 FILLER_30_1818 ();
 b15zdnd11an1n04x5 FILLER_30_1831 ();
 b15zdnd11an1n64x5 FILLER_30_1842 ();
 b15zdnd11an1n64x5 FILLER_30_1906 ();
 b15zdnd11an1n64x5 FILLER_30_1970 ();
 b15zdnd11an1n64x5 FILLER_30_2034 ();
 b15zdnd11an1n32x5 FILLER_30_2098 ();
 b15zdnd11an1n16x5 FILLER_30_2130 ();
 b15zdnd11an1n08x5 FILLER_30_2146 ();
 b15zdnd11an1n64x5 FILLER_30_2162 ();
 b15zdnd11an1n32x5 FILLER_30_2226 ();
 b15zdnd11an1n16x5 FILLER_30_2258 ();
 b15zdnd00an1n02x5 FILLER_30_2274 ();
 b15zdnd11an1n64x5 FILLER_31_0 ();
 b15zdnd11an1n64x5 FILLER_31_64 ();
 b15zdnd11an1n64x5 FILLER_31_128 ();
 b15zdnd11an1n64x5 FILLER_31_192 ();
 b15zdnd11an1n32x5 FILLER_31_256 ();
 b15zdnd00an1n02x5 FILLER_31_288 ();
 b15zdnd11an1n32x5 FILLER_31_299 ();
 b15zdnd11an1n04x5 FILLER_31_331 ();
 b15zdnd11an1n04x5 FILLER_31_338 ();
 b15zdnd11an1n08x5 FILLER_31_347 ();
 b15zdnd11an1n04x5 FILLER_31_359 ();
 b15zdnd11an1n64x5 FILLER_31_405 ();
 b15zdnd11an1n64x5 FILLER_31_469 ();
 b15zdnd11an1n64x5 FILLER_31_533 ();
 b15zdnd11an1n16x5 FILLER_31_597 ();
 b15zdnd11an1n08x5 FILLER_31_613 ();
 b15zdnd11an1n04x5 FILLER_31_621 ();
 b15zdnd11an1n04x5 FILLER_31_667 ();
 b15zdnd11an1n04x5 FILLER_31_677 ();
 b15zdnd11an1n64x5 FILLER_31_723 ();
 b15zdnd11an1n64x5 FILLER_31_787 ();
 b15zdnd11an1n64x5 FILLER_31_851 ();
 b15zdnd11an1n32x5 FILLER_31_915 ();
 b15zdnd11an1n04x5 FILLER_31_947 ();
 b15zdnd11an1n16x5 FILLER_31_955 ();
 b15zdnd00an1n02x5 FILLER_31_971 ();
 b15zdnd11an1n64x5 FILLER_31_987 ();
 b15zdnd11an1n64x5 FILLER_31_1051 ();
 b15zdnd11an1n64x5 FILLER_31_1115 ();
 b15zdnd11an1n64x5 FILLER_31_1179 ();
 b15zdnd11an1n64x5 FILLER_31_1243 ();
 b15zdnd11an1n64x5 FILLER_31_1307 ();
 b15zdnd11an1n64x5 FILLER_31_1371 ();
 b15zdnd11an1n64x5 FILLER_31_1435 ();
 b15zdnd11an1n64x5 FILLER_31_1499 ();
 b15zdnd11an1n64x5 FILLER_31_1563 ();
 b15zdnd11an1n32x5 FILLER_31_1627 ();
 b15zdnd11an1n16x5 FILLER_31_1659 ();
 b15zdnd11an1n04x5 FILLER_31_1675 ();
 b15zdnd00an1n02x5 FILLER_31_1679 ();
 b15zdnd00an1n01x5 FILLER_31_1681 ();
 b15zdnd11an1n32x5 FILLER_31_1734 ();
 b15zdnd11an1n08x5 FILLER_31_1766 ();
 b15zdnd00an1n02x5 FILLER_31_1774 ();
 b15zdnd11an1n32x5 FILLER_31_1782 ();
 b15zdnd11an1n04x5 FILLER_31_1818 ();
 b15zdnd11an1n64x5 FILLER_31_1827 ();
 b15zdnd11an1n64x5 FILLER_31_1891 ();
 b15zdnd11an1n64x5 FILLER_31_1955 ();
 b15zdnd11an1n64x5 FILLER_31_2019 ();
 b15zdnd11an1n64x5 FILLER_31_2083 ();
 b15zdnd11an1n64x5 FILLER_31_2147 ();
 b15zdnd11an1n64x5 FILLER_31_2211 ();
 b15zdnd11an1n08x5 FILLER_31_2275 ();
 b15zdnd00an1n01x5 FILLER_31_2283 ();
 b15zdnd11an1n64x5 FILLER_32_8 ();
 b15zdnd11an1n64x5 FILLER_32_72 ();
 b15zdnd11an1n64x5 FILLER_32_136 ();
 b15zdnd11an1n64x5 FILLER_32_200 ();
 b15zdnd11an1n32x5 FILLER_32_264 ();
 b15zdnd11an1n16x5 FILLER_32_296 ();
 b15zdnd11an1n04x5 FILLER_32_312 ();
 b15zdnd00an1n02x5 FILLER_32_316 ();
 b15zdnd11an1n08x5 FILLER_32_322 ();
 b15zdnd00an1n01x5 FILLER_32_330 ();
 b15zdnd11an1n04x5 FILLER_32_338 ();
 b15zdnd11an1n04x5 FILLER_32_394 ();
 b15zdnd11an1n64x5 FILLER_32_401 ();
 b15zdnd11an1n64x5 FILLER_32_465 ();
 b15zdnd11an1n64x5 FILLER_32_529 ();
 b15zdnd11an1n16x5 FILLER_32_593 ();
 b15zdnd11an1n08x5 FILLER_32_609 ();
 b15zdnd11an1n04x5 FILLER_32_659 ();
 b15zdnd00an1n01x5 FILLER_32_663 ();
 b15zdnd11an1n04x5 FILLER_32_706 ();
 b15zdnd11an1n04x5 FILLER_32_713 ();
 b15zdnd00an1n01x5 FILLER_32_717 ();
 b15zdnd11an1n64x5 FILLER_32_726 ();
 b15zdnd11an1n64x5 FILLER_32_790 ();
 b15zdnd11an1n64x5 FILLER_32_854 ();
 b15zdnd11an1n16x5 FILLER_32_918 ();
 b15zdnd11an1n08x5 FILLER_32_934 ();
 b15zdnd11an1n04x5 FILLER_32_942 ();
 b15zdnd00an1n01x5 FILLER_32_946 ();
 b15zdnd11an1n04x5 FILLER_32_963 ();
 b15zdnd00an1n02x5 FILLER_32_967 ();
 b15zdnd00an1n01x5 FILLER_32_969 ();
 b15zdnd11an1n64x5 FILLER_32_987 ();
 b15zdnd11an1n64x5 FILLER_32_1051 ();
 b15zdnd11an1n64x5 FILLER_32_1115 ();
 b15zdnd11an1n64x5 FILLER_32_1179 ();
 b15zdnd11an1n64x5 FILLER_32_1243 ();
 b15zdnd11an1n64x5 FILLER_32_1307 ();
 b15zdnd11an1n64x5 FILLER_32_1371 ();
 b15zdnd11an1n64x5 FILLER_32_1435 ();
 b15zdnd00an1n01x5 FILLER_32_1499 ();
 b15zdnd11an1n32x5 FILLER_32_1506 ();
 b15zdnd11an1n08x5 FILLER_32_1538 ();
 b15zdnd11an1n04x5 FILLER_32_1546 ();
 b15zdnd00an1n02x5 FILLER_32_1550 ();
 b15zdnd00an1n01x5 FILLER_32_1552 ();
 b15zdnd11an1n64x5 FILLER_32_1558 ();
 b15zdnd11an1n64x5 FILLER_32_1622 ();
 b15zdnd11an1n08x5 FILLER_32_1686 ();
 b15zdnd11an1n04x5 FILLER_32_1694 ();
 b15zdnd00an1n02x5 FILLER_32_1698 ();
 b15zdnd11an1n04x5 FILLER_32_1703 ();
 b15zdnd11an1n16x5 FILLER_32_1710 ();
 b15zdnd11an1n04x5 FILLER_32_1726 ();
 b15zdnd00an1n02x5 FILLER_32_1730 ();
 b15zdnd00an1n01x5 FILLER_32_1732 ();
 b15zdnd11an1n32x5 FILLER_32_1775 ();
 b15zdnd11an1n08x5 FILLER_32_1807 ();
 b15zdnd00an1n02x5 FILLER_32_1815 ();
 b15zdnd11an1n04x5 FILLER_32_1826 ();
 b15zdnd11an1n64x5 FILLER_32_1834 ();
 b15zdnd11an1n64x5 FILLER_32_1898 ();
 b15zdnd11an1n64x5 FILLER_32_1962 ();
 b15zdnd11an1n64x5 FILLER_32_2026 ();
 b15zdnd11an1n64x5 FILLER_32_2090 ();
 b15zdnd11an1n64x5 FILLER_32_2162 ();
 b15zdnd11an1n32x5 FILLER_32_2226 ();
 b15zdnd11an1n16x5 FILLER_32_2258 ();
 b15zdnd00an1n02x5 FILLER_32_2274 ();
 b15zdnd11an1n64x5 FILLER_33_0 ();
 b15zdnd11an1n64x5 FILLER_33_64 ();
 b15zdnd11an1n64x5 FILLER_33_128 ();
 b15zdnd11an1n64x5 FILLER_33_192 ();
 b15zdnd11an1n64x5 FILLER_33_256 ();
 b15zdnd11an1n32x5 FILLER_33_320 ();
 b15zdnd00an1n02x5 FILLER_33_352 ();
 b15zdnd11an1n64x5 FILLER_33_396 ();
 b15zdnd11an1n64x5 FILLER_33_460 ();
 b15zdnd11an1n64x5 FILLER_33_524 ();
 b15zdnd11an1n64x5 FILLER_33_588 ();
 b15zdnd00an1n02x5 FILLER_33_652 ();
 b15zdnd00an1n01x5 FILLER_33_654 ();
 b15zdnd11an1n04x5 FILLER_33_665 ();
 b15zdnd11an1n08x5 FILLER_33_679 ();
 b15zdnd11an1n64x5 FILLER_33_729 ();
 b15zdnd11an1n64x5 FILLER_33_793 ();
 b15zdnd11an1n64x5 FILLER_33_857 ();
 b15zdnd11an1n32x5 FILLER_33_921 ();
 b15zdnd11an1n04x5 FILLER_33_953 ();
 b15zdnd00an1n02x5 FILLER_33_957 ();
 b15zdnd00an1n01x5 FILLER_33_959 ();
 b15zdnd11an1n08x5 FILLER_33_963 ();
 b15zdnd00an1n02x5 FILLER_33_971 ();
 b15zdnd11an1n04x5 FILLER_33_977 ();
 b15zdnd00an1n02x5 FILLER_33_981 ();
 b15zdnd00an1n01x5 FILLER_33_983 ();
 b15zdnd11an1n64x5 FILLER_33_987 ();
 b15zdnd11an1n32x5 FILLER_33_1051 ();
 b15zdnd11an1n08x5 FILLER_33_1083 ();
 b15zdnd11an1n04x5 FILLER_33_1091 ();
 b15zdnd00an1n02x5 FILLER_33_1095 ();
 b15zdnd11an1n64x5 FILLER_33_1107 ();
 b15zdnd11an1n08x5 FILLER_33_1171 ();
 b15zdnd00an1n02x5 FILLER_33_1179 ();
 b15zdnd00an1n01x5 FILLER_33_1181 ();
 b15zdnd11an1n64x5 FILLER_33_1197 ();
 b15zdnd11an1n64x5 FILLER_33_1261 ();
 b15zdnd11an1n64x5 FILLER_33_1325 ();
 b15zdnd11an1n64x5 FILLER_33_1389 ();
 b15zdnd11an1n32x5 FILLER_33_1453 ();
 b15zdnd11an1n08x5 FILLER_33_1485 ();
 b15zdnd11an1n04x5 FILLER_33_1493 ();
 b15zdnd00an1n02x5 FILLER_33_1497 ();
 b15zdnd11an1n64x5 FILLER_33_1512 ();
 b15zdnd11an1n64x5 FILLER_33_1576 ();
 b15zdnd11an1n16x5 FILLER_33_1640 ();
 b15zdnd11an1n08x5 FILLER_33_1656 ();
 b15zdnd00an1n02x5 FILLER_33_1664 ();
 b15zdnd11an1n04x5 FILLER_33_1669 ();
 b15zdnd00an1n01x5 FILLER_33_1673 ();
 b15zdnd11an1n16x5 FILLER_33_1677 ();
 b15zdnd11an1n08x5 FILLER_33_1693 ();
 b15zdnd11an1n04x5 FILLER_33_1701 ();
 b15zdnd11an1n16x5 FILLER_33_1708 ();
 b15zdnd11an1n08x5 FILLER_33_1724 ();
 b15zdnd11an1n64x5 FILLER_33_1750 ();
 b15zdnd11an1n64x5 FILLER_33_1814 ();
 b15zdnd11an1n64x5 FILLER_33_1878 ();
 b15zdnd11an1n64x5 FILLER_33_1942 ();
 b15zdnd11an1n64x5 FILLER_33_2006 ();
 b15zdnd11an1n64x5 FILLER_33_2070 ();
 b15zdnd11an1n64x5 FILLER_33_2134 ();
 b15zdnd11an1n64x5 FILLER_33_2198 ();
 b15zdnd11an1n16x5 FILLER_33_2262 ();
 b15zdnd11an1n04x5 FILLER_33_2278 ();
 b15zdnd00an1n02x5 FILLER_33_2282 ();
 b15zdnd11an1n64x5 FILLER_34_8 ();
 b15zdnd11an1n64x5 FILLER_34_72 ();
 b15zdnd11an1n64x5 FILLER_34_136 ();
 b15zdnd11an1n64x5 FILLER_34_200 ();
 b15zdnd11an1n64x5 FILLER_34_264 ();
 b15zdnd11an1n04x5 FILLER_34_328 ();
 b15zdnd11an1n04x5 FILLER_34_374 ();
 b15zdnd00an1n02x5 FILLER_34_378 ();
 b15zdnd00an1n01x5 FILLER_34_380 ();
 b15zdnd11an1n64x5 FILLER_34_384 ();
 b15zdnd11an1n64x5 FILLER_34_448 ();
 b15zdnd11an1n64x5 FILLER_34_512 ();
 b15zdnd11an1n64x5 FILLER_34_576 ();
 b15zdnd11an1n16x5 FILLER_34_640 ();
 b15zdnd00an1n02x5 FILLER_34_656 ();
 b15zdnd00an1n01x5 FILLER_34_658 ();
 b15zdnd11an1n04x5 FILLER_34_669 ();
 b15zdnd11an1n04x5 FILLER_34_680 ();
 b15zdnd11an1n04x5 FILLER_34_688 ();
 b15zdnd11an1n16x5 FILLER_34_695 ();
 b15zdnd11an1n04x5 FILLER_34_711 ();
 b15zdnd00an1n02x5 FILLER_34_715 ();
 b15zdnd00an1n01x5 FILLER_34_717 ();
 b15zdnd11an1n64x5 FILLER_34_726 ();
 b15zdnd11an1n64x5 FILLER_34_790 ();
 b15zdnd11an1n64x5 FILLER_34_854 ();
 b15zdnd11an1n32x5 FILLER_34_918 ();
 b15zdnd11an1n08x5 FILLER_34_950 ();
 b15zdnd11an1n04x5 FILLER_34_958 ();
 b15zdnd00an1n02x5 FILLER_34_962 ();
 b15zdnd11an1n64x5 FILLER_34_974 ();
 b15zdnd11an1n32x5 FILLER_34_1038 ();
 b15zdnd11an1n08x5 FILLER_34_1070 ();
 b15zdnd00an1n02x5 FILLER_34_1078 ();
 b15zdnd00an1n01x5 FILLER_34_1080 ();
 b15zdnd11an1n64x5 FILLER_34_1088 ();
 b15zdnd11an1n64x5 FILLER_34_1152 ();
 b15zdnd11an1n64x5 FILLER_34_1216 ();
 b15zdnd11an1n64x5 FILLER_34_1280 ();
 b15zdnd11an1n64x5 FILLER_34_1344 ();
 b15zdnd11an1n64x5 FILLER_34_1408 ();
 b15zdnd11an1n16x5 FILLER_34_1472 ();
 b15zdnd11an1n08x5 FILLER_34_1488 ();
 b15zdnd00an1n02x5 FILLER_34_1496 ();
 b15zdnd11an1n04x5 FILLER_34_1507 ();
 b15zdnd11an1n04x5 FILLER_34_1515 ();
 b15zdnd00an1n01x5 FILLER_34_1519 ();
 b15zdnd11an1n64x5 FILLER_34_1529 ();
 b15zdnd11an1n32x5 FILLER_34_1593 ();
 b15zdnd11an1n08x5 FILLER_34_1625 ();
 b15zdnd00an1n02x5 FILLER_34_1633 ();
 b15zdnd11an1n64x5 FILLER_34_1675 ();
 b15zdnd11an1n64x5 FILLER_34_1739 ();
 b15zdnd11an1n64x5 FILLER_34_1803 ();
 b15zdnd11an1n64x5 FILLER_34_1867 ();
 b15zdnd11an1n64x5 FILLER_34_1931 ();
 b15zdnd11an1n64x5 FILLER_34_1995 ();
 b15zdnd11an1n64x5 FILLER_34_2059 ();
 b15zdnd11an1n16x5 FILLER_34_2123 ();
 b15zdnd11an1n08x5 FILLER_34_2139 ();
 b15zdnd11an1n04x5 FILLER_34_2147 ();
 b15zdnd00an1n02x5 FILLER_34_2151 ();
 b15zdnd00an1n01x5 FILLER_34_2153 ();
 b15zdnd11an1n64x5 FILLER_34_2162 ();
 b15zdnd11an1n32x5 FILLER_34_2226 ();
 b15zdnd11an1n16x5 FILLER_34_2258 ();
 b15zdnd00an1n02x5 FILLER_34_2274 ();
 b15zdnd11an1n64x5 FILLER_35_0 ();
 b15zdnd11an1n64x5 FILLER_35_64 ();
 b15zdnd11an1n64x5 FILLER_35_128 ();
 b15zdnd11an1n64x5 FILLER_35_192 ();
 b15zdnd11an1n32x5 FILLER_35_256 ();
 b15zdnd11an1n04x5 FILLER_35_288 ();
 b15zdnd00an1n02x5 FILLER_35_292 ();
 b15zdnd00an1n01x5 FILLER_35_294 ();
 b15zdnd11an1n16x5 FILLER_35_301 ();
 b15zdnd11an1n04x5 FILLER_35_317 ();
 b15zdnd11an1n08x5 FILLER_35_363 ();
 b15zdnd11an1n64x5 FILLER_35_374 ();
 b15zdnd11an1n64x5 FILLER_35_438 ();
 b15zdnd11an1n64x5 FILLER_35_502 ();
 b15zdnd11an1n64x5 FILLER_35_566 ();
 b15zdnd11an1n16x5 FILLER_35_630 ();
 b15zdnd11an1n04x5 FILLER_35_646 ();
 b15zdnd00an1n02x5 FILLER_35_650 ();
 b15zdnd00an1n01x5 FILLER_35_652 ();
 b15zdnd11an1n04x5 FILLER_35_663 ();
 b15zdnd11an1n64x5 FILLER_35_672 ();
 b15zdnd11an1n64x5 FILLER_35_736 ();
 b15zdnd11an1n64x5 FILLER_35_800 ();
 b15zdnd11an1n64x5 FILLER_35_864 ();
 b15zdnd11an1n64x5 FILLER_35_928 ();
 b15zdnd11an1n64x5 FILLER_35_992 ();
 b15zdnd11an1n64x5 FILLER_35_1056 ();
 b15zdnd11an1n64x5 FILLER_35_1120 ();
 b15zdnd11an1n64x5 FILLER_35_1184 ();
 b15zdnd11an1n64x5 FILLER_35_1248 ();
 b15zdnd11an1n64x5 FILLER_35_1312 ();
 b15zdnd11an1n32x5 FILLER_35_1376 ();
 b15zdnd11an1n08x5 FILLER_35_1408 ();
 b15zdnd11an1n04x5 FILLER_35_1416 ();
 b15zdnd00an1n02x5 FILLER_35_1420 ();
 b15zdnd00an1n01x5 FILLER_35_1422 ();
 b15zdnd11an1n64x5 FILLER_35_1432 ();
 b15zdnd11an1n04x5 FILLER_35_1496 ();
 b15zdnd00an1n01x5 FILLER_35_1500 ();
 b15zdnd11an1n64x5 FILLER_35_1515 ();
 b15zdnd11an1n64x5 FILLER_35_1579 ();
 b15zdnd11an1n64x5 FILLER_35_1643 ();
 b15zdnd11an1n64x5 FILLER_35_1707 ();
 b15zdnd11an1n64x5 FILLER_35_1771 ();
 b15zdnd11an1n64x5 FILLER_35_1835 ();
 b15zdnd11an1n64x5 FILLER_35_1899 ();
 b15zdnd11an1n64x5 FILLER_35_1963 ();
 b15zdnd11an1n64x5 FILLER_35_2027 ();
 b15zdnd11an1n64x5 FILLER_35_2091 ();
 b15zdnd11an1n64x5 FILLER_35_2155 ();
 b15zdnd11an1n64x5 FILLER_35_2219 ();
 b15zdnd00an1n01x5 FILLER_35_2283 ();
 b15zdnd11an1n64x5 FILLER_36_8 ();
 b15zdnd11an1n64x5 FILLER_36_72 ();
 b15zdnd11an1n64x5 FILLER_36_136 ();
 b15zdnd11an1n64x5 FILLER_36_200 ();
 b15zdnd11an1n16x5 FILLER_36_264 ();
 b15zdnd11an1n08x5 FILLER_36_280 ();
 b15zdnd00an1n02x5 FILLER_36_288 ();
 b15zdnd00an1n01x5 FILLER_36_290 ();
 b15zdnd11an1n64x5 FILLER_36_297 ();
 b15zdnd11an1n64x5 FILLER_36_361 ();
 b15zdnd11an1n64x5 FILLER_36_425 ();
 b15zdnd11an1n32x5 FILLER_36_489 ();
 b15zdnd11an1n16x5 FILLER_36_521 ();
 b15zdnd00an1n01x5 FILLER_36_537 ();
 b15zdnd11an1n64x5 FILLER_36_580 ();
 b15zdnd11an1n16x5 FILLER_36_644 ();
 b15zdnd11an1n08x5 FILLER_36_660 ();
 b15zdnd00an1n02x5 FILLER_36_668 ();
 b15zdnd11an1n32x5 FILLER_36_676 ();
 b15zdnd11an1n08x5 FILLER_36_708 ();
 b15zdnd00an1n02x5 FILLER_36_716 ();
 b15zdnd11an1n64x5 FILLER_36_726 ();
 b15zdnd11an1n64x5 FILLER_36_790 ();
 b15zdnd11an1n64x5 FILLER_36_854 ();
 b15zdnd11an1n64x5 FILLER_36_918 ();
 b15zdnd11an1n64x5 FILLER_36_982 ();
 b15zdnd11an1n64x5 FILLER_36_1046 ();
 b15zdnd11an1n16x5 FILLER_36_1110 ();
 b15zdnd11an1n08x5 FILLER_36_1126 ();
 b15zdnd11an1n04x5 FILLER_36_1134 ();
 b15zdnd00an1n02x5 FILLER_36_1138 ();
 b15zdnd00an1n01x5 FILLER_36_1140 ();
 b15zdnd11an1n64x5 FILLER_36_1146 ();
 b15zdnd11an1n64x5 FILLER_36_1210 ();
 b15zdnd11an1n16x5 FILLER_36_1274 ();
 b15zdnd11an1n08x5 FILLER_36_1290 ();
 b15zdnd00an1n02x5 FILLER_36_1298 ();
 b15zdnd11an1n32x5 FILLER_36_1305 ();
 b15zdnd11an1n08x5 FILLER_36_1337 ();
 b15zdnd11an1n04x5 FILLER_36_1345 ();
 b15zdnd00an1n01x5 FILLER_36_1349 ();
 b15zdnd11an1n64x5 FILLER_36_1359 ();
 b15zdnd11an1n64x5 FILLER_36_1423 ();
 b15zdnd11an1n16x5 FILLER_36_1487 ();
 b15zdnd11an1n04x5 FILLER_36_1506 ();
 b15zdnd11an1n64x5 FILLER_36_1520 ();
 b15zdnd11an1n64x5 FILLER_36_1584 ();
 b15zdnd11an1n64x5 FILLER_36_1648 ();
 b15zdnd11an1n64x5 FILLER_36_1712 ();
 b15zdnd11an1n64x5 FILLER_36_1776 ();
 b15zdnd11an1n64x5 FILLER_36_1840 ();
 b15zdnd11an1n64x5 FILLER_36_1904 ();
 b15zdnd11an1n64x5 FILLER_36_1968 ();
 b15zdnd11an1n64x5 FILLER_36_2032 ();
 b15zdnd11an1n32x5 FILLER_36_2096 ();
 b15zdnd11an1n16x5 FILLER_36_2128 ();
 b15zdnd11an1n08x5 FILLER_36_2144 ();
 b15zdnd00an1n02x5 FILLER_36_2152 ();
 b15zdnd11an1n64x5 FILLER_36_2162 ();
 b15zdnd11an1n32x5 FILLER_36_2226 ();
 b15zdnd11an1n16x5 FILLER_36_2258 ();
 b15zdnd00an1n02x5 FILLER_36_2274 ();
 b15zdnd11an1n64x5 FILLER_37_0 ();
 b15zdnd11an1n64x5 FILLER_37_64 ();
 b15zdnd11an1n64x5 FILLER_37_128 ();
 b15zdnd11an1n64x5 FILLER_37_192 ();
 b15zdnd11an1n32x5 FILLER_37_256 ();
 b15zdnd00an1n01x5 FILLER_37_288 ();
 b15zdnd11an1n04x5 FILLER_37_292 ();
 b15zdnd11an1n04x5 FILLER_37_300 ();
 b15zdnd00an1n01x5 FILLER_37_304 ();
 b15zdnd11an1n64x5 FILLER_37_310 ();
 b15zdnd11an1n64x5 FILLER_37_374 ();
 b15zdnd11an1n64x5 FILLER_37_438 ();
 b15zdnd11an1n64x5 FILLER_37_502 ();
 b15zdnd11an1n64x5 FILLER_37_566 ();
 b15zdnd11an1n64x5 FILLER_37_630 ();
 b15zdnd11an1n64x5 FILLER_37_694 ();
 b15zdnd11an1n08x5 FILLER_37_758 ();
 b15zdnd00an1n02x5 FILLER_37_766 ();
 b15zdnd11an1n64x5 FILLER_37_793 ();
 b15zdnd11an1n64x5 FILLER_37_857 ();
 b15zdnd11an1n32x5 FILLER_37_921 ();
 b15zdnd00an1n02x5 FILLER_37_953 ();
 b15zdnd00an1n01x5 FILLER_37_955 ();
 b15zdnd11an1n04x5 FILLER_37_998 ();
 b15zdnd00an1n02x5 FILLER_37_1002 ();
 b15zdnd00an1n01x5 FILLER_37_1004 ();
 b15zdnd11an1n64x5 FILLER_37_1047 ();
 b15zdnd11an1n64x5 FILLER_37_1111 ();
 b15zdnd11an1n64x5 FILLER_37_1175 ();
 b15zdnd11an1n64x5 FILLER_37_1239 ();
 b15zdnd11an1n64x5 FILLER_37_1303 ();
 b15zdnd11an1n64x5 FILLER_37_1367 ();
 b15zdnd11an1n64x5 FILLER_37_1431 ();
 b15zdnd11an1n08x5 FILLER_37_1495 ();
 b15zdnd00an1n02x5 FILLER_37_1503 ();
 b15zdnd00an1n01x5 FILLER_37_1505 ();
 b15zdnd11an1n64x5 FILLER_37_1511 ();
 b15zdnd11an1n64x5 FILLER_37_1575 ();
 b15zdnd11an1n64x5 FILLER_37_1639 ();
 b15zdnd11an1n64x5 FILLER_37_1703 ();
 b15zdnd11an1n64x5 FILLER_37_1767 ();
 b15zdnd11an1n64x5 FILLER_37_1831 ();
 b15zdnd11an1n64x5 FILLER_37_1895 ();
 b15zdnd11an1n64x5 FILLER_37_1959 ();
 b15zdnd11an1n64x5 FILLER_37_2023 ();
 b15zdnd11an1n64x5 FILLER_37_2087 ();
 b15zdnd11an1n64x5 FILLER_37_2151 ();
 b15zdnd11an1n64x5 FILLER_37_2215 ();
 b15zdnd11an1n04x5 FILLER_37_2279 ();
 b15zdnd00an1n01x5 FILLER_37_2283 ();
 b15zdnd11an1n64x5 FILLER_38_8 ();
 b15zdnd11an1n64x5 FILLER_38_72 ();
 b15zdnd11an1n64x5 FILLER_38_136 ();
 b15zdnd11an1n64x5 FILLER_38_200 ();
 b15zdnd11an1n16x5 FILLER_38_264 ();
 b15zdnd11an1n08x5 FILLER_38_280 ();
 b15zdnd11an1n04x5 FILLER_38_288 ();
 b15zdnd00an1n02x5 FILLER_38_292 ();
 b15zdnd00an1n01x5 FILLER_38_294 ();
 b15zdnd11an1n64x5 FILLER_38_337 ();
 b15zdnd11an1n64x5 FILLER_38_401 ();
 b15zdnd11an1n32x5 FILLER_38_465 ();
 b15zdnd11an1n08x5 FILLER_38_497 ();
 b15zdnd11an1n64x5 FILLER_38_508 ();
 b15zdnd11an1n64x5 FILLER_38_572 ();
 b15zdnd11an1n64x5 FILLER_38_636 ();
 b15zdnd11an1n16x5 FILLER_38_700 ();
 b15zdnd00an1n02x5 FILLER_38_716 ();
 b15zdnd11an1n64x5 FILLER_38_726 ();
 b15zdnd11an1n64x5 FILLER_38_790 ();
 b15zdnd11an1n64x5 FILLER_38_854 ();
 b15zdnd11an1n64x5 FILLER_38_918 ();
 b15zdnd11an1n64x5 FILLER_38_982 ();
 b15zdnd11an1n32x5 FILLER_38_1046 ();
 b15zdnd11an1n16x5 FILLER_38_1078 ();
 b15zdnd00an1n02x5 FILLER_38_1094 ();
 b15zdnd11an1n64x5 FILLER_38_1108 ();
 b15zdnd11an1n64x5 FILLER_38_1172 ();
 b15zdnd11an1n64x5 FILLER_38_1236 ();
 b15zdnd11an1n08x5 FILLER_38_1300 ();
 b15zdnd00an1n02x5 FILLER_38_1308 ();
 b15zdnd00an1n01x5 FILLER_38_1310 ();
 b15zdnd11an1n32x5 FILLER_38_1316 ();
 b15zdnd11an1n08x5 FILLER_38_1348 ();
 b15zdnd11an1n04x5 FILLER_38_1356 ();
 b15zdnd00an1n01x5 FILLER_38_1360 ();
 b15zdnd11an1n64x5 FILLER_38_1369 ();
 b15zdnd11an1n64x5 FILLER_38_1433 ();
 b15zdnd11an1n08x5 FILLER_38_1497 ();
 b15zdnd11an1n04x5 FILLER_38_1505 ();
 b15zdnd00an1n01x5 FILLER_38_1509 ();
 b15zdnd11an1n64x5 FILLER_38_1516 ();
 b15zdnd11an1n64x5 FILLER_38_1580 ();
 b15zdnd11an1n64x5 FILLER_38_1644 ();
 b15zdnd11an1n64x5 FILLER_38_1708 ();
 b15zdnd11an1n32x5 FILLER_38_1772 ();
 b15zdnd11an1n08x5 FILLER_38_1804 ();
 b15zdnd00an1n02x5 FILLER_38_1812 ();
 b15zdnd00an1n01x5 FILLER_38_1814 ();
 b15zdnd11an1n64x5 FILLER_38_1820 ();
 b15zdnd11an1n64x5 FILLER_38_1884 ();
 b15zdnd11an1n64x5 FILLER_38_1948 ();
 b15zdnd11an1n64x5 FILLER_38_2012 ();
 b15zdnd11an1n64x5 FILLER_38_2076 ();
 b15zdnd11an1n08x5 FILLER_38_2140 ();
 b15zdnd11an1n04x5 FILLER_38_2148 ();
 b15zdnd00an1n02x5 FILLER_38_2152 ();
 b15zdnd11an1n64x5 FILLER_38_2162 ();
 b15zdnd11an1n32x5 FILLER_38_2226 ();
 b15zdnd11an1n16x5 FILLER_38_2258 ();
 b15zdnd00an1n02x5 FILLER_38_2274 ();
 b15zdnd11an1n64x5 FILLER_39_0 ();
 b15zdnd11an1n64x5 FILLER_39_64 ();
 b15zdnd11an1n64x5 FILLER_39_128 ();
 b15zdnd11an1n64x5 FILLER_39_192 ();
 b15zdnd11an1n32x5 FILLER_39_256 ();
 b15zdnd00an1n02x5 FILLER_39_288 ();
 b15zdnd00an1n01x5 FILLER_39_290 ();
 b15zdnd11an1n64x5 FILLER_39_294 ();
 b15zdnd11an1n64x5 FILLER_39_358 ();
 b15zdnd11an1n32x5 FILLER_39_422 ();
 b15zdnd11an1n16x5 FILLER_39_454 ();
 b15zdnd11an1n08x5 FILLER_39_470 ();
 b15zdnd11an1n64x5 FILLER_39_530 ();
 b15zdnd11an1n64x5 FILLER_39_594 ();
 b15zdnd11an1n64x5 FILLER_39_658 ();
 b15zdnd11an1n64x5 FILLER_39_722 ();
 b15zdnd11an1n64x5 FILLER_39_786 ();
 b15zdnd11an1n64x5 FILLER_39_850 ();
 b15zdnd11an1n64x5 FILLER_39_914 ();
 b15zdnd11an1n64x5 FILLER_39_978 ();
 b15zdnd11an1n64x5 FILLER_39_1042 ();
 b15zdnd11an1n64x5 FILLER_39_1106 ();
 b15zdnd11an1n64x5 FILLER_39_1170 ();
 b15zdnd11an1n64x5 FILLER_39_1234 ();
 b15zdnd11an1n32x5 FILLER_39_1298 ();
 b15zdnd11an1n08x5 FILLER_39_1330 ();
 b15zdnd00an1n01x5 FILLER_39_1338 ();
 b15zdnd11an1n64x5 FILLER_39_1381 ();
 b15zdnd11an1n32x5 FILLER_39_1445 ();
 b15zdnd11an1n16x5 FILLER_39_1477 ();
 b15zdnd11an1n08x5 FILLER_39_1493 ();
 b15zdnd00an1n02x5 FILLER_39_1501 ();
 b15zdnd00an1n01x5 FILLER_39_1503 ();
 b15zdnd11an1n64x5 FILLER_39_1508 ();
 b15zdnd11an1n64x5 FILLER_39_1572 ();
 b15zdnd11an1n64x5 FILLER_39_1636 ();
 b15zdnd11an1n64x5 FILLER_39_1700 ();
 b15zdnd11an1n64x5 FILLER_39_1764 ();
 b15zdnd11an1n64x5 FILLER_39_1828 ();
 b15zdnd11an1n64x5 FILLER_39_1892 ();
 b15zdnd11an1n64x5 FILLER_39_1956 ();
 b15zdnd11an1n64x5 FILLER_39_2020 ();
 b15zdnd11an1n64x5 FILLER_39_2084 ();
 b15zdnd11an1n64x5 FILLER_39_2148 ();
 b15zdnd11an1n64x5 FILLER_39_2212 ();
 b15zdnd11an1n08x5 FILLER_39_2276 ();
 b15zdnd11an1n64x5 FILLER_40_8 ();
 b15zdnd11an1n64x5 FILLER_40_72 ();
 b15zdnd11an1n64x5 FILLER_40_136 ();
 b15zdnd11an1n64x5 FILLER_40_200 ();
 b15zdnd11an1n16x5 FILLER_40_264 ();
 b15zdnd11an1n08x5 FILLER_40_280 ();
 b15zdnd11an1n04x5 FILLER_40_295 ();
 b15zdnd11an1n64x5 FILLER_40_305 ();
 b15zdnd11an1n64x5 FILLER_40_369 ();
 b15zdnd11an1n32x5 FILLER_40_433 ();
 b15zdnd11an1n16x5 FILLER_40_465 ();
 b15zdnd11an1n08x5 FILLER_40_481 ();
 b15zdnd11an1n04x5 FILLER_40_489 ();
 b15zdnd00an1n02x5 FILLER_40_493 ();
 b15zdnd00an1n01x5 FILLER_40_495 ();
 b15zdnd11an1n04x5 FILLER_40_499 ();
 b15zdnd11an1n04x5 FILLER_40_506 ();
 b15zdnd00an1n02x5 FILLER_40_510 ();
 b15zdnd11an1n64x5 FILLER_40_519 ();
 b15zdnd11an1n64x5 FILLER_40_583 ();
 b15zdnd11an1n64x5 FILLER_40_647 ();
 b15zdnd11an1n04x5 FILLER_40_711 ();
 b15zdnd00an1n02x5 FILLER_40_715 ();
 b15zdnd00an1n01x5 FILLER_40_717 ();
 b15zdnd11an1n32x5 FILLER_40_726 ();
 b15zdnd11an1n08x5 FILLER_40_758 ();
 b15zdnd00an1n02x5 FILLER_40_766 ();
 b15zdnd11an1n64x5 FILLER_40_775 ();
 b15zdnd11an1n64x5 FILLER_40_839 ();
 b15zdnd11an1n64x5 FILLER_40_903 ();
 b15zdnd11an1n64x5 FILLER_40_967 ();
 b15zdnd11an1n64x5 FILLER_40_1031 ();
 b15zdnd11an1n64x5 FILLER_40_1095 ();
 b15zdnd11an1n64x5 FILLER_40_1159 ();
 b15zdnd11an1n64x5 FILLER_40_1223 ();
 b15zdnd11an1n32x5 FILLER_40_1287 ();
 b15zdnd11an1n08x5 FILLER_40_1319 ();
 b15zdnd11an1n04x5 FILLER_40_1327 ();
 b15zdnd00an1n02x5 FILLER_40_1331 ();
 b15zdnd00an1n01x5 FILLER_40_1333 ();
 b15zdnd11an1n64x5 FILLER_40_1376 ();
 b15zdnd11an1n64x5 FILLER_40_1440 ();
 b15zdnd11an1n64x5 FILLER_40_1504 ();
 b15zdnd11an1n64x5 FILLER_40_1568 ();
 b15zdnd11an1n64x5 FILLER_40_1632 ();
 b15zdnd11an1n64x5 FILLER_40_1696 ();
 b15zdnd11an1n64x5 FILLER_40_1760 ();
 b15zdnd11an1n64x5 FILLER_40_1824 ();
 b15zdnd11an1n64x5 FILLER_40_1888 ();
 b15zdnd11an1n64x5 FILLER_40_1952 ();
 b15zdnd11an1n64x5 FILLER_40_2016 ();
 b15zdnd11an1n64x5 FILLER_40_2080 ();
 b15zdnd11an1n08x5 FILLER_40_2144 ();
 b15zdnd00an1n02x5 FILLER_40_2152 ();
 b15zdnd11an1n64x5 FILLER_40_2162 ();
 b15zdnd11an1n32x5 FILLER_40_2226 ();
 b15zdnd11an1n16x5 FILLER_40_2258 ();
 b15zdnd00an1n02x5 FILLER_40_2274 ();
 b15zdnd11an1n64x5 FILLER_41_0 ();
 b15zdnd11an1n64x5 FILLER_41_64 ();
 b15zdnd11an1n64x5 FILLER_41_128 ();
 b15zdnd11an1n64x5 FILLER_41_192 ();
 b15zdnd11an1n16x5 FILLER_41_256 ();
 b15zdnd11an1n04x5 FILLER_41_272 ();
 b15zdnd00an1n02x5 FILLER_41_276 ();
 b15zdnd11an1n64x5 FILLER_41_320 ();
 b15zdnd11an1n64x5 FILLER_41_384 ();
 b15zdnd11an1n32x5 FILLER_41_448 ();
 b15zdnd11an1n16x5 FILLER_41_480 ();
 b15zdnd11an1n08x5 FILLER_41_496 ();
 b15zdnd11an1n64x5 FILLER_41_513 ();
 b15zdnd11an1n64x5 FILLER_41_577 ();
 b15zdnd11an1n64x5 FILLER_41_641 ();
 b15zdnd11an1n64x5 FILLER_41_705 ();
 b15zdnd11an1n16x5 FILLER_41_769 ();
 b15zdnd11an1n08x5 FILLER_41_785 ();
 b15zdnd11an1n04x5 FILLER_41_793 ();
 b15zdnd00an1n02x5 FILLER_41_797 ();
 b15zdnd11an1n32x5 FILLER_41_802 ();
 b15zdnd11an1n08x5 FILLER_41_834 ();
 b15zdnd11an1n04x5 FILLER_41_842 ();
 b15zdnd00an1n02x5 FILLER_41_846 ();
 b15zdnd00an1n01x5 FILLER_41_848 ();
 b15zdnd11an1n64x5 FILLER_41_852 ();
 b15zdnd11an1n64x5 FILLER_41_916 ();
 b15zdnd11an1n64x5 FILLER_41_980 ();
 b15zdnd11an1n64x5 FILLER_41_1044 ();
 b15zdnd11an1n32x5 FILLER_41_1108 ();
 b15zdnd11an1n04x5 FILLER_41_1140 ();
 b15zdnd00an1n02x5 FILLER_41_1144 ();
 b15zdnd00an1n01x5 FILLER_41_1146 ();
 b15zdnd11an1n64x5 FILLER_41_1152 ();
 b15zdnd11an1n64x5 FILLER_41_1216 ();
 b15zdnd11an1n16x5 FILLER_41_1280 ();
 b15zdnd00an1n01x5 FILLER_41_1296 ();
 b15zdnd11an1n04x5 FILLER_41_1306 ();
 b15zdnd11an1n64x5 FILLER_41_1315 ();
 b15zdnd11an1n64x5 FILLER_41_1379 ();
 b15zdnd11an1n32x5 FILLER_41_1443 ();
 b15zdnd11an1n08x5 FILLER_41_1475 ();
 b15zdnd11an1n04x5 FILLER_41_1483 ();
 b15zdnd00an1n02x5 FILLER_41_1487 ();
 b15zdnd00an1n01x5 FILLER_41_1489 ();
 b15zdnd11an1n64x5 FILLER_41_1496 ();
 b15zdnd11an1n64x5 FILLER_41_1560 ();
 b15zdnd11an1n64x5 FILLER_41_1624 ();
 b15zdnd11an1n64x5 FILLER_41_1688 ();
 b15zdnd11an1n64x5 FILLER_41_1752 ();
 b15zdnd11an1n64x5 FILLER_41_1816 ();
 b15zdnd11an1n64x5 FILLER_41_1880 ();
 b15zdnd11an1n64x5 FILLER_41_1944 ();
 b15zdnd11an1n64x5 FILLER_41_2008 ();
 b15zdnd11an1n64x5 FILLER_41_2072 ();
 b15zdnd11an1n64x5 FILLER_41_2136 ();
 b15zdnd11an1n64x5 FILLER_41_2200 ();
 b15zdnd11an1n16x5 FILLER_41_2264 ();
 b15zdnd11an1n04x5 FILLER_41_2280 ();
 b15zdnd11an1n64x5 FILLER_42_8 ();
 b15zdnd11an1n64x5 FILLER_42_72 ();
 b15zdnd11an1n64x5 FILLER_42_136 ();
 b15zdnd11an1n64x5 FILLER_42_200 ();
 b15zdnd11an1n32x5 FILLER_42_264 ();
 b15zdnd11an1n64x5 FILLER_42_338 ();
 b15zdnd11an1n64x5 FILLER_42_402 ();
 b15zdnd11an1n64x5 FILLER_42_466 ();
 b15zdnd11an1n64x5 FILLER_42_530 ();
 b15zdnd11an1n64x5 FILLER_42_594 ();
 b15zdnd11an1n32x5 FILLER_42_658 ();
 b15zdnd11an1n16x5 FILLER_42_690 ();
 b15zdnd11an1n08x5 FILLER_42_706 ();
 b15zdnd11an1n04x5 FILLER_42_714 ();
 b15zdnd11an1n32x5 FILLER_42_726 ();
 b15zdnd11an1n04x5 FILLER_42_758 ();
 b15zdnd00an1n01x5 FILLER_42_762 ();
 b15zdnd11an1n16x5 FILLER_42_803 ();
 b15zdnd00an1n02x5 FILLER_42_819 ();
 b15zdnd00an1n01x5 FILLER_42_821 ();
 b15zdnd11an1n64x5 FILLER_42_874 ();
 b15zdnd11an1n64x5 FILLER_42_938 ();
 b15zdnd11an1n64x5 FILLER_42_1002 ();
 b15zdnd11an1n64x5 FILLER_42_1066 ();
 b15zdnd11an1n64x5 FILLER_42_1130 ();
 b15zdnd11an1n64x5 FILLER_42_1194 ();
 b15zdnd11an1n64x5 FILLER_42_1258 ();
 b15zdnd11an1n64x5 FILLER_42_1322 ();
 b15zdnd11an1n64x5 FILLER_42_1386 ();
 b15zdnd11an1n64x5 FILLER_42_1450 ();
 b15zdnd11an1n64x5 FILLER_42_1514 ();
 b15zdnd11an1n64x5 FILLER_42_1578 ();
 b15zdnd11an1n64x5 FILLER_42_1642 ();
 b15zdnd11an1n64x5 FILLER_42_1706 ();
 b15zdnd11an1n64x5 FILLER_42_1770 ();
 b15zdnd11an1n64x5 FILLER_42_1834 ();
 b15zdnd11an1n64x5 FILLER_42_1898 ();
 b15zdnd11an1n64x5 FILLER_42_1962 ();
 b15zdnd11an1n64x5 FILLER_42_2026 ();
 b15zdnd11an1n64x5 FILLER_42_2090 ();
 b15zdnd11an1n64x5 FILLER_42_2162 ();
 b15zdnd11an1n32x5 FILLER_42_2226 ();
 b15zdnd11an1n16x5 FILLER_42_2258 ();
 b15zdnd00an1n02x5 FILLER_42_2274 ();
 b15zdnd11an1n64x5 FILLER_43_0 ();
 b15zdnd11an1n64x5 FILLER_43_64 ();
 b15zdnd11an1n64x5 FILLER_43_128 ();
 b15zdnd11an1n64x5 FILLER_43_192 ();
 b15zdnd11an1n08x5 FILLER_43_256 ();
 b15zdnd11an1n04x5 FILLER_43_264 ();
 b15zdnd00an1n01x5 FILLER_43_268 ();
 b15zdnd11an1n16x5 FILLER_43_272 ();
 b15zdnd11an1n64x5 FILLER_43_330 ();
 b15zdnd11an1n64x5 FILLER_43_394 ();
 b15zdnd11an1n64x5 FILLER_43_458 ();
 b15zdnd11an1n64x5 FILLER_43_522 ();
 b15zdnd11an1n64x5 FILLER_43_586 ();
 b15zdnd11an1n64x5 FILLER_43_650 ();
 b15zdnd11an1n64x5 FILLER_43_714 ();
 b15zdnd11an1n16x5 FILLER_43_778 ();
 b15zdnd11an1n04x5 FILLER_43_794 ();
 b15zdnd00an1n01x5 FILLER_43_798 ();
 b15zdnd11an1n32x5 FILLER_43_802 ();
 b15zdnd11an1n04x5 FILLER_43_834 ();
 b15zdnd00an1n02x5 FILLER_43_838 ();
 b15zdnd00an1n01x5 FILLER_43_840 ();
 b15zdnd11an1n04x5 FILLER_43_844 ();
 b15zdnd11an1n64x5 FILLER_43_851 ();
 b15zdnd11an1n64x5 FILLER_43_915 ();
 b15zdnd11an1n64x5 FILLER_43_979 ();
 b15zdnd11an1n64x5 FILLER_43_1043 ();
 b15zdnd11an1n64x5 FILLER_43_1107 ();
 b15zdnd11an1n64x5 FILLER_43_1171 ();
 b15zdnd11an1n64x5 FILLER_43_1235 ();
 b15zdnd11an1n64x5 FILLER_43_1299 ();
 b15zdnd11an1n64x5 FILLER_43_1363 ();
 b15zdnd11an1n64x5 FILLER_43_1427 ();
 b15zdnd11an1n64x5 FILLER_43_1491 ();
 b15zdnd11an1n64x5 FILLER_43_1555 ();
 b15zdnd11an1n64x5 FILLER_43_1619 ();
 b15zdnd11an1n64x5 FILLER_43_1683 ();
 b15zdnd11an1n64x5 FILLER_43_1747 ();
 b15zdnd11an1n04x5 FILLER_43_1811 ();
 b15zdnd11an1n64x5 FILLER_43_1857 ();
 b15zdnd11an1n64x5 FILLER_43_1921 ();
 b15zdnd11an1n64x5 FILLER_43_1985 ();
 b15zdnd11an1n64x5 FILLER_43_2049 ();
 b15zdnd11an1n64x5 FILLER_43_2113 ();
 b15zdnd11an1n64x5 FILLER_43_2177 ();
 b15zdnd11an1n32x5 FILLER_43_2241 ();
 b15zdnd11an1n08x5 FILLER_43_2273 ();
 b15zdnd00an1n02x5 FILLER_43_2281 ();
 b15zdnd00an1n01x5 FILLER_43_2283 ();
 b15zdnd11an1n64x5 FILLER_44_8 ();
 b15zdnd11an1n64x5 FILLER_44_72 ();
 b15zdnd11an1n64x5 FILLER_44_136 ();
 b15zdnd11an1n32x5 FILLER_44_200 ();
 b15zdnd11an1n08x5 FILLER_44_232 ();
 b15zdnd00an1n02x5 FILLER_44_240 ();
 b15zdnd11an1n64x5 FILLER_44_294 ();
 b15zdnd11an1n64x5 FILLER_44_358 ();
 b15zdnd11an1n64x5 FILLER_44_422 ();
 b15zdnd11an1n64x5 FILLER_44_486 ();
 b15zdnd11an1n64x5 FILLER_44_550 ();
 b15zdnd11an1n64x5 FILLER_44_614 ();
 b15zdnd11an1n32x5 FILLER_44_678 ();
 b15zdnd11an1n08x5 FILLER_44_710 ();
 b15zdnd11an1n64x5 FILLER_44_726 ();
 b15zdnd11an1n64x5 FILLER_44_790 ();
 b15zdnd11an1n64x5 FILLER_44_854 ();
 b15zdnd11an1n64x5 FILLER_44_918 ();
 b15zdnd11an1n64x5 FILLER_44_982 ();
 b15zdnd11an1n64x5 FILLER_44_1046 ();
 b15zdnd11an1n04x5 FILLER_44_1110 ();
 b15zdnd00an1n02x5 FILLER_44_1114 ();
 b15zdnd00an1n01x5 FILLER_44_1116 ();
 b15zdnd11an1n64x5 FILLER_44_1127 ();
 b15zdnd11an1n64x5 FILLER_44_1191 ();
 b15zdnd11an1n64x5 FILLER_44_1255 ();
 b15zdnd11an1n64x5 FILLER_44_1319 ();
 b15zdnd11an1n64x5 FILLER_44_1383 ();
 b15zdnd11an1n64x5 FILLER_44_1447 ();
 b15zdnd11an1n64x5 FILLER_44_1511 ();
 b15zdnd11an1n64x5 FILLER_44_1575 ();
 b15zdnd11an1n64x5 FILLER_44_1639 ();
 b15zdnd11an1n64x5 FILLER_44_1703 ();
 b15zdnd11an1n32x5 FILLER_44_1767 ();
 b15zdnd11an1n04x5 FILLER_44_1799 ();
 b15zdnd00an1n02x5 FILLER_44_1803 ();
 b15zdnd11an1n64x5 FILLER_44_1847 ();
 b15zdnd11an1n64x5 FILLER_44_1911 ();
 b15zdnd11an1n64x5 FILLER_44_1975 ();
 b15zdnd11an1n16x5 FILLER_44_2039 ();
 b15zdnd11an1n08x5 FILLER_44_2055 ();
 b15zdnd00an1n01x5 FILLER_44_2063 ();
 b15zdnd11an1n08x5 FILLER_44_2070 ();
 b15zdnd11an1n04x5 FILLER_44_2078 ();
 b15zdnd00an1n02x5 FILLER_44_2082 ();
 b15zdnd00an1n01x5 FILLER_44_2084 ();
 b15zdnd11an1n04x5 FILLER_44_2088 ();
 b15zdnd11an1n32x5 FILLER_44_2095 ();
 b15zdnd11an1n16x5 FILLER_44_2127 ();
 b15zdnd11an1n08x5 FILLER_44_2143 ();
 b15zdnd00an1n02x5 FILLER_44_2151 ();
 b15zdnd00an1n01x5 FILLER_44_2153 ();
 b15zdnd11an1n64x5 FILLER_44_2162 ();
 b15zdnd11an1n32x5 FILLER_44_2226 ();
 b15zdnd11an1n16x5 FILLER_44_2258 ();
 b15zdnd00an1n02x5 FILLER_44_2274 ();
 b15zdnd11an1n64x5 FILLER_45_0 ();
 b15zdnd11an1n64x5 FILLER_45_64 ();
 b15zdnd11an1n64x5 FILLER_45_128 ();
 b15zdnd11an1n64x5 FILLER_45_192 ();
 b15zdnd11an1n08x5 FILLER_45_256 ();
 b15zdnd11an1n04x5 FILLER_45_264 ();
 b15zdnd11an1n64x5 FILLER_45_271 ();
 b15zdnd11an1n64x5 FILLER_45_335 ();
 b15zdnd11an1n64x5 FILLER_45_399 ();
 b15zdnd11an1n64x5 FILLER_45_463 ();
 b15zdnd11an1n64x5 FILLER_45_527 ();
 b15zdnd11an1n64x5 FILLER_45_591 ();
 b15zdnd11an1n64x5 FILLER_45_655 ();
 b15zdnd11an1n64x5 FILLER_45_719 ();
 b15zdnd11an1n08x5 FILLER_45_783 ();
 b15zdnd00an1n01x5 FILLER_45_791 ();
 b15zdnd11an1n04x5 FILLER_45_803 ();
 b15zdnd11an1n64x5 FILLER_45_846 ();
 b15zdnd11an1n64x5 FILLER_45_910 ();
 b15zdnd11an1n64x5 FILLER_45_974 ();
 b15zdnd11an1n64x5 FILLER_45_1038 ();
 b15zdnd11an1n64x5 FILLER_45_1102 ();
 b15zdnd11an1n16x5 FILLER_45_1166 ();
 b15zdnd11an1n08x5 FILLER_45_1182 ();
 b15zdnd11an1n04x5 FILLER_45_1190 ();
 b15zdnd00an1n01x5 FILLER_45_1194 ();
 b15zdnd11an1n64x5 FILLER_45_1216 ();
 b15zdnd11an1n64x5 FILLER_45_1280 ();
 b15zdnd11an1n64x5 FILLER_45_1344 ();
 b15zdnd11an1n64x5 FILLER_45_1408 ();
 b15zdnd11an1n64x5 FILLER_45_1472 ();
 b15zdnd11an1n64x5 FILLER_45_1536 ();
 b15zdnd11an1n64x5 FILLER_45_1600 ();
 b15zdnd11an1n64x5 FILLER_45_1664 ();
 b15zdnd11an1n64x5 FILLER_45_1728 ();
 b15zdnd11an1n64x5 FILLER_45_1792 ();
 b15zdnd11an1n64x5 FILLER_45_1856 ();
 b15zdnd11an1n64x5 FILLER_45_1920 ();
 b15zdnd11an1n32x5 FILLER_45_1984 ();
 b15zdnd11an1n16x5 FILLER_45_2016 ();
 b15zdnd11an1n04x5 FILLER_45_2032 ();
 b15zdnd11an1n04x5 FILLER_45_2042 ();
 b15zdnd11an1n04x5 FILLER_45_2054 ();
 b15zdnd00an1n02x5 FILLER_45_2058 ();
 b15zdnd11an1n64x5 FILLER_45_2112 ();
 b15zdnd11an1n64x5 FILLER_45_2176 ();
 b15zdnd11an1n32x5 FILLER_45_2240 ();
 b15zdnd11an1n08x5 FILLER_45_2272 ();
 b15zdnd11an1n04x5 FILLER_45_2280 ();
 b15zdnd11an1n64x5 FILLER_46_8 ();
 b15zdnd11an1n64x5 FILLER_46_72 ();
 b15zdnd11an1n64x5 FILLER_46_136 ();
 b15zdnd11an1n64x5 FILLER_46_200 ();
 b15zdnd11an1n04x5 FILLER_46_264 ();
 b15zdnd00an1n01x5 FILLER_46_268 ();
 b15zdnd11an1n64x5 FILLER_46_272 ();
 b15zdnd11an1n64x5 FILLER_46_336 ();
 b15zdnd11an1n64x5 FILLER_46_400 ();
 b15zdnd11an1n64x5 FILLER_46_464 ();
 b15zdnd11an1n64x5 FILLER_46_528 ();
 b15zdnd11an1n64x5 FILLER_46_592 ();
 b15zdnd11an1n32x5 FILLER_46_656 ();
 b15zdnd11an1n16x5 FILLER_46_688 ();
 b15zdnd11an1n08x5 FILLER_46_704 ();
 b15zdnd11an1n04x5 FILLER_46_712 ();
 b15zdnd00an1n02x5 FILLER_46_716 ();
 b15zdnd11an1n64x5 FILLER_46_726 ();
 b15zdnd11an1n16x5 FILLER_46_790 ();
 b15zdnd11an1n08x5 FILLER_46_806 ();
 b15zdnd00an1n01x5 FILLER_46_814 ();
 b15zdnd11an1n64x5 FILLER_46_822 ();
 b15zdnd11an1n64x5 FILLER_46_886 ();
 b15zdnd11an1n64x5 FILLER_46_950 ();
 b15zdnd11an1n64x5 FILLER_46_1014 ();
 b15zdnd11an1n64x5 FILLER_46_1078 ();
 b15zdnd11an1n64x5 FILLER_46_1142 ();
 b15zdnd11an1n64x5 FILLER_46_1206 ();
 b15zdnd11an1n64x5 FILLER_46_1270 ();
 b15zdnd11an1n32x5 FILLER_46_1334 ();
 b15zdnd11an1n04x5 FILLER_46_1366 ();
 b15zdnd00an1n02x5 FILLER_46_1370 ();
 b15zdnd00an1n01x5 FILLER_46_1372 ();
 b15zdnd11an1n64x5 FILLER_46_1383 ();
 b15zdnd11an1n64x5 FILLER_46_1447 ();
 b15zdnd11an1n64x5 FILLER_46_1511 ();
 b15zdnd11an1n64x5 FILLER_46_1575 ();
 b15zdnd11an1n64x5 FILLER_46_1639 ();
 b15zdnd11an1n64x5 FILLER_46_1703 ();
 b15zdnd11an1n64x5 FILLER_46_1767 ();
 b15zdnd11an1n64x5 FILLER_46_1831 ();
 b15zdnd11an1n64x5 FILLER_46_1895 ();
 b15zdnd11an1n32x5 FILLER_46_1959 ();
 b15zdnd11an1n08x5 FILLER_46_1994 ();
 b15zdnd11an1n08x5 FILLER_46_2005 ();
 b15zdnd00an1n01x5 FILLER_46_2013 ();
 b15zdnd11an1n04x5 FILLER_46_2024 ();
 b15zdnd11an1n04x5 FILLER_46_2032 ();
 b15zdnd00an1n02x5 FILLER_46_2036 ();
 b15zdnd11an1n08x5 FILLER_46_2080 ();
 b15zdnd11an1n16x5 FILLER_46_2130 ();
 b15zdnd11an1n08x5 FILLER_46_2146 ();
 b15zdnd11an1n64x5 FILLER_46_2162 ();
 b15zdnd11an1n32x5 FILLER_46_2226 ();
 b15zdnd11an1n16x5 FILLER_46_2258 ();
 b15zdnd00an1n02x5 FILLER_46_2274 ();
 b15zdnd11an1n64x5 FILLER_47_0 ();
 b15zdnd11an1n64x5 FILLER_47_64 ();
 b15zdnd11an1n64x5 FILLER_47_128 ();
 b15zdnd11an1n64x5 FILLER_47_192 ();
 b15zdnd11an1n64x5 FILLER_47_256 ();
 b15zdnd11an1n64x5 FILLER_47_320 ();
 b15zdnd11an1n64x5 FILLER_47_384 ();
 b15zdnd11an1n64x5 FILLER_47_448 ();
 b15zdnd11an1n64x5 FILLER_47_512 ();
 b15zdnd11an1n64x5 FILLER_47_576 ();
 b15zdnd11an1n64x5 FILLER_47_640 ();
 b15zdnd11an1n64x5 FILLER_47_704 ();
 b15zdnd11an1n64x5 FILLER_47_768 ();
 b15zdnd11an1n64x5 FILLER_47_832 ();
 b15zdnd11an1n64x5 FILLER_47_896 ();
 b15zdnd11an1n16x5 FILLER_47_960 ();
 b15zdnd11an1n04x5 FILLER_47_976 ();
 b15zdnd00an1n01x5 FILLER_47_980 ();
 b15zdnd11an1n64x5 FILLER_47_984 ();
 b15zdnd11an1n16x5 FILLER_47_1048 ();
 b15zdnd11an1n08x5 FILLER_47_1064 ();
 b15zdnd11an1n64x5 FILLER_47_1075 ();
 b15zdnd11an1n64x5 FILLER_47_1139 ();
 b15zdnd11an1n64x5 FILLER_47_1203 ();
 b15zdnd11an1n64x5 FILLER_47_1267 ();
 b15zdnd11an1n64x5 FILLER_47_1331 ();
 b15zdnd11an1n64x5 FILLER_47_1395 ();
 b15zdnd11an1n32x5 FILLER_47_1459 ();
 b15zdnd11an1n16x5 FILLER_47_1491 ();
 b15zdnd11an1n08x5 FILLER_47_1507 ();
 b15zdnd11an1n04x5 FILLER_47_1515 ();
 b15zdnd00an1n02x5 FILLER_47_1519 ();
 b15zdnd00an1n01x5 FILLER_47_1521 ();
 b15zdnd11an1n64x5 FILLER_47_1525 ();
 b15zdnd11an1n32x5 FILLER_47_1589 ();
 b15zdnd00an1n02x5 FILLER_47_1621 ();
 b15zdnd11an1n04x5 FILLER_47_1626 ();
 b15zdnd11an1n64x5 FILLER_47_1633 ();
 b15zdnd11an1n32x5 FILLER_47_1697 ();
 b15zdnd11an1n08x5 FILLER_47_1729 ();
 b15zdnd11an1n04x5 FILLER_47_1737 ();
 b15zdnd00an1n02x5 FILLER_47_1741 ();
 b15zdnd00an1n01x5 FILLER_47_1743 ();
 b15zdnd11an1n64x5 FILLER_47_1753 ();
 b15zdnd11an1n64x5 FILLER_47_1817 ();
 b15zdnd11an1n32x5 FILLER_47_1881 ();
 b15zdnd00an1n02x5 FILLER_47_1913 ();
 b15zdnd11an1n64x5 FILLER_47_1918 ();
 b15zdnd11an1n04x5 FILLER_47_1982 ();
 b15zdnd11an1n04x5 FILLER_47_1992 ();
 b15zdnd11an1n04x5 FILLER_47_2005 ();
 b15zdnd11an1n08x5 FILLER_47_2051 ();
 b15zdnd11an1n04x5 FILLER_47_2059 ();
 b15zdnd00an1n02x5 FILLER_47_2063 ();
 b15zdnd11an1n64x5 FILLER_47_2107 ();
 b15zdnd11an1n64x5 FILLER_47_2171 ();
 b15zdnd11an1n32x5 FILLER_47_2235 ();
 b15zdnd11an1n16x5 FILLER_47_2267 ();
 b15zdnd00an1n01x5 FILLER_47_2283 ();
 b15zdnd11an1n64x5 FILLER_48_8 ();
 b15zdnd11an1n64x5 FILLER_48_72 ();
 b15zdnd11an1n64x5 FILLER_48_136 ();
 b15zdnd11an1n64x5 FILLER_48_200 ();
 b15zdnd11an1n64x5 FILLER_48_264 ();
 b15zdnd11an1n64x5 FILLER_48_328 ();
 b15zdnd11an1n04x5 FILLER_48_392 ();
 b15zdnd00an1n02x5 FILLER_48_396 ();
 b15zdnd11an1n64x5 FILLER_48_401 ();
 b15zdnd11an1n64x5 FILLER_48_465 ();
 b15zdnd11an1n64x5 FILLER_48_529 ();
 b15zdnd11an1n64x5 FILLER_48_593 ();
 b15zdnd11an1n32x5 FILLER_48_657 ();
 b15zdnd11an1n16x5 FILLER_48_689 ();
 b15zdnd11an1n08x5 FILLER_48_705 ();
 b15zdnd11an1n04x5 FILLER_48_713 ();
 b15zdnd00an1n01x5 FILLER_48_717 ();
 b15zdnd11an1n64x5 FILLER_48_726 ();
 b15zdnd11an1n64x5 FILLER_48_790 ();
 b15zdnd11an1n64x5 FILLER_48_854 ();
 b15zdnd11an1n32x5 FILLER_48_918 ();
 b15zdnd11an1n04x5 FILLER_48_950 ();
 b15zdnd11an1n32x5 FILLER_48_1006 ();
 b15zdnd11an1n04x5 FILLER_48_1038 ();
 b15zdnd00an1n02x5 FILLER_48_1042 ();
 b15zdnd00an1n01x5 FILLER_48_1044 ();
 b15zdnd11an1n32x5 FILLER_48_1097 ();
 b15zdnd11an1n16x5 FILLER_48_1129 ();
 b15zdnd00an1n02x5 FILLER_48_1145 ();
 b15zdnd11an1n64x5 FILLER_48_1150 ();
 b15zdnd11an1n64x5 FILLER_48_1214 ();
 b15zdnd11an1n32x5 FILLER_48_1278 ();
 b15zdnd11an1n16x5 FILLER_48_1310 ();
 b15zdnd11an1n04x5 FILLER_48_1326 ();
 b15zdnd11an1n04x5 FILLER_48_1333 ();
 b15zdnd11an1n64x5 FILLER_48_1340 ();
 b15zdnd11an1n32x5 FILLER_48_1404 ();
 b15zdnd11an1n08x5 FILLER_48_1436 ();
 b15zdnd00an1n01x5 FILLER_48_1444 ();
 b15zdnd11an1n64x5 FILLER_48_1448 ();
 b15zdnd11an1n08x5 FILLER_48_1512 ();
 b15zdnd00an1n02x5 FILLER_48_1520 ();
 b15zdnd11an1n04x5 FILLER_48_1525 ();
 b15zdnd00an1n02x5 FILLER_48_1529 ();
 b15zdnd11an1n64x5 FILLER_48_1534 ();
 b15zdnd11an1n04x5 FILLER_48_1598 ();
 b15zdnd00an1n02x5 FILLER_48_1602 ();
 b15zdnd00an1n01x5 FILLER_48_1604 ();
 b15zdnd11an1n64x5 FILLER_48_1657 ();
 b15zdnd11an1n64x5 FILLER_48_1721 ();
 b15zdnd00an1n02x5 FILLER_48_1785 ();
 b15zdnd00an1n01x5 FILLER_48_1787 ();
 b15zdnd11an1n64x5 FILLER_48_1791 ();
 b15zdnd11an1n16x5 FILLER_48_1855 ();
 b15zdnd11an1n08x5 FILLER_48_1871 ();
 b15zdnd00an1n02x5 FILLER_48_1879 ();
 b15zdnd11an1n32x5 FILLER_48_1921 ();
 b15zdnd11an1n08x5 FILLER_48_1953 ();
 b15zdnd11an1n04x5 FILLER_48_1961 ();
 b15zdnd00an1n01x5 FILLER_48_1965 ();
 b15zdnd11an1n04x5 FILLER_48_2018 ();
 b15zdnd11an1n32x5 FILLER_48_2028 ();
 b15zdnd11an1n16x5 FILLER_48_2060 ();
 b15zdnd11an1n08x5 FILLER_48_2076 ();
 b15zdnd00an1n01x5 FILLER_48_2084 ();
 b15zdnd11an1n64x5 FILLER_48_2088 ();
 b15zdnd00an1n02x5 FILLER_48_2152 ();
 b15zdnd11an1n64x5 FILLER_48_2162 ();
 b15zdnd11an1n32x5 FILLER_48_2226 ();
 b15zdnd11an1n16x5 FILLER_48_2258 ();
 b15zdnd00an1n02x5 FILLER_48_2274 ();
 b15zdnd11an1n64x5 FILLER_49_0 ();
 b15zdnd11an1n64x5 FILLER_49_64 ();
 b15zdnd11an1n64x5 FILLER_49_128 ();
 b15zdnd11an1n64x5 FILLER_49_192 ();
 b15zdnd11an1n64x5 FILLER_49_256 ();
 b15zdnd11an1n64x5 FILLER_49_320 ();
 b15zdnd11an1n08x5 FILLER_49_384 ();
 b15zdnd11an1n04x5 FILLER_49_392 ();
 b15zdnd11an1n04x5 FILLER_49_399 ();
 b15zdnd00an1n01x5 FILLER_49_403 ();
 b15zdnd11an1n64x5 FILLER_49_407 ();
 b15zdnd11an1n64x5 FILLER_49_471 ();
 b15zdnd11an1n64x5 FILLER_49_535 ();
 b15zdnd11an1n64x5 FILLER_49_599 ();
 b15zdnd11an1n64x5 FILLER_49_663 ();
 b15zdnd11an1n64x5 FILLER_49_727 ();
 b15zdnd11an1n64x5 FILLER_49_791 ();
 b15zdnd11an1n64x5 FILLER_49_855 ();
 b15zdnd11an1n32x5 FILLER_49_919 ();
 b15zdnd11an1n16x5 FILLER_49_951 ();
 b15zdnd11an1n08x5 FILLER_49_967 ();
 b15zdnd11an1n04x5 FILLER_49_975 ();
 b15zdnd00an1n01x5 FILLER_49_979 ();
 b15zdnd11an1n04x5 FILLER_49_983 ();
 b15zdnd11an1n64x5 FILLER_49_990 ();
 b15zdnd11an1n08x5 FILLER_49_1054 ();
 b15zdnd00an1n02x5 FILLER_49_1062 ();
 b15zdnd11an1n04x5 FILLER_49_1067 ();
 b15zdnd11an1n32x5 FILLER_49_1074 ();
 b15zdnd11an1n16x5 FILLER_49_1106 ();
 b15zdnd11an1n16x5 FILLER_49_1174 ();
 b15zdnd11an1n08x5 FILLER_49_1190 ();
 b15zdnd11an1n04x5 FILLER_49_1198 ();
 b15zdnd00an1n02x5 FILLER_49_1202 ();
 b15zdnd00an1n01x5 FILLER_49_1204 ();
 b15zdnd11an1n64x5 FILLER_49_1212 ();
 b15zdnd11an1n32x5 FILLER_49_1276 ();
 b15zdnd11an1n04x5 FILLER_49_1308 ();
 b15zdnd11an1n32x5 FILLER_49_1364 ();
 b15zdnd11an1n04x5 FILLER_49_1396 ();
 b15zdnd00an1n02x5 FILLER_49_1400 ();
 b15zdnd00an1n01x5 FILLER_49_1402 ();
 b15zdnd11an1n04x5 FILLER_49_1410 ();
 b15zdnd11an1n32x5 FILLER_49_1456 ();
 b15zdnd11an1n08x5 FILLER_49_1488 ();
 b15zdnd00an1n02x5 FILLER_49_1496 ();
 b15zdnd00an1n01x5 FILLER_49_1498 ();
 b15zdnd11an1n64x5 FILLER_49_1551 ();
 b15zdnd11an1n08x5 FILLER_49_1615 ();
 b15zdnd11an1n04x5 FILLER_49_1623 ();
 b15zdnd00an1n02x5 FILLER_49_1627 ();
 b15zdnd00an1n01x5 FILLER_49_1629 ();
 b15zdnd11an1n64x5 FILLER_49_1633 ();
 b15zdnd11an1n64x5 FILLER_49_1697 ();
 b15zdnd00an1n01x5 FILLER_49_1761 ();
 b15zdnd11an1n64x5 FILLER_49_1814 ();
 b15zdnd11an1n32x5 FILLER_49_1878 ();
 b15zdnd11an1n04x5 FILLER_49_1910 ();
 b15zdnd00an1n02x5 FILLER_49_1914 ();
 b15zdnd00an1n01x5 FILLER_49_1916 ();
 b15zdnd11an1n32x5 FILLER_49_1920 ();
 b15zdnd11an1n16x5 FILLER_49_1952 ();
 b15zdnd11an1n08x5 FILLER_49_1968 ();
 b15zdnd11an1n04x5 FILLER_49_1976 ();
 b15zdnd11an1n04x5 FILLER_49_1983 ();
 b15zdnd11an1n64x5 FILLER_49_2029 ();
 b15zdnd11an1n64x5 FILLER_49_2093 ();
 b15zdnd11an1n64x5 FILLER_49_2157 ();
 b15zdnd11an1n32x5 FILLER_49_2221 ();
 b15zdnd11an1n16x5 FILLER_49_2253 ();
 b15zdnd11an1n08x5 FILLER_49_2269 ();
 b15zdnd11an1n04x5 FILLER_49_2277 ();
 b15zdnd00an1n02x5 FILLER_49_2281 ();
 b15zdnd00an1n01x5 FILLER_49_2283 ();
 b15zdnd11an1n64x5 FILLER_50_8 ();
 b15zdnd11an1n64x5 FILLER_50_72 ();
 b15zdnd11an1n64x5 FILLER_50_136 ();
 b15zdnd11an1n64x5 FILLER_50_200 ();
 b15zdnd11an1n64x5 FILLER_50_264 ();
 b15zdnd11an1n32x5 FILLER_50_328 ();
 b15zdnd11an1n08x5 FILLER_50_360 ();
 b15zdnd11an1n04x5 FILLER_50_368 ();
 b15zdnd00an1n01x5 FILLER_50_372 ();
 b15zdnd11an1n64x5 FILLER_50_425 ();
 b15zdnd11an1n64x5 FILLER_50_489 ();
 b15zdnd11an1n64x5 FILLER_50_553 ();
 b15zdnd11an1n64x5 FILLER_50_617 ();
 b15zdnd11an1n32x5 FILLER_50_681 ();
 b15zdnd11an1n04x5 FILLER_50_713 ();
 b15zdnd00an1n01x5 FILLER_50_717 ();
 b15zdnd11an1n64x5 FILLER_50_726 ();
 b15zdnd11an1n64x5 FILLER_50_790 ();
 b15zdnd11an1n64x5 FILLER_50_854 ();
 b15zdnd11an1n64x5 FILLER_50_918 ();
 b15zdnd11an1n64x5 FILLER_50_982 ();
 b15zdnd11an1n64x5 FILLER_50_1046 ();
 b15zdnd11an1n16x5 FILLER_50_1110 ();
 b15zdnd11an1n08x5 FILLER_50_1126 ();
 b15zdnd00an1n01x5 FILLER_50_1134 ();
 b15zdnd11an1n04x5 FILLER_50_1138 ();
 b15zdnd11an1n16x5 FILLER_50_1145 ();
 b15zdnd11an1n08x5 FILLER_50_1161 ();
 b15zdnd11an1n04x5 FILLER_50_1169 ();
 b15zdnd11an1n64x5 FILLER_50_1199 ();
 b15zdnd11an1n64x5 FILLER_50_1263 ();
 b15zdnd11an1n08x5 FILLER_50_1327 ();
 b15zdnd00an1n02x5 FILLER_50_1335 ();
 b15zdnd11an1n64x5 FILLER_50_1340 ();
 b15zdnd11an1n16x5 FILLER_50_1404 ();
 b15zdnd11an1n32x5 FILLER_50_1472 ();
 b15zdnd00an1n02x5 FILLER_50_1504 ();
 b15zdnd11an1n64x5 FILLER_50_1510 ();
 b15zdnd11an1n64x5 FILLER_50_1574 ();
 b15zdnd11an1n64x5 FILLER_50_1638 ();
 b15zdnd11an1n64x5 FILLER_50_1702 ();
 b15zdnd11an1n16x5 FILLER_50_1766 ();
 b15zdnd11an1n04x5 FILLER_50_1782 ();
 b15zdnd00an1n01x5 FILLER_50_1786 ();
 b15zdnd11an1n64x5 FILLER_50_1790 ();
 b15zdnd11an1n64x5 FILLER_50_1854 ();
 b15zdnd11an1n64x5 FILLER_50_1918 ();
 b15zdnd11an1n04x5 FILLER_50_1982 ();
 b15zdnd00an1n02x5 FILLER_50_1986 ();
 b15zdnd00an1n01x5 FILLER_50_1988 ();
 b15zdnd11an1n04x5 FILLER_50_1992 ();
 b15zdnd11an1n04x5 FILLER_50_2001 ();
 b15zdnd11an1n64x5 FILLER_50_2010 ();
 b15zdnd11an1n64x5 FILLER_50_2074 ();
 b15zdnd11an1n16x5 FILLER_50_2138 ();
 b15zdnd11an1n64x5 FILLER_50_2162 ();
 b15zdnd11an1n32x5 FILLER_50_2226 ();
 b15zdnd11an1n16x5 FILLER_50_2258 ();
 b15zdnd00an1n02x5 FILLER_50_2274 ();
 b15zdnd11an1n64x5 FILLER_51_0 ();
 b15zdnd11an1n64x5 FILLER_51_64 ();
 b15zdnd11an1n64x5 FILLER_51_128 ();
 b15zdnd11an1n64x5 FILLER_51_192 ();
 b15zdnd11an1n64x5 FILLER_51_256 ();
 b15zdnd11an1n64x5 FILLER_51_320 ();
 b15zdnd11an1n64x5 FILLER_51_384 ();
 b15zdnd11an1n64x5 FILLER_51_448 ();
 b15zdnd11an1n64x5 FILLER_51_512 ();
 b15zdnd11an1n64x5 FILLER_51_576 ();
 b15zdnd11an1n64x5 FILLER_51_640 ();
 b15zdnd11an1n64x5 FILLER_51_704 ();
 b15zdnd11an1n64x5 FILLER_51_768 ();
 b15zdnd11an1n64x5 FILLER_51_832 ();
 b15zdnd11an1n64x5 FILLER_51_896 ();
 b15zdnd11an1n64x5 FILLER_51_960 ();
 b15zdnd11an1n64x5 FILLER_51_1024 ();
 b15zdnd11an1n32x5 FILLER_51_1088 ();
 b15zdnd11an1n16x5 FILLER_51_1120 ();
 b15zdnd11an1n08x5 FILLER_51_1136 ();
 b15zdnd11an1n04x5 FILLER_51_1144 ();
 b15zdnd11an1n04x5 FILLER_51_1155 ();
 b15zdnd11an1n04x5 FILLER_51_1169 ();
 b15zdnd11an1n64x5 FILLER_51_1215 ();
 b15zdnd11an1n64x5 FILLER_51_1279 ();
 b15zdnd11an1n04x5 FILLER_51_1343 ();
 b15zdnd11an1n64x5 FILLER_51_1350 ();
 b15zdnd11an1n04x5 FILLER_51_1414 ();
 b15zdnd11an1n04x5 FILLER_51_1449 ();
 b15zdnd11an1n08x5 FILLER_51_1456 ();
 b15zdnd00an1n02x5 FILLER_51_1464 ();
 b15zdnd11an1n64x5 FILLER_51_1508 ();
 b15zdnd11an1n64x5 FILLER_51_1572 ();
 b15zdnd11an1n16x5 FILLER_51_1636 ();
 b15zdnd11an1n08x5 FILLER_51_1652 ();
 b15zdnd11an1n04x5 FILLER_51_1660 ();
 b15zdnd11an1n04x5 FILLER_51_1670 ();
 b15zdnd00an1n02x5 FILLER_51_1674 ();
 b15zdnd11an1n04x5 FILLER_51_1680 ();
 b15zdnd11an1n64x5 FILLER_51_1687 ();
 b15zdnd11an1n32x5 FILLER_51_1751 ();
 b15zdnd00an1n02x5 FILLER_51_1783 ();
 b15zdnd00an1n01x5 FILLER_51_1785 ();
 b15zdnd11an1n64x5 FILLER_51_1789 ();
 b15zdnd11an1n04x5 FILLER_51_1853 ();
 b15zdnd11an1n04x5 FILLER_51_1899 ();
 b15zdnd00an1n02x5 FILLER_51_1903 ();
 b15zdnd00an1n01x5 FILLER_51_1905 ();
 b15zdnd11an1n64x5 FILLER_51_1910 ();
 b15zdnd11an1n64x5 FILLER_51_1974 ();
 b15zdnd11an1n64x5 FILLER_51_2038 ();
 b15zdnd11an1n64x5 FILLER_51_2102 ();
 b15zdnd11an1n64x5 FILLER_51_2166 ();
 b15zdnd11an1n32x5 FILLER_51_2230 ();
 b15zdnd11an1n16x5 FILLER_51_2262 ();
 b15zdnd11an1n04x5 FILLER_51_2278 ();
 b15zdnd00an1n02x5 FILLER_51_2282 ();
 b15zdnd11an1n64x5 FILLER_52_8 ();
 b15zdnd11an1n64x5 FILLER_52_72 ();
 b15zdnd11an1n64x5 FILLER_52_136 ();
 b15zdnd11an1n64x5 FILLER_52_200 ();
 b15zdnd11an1n64x5 FILLER_52_264 ();
 b15zdnd11an1n64x5 FILLER_52_328 ();
 b15zdnd11an1n64x5 FILLER_52_392 ();
 b15zdnd11an1n32x5 FILLER_52_456 ();
 b15zdnd11an1n16x5 FILLER_52_488 ();
 b15zdnd00an1n01x5 FILLER_52_504 ();
 b15zdnd11an1n04x5 FILLER_52_508 ();
 b15zdnd00an1n01x5 FILLER_52_512 ();
 b15zdnd11an1n64x5 FILLER_52_555 ();
 b15zdnd11an1n64x5 FILLER_52_619 ();
 b15zdnd11an1n32x5 FILLER_52_683 ();
 b15zdnd00an1n02x5 FILLER_52_715 ();
 b15zdnd00an1n01x5 FILLER_52_717 ();
 b15zdnd11an1n64x5 FILLER_52_726 ();
 b15zdnd11an1n64x5 FILLER_52_790 ();
 b15zdnd11an1n64x5 FILLER_52_854 ();
 b15zdnd11an1n64x5 FILLER_52_918 ();
 b15zdnd11an1n64x5 FILLER_52_982 ();
 b15zdnd11an1n64x5 FILLER_52_1046 ();
 b15zdnd11an1n32x5 FILLER_52_1110 ();
 b15zdnd11an1n04x5 FILLER_52_1142 ();
 b15zdnd00an1n02x5 FILLER_52_1146 ();
 b15zdnd00an1n01x5 FILLER_52_1148 ();
 b15zdnd11an1n08x5 FILLER_52_1163 ();
 b15zdnd11an1n04x5 FILLER_52_1175 ();
 b15zdnd11an1n08x5 FILLER_52_1189 ();
 b15zdnd11an1n04x5 FILLER_52_1197 ();
 b15zdnd11an1n04x5 FILLER_52_1225 ();
 b15zdnd11an1n64x5 FILLER_52_1232 ();
 b15zdnd11an1n08x5 FILLER_52_1296 ();
 b15zdnd00an1n01x5 FILLER_52_1304 ();
 b15zdnd11an1n32x5 FILLER_52_1313 ();
 b15zdnd00an1n01x5 FILLER_52_1345 ();
 b15zdnd11an1n32x5 FILLER_52_1373 ();
 b15zdnd11an1n04x5 FILLER_52_1405 ();
 b15zdnd00an1n01x5 FILLER_52_1409 ();
 b15zdnd11an1n16x5 FILLER_52_1427 ();
 b15zdnd00an1n01x5 FILLER_52_1443 ();
 b15zdnd11an1n08x5 FILLER_52_1447 ();
 b15zdnd11an1n04x5 FILLER_52_1455 ();
 b15zdnd00an1n02x5 FILLER_52_1459 ();
 b15zdnd11an1n64x5 FILLER_52_1468 ();
 b15zdnd11an1n64x5 FILLER_52_1532 ();
 b15zdnd11an1n32x5 FILLER_52_1596 ();
 b15zdnd11an1n16x5 FILLER_52_1628 ();
 b15zdnd11an1n08x5 FILLER_52_1644 ();
 b15zdnd11an1n16x5 FILLER_52_1694 ();
 b15zdnd11an1n08x5 FILLER_52_1710 ();
 b15zdnd00an1n02x5 FILLER_52_1718 ();
 b15zdnd00an1n01x5 FILLER_52_1720 ();
 b15zdnd11an1n64x5 FILLER_52_1763 ();
 b15zdnd00an1n02x5 FILLER_52_1827 ();
 b15zdnd11an1n32x5 FILLER_52_1837 ();
 b15zdnd11an1n16x5 FILLER_52_1869 ();
 b15zdnd11an1n04x5 FILLER_52_1885 ();
 b15zdnd11an1n64x5 FILLER_52_1929 ();
 b15zdnd11an1n64x5 FILLER_52_1993 ();
 b15zdnd11an1n64x5 FILLER_52_2057 ();
 b15zdnd11an1n32x5 FILLER_52_2121 ();
 b15zdnd00an1n01x5 FILLER_52_2153 ();
 b15zdnd11an1n64x5 FILLER_52_2162 ();
 b15zdnd11an1n32x5 FILLER_52_2226 ();
 b15zdnd11an1n16x5 FILLER_52_2258 ();
 b15zdnd00an1n02x5 FILLER_52_2274 ();
 b15zdnd11an1n64x5 FILLER_53_0 ();
 b15zdnd11an1n64x5 FILLER_53_64 ();
 b15zdnd11an1n64x5 FILLER_53_128 ();
 b15zdnd11an1n64x5 FILLER_53_192 ();
 b15zdnd11an1n64x5 FILLER_53_256 ();
 b15zdnd11an1n64x5 FILLER_53_320 ();
 b15zdnd11an1n04x5 FILLER_53_384 ();
 b15zdnd11an1n04x5 FILLER_53_394 ();
 b15zdnd11an1n32x5 FILLER_53_440 ();
 b15zdnd11an1n04x5 FILLER_53_472 ();
 b15zdnd00an1n02x5 FILLER_53_476 ();
 b15zdnd11an1n64x5 FILLER_53_530 ();
 b15zdnd11an1n64x5 FILLER_53_594 ();
 b15zdnd11an1n64x5 FILLER_53_658 ();
 b15zdnd11an1n64x5 FILLER_53_722 ();
 b15zdnd11an1n64x5 FILLER_53_786 ();
 b15zdnd11an1n64x5 FILLER_53_850 ();
 b15zdnd11an1n64x5 FILLER_53_914 ();
 b15zdnd11an1n16x5 FILLER_53_978 ();
 b15zdnd11an1n08x5 FILLER_53_994 ();
 b15zdnd11an1n04x5 FILLER_53_1002 ();
 b15zdnd11an1n64x5 FILLER_53_1018 ();
 b15zdnd11an1n64x5 FILLER_53_1082 ();
 b15zdnd11an1n04x5 FILLER_53_1146 ();
 b15zdnd00an1n01x5 FILLER_53_1150 ();
 b15zdnd11an1n04x5 FILLER_53_1158 ();
 b15zdnd11an1n08x5 FILLER_53_1172 ();
 b15zdnd00an1n02x5 FILLER_53_1180 ();
 b15zdnd11an1n04x5 FILLER_53_1193 ();
 b15zdnd00an1n02x5 FILLER_53_1197 ();
 b15zdnd11an1n08x5 FILLER_53_1205 ();
 b15zdnd11an1n04x5 FILLER_53_1213 ();
 b15zdnd00an1n02x5 FILLER_53_1217 ();
 b15zdnd00an1n01x5 FILLER_53_1219 ();
 b15zdnd11an1n64x5 FILLER_53_1226 ();
 b15zdnd11an1n08x5 FILLER_53_1290 ();
 b15zdnd11an1n04x5 FILLER_53_1298 ();
 b15zdnd00an1n01x5 FILLER_53_1302 ();
 b15zdnd11an1n64x5 FILLER_53_1345 ();
 b15zdnd11an1n64x5 FILLER_53_1409 ();
 b15zdnd11an1n64x5 FILLER_53_1473 ();
 b15zdnd11an1n64x5 FILLER_53_1537 ();
 b15zdnd11an1n32x5 FILLER_53_1601 ();
 b15zdnd11an1n16x5 FILLER_53_1633 ();
 b15zdnd11an1n08x5 FILLER_53_1649 ();
 b15zdnd00an1n02x5 FILLER_53_1657 ();
 b15zdnd00an1n01x5 FILLER_53_1659 ();
 b15zdnd11an1n64x5 FILLER_53_1702 ();
 b15zdnd11an1n32x5 FILLER_53_1766 ();
 b15zdnd11an1n08x5 FILLER_53_1798 ();
 b15zdnd00an1n02x5 FILLER_53_1806 ();
 b15zdnd00an1n01x5 FILLER_53_1808 ();
 b15zdnd11an1n64x5 FILLER_53_1836 ();
 b15zdnd11an1n64x5 FILLER_53_1900 ();
 b15zdnd11an1n64x5 FILLER_53_1964 ();
 b15zdnd11an1n64x5 FILLER_53_2028 ();
 b15zdnd11an1n64x5 FILLER_53_2092 ();
 b15zdnd11an1n64x5 FILLER_53_2156 ();
 b15zdnd11an1n64x5 FILLER_53_2220 ();
 b15zdnd11an1n64x5 FILLER_54_8 ();
 b15zdnd11an1n64x5 FILLER_54_72 ();
 b15zdnd11an1n64x5 FILLER_54_136 ();
 b15zdnd11an1n32x5 FILLER_54_200 ();
 b15zdnd00an1n02x5 FILLER_54_232 ();
 b15zdnd00an1n01x5 FILLER_54_234 ();
 b15zdnd11an1n64x5 FILLER_54_238 ();
 b15zdnd11an1n64x5 FILLER_54_302 ();
 b15zdnd11an1n04x5 FILLER_54_369 ();
 b15zdnd11an1n04x5 FILLER_54_383 ();
 b15zdnd11an1n64x5 FILLER_54_429 ();
 b15zdnd11an1n04x5 FILLER_54_493 ();
 b15zdnd11an1n04x5 FILLER_54_500 ();
 b15zdnd11an1n64x5 FILLER_54_507 ();
 b15zdnd11an1n64x5 FILLER_54_571 ();
 b15zdnd11an1n64x5 FILLER_54_635 ();
 b15zdnd11an1n16x5 FILLER_54_699 ();
 b15zdnd00an1n02x5 FILLER_54_715 ();
 b15zdnd00an1n01x5 FILLER_54_717 ();
 b15zdnd11an1n64x5 FILLER_54_726 ();
 b15zdnd11an1n04x5 FILLER_54_790 ();
 b15zdnd11an1n64x5 FILLER_54_798 ();
 b15zdnd11an1n64x5 FILLER_54_862 ();
 b15zdnd11an1n32x5 FILLER_54_926 ();
 b15zdnd11an1n08x5 FILLER_54_958 ();
 b15zdnd11an1n04x5 FILLER_54_966 ();
 b15zdnd00an1n01x5 FILLER_54_970 ();
 b15zdnd11an1n08x5 FILLER_54_976 ();
 b15zdnd11an1n04x5 FILLER_54_984 ();
 b15zdnd11an1n64x5 FILLER_54_997 ();
 b15zdnd11an1n64x5 FILLER_54_1061 ();
 b15zdnd11an1n64x5 FILLER_54_1125 ();
 b15zdnd11an1n64x5 FILLER_54_1189 ();
 b15zdnd11an1n32x5 FILLER_54_1253 ();
 b15zdnd11an1n08x5 FILLER_54_1285 ();
 b15zdnd00an1n01x5 FILLER_54_1293 ();
 b15zdnd11an1n16x5 FILLER_54_1336 ();
 b15zdnd11an1n04x5 FILLER_54_1355 ();
 b15zdnd11an1n64x5 FILLER_54_1362 ();
 b15zdnd11an1n64x5 FILLER_54_1426 ();
 b15zdnd11an1n64x5 FILLER_54_1490 ();
 b15zdnd11an1n64x5 FILLER_54_1554 ();
 b15zdnd11an1n32x5 FILLER_54_1618 ();
 b15zdnd11an1n16x5 FILLER_54_1650 ();
 b15zdnd11an1n08x5 FILLER_54_1666 ();
 b15zdnd11an1n04x5 FILLER_54_1674 ();
 b15zdnd11an1n16x5 FILLER_54_1687 ();
 b15zdnd11an1n04x5 FILLER_54_1703 ();
 b15zdnd00an1n02x5 FILLER_54_1707 ();
 b15zdnd11an1n64x5 FILLER_54_1751 ();
 b15zdnd11an1n64x5 FILLER_54_1815 ();
 b15zdnd11an1n64x5 FILLER_54_1879 ();
 b15zdnd11an1n64x5 FILLER_54_1943 ();
 b15zdnd11an1n64x5 FILLER_54_2007 ();
 b15zdnd11an1n64x5 FILLER_54_2071 ();
 b15zdnd11an1n16x5 FILLER_54_2135 ();
 b15zdnd00an1n02x5 FILLER_54_2151 ();
 b15zdnd00an1n01x5 FILLER_54_2153 ();
 b15zdnd11an1n64x5 FILLER_54_2162 ();
 b15zdnd11an1n32x5 FILLER_54_2226 ();
 b15zdnd11an1n16x5 FILLER_54_2258 ();
 b15zdnd00an1n02x5 FILLER_54_2274 ();
 b15zdnd11an1n64x5 FILLER_55_0 ();
 b15zdnd11an1n64x5 FILLER_55_64 ();
 b15zdnd11an1n64x5 FILLER_55_128 ();
 b15zdnd11an1n16x5 FILLER_55_192 ();
 b15zdnd11an1n64x5 FILLER_55_260 ();
 b15zdnd11an1n32x5 FILLER_55_324 ();
 b15zdnd00an1n02x5 FILLER_55_356 ();
 b15zdnd00an1n01x5 FILLER_55_358 ();
 b15zdnd11an1n04x5 FILLER_55_368 ();
 b15zdnd00an1n01x5 FILLER_55_372 ();
 b15zdnd11an1n08x5 FILLER_55_387 ();
 b15zdnd11an1n64x5 FILLER_55_437 ();
 b15zdnd11an1n64x5 FILLER_55_501 ();
 b15zdnd11an1n64x5 FILLER_55_565 ();
 b15zdnd11an1n64x5 FILLER_55_629 ();
 b15zdnd11an1n64x5 FILLER_55_693 ();
 b15zdnd00an1n02x5 FILLER_55_757 ();
 b15zdnd00an1n01x5 FILLER_55_759 ();
 b15zdnd11an1n04x5 FILLER_55_764 ();
 b15zdnd00an1n01x5 FILLER_55_768 ();
 b15zdnd11an1n64x5 FILLER_55_773 ();
 b15zdnd11an1n64x5 FILLER_55_837 ();
 b15zdnd11an1n64x5 FILLER_55_901 ();
 b15zdnd11an1n64x5 FILLER_55_965 ();
 b15zdnd11an1n64x5 FILLER_55_1029 ();
 b15zdnd11an1n16x5 FILLER_55_1093 ();
 b15zdnd11an1n08x5 FILLER_55_1109 ();
 b15zdnd11an1n04x5 FILLER_55_1117 ();
 b15zdnd11an1n64x5 FILLER_55_1166 ();
 b15zdnd11an1n64x5 FILLER_55_1230 ();
 b15zdnd11an1n32x5 FILLER_55_1294 ();
 b15zdnd11an1n08x5 FILLER_55_1326 ();
 b15zdnd11an1n64x5 FILLER_55_1386 ();
 b15zdnd11an1n64x5 FILLER_55_1450 ();
 b15zdnd11an1n64x5 FILLER_55_1514 ();
 b15zdnd11an1n64x5 FILLER_55_1578 ();
 b15zdnd11an1n16x5 FILLER_55_1642 ();
 b15zdnd11an1n08x5 FILLER_55_1658 ();
 b15zdnd00an1n02x5 FILLER_55_1666 ();
 b15zdnd00an1n01x5 FILLER_55_1668 ();
 b15zdnd11an1n04x5 FILLER_55_1675 ();
 b15zdnd11an1n04x5 FILLER_55_1721 ();
 b15zdnd11an1n04x5 FILLER_55_1728 ();
 b15zdnd11an1n64x5 FILLER_55_1735 ();
 b15zdnd11an1n64x5 FILLER_55_1799 ();
 b15zdnd11an1n64x5 FILLER_55_1863 ();
 b15zdnd11an1n64x5 FILLER_55_1927 ();
 b15zdnd11an1n64x5 FILLER_55_1991 ();
 b15zdnd11an1n64x5 FILLER_55_2055 ();
 b15zdnd11an1n64x5 FILLER_55_2119 ();
 b15zdnd11an1n64x5 FILLER_55_2183 ();
 b15zdnd11an1n32x5 FILLER_55_2247 ();
 b15zdnd11an1n04x5 FILLER_55_2279 ();
 b15zdnd00an1n01x5 FILLER_55_2283 ();
 b15zdnd11an1n64x5 FILLER_56_8 ();
 b15zdnd11an1n64x5 FILLER_56_72 ();
 b15zdnd11an1n64x5 FILLER_56_136 ();
 b15zdnd11an1n16x5 FILLER_56_200 ();
 b15zdnd11an1n08x5 FILLER_56_216 ();
 b15zdnd00an1n02x5 FILLER_56_224 ();
 b15zdnd00an1n01x5 FILLER_56_226 ();
 b15zdnd11an1n04x5 FILLER_56_230 ();
 b15zdnd11an1n64x5 FILLER_56_237 ();
 b15zdnd11an1n64x5 FILLER_56_301 ();
 b15zdnd00an1n01x5 FILLER_56_365 ();
 b15zdnd11an1n04x5 FILLER_56_369 ();
 b15zdnd00an1n02x5 FILLER_56_373 ();
 b15zdnd00an1n01x5 FILLER_56_375 ();
 b15zdnd11an1n08x5 FILLER_56_381 ();
 b15zdnd00an1n02x5 FILLER_56_389 ();
 b15zdnd11an1n64x5 FILLER_56_398 ();
 b15zdnd11an1n16x5 FILLER_56_462 ();
 b15zdnd00an1n02x5 FILLER_56_478 ();
 b15zdnd11an1n64x5 FILLER_56_522 ();
 b15zdnd11an1n64x5 FILLER_56_586 ();
 b15zdnd11an1n64x5 FILLER_56_650 ();
 b15zdnd11an1n04x5 FILLER_56_714 ();
 b15zdnd11an1n32x5 FILLER_56_726 ();
 b15zdnd11an1n08x5 FILLER_56_758 ();
 b15zdnd00an1n02x5 FILLER_56_766 ();
 b15zdnd11an1n64x5 FILLER_56_772 ();
 b15zdnd11an1n64x5 FILLER_56_836 ();
 b15zdnd11an1n64x5 FILLER_56_900 ();
 b15zdnd11an1n64x5 FILLER_56_964 ();
 b15zdnd11an1n64x5 FILLER_56_1028 ();
 b15zdnd11an1n64x5 FILLER_56_1092 ();
 b15zdnd11an1n64x5 FILLER_56_1156 ();
 b15zdnd11an1n64x5 FILLER_56_1220 ();
 b15zdnd11an1n64x5 FILLER_56_1284 ();
 b15zdnd11an1n08x5 FILLER_56_1348 ();
 b15zdnd11an1n04x5 FILLER_56_1356 ();
 b15zdnd11an1n64x5 FILLER_56_1363 ();
 b15zdnd11an1n64x5 FILLER_56_1427 ();
 b15zdnd11an1n64x5 FILLER_56_1491 ();
 b15zdnd11an1n64x5 FILLER_56_1555 ();
 b15zdnd11an1n32x5 FILLER_56_1619 ();
 b15zdnd11an1n08x5 FILLER_56_1651 ();
 b15zdnd00an1n02x5 FILLER_56_1659 ();
 b15zdnd00an1n01x5 FILLER_56_1661 ();
 b15zdnd11an1n04x5 FILLER_56_1672 ();
 b15zdnd11an1n16x5 FILLER_56_1686 ();
 b15zdnd11an1n04x5 FILLER_56_1702 ();
 b15zdnd11an1n64x5 FILLER_56_1758 ();
 b15zdnd11an1n64x5 FILLER_56_1822 ();
 b15zdnd11an1n64x5 FILLER_56_1886 ();
 b15zdnd11an1n64x5 FILLER_56_1950 ();
 b15zdnd11an1n64x5 FILLER_56_2014 ();
 b15zdnd11an1n64x5 FILLER_56_2078 ();
 b15zdnd11an1n08x5 FILLER_56_2142 ();
 b15zdnd11an1n04x5 FILLER_56_2150 ();
 b15zdnd11an1n64x5 FILLER_56_2162 ();
 b15zdnd11an1n32x5 FILLER_56_2226 ();
 b15zdnd11an1n16x5 FILLER_56_2258 ();
 b15zdnd00an1n02x5 FILLER_56_2274 ();
 b15zdnd11an1n64x5 FILLER_57_0 ();
 b15zdnd11an1n64x5 FILLER_57_64 ();
 b15zdnd11an1n64x5 FILLER_57_128 ();
 b15zdnd11an1n64x5 FILLER_57_192 ();
 b15zdnd11an1n64x5 FILLER_57_256 ();
 b15zdnd11an1n32x5 FILLER_57_320 ();
 b15zdnd11an1n16x5 FILLER_57_352 ();
 b15zdnd11an1n04x5 FILLER_57_368 ();
 b15zdnd11an1n04x5 FILLER_57_382 ();
 b15zdnd11an1n64x5 FILLER_57_390 ();
 b15zdnd11an1n04x5 FILLER_57_454 ();
 b15zdnd00an1n02x5 FILLER_57_458 ();
 b15zdnd00an1n01x5 FILLER_57_460 ();
 b15zdnd11an1n64x5 FILLER_57_486 ();
 b15zdnd11an1n64x5 FILLER_57_550 ();
 b15zdnd11an1n64x5 FILLER_57_614 ();
 b15zdnd11an1n64x5 FILLER_57_678 ();
 b15zdnd11an1n64x5 FILLER_57_742 ();
 b15zdnd11an1n64x5 FILLER_57_806 ();
 b15zdnd11an1n64x5 FILLER_57_870 ();
 b15zdnd11an1n64x5 FILLER_57_934 ();
 b15zdnd11an1n64x5 FILLER_57_998 ();
 b15zdnd11an1n64x5 FILLER_57_1062 ();
 b15zdnd11an1n64x5 FILLER_57_1126 ();
 b15zdnd11an1n64x5 FILLER_57_1190 ();
 b15zdnd11an1n64x5 FILLER_57_1254 ();
 b15zdnd11an1n64x5 FILLER_57_1318 ();
 b15zdnd11an1n64x5 FILLER_57_1382 ();
 b15zdnd11an1n64x5 FILLER_57_1446 ();
 b15zdnd11an1n64x5 FILLER_57_1510 ();
 b15zdnd11an1n64x5 FILLER_57_1574 ();
 b15zdnd11an1n32x5 FILLER_57_1638 ();
 b15zdnd00an1n02x5 FILLER_57_1670 ();
 b15zdnd00an1n01x5 FILLER_57_1672 ();
 b15zdnd11an1n08x5 FILLER_57_1682 ();
 b15zdnd11an1n04x5 FILLER_57_1690 ();
 b15zdnd00an1n02x5 FILLER_57_1694 ();
 b15zdnd11an1n04x5 FILLER_57_1738 ();
 b15zdnd11an1n64x5 FILLER_57_1745 ();
 b15zdnd11an1n64x5 FILLER_57_1809 ();
 b15zdnd11an1n64x5 FILLER_57_1873 ();
 b15zdnd11an1n64x5 FILLER_57_1937 ();
 b15zdnd11an1n64x5 FILLER_57_2001 ();
 b15zdnd11an1n64x5 FILLER_57_2065 ();
 b15zdnd11an1n64x5 FILLER_57_2129 ();
 b15zdnd11an1n64x5 FILLER_57_2193 ();
 b15zdnd11an1n16x5 FILLER_57_2257 ();
 b15zdnd11an1n08x5 FILLER_57_2273 ();
 b15zdnd00an1n02x5 FILLER_57_2281 ();
 b15zdnd00an1n01x5 FILLER_57_2283 ();
 b15zdnd11an1n64x5 FILLER_58_8 ();
 b15zdnd11an1n64x5 FILLER_58_72 ();
 b15zdnd11an1n64x5 FILLER_58_136 ();
 b15zdnd11an1n64x5 FILLER_58_200 ();
 b15zdnd11an1n64x5 FILLER_58_264 ();
 b15zdnd11an1n32x5 FILLER_58_328 ();
 b15zdnd11an1n08x5 FILLER_58_360 ();
 b15zdnd00an1n02x5 FILLER_58_368 ();
 b15zdnd00an1n01x5 FILLER_58_370 ();
 b15zdnd11an1n64x5 FILLER_58_381 ();
 b15zdnd11an1n64x5 FILLER_58_445 ();
 b15zdnd11an1n64x5 FILLER_58_509 ();
 b15zdnd11an1n64x5 FILLER_58_573 ();
 b15zdnd11an1n64x5 FILLER_58_637 ();
 b15zdnd11an1n16x5 FILLER_58_701 ();
 b15zdnd00an1n01x5 FILLER_58_717 ();
 b15zdnd11an1n64x5 FILLER_58_726 ();
 b15zdnd11an1n16x5 FILLER_58_790 ();
 b15zdnd11an1n08x5 FILLER_58_806 ();
 b15zdnd11an1n04x5 FILLER_58_814 ();
 b15zdnd11an1n64x5 FILLER_58_860 ();
 b15zdnd11an1n64x5 FILLER_58_924 ();
 b15zdnd11an1n64x5 FILLER_58_988 ();
 b15zdnd11an1n64x5 FILLER_58_1052 ();
 b15zdnd11an1n64x5 FILLER_58_1116 ();
 b15zdnd11an1n64x5 FILLER_58_1180 ();
 b15zdnd11an1n64x5 FILLER_58_1244 ();
 b15zdnd11an1n64x5 FILLER_58_1308 ();
 b15zdnd11an1n64x5 FILLER_58_1372 ();
 b15zdnd11an1n64x5 FILLER_58_1436 ();
 b15zdnd11an1n64x5 FILLER_58_1500 ();
 b15zdnd11an1n64x5 FILLER_58_1564 ();
 b15zdnd11an1n16x5 FILLER_58_1628 ();
 b15zdnd11an1n08x5 FILLER_58_1644 ();
 b15zdnd11an1n04x5 FILLER_58_1652 ();
 b15zdnd00an1n02x5 FILLER_58_1656 ();
 b15zdnd11an1n04x5 FILLER_58_1668 ();
 b15zdnd11an1n32x5 FILLER_58_1682 ();
 b15zdnd11an1n04x5 FILLER_58_1714 ();
 b15zdnd00an1n02x5 FILLER_58_1718 ();
 b15zdnd00an1n01x5 FILLER_58_1720 ();
 b15zdnd11an1n64x5 FILLER_58_1763 ();
 b15zdnd11an1n64x5 FILLER_58_1827 ();
 b15zdnd11an1n64x5 FILLER_58_1891 ();
 b15zdnd11an1n64x5 FILLER_58_1955 ();
 b15zdnd11an1n64x5 FILLER_58_2019 ();
 b15zdnd11an1n64x5 FILLER_58_2083 ();
 b15zdnd11an1n04x5 FILLER_58_2147 ();
 b15zdnd00an1n02x5 FILLER_58_2151 ();
 b15zdnd00an1n01x5 FILLER_58_2153 ();
 b15zdnd11an1n64x5 FILLER_58_2162 ();
 b15zdnd11an1n32x5 FILLER_58_2226 ();
 b15zdnd11an1n16x5 FILLER_58_2258 ();
 b15zdnd00an1n02x5 FILLER_58_2274 ();
 b15zdnd11an1n64x5 FILLER_59_0 ();
 b15zdnd11an1n64x5 FILLER_59_64 ();
 b15zdnd11an1n64x5 FILLER_59_128 ();
 b15zdnd11an1n64x5 FILLER_59_192 ();
 b15zdnd11an1n64x5 FILLER_59_256 ();
 b15zdnd11an1n64x5 FILLER_59_320 ();
 b15zdnd11an1n64x5 FILLER_59_384 ();
 b15zdnd11an1n64x5 FILLER_59_448 ();
 b15zdnd11an1n64x5 FILLER_59_512 ();
 b15zdnd11an1n64x5 FILLER_59_576 ();
 b15zdnd11an1n64x5 FILLER_59_640 ();
 b15zdnd11an1n64x5 FILLER_59_704 ();
 b15zdnd11an1n64x5 FILLER_59_768 ();
 b15zdnd11an1n64x5 FILLER_59_832 ();
 b15zdnd11an1n64x5 FILLER_59_896 ();
 b15zdnd11an1n64x5 FILLER_59_960 ();
 b15zdnd11an1n64x5 FILLER_59_1024 ();
 b15zdnd11an1n32x5 FILLER_59_1088 ();
 b15zdnd11an1n08x5 FILLER_59_1120 ();
 b15zdnd11an1n04x5 FILLER_59_1128 ();
 b15zdnd11an1n64x5 FILLER_59_1152 ();
 b15zdnd11an1n64x5 FILLER_59_1216 ();
 b15zdnd11an1n32x5 FILLER_59_1280 ();
 b15zdnd11an1n16x5 FILLER_59_1312 ();
 b15zdnd11an1n08x5 FILLER_59_1328 ();
 b15zdnd11an1n04x5 FILLER_59_1336 ();
 b15zdnd00an1n02x5 FILLER_59_1340 ();
 b15zdnd11an1n64x5 FILLER_59_1384 ();
 b15zdnd11an1n16x5 FILLER_59_1448 ();
 b15zdnd11an1n04x5 FILLER_59_1464 ();
 b15zdnd00an1n02x5 FILLER_59_1468 ();
 b15zdnd00an1n01x5 FILLER_59_1470 ();
 b15zdnd11an1n64x5 FILLER_59_1491 ();
 b15zdnd11an1n64x5 FILLER_59_1555 ();
 b15zdnd11an1n32x5 FILLER_59_1619 ();
 b15zdnd11an1n04x5 FILLER_59_1651 ();
 b15zdnd00an1n02x5 FILLER_59_1655 ();
 b15zdnd00an1n01x5 FILLER_59_1657 ();
 b15zdnd11an1n04x5 FILLER_59_1663 ();
 b15zdnd11an1n64x5 FILLER_59_1670 ();
 b15zdnd11an1n64x5 FILLER_59_1734 ();
 b15zdnd11an1n64x5 FILLER_59_1798 ();
 b15zdnd11an1n64x5 FILLER_59_1862 ();
 b15zdnd11an1n64x5 FILLER_59_1926 ();
 b15zdnd11an1n64x5 FILLER_59_1990 ();
 b15zdnd11an1n64x5 FILLER_59_2054 ();
 b15zdnd11an1n64x5 FILLER_59_2118 ();
 b15zdnd11an1n64x5 FILLER_59_2182 ();
 b15zdnd11an1n32x5 FILLER_59_2246 ();
 b15zdnd11an1n04x5 FILLER_59_2278 ();
 b15zdnd00an1n02x5 FILLER_59_2282 ();
 b15zdnd11an1n64x5 FILLER_60_8 ();
 b15zdnd11an1n64x5 FILLER_60_72 ();
 b15zdnd11an1n64x5 FILLER_60_136 ();
 b15zdnd11an1n64x5 FILLER_60_200 ();
 b15zdnd11an1n64x5 FILLER_60_264 ();
 b15zdnd11an1n32x5 FILLER_60_328 ();
 b15zdnd11an1n16x5 FILLER_60_360 ();
 b15zdnd11an1n04x5 FILLER_60_376 ();
 b15zdnd00an1n01x5 FILLER_60_380 ();
 b15zdnd11an1n64x5 FILLER_60_388 ();
 b15zdnd11an1n64x5 FILLER_60_452 ();
 b15zdnd11an1n64x5 FILLER_60_516 ();
 b15zdnd11an1n64x5 FILLER_60_580 ();
 b15zdnd11an1n64x5 FILLER_60_644 ();
 b15zdnd11an1n08x5 FILLER_60_708 ();
 b15zdnd00an1n02x5 FILLER_60_716 ();
 b15zdnd11an1n64x5 FILLER_60_726 ();
 b15zdnd11an1n64x5 FILLER_60_790 ();
 b15zdnd11an1n64x5 FILLER_60_854 ();
 b15zdnd11an1n64x5 FILLER_60_918 ();
 b15zdnd11an1n64x5 FILLER_60_982 ();
 b15zdnd11an1n64x5 FILLER_60_1046 ();
 b15zdnd11an1n64x5 FILLER_60_1110 ();
 b15zdnd11an1n64x5 FILLER_60_1174 ();
 b15zdnd11an1n64x5 FILLER_60_1238 ();
 b15zdnd11an1n64x5 FILLER_60_1302 ();
 b15zdnd11an1n64x5 FILLER_60_1366 ();
 b15zdnd11an1n64x5 FILLER_60_1430 ();
 b15zdnd11an1n64x5 FILLER_60_1494 ();
 b15zdnd11an1n64x5 FILLER_60_1558 ();
 b15zdnd11an1n64x5 FILLER_60_1622 ();
 b15zdnd11an1n64x5 FILLER_60_1686 ();
 b15zdnd11an1n64x5 FILLER_60_1750 ();
 b15zdnd11an1n64x5 FILLER_60_1814 ();
 b15zdnd11an1n32x5 FILLER_60_1878 ();
 b15zdnd11an1n04x5 FILLER_60_1910 ();
 b15zdnd11an1n64x5 FILLER_60_1956 ();
 b15zdnd11an1n64x5 FILLER_60_2020 ();
 b15zdnd11an1n64x5 FILLER_60_2084 ();
 b15zdnd11an1n04x5 FILLER_60_2148 ();
 b15zdnd00an1n02x5 FILLER_60_2152 ();
 b15zdnd11an1n64x5 FILLER_60_2162 ();
 b15zdnd11an1n32x5 FILLER_60_2226 ();
 b15zdnd11an1n16x5 FILLER_60_2258 ();
 b15zdnd00an1n02x5 FILLER_60_2274 ();
 b15zdnd11an1n64x5 FILLER_61_0 ();
 b15zdnd11an1n64x5 FILLER_61_64 ();
 b15zdnd11an1n64x5 FILLER_61_128 ();
 b15zdnd11an1n64x5 FILLER_61_192 ();
 b15zdnd11an1n64x5 FILLER_61_256 ();
 b15zdnd11an1n64x5 FILLER_61_320 ();
 b15zdnd00an1n02x5 FILLER_61_384 ();
 b15zdnd11an1n64x5 FILLER_61_428 ();
 b15zdnd11an1n64x5 FILLER_61_492 ();
 b15zdnd11an1n64x5 FILLER_61_556 ();
 b15zdnd11an1n64x5 FILLER_61_620 ();
 b15zdnd11an1n64x5 FILLER_61_684 ();
 b15zdnd11an1n64x5 FILLER_61_748 ();
 b15zdnd11an1n64x5 FILLER_61_812 ();
 b15zdnd11an1n64x5 FILLER_61_876 ();
 b15zdnd11an1n64x5 FILLER_61_940 ();
 b15zdnd11an1n64x5 FILLER_61_1004 ();
 b15zdnd11an1n64x5 FILLER_61_1068 ();
 b15zdnd11an1n64x5 FILLER_61_1132 ();
 b15zdnd11an1n64x5 FILLER_61_1196 ();
 b15zdnd11an1n08x5 FILLER_61_1260 ();
 b15zdnd00an1n01x5 FILLER_61_1268 ();
 b15zdnd11an1n64x5 FILLER_61_1286 ();
 b15zdnd11an1n64x5 FILLER_61_1350 ();
 b15zdnd11an1n64x5 FILLER_61_1414 ();
 b15zdnd11an1n64x5 FILLER_61_1478 ();
 b15zdnd11an1n64x5 FILLER_61_1542 ();
 b15zdnd11an1n64x5 FILLER_61_1606 ();
 b15zdnd11an1n64x5 FILLER_61_1670 ();
 b15zdnd11an1n64x5 FILLER_61_1734 ();
 b15zdnd11an1n64x5 FILLER_61_1798 ();
 b15zdnd11an1n32x5 FILLER_61_1862 ();
 b15zdnd00an1n02x5 FILLER_61_1894 ();
 b15zdnd00an1n01x5 FILLER_61_1896 ();
 b15zdnd11an1n64x5 FILLER_61_1939 ();
 b15zdnd11an1n64x5 FILLER_61_2003 ();
 b15zdnd11an1n64x5 FILLER_61_2067 ();
 b15zdnd11an1n64x5 FILLER_61_2131 ();
 b15zdnd11an1n64x5 FILLER_61_2195 ();
 b15zdnd11an1n16x5 FILLER_61_2259 ();
 b15zdnd11an1n08x5 FILLER_61_2275 ();
 b15zdnd00an1n01x5 FILLER_61_2283 ();
 b15zdnd11an1n64x5 FILLER_62_8 ();
 b15zdnd11an1n64x5 FILLER_62_72 ();
 b15zdnd11an1n64x5 FILLER_62_136 ();
 b15zdnd11an1n64x5 FILLER_62_200 ();
 b15zdnd11an1n64x5 FILLER_62_264 ();
 b15zdnd11an1n64x5 FILLER_62_328 ();
 b15zdnd11an1n64x5 FILLER_62_392 ();
 b15zdnd11an1n64x5 FILLER_62_456 ();
 b15zdnd11an1n64x5 FILLER_62_520 ();
 b15zdnd11an1n64x5 FILLER_62_584 ();
 b15zdnd11an1n64x5 FILLER_62_648 ();
 b15zdnd11an1n04x5 FILLER_62_712 ();
 b15zdnd00an1n02x5 FILLER_62_716 ();
 b15zdnd11an1n64x5 FILLER_62_726 ();
 b15zdnd11an1n64x5 FILLER_62_790 ();
 b15zdnd11an1n64x5 FILLER_62_854 ();
 b15zdnd11an1n64x5 FILLER_62_918 ();
 b15zdnd11an1n64x5 FILLER_62_982 ();
 b15zdnd11an1n64x5 FILLER_62_1046 ();
 b15zdnd11an1n64x5 FILLER_62_1110 ();
 b15zdnd11an1n64x5 FILLER_62_1174 ();
 b15zdnd11an1n64x5 FILLER_62_1238 ();
 b15zdnd11an1n64x5 FILLER_62_1302 ();
 b15zdnd11an1n64x5 FILLER_62_1366 ();
 b15zdnd11an1n64x5 FILLER_62_1430 ();
 b15zdnd11an1n08x5 FILLER_62_1494 ();
 b15zdnd11an1n04x5 FILLER_62_1502 ();
 b15zdnd11an1n04x5 FILLER_62_1537 ();
 b15zdnd11an1n04x5 FILLER_62_1593 ();
 b15zdnd00an1n02x5 FILLER_62_1597 ();
 b15zdnd00an1n01x5 FILLER_62_1599 ();
 b15zdnd11an1n08x5 FILLER_62_1605 ();
 b15zdnd00an1n02x5 FILLER_62_1613 ();
 b15zdnd11an1n64x5 FILLER_62_1626 ();
 b15zdnd11an1n64x5 FILLER_62_1690 ();
 b15zdnd11an1n64x5 FILLER_62_1754 ();
 b15zdnd11an1n64x5 FILLER_62_1818 ();
 b15zdnd11an1n64x5 FILLER_62_1882 ();
 b15zdnd11an1n64x5 FILLER_62_1946 ();
 b15zdnd11an1n64x5 FILLER_62_2010 ();
 b15zdnd11an1n64x5 FILLER_62_2074 ();
 b15zdnd11an1n16x5 FILLER_62_2138 ();
 b15zdnd11an1n64x5 FILLER_62_2162 ();
 b15zdnd11an1n32x5 FILLER_62_2226 ();
 b15zdnd11an1n16x5 FILLER_62_2258 ();
 b15zdnd00an1n02x5 FILLER_62_2274 ();
 b15zdnd11an1n64x5 FILLER_63_0 ();
 b15zdnd11an1n64x5 FILLER_63_64 ();
 b15zdnd11an1n64x5 FILLER_63_128 ();
 b15zdnd11an1n64x5 FILLER_63_192 ();
 b15zdnd11an1n04x5 FILLER_63_256 ();
 b15zdnd11an1n64x5 FILLER_63_302 ();
 b15zdnd11an1n64x5 FILLER_63_366 ();
 b15zdnd11an1n64x5 FILLER_63_430 ();
 b15zdnd11an1n64x5 FILLER_63_494 ();
 b15zdnd11an1n64x5 FILLER_63_558 ();
 b15zdnd11an1n64x5 FILLER_63_622 ();
 b15zdnd11an1n64x5 FILLER_63_686 ();
 b15zdnd11an1n64x5 FILLER_63_750 ();
 b15zdnd11an1n64x5 FILLER_63_814 ();
 b15zdnd11an1n64x5 FILLER_63_878 ();
 b15zdnd11an1n64x5 FILLER_63_942 ();
 b15zdnd11an1n64x5 FILLER_63_1006 ();
 b15zdnd11an1n64x5 FILLER_63_1070 ();
 b15zdnd11an1n64x5 FILLER_63_1134 ();
 b15zdnd11an1n32x5 FILLER_63_1198 ();
 b15zdnd11an1n08x5 FILLER_63_1230 ();
 b15zdnd00an1n01x5 FILLER_63_1238 ();
 b15zdnd11an1n08x5 FILLER_63_1242 ();
 b15zdnd00an1n01x5 FILLER_63_1250 ();
 b15zdnd11an1n64x5 FILLER_63_1254 ();
 b15zdnd11an1n64x5 FILLER_63_1318 ();
 b15zdnd11an1n64x5 FILLER_63_1382 ();
 b15zdnd11an1n64x5 FILLER_63_1446 ();
 b15zdnd11an1n32x5 FILLER_63_1510 ();
 b15zdnd11an1n16x5 FILLER_63_1542 ();
 b15zdnd00an1n02x5 FILLER_63_1558 ();
 b15zdnd11an1n04x5 FILLER_63_1563 ();
 b15zdnd11an1n32x5 FILLER_63_1570 ();
 b15zdnd11an1n64x5 FILLER_63_1644 ();
 b15zdnd11an1n64x5 FILLER_63_1708 ();
 b15zdnd11an1n64x5 FILLER_63_1772 ();
 b15zdnd11an1n64x5 FILLER_63_1836 ();
 b15zdnd11an1n64x5 FILLER_63_1900 ();
 b15zdnd11an1n64x5 FILLER_63_1964 ();
 b15zdnd11an1n64x5 FILLER_63_2028 ();
 b15zdnd11an1n64x5 FILLER_63_2092 ();
 b15zdnd11an1n64x5 FILLER_63_2156 ();
 b15zdnd11an1n64x5 FILLER_63_2220 ();
 b15zdnd11an1n64x5 FILLER_64_8 ();
 b15zdnd11an1n64x5 FILLER_64_72 ();
 b15zdnd11an1n64x5 FILLER_64_136 ();
 b15zdnd11an1n64x5 FILLER_64_200 ();
 b15zdnd11an1n64x5 FILLER_64_264 ();
 b15zdnd11an1n16x5 FILLER_64_328 ();
 b15zdnd11an1n04x5 FILLER_64_344 ();
 b15zdnd00an1n01x5 FILLER_64_348 ();
 b15zdnd11an1n64x5 FILLER_64_401 ();
 b15zdnd11an1n16x5 FILLER_64_465 ();
 b15zdnd11an1n04x5 FILLER_64_481 ();
 b15zdnd00an1n02x5 FILLER_64_485 ();
 b15zdnd11an1n04x5 FILLER_64_491 ();
 b15zdnd11an1n64x5 FILLER_64_537 ();
 b15zdnd11an1n64x5 FILLER_64_601 ();
 b15zdnd11an1n32x5 FILLER_64_665 ();
 b15zdnd11an1n16x5 FILLER_64_697 ();
 b15zdnd11an1n04x5 FILLER_64_713 ();
 b15zdnd00an1n01x5 FILLER_64_717 ();
 b15zdnd11an1n64x5 FILLER_64_726 ();
 b15zdnd11an1n64x5 FILLER_64_790 ();
 b15zdnd11an1n64x5 FILLER_64_854 ();
 b15zdnd11an1n64x5 FILLER_64_918 ();
 b15zdnd11an1n64x5 FILLER_64_982 ();
 b15zdnd11an1n64x5 FILLER_64_1046 ();
 b15zdnd11an1n64x5 FILLER_64_1110 ();
 b15zdnd11an1n32x5 FILLER_64_1174 ();
 b15zdnd11an1n08x5 FILLER_64_1206 ();
 b15zdnd11an1n04x5 FILLER_64_1214 ();
 b15zdnd00an1n01x5 FILLER_64_1218 ();
 b15zdnd11an1n64x5 FILLER_64_1271 ();
 b15zdnd11an1n64x5 FILLER_64_1335 ();
 b15zdnd11an1n64x5 FILLER_64_1399 ();
 b15zdnd11an1n04x5 FILLER_64_1463 ();
 b15zdnd00an1n02x5 FILLER_64_1467 ();
 b15zdnd00an1n01x5 FILLER_64_1469 ();
 b15zdnd11an1n64x5 FILLER_64_1477 ();
 b15zdnd11an1n16x5 FILLER_64_1541 ();
 b15zdnd11an1n08x5 FILLER_64_1557 ();
 b15zdnd00an1n02x5 FILLER_64_1565 ();
 b15zdnd11an1n16x5 FILLER_64_1570 ();
 b15zdnd11an1n64x5 FILLER_64_1625 ();
 b15zdnd11an1n64x5 FILLER_64_1689 ();
 b15zdnd11an1n64x5 FILLER_64_1753 ();
 b15zdnd11an1n64x5 FILLER_64_1817 ();
 b15zdnd11an1n64x5 FILLER_64_1881 ();
 b15zdnd11an1n64x5 FILLER_64_1945 ();
 b15zdnd11an1n64x5 FILLER_64_2009 ();
 b15zdnd11an1n64x5 FILLER_64_2073 ();
 b15zdnd11an1n16x5 FILLER_64_2137 ();
 b15zdnd00an1n01x5 FILLER_64_2153 ();
 b15zdnd11an1n64x5 FILLER_64_2162 ();
 b15zdnd11an1n32x5 FILLER_64_2226 ();
 b15zdnd11an1n16x5 FILLER_64_2258 ();
 b15zdnd00an1n02x5 FILLER_64_2274 ();
 b15zdnd11an1n64x5 FILLER_65_0 ();
 b15zdnd11an1n64x5 FILLER_65_64 ();
 b15zdnd11an1n64x5 FILLER_65_128 ();
 b15zdnd11an1n64x5 FILLER_65_192 ();
 b15zdnd11an1n64x5 FILLER_65_256 ();
 b15zdnd11an1n32x5 FILLER_65_320 ();
 b15zdnd11an1n08x5 FILLER_65_352 ();
 b15zdnd00an1n02x5 FILLER_65_360 ();
 b15zdnd11an1n08x5 FILLER_65_365 ();
 b15zdnd00an1n01x5 FILLER_65_373 ();
 b15zdnd11an1n64x5 FILLER_65_377 ();
 b15zdnd11an1n64x5 FILLER_65_441 ();
 b15zdnd11an1n64x5 FILLER_65_505 ();
 b15zdnd11an1n64x5 FILLER_65_569 ();
 b15zdnd11an1n64x5 FILLER_65_633 ();
 b15zdnd11an1n64x5 FILLER_65_697 ();
 b15zdnd11an1n64x5 FILLER_65_761 ();
 b15zdnd11an1n64x5 FILLER_65_825 ();
 b15zdnd11an1n64x5 FILLER_65_889 ();
 b15zdnd11an1n64x5 FILLER_65_953 ();
 b15zdnd11an1n64x5 FILLER_65_1017 ();
 b15zdnd11an1n64x5 FILLER_65_1081 ();
 b15zdnd11an1n64x5 FILLER_65_1145 ();
 b15zdnd11an1n64x5 FILLER_65_1209 ();
 b15zdnd11an1n64x5 FILLER_65_1273 ();
 b15zdnd11an1n64x5 FILLER_65_1337 ();
 b15zdnd11an1n64x5 FILLER_65_1401 ();
 b15zdnd11an1n64x5 FILLER_65_1465 ();
 b15zdnd11an1n64x5 FILLER_65_1529 ();
 b15zdnd11an1n08x5 FILLER_65_1593 ();
 b15zdnd11an1n04x5 FILLER_65_1601 ();
 b15zdnd11an1n64x5 FILLER_65_1620 ();
 b15zdnd11an1n64x5 FILLER_65_1684 ();
 b15zdnd11an1n64x5 FILLER_65_1748 ();
 b15zdnd11an1n64x5 FILLER_65_1812 ();
 b15zdnd11an1n64x5 FILLER_65_1876 ();
 b15zdnd11an1n64x5 FILLER_65_1940 ();
 b15zdnd11an1n64x5 FILLER_65_2004 ();
 b15zdnd11an1n64x5 FILLER_65_2068 ();
 b15zdnd11an1n64x5 FILLER_65_2132 ();
 b15zdnd11an1n64x5 FILLER_65_2196 ();
 b15zdnd11an1n16x5 FILLER_65_2260 ();
 b15zdnd11an1n08x5 FILLER_65_2276 ();
 b15zdnd11an1n64x5 FILLER_66_8 ();
 b15zdnd11an1n64x5 FILLER_66_72 ();
 b15zdnd11an1n64x5 FILLER_66_136 ();
 b15zdnd11an1n64x5 FILLER_66_200 ();
 b15zdnd11an1n64x5 FILLER_66_264 ();
 b15zdnd11an1n32x5 FILLER_66_328 ();
 b15zdnd11an1n08x5 FILLER_66_360 ();
 b15zdnd11an1n04x5 FILLER_66_368 ();
 b15zdnd11an1n64x5 FILLER_66_375 ();
 b15zdnd11an1n64x5 FILLER_66_439 ();
 b15zdnd00an1n01x5 FILLER_66_503 ();
 b15zdnd11an1n64x5 FILLER_66_507 ();
 b15zdnd11an1n64x5 FILLER_66_571 ();
 b15zdnd11an1n64x5 FILLER_66_635 ();
 b15zdnd11an1n16x5 FILLER_66_699 ();
 b15zdnd00an1n02x5 FILLER_66_715 ();
 b15zdnd00an1n01x5 FILLER_66_717 ();
 b15zdnd11an1n64x5 FILLER_66_726 ();
 b15zdnd11an1n64x5 FILLER_66_790 ();
 b15zdnd11an1n64x5 FILLER_66_854 ();
 b15zdnd11an1n64x5 FILLER_66_918 ();
 b15zdnd11an1n64x5 FILLER_66_982 ();
 b15zdnd11an1n64x5 FILLER_66_1046 ();
 b15zdnd11an1n04x5 FILLER_66_1110 ();
 b15zdnd00an1n01x5 FILLER_66_1114 ();
 b15zdnd11an1n64x5 FILLER_66_1129 ();
 b15zdnd11an1n32x5 FILLER_66_1193 ();
 b15zdnd11an1n16x5 FILLER_66_1225 ();
 b15zdnd11an1n04x5 FILLER_66_1241 ();
 b15zdnd00an1n01x5 FILLER_66_1245 ();
 b15zdnd11an1n64x5 FILLER_66_1249 ();
 b15zdnd11an1n64x5 FILLER_66_1313 ();
 b15zdnd11an1n64x5 FILLER_66_1377 ();
 b15zdnd11an1n64x5 FILLER_66_1441 ();
 b15zdnd11an1n64x5 FILLER_66_1505 ();
 b15zdnd11an1n32x5 FILLER_66_1569 ();
 b15zdnd00an1n01x5 FILLER_66_1601 ();
 b15zdnd11an1n64x5 FILLER_66_1609 ();
 b15zdnd11an1n64x5 FILLER_66_1673 ();
 b15zdnd11an1n64x5 FILLER_66_1737 ();
 b15zdnd11an1n64x5 FILLER_66_1801 ();
 b15zdnd11an1n64x5 FILLER_66_1865 ();
 b15zdnd11an1n64x5 FILLER_66_1929 ();
 b15zdnd11an1n64x5 FILLER_66_1993 ();
 b15zdnd11an1n64x5 FILLER_66_2057 ();
 b15zdnd11an1n32x5 FILLER_66_2121 ();
 b15zdnd00an1n01x5 FILLER_66_2153 ();
 b15zdnd11an1n64x5 FILLER_66_2162 ();
 b15zdnd11an1n32x5 FILLER_66_2226 ();
 b15zdnd11an1n16x5 FILLER_66_2258 ();
 b15zdnd00an1n02x5 FILLER_66_2274 ();
 b15zdnd11an1n64x5 FILLER_67_0 ();
 b15zdnd11an1n64x5 FILLER_67_64 ();
 b15zdnd11an1n64x5 FILLER_67_128 ();
 b15zdnd11an1n64x5 FILLER_67_192 ();
 b15zdnd11an1n64x5 FILLER_67_256 ();
 b15zdnd11an1n64x5 FILLER_67_320 ();
 b15zdnd11an1n64x5 FILLER_67_384 ();
 b15zdnd11an1n16x5 FILLER_67_448 ();
 b15zdnd11an1n04x5 FILLER_67_464 ();
 b15zdnd11an1n04x5 FILLER_67_508 ();
 b15zdnd11an1n64x5 FILLER_67_515 ();
 b15zdnd11an1n64x5 FILLER_67_579 ();
 b15zdnd11an1n64x5 FILLER_67_643 ();
 b15zdnd11an1n64x5 FILLER_67_707 ();
 b15zdnd11an1n32x5 FILLER_67_771 ();
 b15zdnd11an1n16x5 FILLER_67_803 ();
 b15zdnd00an1n02x5 FILLER_67_819 ();
 b15zdnd11an1n64x5 FILLER_67_829 ();
 b15zdnd11an1n64x5 FILLER_67_893 ();
 b15zdnd11an1n64x5 FILLER_67_957 ();
 b15zdnd11an1n64x5 FILLER_67_1021 ();
 b15zdnd11an1n64x5 FILLER_67_1085 ();
 b15zdnd11an1n64x5 FILLER_67_1149 ();
 b15zdnd11an1n64x5 FILLER_67_1213 ();
 b15zdnd11an1n08x5 FILLER_67_1277 ();
 b15zdnd11an1n04x5 FILLER_67_1285 ();
 b15zdnd00an1n02x5 FILLER_67_1289 ();
 b15zdnd00an1n01x5 FILLER_67_1291 ();
 b15zdnd11an1n64x5 FILLER_67_1303 ();
 b15zdnd11an1n64x5 FILLER_67_1367 ();
 b15zdnd11an1n64x5 FILLER_67_1431 ();
 b15zdnd11an1n64x5 FILLER_67_1495 ();
 b15zdnd11an1n64x5 FILLER_67_1559 ();
 b15zdnd11an1n64x5 FILLER_67_1623 ();
 b15zdnd11an1n64x5 FILLER_67_1687 ();
 b15zdnd11an1n64x5 FILLER_67_1751 ();
 b15zdnd11an1n64x5 FILLER_67_1815 ();
 b15zdnd11an1n64x5 FILLER_67_1879 ();
 b15zdnd11an1n64x5 FILLER_67_1943 ();
 b15zdnd11an1n64x5 FILLER_67_2007 ();
 b15zdnd11an1n64x5 FILLER_67_2071 ();
 b15zdnd11an1n64x5 FILLER_67_2135 ();
 b15zdnd11an1n64x5 FILLER_67_2199 ();
 b15zdnd11an1n16x5 FILLER_67_2263 ();
 b15zdnd11an1n04x5 FILLER_67_2279 ();
 b15zdnd00an1n01x5 FILLER_67_2283 ();
 b15zdnd11an1n64x5 FILLER_68_8 ();
 b15zdnd11an1n64x5 FILLER_68_72 ();
 b15zdnd11an1n64x5 FILLER_68_136 ();
 b15zdnd11an1n64x5 FILLER_68_200 ();
 b15zdnd11an1n64x5 FILLER_68_264 ();
 b15zdnd11an1n64x5 FILLER_68_328 ();
 b15zdnd11an1n64x5 FILLER_68_392 ();
 b15zdnd11an1n64x5 FILLER_68_456 ();
 b15zdnd11an1n64x5 FILLER_68_520 ();
 b15zdnd11an1n64x5 FILLER_68_584 ();
 b15zdnd11an1n64x5 FILLER_68_648 ();
 b15zdnd11an1n04x5 FILLER_68_712 ();
 b15zdnd00an1n02x5 FILLER_68_716 ();
 b15zdnd11an1n64x5 FILLER_68_726 ();
 b15zdnd11an1n64x5 FILLER_68_790 ();
 b15zdnd11an1n64x5 FILLER_68_854 ();
 b15zdnd11an1n32x5 FILLER_68_918 ();
 b15zdnd11an1n16x5 FILLER_68_950 ();
 b15zdnd11an1n08x5 FILLER_68_966 ();
 b15zdnd11an1n04x5 FILLER_68_974 ();
 b15zdnd00an1n02x5 FILLER_68_978 ();
 b15zdnd00an1n01x5 FILLER_68_980 ();
 b15zdnd11an1n64x5 FILLER_68_990 ();
 b15zdnd11an1n64x5 FILLER_68_1054 ();
 b15zdnd11an1n64x5 FILLER_68_1118 ();
 b15zdnd11an1n64x5 FILLER_68_1182 ();
 b15zdnd11an1n64x5 FILLER_68_1246 ();
 b15zdnd11an1n64x5 FILLER_68_1310 ();
 b15zdnd11an1n64x5 FILLER_68_1374 ();
 b15zdnd11an1n64x5 FILLER_68_1438 ();
 b15zdnd11an1n64x5 FILLER_68_1502 ();
 b15zdnd11an1n64x5 FILLER_68_1566 ();
 b15zdnd11an1n64x5 FILLER_68_1630 ();
 b15zdnd11an1n64x5 FILLER_68_1694 ();
 b15zdnd11an1n64x5 FILLER_68_1758 ();
 b15zdnd11an1n64x5 FILLER_68_1822 ();
 b15zdnd11an1n64x5 FILLER_68_1886 ();
 b15zdnd11an1n64x5 FILLER_68_1950 ();
 b15zdnd11an1n08x5 FILLER_68_2014 ();
 b15zdnd11an1n04x5 FILLER_68_2026 ();
 b15zdnd11an1n04x5 FILLER_68_2035 ();
 b15zdnd11an1n32x5 FILLER_68_2044 ();
 b15zdnd11an1n08x5 FILLER_68_2076 ();
 b15zdnd11an1n64x5 FILLER_68_2087 ();
 b15zdnd00an1n02x5 FILLER_68_2151 ();
 b15zdnd00an1n01x5 FILLER_68_2153 ();
 b15zdnd11an1n64x5 FILLER_68_2162 ();
 b15zdnd11an1n32x5 FILLER_68_2226 ();
 b15zdnd11an1n16x5 FILLER_68_2258 ();
 b15zdnd00an1n02x5 FILLER_68_2274 ();
 b15zdnd11an1n64x5 FILLER_69_0 ();
 b15zdnd11an1n64x5 FILLER_69_64 ();
 b15zdnd11an1n64x5 FILLER_69_128 ();
 b15zdnd11an1n64x5 FILLER_69_192 ();
 b15zdnd11an1n04x5 FILLER_69_256 ();
 b15zdnd00an1n02x5 FILLER_69_260 ();
 b15zdnd11an1n64x5 FILLER_69_267 ();
 b15zdnd11an1n64x5 FILLER_69_331 ();
 b15zdnd11an1n64x5 FILLER_69_395 ();
 b15zdnd11an1n32x5 FILLER_69_459 ();
 b15zdnd11an1n04x5 FILLER_69_491 ();
 b15zdnd00an1n02x5 FILLER_69_495 ();
 b15zdnd11an1n64x5 FILLER_69_513 ();
 b15zdnd11an1n64x5 FILLER_69_577 ();
 b15zdnd11an1n64x5 FILLER_69_641 ();
 b15zdnd11an1n32x5 FILLER_69_705 ();
 b15zdnd11an1n16x5 FILLER_69_737 ();
 b15zdnd11an1n08x5 FILLER_69_753 ();
 b15zdnd11an1n04x5 FILLER_69_761 ();
 b15zdnd00an1n02x5 FILLER_69_765 ();
 b15zdnd00an1n01x5 FILLER_69_767 ();
 b15zdnd11an1n64x5 FILLER_69_771 ();
 b15zdnd11an1n64x5 FILLER_69_835 ();
 b15zdnd11an1n64x5 FILLER_69_899 ();
 b15zdnd11an1n64x5 FILLER_69_963 ();
 b15zdnd11an1n64x5 FILLER_69_1027 ();
 b15zdnd11an1n64x5 FILLER_69_1091 ();
 b15zdnd11an1n64x5 FILLER_69_1155 ();
 b15zdnd11an1n16x5 FILLER_69_1219 ();
 b15zdnd11an1n08x5 FILLER_69_1235 ();
 b15zdnd11an1n04x5 FILLER_69_1243 ();
 b15zdnd11an1n64x5 FILLER_69_1289 ();
 b15zdnd11an1n64x5 FILLER_69_1353 ();
 b15zdnd11an1n32x5 FILLER_69_1417 ();
 b15zdnd11an1n08x5 FILLER_69_1449 ();
 b15zdnd11an1n04x5 FILLER_69_1457 ();
 b15zdnd00an1n02x5 FILLER_69_1461 ();
 b15zdnd11an1n64x5 FILLER_69_1471 ();
 b15zdnd11an1n64x5 FILLER_69_1535 ();
 b15zdnd11an1n64x5 FILLER_69_1599 ();
 b15zdnd11an1n64x5 FILLER_69_1663 ();
 b15zdnd11an1n64x5 FILLER_69_1727 ();
 b15zdnd11an1n64x5 FILLER_69_1791 ();
 b15zdnd11an1n32x5 FILLER_69_1855 ();
 b15zdnd11an1n16x5 FILLER_69_1887 ();
 b15zdnd11an1n08x5 FILLER_69_1903 ();
 b15zdnd11an1n04x5 FILLER_69_1911 ();
 b15zdnd00an1n01x5 FILLER_69_1915 ();
 b15zdnd11an1n04x5 FILLER_69_1919 ();
 b15zdnd11an1n08x5 FILLER_69_1926 ();
 b15zdnd00an1n02x5 FILLER_69_1934 ();
 b15zdnd00an1n01x5 FILLER_69_1936 ();
 b15zdnd11an1n64x5 FILLER_69_1940 ();
 b15zdnd11an1n16x5 FILLER_69_2004 ();
 b15zdnd00an1n02x5 FILLER_69_2020 ();
 b15zdnd11an1n04x5 FILLER_69_2033 ();
 b15zdnd11an1n04x5 FILLER_69_2050 ();
 b15zdnd11an1n08x5 FILLER_69_2057 ();
 b15zdnd00an1n01x5 FILLER_69_2065 ();
 b15zdnd11an1n64x5 FILLER_69_2118 ();
 b15zdnd11an1n64x5 FILLER_69_2182 ();
 b15zdnd11an1n32x5 FILLER_69_2246 ();
 b15zdnd11an1n04x5 FILLER_69_2278 ();
 b15zdnd00an1n02x5 FILLER_69_2282 ();
 b15zdnd11an1n64x5 FILLER_70_8 ();
 b15zdnd11an1n64x5 FILLER_70_72 ();
 b15zdnd11an1n64x5 FILLER_70_136 ();
 b15zdnd11an1n32x5 FILLER_70_200 ();
 b15zdnd11an1n08x5 FILLER_70_232 ();
 b15zdnd11an1n04x5 FILLER_70_240 ();
 b15zdnd11an1n04x5 FILLER_70_253 ();
 b15zdnd11an1n04x5 FILLER_70_267 ();
 b15zdnd11an1n64x5 FILLER_70_278 ();
 b15zdnd11an1n64x5 FILLER_70_342 ();
 b15zdnd11an1n64x5 FILLER_70_406 ();
 b15zdnd11an1n08x5 FILLER_70_470 ();
 b15zdnd00an1n02x5 FILLER_70_478 ();
 b15zdnd00an1n01x5 FILLER_70_480 ();
 b15zdnd11an1n64x5 FILLER_70_508 ();
 b15zdnd11an1n64x5 FILLER_70_572 ();
 b15zdnd11an1n08x5 FILLER_70_636 ();
 b15zdnd11an1n64x5 FILLER_70_647 ();
 b15zdnd11an1n04x5 FILLER_70_711 ();
 b15zdnd00an1n02x5 FILLER_70_715 ();
 b15zdnd00an1n01x5 FILLER_70_717 ();
 b15zdnd11an1n32x5 FILLER_70_726 ();
 b15zdnd00an1n02x5 FILLER_70_758 ();
 b15zdnd00an1n01x5 FILLER_70_760 ();
 b15zdnd11an1n04x5 FILLER_70_764 ();
 b15zdnd11an1n08x5 FILLER_70_771 ();
 b15zdnd00an1n02x5 FILLER_70_779 ();
 b15zdnd00an1n01x5 FILLER_70_781 ();
 b15zdnd11an1n04x5 FILLER_70_785 ();
 b15zdnd11an1n64x5 FILLER_70_792 ();
 b15zdnd11an1n64x5 FILLER_70_856 ();
 b15zdnd11an1n64x5 FILLER_70_920 ();
 b15zdnd11an1n04x5 FILLER_70_984 ();
 b15zdnd00an1n02x5 FILLER_70_988 ();
 b15zdnd00an1n01x5 FILLER_70_990 ();
 b15zdnd11an1n64x5 FILLER_70_1036 ();
 b15zdnd11an1n64x5 FILLER_70_1100 ();
 b15zdnd11an1n64x5 FILLER_70_1164 ();
 b15zdnd11an1n64x5 FILLER_70_1228 ();
 b15zdnd11an1n64x5 FILLER_70_1292 ();
 b15zdnd11an1n08x5 FILLER_70_1356 ();
 b15zdnd11an1n04x5 FILLER_70_1364 ();
 b15zdnd00an1n02x5 FILLER_70_1368 ();
 b15zdnd00an1n01x5 FILLER_70_1370 ();
 b15zdnd11an1n32x5 FILLER_70_1396 ();
 b15zdnd00an1n02x5 FILLER_70_1428 ();
 b15zdnd00an1n01x5 FILLER_70_1430 ();
 b15zdnd11an1n04x5 FILLER_70_1434 ();
 b15zdnd11an1n64x5 FILLER_70_1441 ();
 b15zdnd11an1n64x5 FILLER_70_1505 ();
 b15zdnd11an1n64x5 FILLER_70_1569 ();
 b15zdnd11an1n64x5 FILLER_70_1633 ();
 b15zdnd11an1n64x5 FILLER_70_1697 ();
 b15zdnd11an1n64x5 FILLER_70_1761 ();
 b15zdnd11an1n64x5 FILLER_70_1825 ();
 b15zdnd00an1n02x5 FILLER_70_1889 ();
 b15zdnd11an1n64x5 FILLER_70_1943 ();
 b15zdnd11an1n08x5 FILLER_70_2007 ();
 b15zdnd00an1n02x5 FILLER_70_2015 ();
 b15zdnd00an1n01x5 FILLER_70_2017 ();
 b15zdnd11an1n04x5 FILLER_70_2028 ();
 b15zdnd11an1n16x5 FILLER_70_2045 ();
 b15zdnd00an1n02x5 FILLER_70_2061 ();
 b15zdnd11an1n04x5 FILLER_70_2105 ();
 b15zdnd11an1n32x5 FILLER_70_2112 ();
 b15zdnd11an1n08x5 FILLER_70_2144 ();
 b15zdnd00an1n02x5 FILLER_70_2152 ();
 b15zdnd11an1n64x5 FILLER_70_2162 ();
 b15zdnd11an1n32x5 FILLER_70_2226 ();
 b15zdnd11an1n16x5 FILLER_70_2258 ();
 b15zdnd00an1n02x5 FILLER_70_2274 ();
 b15zdnd11an1n64x5 FILLER_71_0 ();
 b15zdnd11an1n64x5 FILLER_71_64 ();
 b15zdnd11an1n64x5 FILLER_71_128 ();
 b15zdnd11an1n32x5 FILLER_71_192 ();
 b15zdnd11an1n08x5 FILLER_71_224 ();
 b15zdnd11an1n04x5 FILLER_71_232 ();
 b15zdnd00an1n02x5 FILLER_71_236 ();
 b15zdnd00an1n01x5 FILLER_71_238 ();
 b15zdnd11an1n64x5 FILLER_71_281 ();
 b15zdnd11an1n64x5 FILLER_71_345 ();
 b15zdnd11an1n64x5 FILLER_71_409 ();
 b15zdnd11an1n64x5 FILLER_71_473 ();
 b15zdnd11an1n64x5 FILLER_71_537 ();
 b15zdnd11an1n32x5 FILLER_71_601 ();
 b15zdnd00an1n02x5 FILLER_71_633 ();
 b15zdnd00an1n01x5 FILLER_71_635 ();
 b15zdnd11an1n04x5 FILLER_71_639 ();
 b15zdnd11an1n64x5 FILLER_71_646 ();
 b15zdnd11an1n32x5 FILLER_71_710 ();
 b15zdnd00an1n01x5 FILLER_71_742 ();
 b15zdnd11an1n04x5 FILLER_71_795 ();
 b15zdnd11an1n64x5 FILLER_71_802 ();
 b15zdnd11an1n64x5 FILLER_71_866 ();
 b15zdnd00an1n01x5 FILLER_71_930 ();
 b15zdnd11an1n04x5 FILLER_71_934 ();
 b15zdnd00an1n02x5 FILLER_71_938 ();
 b15zdnd00an1n01x5 FILLER_71_940 ();
 b15zdnd11an1n64x5 FILLER_71_944 ();
 b15zdnd11an1n32x5 FILLER_71_1008 ();
 b15zdnd11an1n16x5 FILLER_71_1040 ();
 b15zdnd11an1n08x5 FILLER_71_1056 ();
 b15zdnd11an1n04x5 FILLER_71_1064 ();
 b15zdnd00an1n02x5 FILLER_71_1068 ();
 b15zdnd00an1n01x5 FILLER_71_1070 ();
 b15zdnd11an1n04x5 FILLER_71_1074 ();
 b15zdnd11an1n04x5 FILLER_71_1081 ();
 b15zdnd11an1n16x5 FILLER_71_1088 ();
 b15zdnd00an1n02x5 FILLER_71_1104 ();
 b15zdnd00an1n01x5 FILLER_71_1106 ();
 b15zdnd11an1n16x5 FILLER_71_1118 ();
 b15zdnd00an1n02x5 FILLER_71_1134 ();
 b15zdnd00an1n01x5 FILLER_71_1136 ();
 b15zdnd11an1n64x5 FILLER_71_1145 ();
 b15zdnd11an1n64x5 FILLER_71_1209 ();
 b15zdnd11an1n64x5 FILLER_71_1273 ();
 b15zdnd11an1n04x5 FILLER_71_1337 ();
 b15zdnd11an1n04x5 FILLER_71_1350 ();
 b15zdnd00an1n02x5 FILLER_71_1354 ();
 b15zdnd11an1n04x5 FILLER_71_1395 ();
 b15zdnd11an1n64x5 FILLER_71_1439 ();
 b15zdnd11an1n64x5 FILLER_71_1503 ();
 b15zdnd11an1n64x5 FILLER_71_1567 ();
 b15zdnd11an1n64x5 FILLER_71_1631 ();
 b15zdnd11an1n64x5 FILLER_71_1695 ();
 b15zdnd11an1n64x5 FILLER_71_1759 ();
 b15zdnd11an1n64x5 FILLER_71_1823 ();
 b15zdnd11an1n16x5 FILLER_71_1887 ();
 b15zdnd11an1n04x5 FILLER_71_1903 ();
 b15zdnd00an1n02x5 FILLER_71_1907 ();
 b15zdnd00an1n01x5 FILLER_71_1909 ();
 b15zdnd11an1n32x5 FILLER_71_1962 ();
 b15zdnd11an1n04x5 FILLER_71_1994 ();
 b15zdnd00an1n01x5 FILLER_71_1998 ();
 b15zdnd11an1n08x5 FILLER_71_2041 ();
 b15zdnd11an1n08x5 FILLER_71_2060 ();
 b15zdnd11an1n04x5 FILLER_71_2068 ();
 b15zdnd00an1n02x5 FILLER_71_2072 ();
 b15zdnd00an1n01x5 FILLER_71_2074 ();
 b15zdnd11an1n64x5 FILLER_71_2117 ();
 b15zdnd11an1n64x5 FILLER_71_2181 ();
 b15zdnd11an1n32x5 FILLER_71_2245 ();
 b15zdnd11an1n04x5 FILLER_71_2277 ();
 b15zdnd00an1n02x5 FILLER_71_2281 ();
 b15zdnd00an1n01x5 FILLER_71_2283 ();
 b15zdnd11an1n64x5 FILLER_72_8 ();
 b15zdnd11an1n64x5 FILLER_72_72 ();
 b15zdnd11an1n64x5 FILLER_72_136 ();
 b15zdnd11an1n16x5 FILLER_72_200 ();
 b15zdnd11an1n08x5 FILLER_72_216 ();
 b15zdnd11an1n08x5 FILLER_72_227 ();
 b15zdnd00an1n02x5 FILLER_72_235 ();
 b15zdnd11an1n04x5 FILLER_72_244 ();
 b15zdnd11an1n64x5 FILLER_72_290 ();
 b15zdnd11an1n64x5 FILLER_72_354 ();
 b15zdnd11an1n64x5 FILLER_72_418 ();
 b15zdnd11an1n64x5 FILLER_72_482 ();
 b15zdnd11an1n64x5 FILLER_72_546 ();
 b15zdnd11an1n08x5 FILLER_72_610 ();
 b15zdnd00an1n01x5 FILLER_72_618 ();
 b15zdnd11an1n32x5 FILLER_72_671 ();
 b15zdnd11an1n08x5 FILLER_72_703 ();
 b15zdnd11an1n04x5 FILLER_72_711 ();
 b15zdnd00an1n02x5 FILLER_72_715 ();
 b15zdnd00an1n01x5 FILLER_72_717 ();
 b15zdnd11an1n08x5 FILLER_72_726 ();
 b15zdnd11an1n04x5 FILLER_72_734 ();
 b15zdnd11an1n04x5 FILLER_72_747 ();
 b15zdnd11an1n04x5 FILLER_72_757 ();
 b15zdnd11an1n04x5 FILLER_72_813 ();
 b15zdnd11an1n64x5 FILLER_72_824 ();
 b15zdnd11an1n32x5 FILLER_72_888 ();
 b15zdnd11an1n04x5 FILLER_72_923 ();
 b15zdnd00an1n01x5 FILLER_72_927 ();
 b15zdnd11an1n04x5 FILLER_72_931 ();
 b15zdnd11an1n04x5 FILLER_72_938 ();
 b15zdnd11an1n04x5 FILLER_72_945 ();
 b15zdnd11an1n08x5 FILLER_72_952 ();
 b15zdnd11an1n64x5 FILLER_72_969 ();
 b15zdnd11an1n16x5 FILLER_72_1033 ();
 b15zdnd00an1n02x5 FILLER_72_1049 ();
 b15zdnd11an1n64x5 FILLER_72_1103 ();
 b15zdnd11an1n64x5 FILLER_72_1167 ();
 b15zdnd11an1n64x5 FILLER_72_1231 ();
 b15zdnd11an1n64x5 FILLER_72_1295 ();
 b15zdnd11an1n64x5 FILLER_72_1359 ();
 b15zdnd11an1n64x5 FILLER_72_1423 ();
 b15zdnd11an1n64x5 FILLER_72_1487 ();
 b15zdnd11an1n64x5 FILLER_72_1551 ();
 b15zdnd11an1n64x5 FILLER_72_1615 ();
 b15zdnd11an1n64x5 FILLER_72_1679 ();
 b15zdnd11an1n64x5 FILLER_72_1743 ();
 b15zdnd11an1n16x5 FILLER_72_1807 ();
 b15zdnd00an1n02x5 FILLER_72_1823 ();
 b15zdnd11an1n64x5 FILLER_72_1828 ();
 b15zdnd11an1n16x5 FILLER_72_1892 ();
 b15zdnd11an1n08x5 FILLER_72_1908 ();
 b15zdnd00an1n01x5 FILLER_72_1916 ();
 b15zdnd11an1n08x5 FILLER_72_1920 ();
 b15zdnd11an1n04x5 FILLER_72_1931 ();
 b15zdnd00an1n01x5 FILLER_72_1935 ();
 b15zdnd11an1n64x5 FILLER_72_1978 ();
 b15zdnd11an1n32x5 FILLER_72_2042 ();
 b15zdnd11an1n08x5 FILLER_72_2074 ();
 b15zdnd11an1n04x5 FILLER_72_2082 ();
 b15zdnd00an1n02x5 FILLER_72_2086 ();
 b15zdnd00an1n01x5 FILLER_72_2088 ();
 b15zdnd11an1n32x5 FILLER_72_2092 ();
 b15zdnd11an1n16x5 FILLER_72_2124 ();
 b15zdnd11an1n08x5 FILLER_72_2140 ();
 b15zdnd11an1n04x5 FILLER_72_2148 ();
 b15zdnd00an1n02x5 FILLER_72_2152 ();
 b15zdnd11an1n64x5 FILLER_72_2162 ();
 b15zdnd11an1n32x5 FILLER_72_2226 ();
 b15zdnd11an1n16x5 FILLER_72_2258 ();
 b15zdnd00an1n02x5 FILLER_72_2274 ();
 b15zdnd11an1n64x5 FILLER_73_0 ();
 b15zdnd11an1n64x5 FILLER_73_64 ();
 b15zdnd11an1n64x5 FILLER_73_128 ();
 b15zdnd11an1n08x5 FILLER_73_192 ();
 b15zdnd00an1n02x5 FILLER_73_200 ();
 b15zdnd11an1n04x5 FILLER_73_254 ();
 b15zdnd11an1n04x5 FILLER_73_265 ();
 b15zdnd11an1n64x5 FILLER_73_311 ();
 b15zdnd11an1n64x5 FILLER_73_375 ();
 b15zdnd11an1n64x5 FILLER_73_439 ();
 b15zdnd11an1n64x5 FILLER_73_503 ();
 b15zdnd11an1n16x5 FILLER_73_567 ();
 b15zdnd11an1n04x5 FILLER_73_583 ();
 b15zdnd00an1n02x5 FILLER_73_587 ();
 b15zdnd11an1n32x5 FILLER_73_596 ();
 b15zdnd11an1n04x5 FILLER_73_628 ();
 b15zdnd00an1n02x5 FILLER_73_632 ();
 b15zdnd11an1n08x5 FILLER_73_637 ();
 b15zdnd00an1n02x5 FILLER_73_645 ();
 b15zdnd11an1n08x5 FILLER_73_674 ();
 b15zdnd11an1n32x5 FILLER_73_691 ();
 b15zdnd11an1n16x5 FILLER_73_723 ();
 b15zdnd00an1n02x5 FILLER_73_739 ();
 b15zdnd11an1n16x5 FILLER_73_793 ();
 b15zdnd00an1n01x5 FILLER_73_809 ();
 b15zdnd11an1n64x5 FILLER_73_818 ();
 b15zdnd11an1n32x5 FILLER_73_882 ();
 b15zdnd11an1n04x5 FILLER_73_914 ();
 b15zdnd11an1n32x5 FILLER_73_970 ();
 b15zdnd11an1n08x5 FILLER_73_1002 ();
 b15zdnd11an1n04x5 FILLER_73_1010 ();
 b15zdnd00an1n02x5 FILLER_73_1014 ();
 b15zdnd11an1n16x5 FILLER_73_1025 ();
 b15zdnd11an1n08x5 FILLER_73_1041 ();
 b15zdnd00an1n02x5 FILLER_73_1049 ();
 b15zdnd11an1n16x5 FILLER_73_1103 ();
 b15zdnd11an1n08x5 FILLER_73_1119 ();
 b15zdnd11an1n08x5 FILLER_73_1131 ();
 b15zdnd11an1n16x5 FILLER_73_1143 ();
 b15zdnd11an1n16x5 FILLER_73_1165 ();
 b15zdnd00an1n01x5 FILLER_73_1181 ();
 b15zdnd11an1n64x5 FILLER_73_1186 ();
 b15zdnd11an1n64x5 FILLER_73_1250 ();
 b15zdnd11an1n64x5 FILLER_73_1314 ();
 b15zdnd11an1n64x5 FILLER_73_1378 ();
 b15zdnd11an1n64x5 FILLER_73_1442 ();
 b15zdnd11an1n64x5 FILLER_73_1506 ();
 b15zdnd11an1n64x5 FILLER_73_1570 ();
 b15zdnd11an1n64x5 FILLER_73_1634 ();
 b15zdnd11an1n64x5 FILLER_73_1698 ();
 b15zdnd11an1n32x5 FILLER_73_1762 ();
 b15zdnd11an1n04x5 FILLER_73_1794 ();
 b15zdnd00an1n01x5 FILLER_73_1798 ();
 b15zdnd11an1n64x5 FILLER_73_1851 ();
 b15zdnd11an1n16x5 FILLER_73_1915 ();
 b15zdnd11an1n04x5 FILLER_73_1931 ();
 b15zdnd11an1n64x5 FILLER_73_1938 ();
 b15zdnd11an1n64x5 FILLER_73_2002 ();
 b15zdnd11an1n64x5 FILLER_73_2066 ();
 b15zdnd11an1n64x5 FILLER_73_2130 ();
 b15zdnd11an1n64x5 FILLER_73_2194 ();
 b15zdnd11an1n16x5 FILLER_73_2258 ();
 b15zdnd11an1n08x5 FILLER_73_2274 ();
 b15zdnd00an1n02x5 FILLER_73_2282 ();
 b15zdnd11an1n64x5 FILLER_74_8 ();
 b15zdnd11an1n64x5 FILLER_74_72 ();
 b15zdnd11an1n64x5 FILLER_74_136 ();
 b15zdnd11an1n16x5 FILLER_74_200 ();
 b15zdnd11an1n08x5 FILLER_74_216 ();
 b15zdnd11an1n04x5 FILLER_74_224 ();
 b15zdnd11an1n16x5 FILLER_74_231 ();
 b15zdnd11an1n08x5 FILLER_74_247 ();
 b15zdnd00an1n02x5 FILLER_74_255 ();
 b15zdnd00an1n01x5 FILLER_74_257 ();
 b15zdnd11an1n04x5 FILLER_74_263 ();
 b15zdnd00an1n02x5 FILLER_74_267 ();
 b15zdnd11an1n04x5 FILLER_74_273 ();
 b15zdnd00an1n02x5 FILLER_74_277 ();
 b15zdnd11an1n64x5 FILLER_74_289 ();
 b15zdnd11an1n04x5 FILLER_74_353 ();
 b15zdnd00an1n02x5 FILLER_74_357 ();
 b15zdnd00an1n01x5 FILLER_74_359 ();
 b15zdnd11an1n64x5 FILLER_74_391 ();
 b15zdnd11an1n64x5 FILLER_74_455 ();
 b15zdnd11an1n16x5 FILLER_74_519 ();
 b15zdnd11an1n04x5 FILLER_74_535 ();
 b15zdnd11an1n32x5 FILLER_74_543 ();
 b15zdnd11an1n16x5 FILLER_74_575 ();
 b15zdnd11an1n08x5 FILLER_74_591 ();
 b15zdnd11an1n04x5 FILLER_74_599 ();
 b15zdnd11an1n04x5 FILLER_74_611 ();
 b15zdnd11an1n04x5 FILLER_74_667 ();
 b15zdnd11an1n16x5 FILLER_74_674 ();
 b15zdnd11an1n08x5 FILLER_74_690 ();
 b15zdnd00an1n01x5 FILLER_74_698 ();
 b15zdnd11an1n08x5 FILLER_74_706 ();
 b15zdnd11an1n04x5 FILLER_74_714 ();
 b15zdnd11an1n16x5 FILLER_74_726 ();
 b15zdnd11an1n64x5 FILLER_74_794 ();
 b15zdnd11an1n32x5 FILLER_74_858 ();
 b15zdnd11an1n16x5 FILLER_74_890 ();
 b15zdnd11an1n04x5 FILLER_74_958 ();
 b15zdnd11an1n64x5 FILLER_74_965 ();
 b15zdnd11an1n32x5 FILLER_74_1029 ();
 b15zdnd11an1n08x5 FILLER_74_1061 ();
 b15zdnd00an1n02x5 FILLER_74_1069 ();
 b15zdnd11an1n04x5 FILLER_74_1074 ();
 b15zdnd11an1n04x5 FILLER_74_1081 ();
 b15zdnd11an1n64x5 FILLER_74_1088 ();
 b15zdnd00an1n02x5 FILLER_74_1152 ();
 b15zdnd11an1n04x5 FILLER_74_1162 ();
 b15zdnd00an1n01x5 FILLER_74_1166 ();
 b15zdnd11an1n32x5 FILLER_74_1171 ();
 b15zdnd11an1n16x5 FILLER_74_1203 ();
 b15zdnd11an1n04x5 FILLER_74_1219 ();
 b15zdnd00an1n01x5 FILLER_74_1223 ();
 b15zdnd11an1n64x5 FILLER_74_1236 ();
 b15zdnd11an1n64x5 FILLER_74_1300 ();
 b15zdnd11an1n64x5 FILLER_74_1364 ();
 b15zdnd11an1n64x5 FILLER_74_1428 ();
 b15zdnd11an1n64x5 FILLER_74_1492 ();
 b15zdnd11an1n64x5 FILLER_74_1556 ();
 b15zdnd11an1n64x5 FILLER_74_1620 ();
 b15zdnd11an1n64x5 FILLER_74_1684 ();
 b15zdnd11an1n08x5 FILLER_74_1748 ();
 b15zdnd11an1n04x5 FILLER_74_1756 ();
 b15zdnd00an1n02x5 FILLER_74_1760 ();
 b15zdnd11an1n04x5 FILLER_74_1780 ();
 b15zdnd11an1n04x5 FILLER_74_1826 ();
 b15zdnd11an1n64x5 FILLER_74_1833 ();
 b15zdnd11an1n64x5 FILLER_74_1897 ();
 b15zdnd11an1n64x5 FILLER_74_1961 ();
 b15zdnd11an1n64x5 FILLER_74_2025 ();
 b15zdnd11an1n64x5 FILLER_74_2089 ();
 b15zdnd00an1n01x5 FILLER_74_2153 ();
 b15zdnd11an1n64x5 FILLER_74_2162 ();
 b15zdnd11an1n32x5 FILLER_74_2226 ();
 b15zdnd11an1n16x5 FILLER_74_2258 ();
 b15zdnd00an1n02x5 FILLER_74_2274 ();
 b15zdnd11an1n64x5 FILLER_75_0 ();
 b15zdnd11an1n64x5 FILLER_75_64 ();
 b15zdnd11an1n64x5 FILLER_75_128 ();
 b15zdnd11an1n16x5 FILLER_75_192 ();
 b15zdnd11an1n08x5 FILLER_75_208 ();
 b15zdnd11an1n04x5 FILLER_75_216 ();
 b15zdnd00an1n02x5 FILLER_75_220 ();
 b15zdnd11an1n32x5 FILLER_75_225 ();
 b15zdnd11an1n16x5 FILLER_75_257 ();
 b15zdnd11an1n64x5 FILLER_75_315 ();
 b15zdnd11an1n64x5 FILLER_75_379 ();
 b15zdnd11an1n64x5 FILLER_75_443 ();
 b15zdnd11an1n16x5 FILLER_75_507 ();
 b15zdnd11an1n08x5 FILLER_75_523 ();
 b15zdnd11an1n64x5 FILLER_75_541 ();
 b15zdnd11an1n16x5 FILLER_75_605 ();
 b15zdnd11an1n08x5 FILLER_75_621 ();
 b15zdnd00an1n02x5 FILLER_75_629 ();
 b15zdnd00an1n01x5 FILLER_75_631 ();
 b15zdnd11an1n04x5 FILLER_75_635 ();
 b15zdnd11an1n04x5 FILLER_75_642 ();
 b15zdnd11an1n04x5 FILLER_75_649 ();
 b15zdnd11an1n64x5 FILLER_75_656 ();
 b15zdnd11an1n08x5 FILLER_75_729 ();
 b15zdnd11an1n04x5 FILLER_75_737 ();
 b15zdnd00an1n02x5 FILLER_75_741 ();
 b15zdnd00an1n01x5 FILLER_75_743 ();
 b15zdnd11an1n08x5 FILLER_75_751 ();
 b15zdnd00an1n02x5 FILLER_75_759 ();
 b15zdnd00an1n01x5 FILLER_75_761 ();
 b15zdnd11an1n04x5 FILLER_75_765 ();
 b15zdnd11an1n04x5 FILLER_75_772 ();
 b15zdnd11an1n04x5 FILLER_75_779 ();
 b15zdnd11an1n64x5 FILLER_75_786 ();
 b15zdnd11an1n32x5 FILLER_75_850 ();
 b15zdnd11an1n16x5 FILLER_75_882 ();
 b15zdnd11an1n08x5 FILLER_75_898 ();
 b15zdnd11an1n04x5 FILLER_75_906 ();
 b15zdnd11an1n04x5 FILLER_75_962 ();
 b15zdnd11an1n32x5 FILLER_75_969 ();
 b15zdnd11an1n04x5 FILLER_75_1001 ();
 b15zdnd00an1n02x5 FILLER_75_1005 ();
 b15zdnd00an1n01x5 FILLER_75_1007 ();
 b15zdnd11an1n16x5 FILLER_75_1017 ();
 b15zdnd11an1n08x5 FILLER_75_1033 ();
 b15zdnd00an1n02x5 FILLER_75_1041 ();
 b15zdnd00an1n01x5 FILLER_75_1043 ();
 b15zdnd11an1n16x5 FILLER_75_1052 ();
 b15zdnd11an1n08x5 FILLER_75_1068 ();
 b15zdnd00an1n02x5 FILLER_75_1076 ();
 b15zdnd00an1n01x5 FILLER_75_1078 ();
 b15zdnd11an1n32x5 FILLER_75_1082 ();
 b15zdnd00an1n02x5 FILLER_75_1114 ();
 b15zdnd00an1n01x5 FILLER_75_1116 ();
 b15zdnd11an1n32x5 FILLER_75_1128 ();
 b15zdnd11an1n16x5 FILLER_75_1160 ();
 b15zdnd11an1n08x5 FILLER_75_1176 ();
 b15zdnd11an1n04x5 FILLER_75_1187 ();
 b15zdnd00an1n02x5 FILLER_75_1191 ();
 b15zdnd11an1n64x5 FILLER_75_1204 ();
 b15zdnd11an1n64x5 FILLER_75_1268 ();
 b15zdnd11an1n64x5 FILLER_75_1332 ();
 b15zdnd11an1n32x5 FILLER_75_1396 ();
 b15zdnd11an1n04x5 FILLER_75_1428 ();
 b15zdnd11an1n64x5 FILLER_75_1452 ();
 b15zdnd11an1n64x5 FILLER_75_1516 ();
 b15zdnd11an1n64x5 FILLER_75_1580 ();
 b15zdnd11an1n64x5 FILLER_75_1644 ();
 b15zdnd11an1n32x5 FILLER_75_1708 ();
 b15zdnd11an1n04x5 FILLER_75_1740 ();
 b15zdnd00an1n02x5 FILLER_75_1744 ();
 b15zdnd00an1n01x5 FILLER_75_1746 ();
 b15zdnd11an1n64x5 FILLER_75_1750 ();
 b15zdnd11an1n08x5 FILLER_75_1814 ();
 b15zdnd00an1n02x5 FILLER_75_1822 ();
 b15zdnd00an1n01x5 FILLER_75_1824 ();
 b15zdnd11an1n64x5 FILLER_75_1828 ();
 b15zdnd11an1n08x5 FILLER_75_1892 ();
 b15zdnd11an1n04x5 FILLER_75_1900 ();
 b15zdnd00an1n01x5 FILLER_75_1904 ();
 b15zdnd11an1n64x5 FILLER_75_1919 ();
 b15zdnd11an1n64x5 FILLER_75_1983 ();
 b15zdnd11an1n64x5 FILLER_75_2047 ();
 b15zdnd11an1n64x5 FILLER_75_2111 ();
 b15zdnd11an1n64x5 FILLER_75_2175 ();
 b15zdnd11an1n32x5 FILLER_75_2239 ();
 b15zdnd11an1n08x5 FILLER_75_2271 ();
 b15zdnd11an1n04x5 FILLER_75_2279 ();
 b15zdnd00an1n01x5 FILLER_75_2283 ();
 b15zdnd11an1n64x5 FILLER_76_8 ();
 b15zdnd11an1n64x5 FILLER_76_72 ();
 b15zdnd11an1n64x5 FILLER_76_136 ();
 b15zdnd11an1n64x5 FILLER_76_200 ();
 b15zdnd11an1n16x5 FILLER_76_264 ();
 b15zdnd00an1n02x5 FILLER_76_280 ();
 b15zdnd00an1n01x5 FILLER_76_282 ();
 b15zdnd11an1n64x5 FILLER_76_287 ();
 b15zdnd11an1n64x5 FILLER_76_351 ();
 b15zdnd11an1n64x5 FILLER_76_415 ();
 b15zdnd11an1n64x5 FILLER_76_479 ();
 b15zdnd11an1n64x5 FILLER_76_543 ();
 b15zdnd11an1n08x5 FILLER_76_607 ();
 b15zdnd00an1n01x5 FILLER_76_615 ();
 b15zdnd11an1n32x5 FILLER_76_668 ();
 b15zdnd11an1n16x5 FILLER_76_700 ();
 b15zdnd00an1n02x5 FILLER_76_716 ();
 b15zdnd11an1n16x5 FILLER_76_726 ();
 b15zdnd00an1n01x5 FILLER_76_742 ();
 b15zdnd11an1n08x5 FILLER_76_750 ();
 b15zdnd00an1n02x5 FILLER_76_758 ();
 b15zdnd00an1n01x5 FILLER_76_760 ();
 b15zdnd11an1n04x5 FILLER_76_764 ();
 b15zdnd11an1n32x5 FILLER_76_771 ();
 b15zdnd11an1n08x5 FILLER_76_803 ();
 b15zdnd11an1n04x5 FILLER_76_811 ();
 b15zdnd00an1n01x5 FILLER_76_815 ();
 b15zdnd11an1n64x5 FILLER_76_822 ();
 b15zdnd11an1n08x5 FILLER_76_886 ();
 b15zdnd11an1n04x5 FILLER_76_894 ();
 b15zdnd00an1n02x5 FILLER_76_898 ();
 b15zdnd11an1n04x5 FILLER_76_903 ();
 b15zdnd11an1n64x5 FILLER_76_959 ();
 b15zdnd11an1n16x5 FILLER_76_1023 ();
 b15zdnd11an1n08x5 FILLER_76_1039 ();
 b15zdnd11an1n04x5 FILLER_76_1047 ();
 b15zdnd00an1n01x5 FILLER_76_1051 ();
 b15zdnd11an1n64x5 FILLER_76_1104 ();
 b15zdnd11an1n16x5 FILLER_76_1168 ();
 b15zdnd11an1n64x5 FILLER_76_1199 ();
 b15zdnd11an1n64x5 FILLER_76_1263 ();
 b15zdnd11an1n32x5 FILLER_76_1327 ();
 b15zdnd11an1n08x5 FILLER_76_1359 ();
 b15zdnd00an1n01x5 FILLER_76_1367 ();
 b15zdnd11an1n64x5 FILLER_76_1371 ();
 b15zdnd11an1n08x5 FILLER_76_1435 ();
 b15zdnd11an1n04x5 FILLER_76_1443 ();
 b15zdnd11an1n64x5 FILLER_76_1454 ();
 b15zdnd11an1n64x5 FILLER_76_1518 ();
 b15zdnd11an1n64x5 FILLER_76_1582 ();
 b15zdnd11an1n64x5 FILLER_76_1646 ();
 b15zdnd11an1n32x5 FILLER_76_1710 ();
 b15zdnd11an1n04x5 FILLER_76_1742 ();
 b15zdnd00an1n02x5 FILLER_76_1746 ();
 b15zdnd11an1n04x5 FILLER_76_1751 ();
 b15zdnd11an1n64x5 FILLER_76_1758 ();
 b15zdnd11an1n64x5 FILLER_76_1822 ();
 b15zdnd11an1n64x5 FILLER_76_1886 ();
 b15zdnd11an1n32x5 FILLER_76_1950 ();
 b15zdnd11an1n16x5 FILLER_76_1982 ();
 b15zdnd11an1n04x5 FILLER_76_1998 ();
 b15zdnd00an1n02x5 FILLER_76_2002 ();
 b15zdnd11an1n64x5 FILLER_76_2008 ();
 b15zdnd11an1n64x5 FILLER_76_2072 ();
 b15zdnd11an1n16x5 FILLER_76_2136 ();
 b15zdnd00an1n02x5 FILLER_76_2152 ();
 b15zdnd11an1n64x5 FILLER_76_2162 ();
 b15zdnd11an1n32x5 FILLER_76_2226 ();
 b15zdnd11an1n16x5 FILLER_76_2258 ();
 b15zdnd00an1n02x5 FILLER_76_2274 ();
 b15zdnd11an1n64x5 FILLER_77_0 ();
 b15zdnd11an1n64x5 FILLER_77_64 ();
 b15zdnd11an1n64x5 FILLER_77_128 ();
 b15zdnd11an1n64x5 FILLER_77_192 ();
 b15zdnd11an1n32x5 FILLER_77_256 ();
 b15zdnd11an1n04x5 FILLER_77_288 ();
 b15zdnd00an1n01x5 FILLER_77_292 ();
 b15zdnd11an1n64x5 FILLER_77_296 ();
 b15zdnd11an1n64x5 FILLER_77_360 ();
 b15zdnd11an1n64x5 FILLER_77_424 ();
 b15zdnd11an1n64x5 FILLER_77_488 ();
 b15zdnd11an1n64x5 FILLER_77_552 ();
 b15zdnd00an1n02x5 FILLER_77_616 ();
 b15zdnd00an1n01x5 FILLER_77_618 ();
 b15zdnd11an1n08x5 FILLER_77_671 ();
 b15zdnd11an1n04x5 FILLER_77_679 ();
 b15zdnd00an1n02x5 FILLER_77_683 ();
 b15zdnd11an1n64x5 FILLER_77_691 ();
 b15zdnd11an1n64x5 FILLER_77_755 ();
 b15zdnd11an1n64x5 FILLER_77_819 ();
 b15zdnd11an1n16x5 FILLER_77_883 ();
 b15zdnd11an1n04x5 FILLER_77_899 ();
 b15zdnd00an1n02x5 FILLER_77_903 ();
 b15zdnd11an1n04x5 FILLER_77_919 ();
 b15zdnd11an1n04x5 FILLER_77_926 ();
 b15zdnd11an1n64x5 FILLER_77_957 ();
 b15zdnd11an1n32x5 FILLER_77_1021 ();
 b15zdnd11an1n64x5 FILLER_77_1105 ();
 b15zdnd11an1n64x5 FILLER_77_1169 ();
 b15zdnd11an1n64x5 FILLER_77_1233 ();
 b15zdnd11an1n32x5 FILLER_77_1297 ();
 b15zdnd11an1n08x5 FILLER_77_1329 ();
 b15zdnd11an1n04x5 FILLER_77_1337 ();
 b15zdnd00an1n01x5 FILLER_77_1341 ();
 b15zdnd11an1n32x5 FILLER_77_1394 ();
 b15zdnd11an1n16x5 FILLER_77_1426 ();
 b15zdnd00an1n01x5 FILLER_77_1442 ();
 b15zdnd11an1n64x5 FILLER_77_1468 ();
 b15zdnd11an1n64x5 FILLER_77_1532 ();
 b15zdnd11an1n64x5 FILLER_77_1596 ();
 b15zdnd11an1n32x5 FILLER_77_1660 ();
 b15zdnd11an1n16x5 FILLER_77_1692 ();
 b15zdnd00an1n02x5 FILLER_77_1708 ();
 b15zdnd00an1n01x5 FILLER_77_1710 ();
 b15zdnd11an1n08x5 FILLER_77_1715 ();
 b15zdnd11an1n64x5 FILLER_77_1775 ();
 b15zdnd11an1n64x5 FILLER_77_1839 ();
 b15zdnd11an1n64x5 FILLER_77_1903 ();
 b15zdnd11an1n32x5 FILLER_77_1967 ();
 b15zdnd11an1n16x5 FILLER_77_1999 ();
 b15zdnd11an1n08x5 FILLER_77_2015 ();
 b15zdnd11an1n04x5 FILLER_77_2023 ();
 b15zdnd00an1n01x5 FILLER_77_2027 ();
 b15zdnd11an1n08x5 FILLER_77_2033 ();
 b15zdnd11an1n04x5 FILLER_77_2041 ();
 b15zdnd00an1n01x5 FILLER_77_2045 ();
 b15zdnd11an1n64x5 FILLER_77_2088 ();
 b15zdnd11an1n64x5 FILLER_77_2152 ();
 b15zdnd11an1n64x5 FILLER_77_2216 ();
 b15zdnd11an1n04x5 FILLER_77_2280 ();
 b15zdnd11an1n64x5 FILLER_78_8 ();
 b15zdnd11an1n64x5 FILLER_78_72 ();
 b15zdnd11an1n64x5 FILLER_78_136 ();
 b15zdnd11an1n64x5 FILLER_78_200 ();
 b15zdnd11an1n16x5 FILLER_78_264 ();
 b15zdnd11an1n08x5 FILLER_78_280 ();
 b15zdnd11an1n04x5 FILLER_78_288 ();
 b15zdnd00an1n02x5 FILLER_78_292 ();
 b15zdnd11an1n32x5 FILLER_78_300 ();
 b15zdnd11an1n16x5 FILLER_78_332 ();
 b15zdnd00an1n02x5 FILLER_78_348 ();
 b15zdnd00an1n01x5 FILLER_78_350 ();
 b15zdnd11an1n64x5 FILLER_78_393 ();
 b15zdnd11an1n64x5 FILLER_78_457 ();
 b15zdnd11an1n32x5 FILLER_78_521 ();
 b15zdnd11an1n16x5 FILLER_78_553 ();
 b15zdnd11an1n04x5 FILLER_78_569 ();
 b15zdnd11an1n32x5 FILLER_78_584 ();
 b15zdnd11an1n16x5 FILLER_78_616 ();
 b15zdnd00an1n02x5 FILLER_78_632 ();
 b15zdnd00an1n01x5 FILLER_78_634 ();
 b15zdnd11an1n04x5 FILLER_78_638 ();
 b15zdnd11an1n04x5 FILLER_78_645 ();
 b15zdnd11an1n16x5 FILLER_78_652 ();
 b15zdnd11an1n04x5 FILLER_78_668 ();
 b15zdnd00an1n01x5 FILLER_78_672 ();
 b15zdnd11an1n32x5 FILLER_78_680 ();
 b15zdnd11an1n04x5 FILLER_78_712 ();
 b15zdnd00an1n02x5 FILLER_78_716 ();
 b15zdnd11an1n64x5 FILLER_78_726 ();
 b15zdnd11an1n64x5 FILLER_78_790 ();
 b15zdnd11an1n64x5 FILLER_78_854 ();
 b15zdnd11an1n08x5 FILLER_78_918 ();
 b15zdnd11an1n04x5 FILLER_78_929 ();
 b15zdnd11an1n64x5 FILLER_78_936 ();
 b15zdnd11an1n64x5 FILLER_78_1000 ();
 b15zdnd11an1n08x5 FILLER_78_1064 ();
 b15zdnd00an1n01x5 FILLER_78_1072 ();
 b15zdnd11an1n04x5 FILLER_78_1076 ();
 b15zdnd11an1n04x5 FILLER_78_1083 ();
 b15zdnd11an1n64x5 FILLER_78_1090 ();
 b15zdnd11an1n64x5 FILLER_78_1154 ();
 b15zdnd11an1n64x5 FILLER_78_1218 ();
 b15zdnd11an1n64x5 FILLER_78_1282 ();
 b15zdnd11an1n16x5 FILLER_78_1346 ();
 b15zdnd11an1n04x5 FILLER_78_1362 ();
 b15zdnd00an1n01x5 FILLER_78_1366 ();
 b15zdnd11an1n04x5 FILLER_78_1370 ();
 b15zdnd11an1n64x5 FILLER_78_1377 ();
 b15zdnd11an1n64x5 FILLER_78_1441 ();
 b15zdnd11an1n64x5 FILLER_78_1505 ();
 b15zdnd11an1n64x5 FILLER_78_1569 ();
 b15zdnd11an1n64x5 FILLER_78_1633 ();
 b15zdnd11an1n08x5 FILLER_78_1697 ();
 b15zdnd11an1n04x5 FILLER_78_1705 ();
 b15zdnd00an1n02x5 FILLER_78_1709 ();
 b15zdnd11an1n04x5 FILLER_78_1721 ();
 b15zdnd11an1n04x5 FILLER_78_1767 ();
 b15zdnd11an1n64x5 FILLER_78_1813 ();
 b15zdnd11an1n64x5 FILLER_78_1877 ();
 b15zdnd11an1n64x5 FILLER_78_1941 ();
 b15zdnd11an1n64x5 FILLER_78_2005 ();
 b15zdnd11an1n64x5 FILLER_78_2069 ();
 b15zdnd11an1n16x5 FILLER_78_2133 ();
 b15zdnd11an1n04x5 FILLER_78_2149 ();
 b15zdnd00an1n01x5 FILLER_78_2153 ();
 b15zdnd11an1n64x5 FILLER_78_2162 ();
 b15zdnd11an1n32x5 FILLER_78_2226 ();
 b15zdnd11an1n16x5 FILLER_78_2258 ();
 b15zdnd00an1n02x5 FILLER_78_2274 ();
 b15zdnd11an1n16x5 FILLER_79_0 ();
 b15zdnd11an1n08x5 FILLER_79_16 ();
 b15zdnd11an1n04x5 FILLER_79_24 ();
 b15zdnd00an1n01x5 FILLER_79_28 ();
 b15zdnd11an1n64x5 FILLER_79_34 ();
 b15zdnd11an1n64x5 FILLER_79_98 ();
 b15zdnd11an1n64x5 FILLER_79_162 ();
 b15zdnd11an1n64x5 FILLER_79_226 ();
 b15zdnd11an1n64x5 FILLER_79_290 ();
 b15zdnd11an1n08x5 FILLER_79_354 ();
 b15zdnd11an1n04x5 FILLER_79_362 ();
 b15zdnd11an1n64x5 FILLER_79_369 ();
 b15zdnd11an1n64x5 FILLER_79_433 ();
 b15zdnd11an1n64x5 FILLER_79_497 ();
 b15zdnd11an1n64x5 FILLER_79_561 ();
 b15zdnd11an1n08x5 FILLER_79_625 ();
 b15zdnd11an1n04x5 FILLER_79_633 ();
 b15zdnd00an1n01x5 FILLER_79_637 ();
 b15zdnd11an1n04x5 FILLER_79_641 ();
 b15zdnd11an1n04x5 FILLER_79_653 ();
 b15zdnd00an1n01x5 FILLER_79_657 ();
 b15zdnd11an1n04x5 FILLER_79_665 ();
 b15zdnd00an1n02x5 FILLER_79_669 ();
 b15zdnd11an1n64x5 FILLER_79_691 ();
 b15zdnd11an1n64x5 FILLER_79_755 ();
 b15zdnd11an1n64x5 FILLER_79_819 ();
 b15zdnd11an1n16x5 FILLER_79_883 ();
 b15zdnd11an1n04x5 FILLER_79_899 ();
 b15zdnd00an1n02x5 FILLER_79_903 ();
 b15zdnd00an1n01x5 FILLER_79_905 ();
 b15zdnd11an1n64x5 FILLER_79_915 ();
 b15zdnd11an1n64x5 FILLER_79_979 ();
 b15zdnd11an1n32x5 FILLER_79_1043 ();
 b15zdnd00an1n02x5 FILLER_79_1075 ();
 b15zdnd00an1n01x5 FILLER_79_1077 ();
 b15zdnd11an1n04x5 FILLER_79_1081 ();
 b15zdnd11an1n64x5 FILLER_79_1088 ();
 b15zdnd11an1n64x5 FILLER_79_1152 ();
 b15zdnd11an1n64x5 FILLER_79_1216 ();
 b15zdnd11an1n64x5 FILLER_79_1280 ();
 b15zdnd11an1n64x5 FILLER_79_1344 ();
 b15zdnd11an1n32x5 FILLER_79_1408 ();
 b15zdnd00an1n01x5 FILLER_79_1440 ();
 b15zdnd11an1n04x5 FILLER_79_1480 ();
 b15zdnd11an1n64x5 FILLER_79_1489 ();
 b15zdnd11an1n64x5 FILLER_79_1553 ();
 b15zdnd11an1n16x5 FILLER_79_1617 ();
 b15zdnd00an1n02x5 FILLER_79_1633 ();
 b15zdnd00an1n01x5 FILLER_79_1635 ();
 b15zdnd11an1n64x5 FILLER_79_1640 ();
 b15zdnd11an1n08x5 FILLER_79_1704 ();
 b15zdnd11an1n04x5 FILLER_79_1712 ();
 b15zdnd11an1n08x5 FILLER_79_1723 ();
 b15zdnd11an1n64x5 FILLER_79_1773 ();
 b15zdnd11an1n08x5 FILLER_79_1837 ();
 b15zdnd11an1n64x5 FILLER_79_1855 ();
 b15zdnd11an1n64x5 FILLER_79_1919 ();
 b15zdnd11an1n64x5 FILLER_79_1983 ();
 b15zdnd11an1n64x5 FILLER_79_2047 ();
 b15zdnd11an1n64x5 FILLER_79_2111 ();
 b15zdnd11an1n64x5 FILLER_79_2175 ();
 b15zdnd11an1n32x5 FILLER_79_2239 ();
 b15zdnd11an1n08x5 FILLER_79_2271 ();
 b15zdnd11an1n04x5 FILLER_79_2279 ();
 b15zdnd00an1n01x5 FILLER_79_2283 ();
 b15zdnd11an1n64x5 FILLER_80_8 ();
 b15zdnd11an1n64x5 FILLER_80_72 ();
 b15zdnd11an1n64x5 FILLER_80_136 ();
 b15zdnd11an1n64x5 FILLER_80_200 ();
 b15zdnd11an1n32x5 FILLER_80_264 ();
 b15zdnd11an1n16x5 FILLER_80_296 ();
 b15zdnd11an1n08x5 FILLER_80_312 ();
 b15zdnd00an1n01x5 FILLER_80_320 ();
 b15zdnd11an1n08x5 FILLER_80_363 ();
 b15zdnd00an1n02x5 FILLER_80_371 ();
 b15zdnd11an1n64x5 FILLER_80_376 ();
 b15zdnd11an1n64x5 FILLER_80_440 ();
 b15zdnd11an1n64x5 FILLER_80_504 ();
 b15zdnd11an1n64x5 FILLER_80_568 ();
 b15zdnd11an1n64x5 FILLER_80_632 ();
 b15zdnd11an1n16x5 FILLER_80_696 ();
 b15zdnd11an1n04x5 FILLER_80_712 ();
 b15zdnd00an1n02x5 FILLER_80_716 ();
 b15zdnd11an1n64x5 FILLER_80_726 ();
 b15zdnd11an1n64x5 FILLER_80_790 ();
 b15zdnd11an1n64x5 FILLER_80_854 ();
 b15zdnd11an1n64x5 FILLER_80_918 ();
 b15zdnd11an1n64x5 FILLER_80_982 ();
 b15zdnd11an1n64x5 FILLER_80_1046 ();
 b15zdnd11an1n16x5 FILLER_80_1110 ();
 b15zdnd11an1n08x5 FILLER_80_1126 ();
 b15zdnd11an1n04x5 FILLER_80_1134 ();
 b15zdnd00an1n02x5 FILLER_80_1138 ();
 b15zdnd11an1n64x5 FILLER_80_1162 ();
 b15zdnd11an1n64x5 FILLER_80_1226 ();
 b15zdnd11an1n32x5 FILLER_80_1290 ();
 b15zdnd11an1n16x5 FILLER_80_1322 ();
 b15zdnd11an1n08x5 FILLER_80_1338 ();
 b15zdnd00an1n02x5 FILLER_80_1346 ();
 b15zdnd11an1n64x5 FILLER_80_1390 ();
 b15zdnd11an1n04x5 FILLER_80_1454 ();
 b15zdnd00an1n02x5 FILLER_80_1458 ();
 b15zdnd11an1n16x5 FILLER_80_1468 ();
 b15zdnd11an1n08x5 FILLER_80_1484 ();
 b15zdnd11an1n04x5 FILLER_80_1495 ();
 b15zdnd11an1n08x5 FILLER_80_1502 ();
 b15zdnd00an1n02x5 FILLER_80_1510 ();
 b15zdnd11an1n64x5 FILLER_80_1515 ();
 b15zdnd11an1n16x5 FILLER_80_1579 ();
 b15zdnd11an1n08x5 FILLER_80_1595 ();
 b15zdnd11an1n04x5 FILLER_80_1603 ();
 b15zdnd00an1n01x5 FILLER_80_1607 ();
 b15zdnd11an1n04x5 FILLER_80_1614 ();
 b15zdnd11an1n32x5 FILLER_80_1658 ();
 b15zdnd11an1n16x5 FILLER_80_1690 ();
 b15zdnd11an1n08x5 FILLER_80_1706 ();
 b15zdnd00an1n02x5 FILLER_80_1714 ();
 b15zdnd00an1n01x5 FILLER_80_1716 ();
 b15zdnd11an1n04x5 FILLER_80_1722 ();
 b15zdnd11an1n64x5 FILLER_80_1768 ();
 b15zdnd11an1n64x5 FILLER_80_1832 ();
 b15zdnd11an1n64x5 FILLER_80_1896 ();
 b15zdnd11an1n32x5 FILLER_80_1960 ();
 b15zdnd11an1n08x5 FILLER_80_1992 ();
 b15zdnd11an1n04x5 FILLER_80_2000 ();
 b15zdnd11an1n64x5 FILLER_80_2008 ();
 b15zdnd11an1n64x5 FILLER_80_2072 ();
 b15zdnd11an1n16x5 FILLER_80_2136 ();
 b15zdnd00an1n02x5 FILLER_80_2152 ();
 b15zdnd11an1n64x5 FILLER_80_2162 ();
 b15zdnd11an1n32x5 FILLER_80_2226 ();
 b15zdnd11an1n16x5 FILLER_80_2258 ();
 b15zdnd00an1n02x5 FILLER_80_2274 ();
 b15zdnd11an1n64x5 FILLER_81_0 ();
 b15zdnd11an1n64x5 FILLER_81_64 ();
 b15zdnd11an1n64x5 FILLER_81_128 ();
 b15zdnd11an1n64x5 FILLER_81_192 ();
 b15zdnd11an1n64x5 FILLER_81_256 ();
 b15zdnd11an1n08x5 FILLER_81_320 ();
 b15zdnd11an1n04x5 FILLER_81_328 ();
 b15zdnd00an1n02x5 FILLER_81_332 ();
 b15zdnd11an1n04x5 FILLER_81_374 ();
 b15zdnd11an1n16x5 FILLER_81_381 ();
 b15zdnd11an1n64x5 FILLER_81_422 ();
 b15zdnd11an1n64x5 FILLER_81_486 ();
 b15zdnd11an1n64x5 FILLER_81_550 ();
 b15zdnd11an1n64x5 FILLER_81_614 ();
 b15zdnd11an1n64x5 FILLER_81_678 ();
 b15zdnd11an1n64x5 FILLER_81_742 ();
 b15zdnd11an1n64x5 FILLER_81_806 ();
 b15zdnd11an1n64x5 FILLER_81_870 ();
 b15zdnd11an1n64x5 FILLER_81_934 ();
 b15zdnd11an1n64x5 FILLER_81_998 ();
 b15zdnd11an1n64x5 FILLER_81_1062 ();
 b15zdnd11an1n64x5 FILLER_81_1126 ();
 b15zdnd11an1n64x5 FILLER_81_1190 ();
 b15zdnd11an1n64x5 FILLER_81_1254 ();
 b15zdnd11an1n64x5 FILLER_81_1318 ();
 b15zdnd11an1n64x5 FILLER_81_1382 ();
 b15zdnd11an1n08x5 FILLER_81_1446 ();
 b15zdnd11an1n04x5 FILLER_81_1454 ();
 b15zdnd00an1n02x5 FILLER_81_1458 ();
 b15zdnd11an1n08x5 FILLER_81_1500 ();
 b15zdnd00an1n02x5 FILLER_81_1508 ();
 b15zdnd00an1n01x5 FILLER_81_1510 ();
 b15zdnd11an1n64x5 FILLER_81_1514 ();
 b15zdnd11an1n08x5 FILLER_81_1578 ();
 b15zdnd00an1n01x5 FILLER_81_1586 ();
 b15zdnd11an1n04x5 FILLER_81_1614 ();
 b15zdnd11an1n04x5 FILLER_81_1660 ();
 b15zdnd11an1n32x5 FILLER_81_1667 ();
 b15zdnd11an1n04x5 FILLER_81_1699 ();
 b15zdnd00an1n02x5 FILLER_81_1703 ();
 b15zdnd11an1n08x5 FILLER_81_1709 ();
 b15zdnd11an1n08x5 FILLER_81_1730 ();
 b15zdnd11an1n04x5 FILLER_81_1738 ();
 b15zdnd00an1n02x5 FILLER_81_1742 ();
 b15zdnd11an1n64x5 FILLER_81_1786 ();
 b15zdnd00an1n02x5 FILLER_81_1850 ();
 b15zdnd11an1n64x5 FILLER_81_1894 ();
 b15zdnd11an1n64x5 FILLER_81_1958 ();
 b15zdnd11an1n64x5 FILLER_81_2022 ();
 b15zdnd11an1n64x5 FILLER_81_2086 ();
 b15zdnd11an1n64x5 FILLER_81_2150 ();
 b15zdnd11an1n64x5 FILLER_81_2214 ();
 b15zdnd11an1n04x5 FILLER_81_2278 ();
 b15zdnd00an1n02x5 FILLER_81_2282 ();
 b15zdnd11an1n64x5 FILLER_82_8 ();
 b15zdnd11an1n64x5 FILLER_82_72 ();
 b15zdnd11an1n64x5 FILLER_82_136 ();
 b15zdnd11an1n64x5 FILLER_82_200 ();
 b15zdnd11an1n64x5 FILLER_82_264 ();
 b15zdnd11an1n16x5 FILLER_82_328 ();
 b15zdnd11an1n08x5 FILLER_82_344 ();
 b15zdnd00an1n02x5 FILLER_82_352 ();
 b15zdnd00an1n01x5 FILLER_82_354 ();
 b15zdnd11an1n04x5 FILLER_82_407 ();
 b15zdnd11an1n16x5 FILLER_82_453 ();
 b15zdnd11an1n04x5 FILLER_82_469 ();
 b15zdnd00an1n02x5 FILLER_82_473 ();
 b15zdnd11an1n64x5 FILLER_82_483 ();
 b15zdnd11an1n64x5 FILLER_82_547 ();
 b15zdnd11an1n64x5 FILLER_82_611 ();
 b15zdnd11an1n32x5 FILLER_82_675 ();
 b15zdnd11an1n08x5 FILLER_82_707 ();
 b15zdnd00an1n02x5 FILLER_82_715 ();
 b15zdnd00an1n01x5 FILLER_82_717 ();
 b15zdnd11an1n64x5 FILLER_82_726 ();
 b15zdnd11an1n64x5 FILLER_82_790 ();
 b15zdnd11an1n64x5 FILLER_82_854 ();
 b15zdnd11an1n64x5 FILLER_82_918 ();
 b15zdnd11an1n64x5 FILLER_82_982 ();
 b15zdnd11an1n64x5 FILLER_82_1046 ();
 b15zdnd11an1n64x5 FILLER_82_1110 ();
 b15zdnd11an1n64x5 FILLER_82_1174 ();
 b15zdnd11an1n64x5 FILLER_82_1238 ();
 b15zdnd00an1n01x5 FILLER_82_1302 ();
 b15zdnd11an1n64x5 FILLER_82_1315 ();
 b15zdnd11an1n64x5 FILLER_82_1379 ();
 b15zdnd11an1n32x5 FILLER_82_1443 ();
 b15zdnd11an1n08x5 FILLER_82_1475 ();
 b15zdnd11an1n04x5 FILLER_82_1483 ();
 b15zdnd11an1n32x5 FILLER_82_1539 ();
 b15zdnd11an1n08x5 FILLER_82_1571 ();
 b15zdnd00an1n02x5 FILLER_82_1579 ();
 b15zdnd00an1n01x5 FILLER_82_1581 ();
 b15zdnd11an1n64x5 FILLER_82_1588 ();
 b15zdnd00an1n02x5 FILLER_82_1652 ();
 b15zdnd00an1n01x5 FILLER_82_1654 ();
 b15zdnd11an1n32x5 FILLER_82_1658 ();
 b15zdnd11an1n08x5 FILLER_82_1690 ();
 b15zdnd11an1n04x5 FILLER_82_1698 ();
 b15zdnd00an1n02x5 FILLER_82_1702 ();
 b15zdnd11an1n04x5 FILLER_82_1709 ();
 b15zdnd11an1n08x5 FILLER_82_1726 ();
 b15zdnd11an1n04x5 FILLER_82_1741 ();
 b15zdnd11an1n64x5 FILLER_82_1748 ();
 b15zdnd11an1n16x5 FILLER_82_1812 ();
 b15zdnd11an1n64x5 FILLER_82_1870 ();
 b15zdnd11an1n64x5 FILLER_82_1934 ();
 b15zdnd11an1n16x5 FILLER_82_1998 ();
 b15zdnd11an1n08x5 FILLER_82_2014 ();
 b15zdnd11an1n64x5 FILLER_82_2025 ();
 b15zdnd11an1n64x5 FILLER_82_2089 ();
 b15zdnd00an1n01x5 FILLER_82_2153 ();
 b15zdnd11an1n64x5 FILLER_82_2162 ();
 b15zdnd11an1n32x5 FILLER_82_2226 ();
 b15zdnd11an1n16x5 FILLER_82_2258 ();
 b15zdnd00an1n02x5 FILLER_82_2274 ();
 b15zdnd11an1n64x5 FILLER_83_0 ();
 b15zdnd11an1n64x5 FILLER_83_64 ();
 b15zdnd11an1n64x5 FILLER_83_128 ();
 b15zdnd11an1n64x5 FILLER_83_192 ();
 b15zdnd11an1n64x5 FILLER_83_256 ();
 b15zdnd11an1n32x5 FILLER_83_320 ();
 b15zdnd11an1n16x5 FILLER_83_352 ();
 b15zdnd11an1n04x5 FILLER_83_368 ();
 b15zdnd00an1n02x5 FILLER_83_372 ();
 b15zdnd11an1n04x5 FILLER_83_377 ();
 b15zdnd11an1n64x5 FILLER_83_384 ();
 b15zdnd11an1n64x5 FILLER_83_448 ();
 b15zdnd11an1n64x5 FILLER_83_512 ();
 b15zdnd11an1n64x5 FILLER_83_576 ();
 b15zdnd11an1n64x5 FILLER_83_640 ();
 b15zdnd11an1n64x5 FILLER_83_704 ();
 b15zdnd11an1n64x5 FILLER_83_768 ();
 b15zdnd11an1n64x5 FILLER_83_832 ();
 b15zdnd11an1n64x5 FILLER_83_896 ();
 b15zdnd11an1n64x5 FILLER_83_960 ();
 b15zdnd11an1n64x5 FILLER_83_1024 ();
 b15zdnd11an1n64x5 FILLER_83_1088 ();
 b15zdnd11an1n64x5 FILLER_83_1152 ();
 b15zdnd11an1n32x5 FILLER_83_1216 ();
 b15zdnd11an1n16x5 FILLER_83_1248 ();
 b15zdnd11an1n08x5 FILLER_83_1264 ();
 b15zdnd11an1n64x5 FILLER_83_1283 ();
 b15zdnd11an1n64x5 FILLER_83_1347 ();
 b15zdnd11an1n32x5 FILLER_83_1411 ();
 b15zdnd11an1n16x5 FILLER_83_1443 ();
 b15zdnd00an1n01x5 FILLER_83_1459 ();
 b15zdnd11an1n32x5 FILLER_83_1471 ();
 b15zdnd11an1n08x5 FILLER_83_1503 ();
 b15zdnd00an1n01x5 FILLER_83_1511 ();
 b15zdnd11an1n16x5 FILLER_83_1515 ();
 b15zdnd11an1n04x5 FILLER_83_1531 ();
 b15zdnd00an1n01x5 FILLER_83_1535 ();
 b15zdnd11an1n04x5 FILLER_83_1578 ();
 b15zdnd11an1n04x5 FILLER_83_1585 ();
 b15zdnd11an1n32x5 FILLER_83_1592 ();
 b15zdnd11an1n16x5 FILLER_83_1624 ();
 b15zdnd11an1n08x5 FILLER_83_1640 ();
 b15zdnd11an1n04x5 FILLER_83_1648 ();
 b15zdnd00an1n02x5 FILLER_83_1652 ();
 b15zdnd11an1n64x5 FILLER_83_1696 ();
 b15zdnd11an1n64x5 FILLER_83_1760 ();
 b15zdnd11an1n64x5 FILLER_83_1824 ();
 b15zdnd11an1n64x5 FILLER_83_1888 ();
 b15zdnd11an1n32x5 FILLER_83_1952 ();
 b15zdnd11an1n16x5 FILLER_83_1984 ();
 b15zdnd00an1n02x5 FILLER_83_2000 ();
 b15zdnd11an1n04x5 FILLER_83_2044 ();
 b15zdnd11an1n64x5 FILLER_83_2066 ();
 b15zdnd11an1n64x5 FILLER_83_2130 ();
 b15zdnd11an1n64x5 FILLER_83_2194 ();
 b15zdnd11an1n16x5 FILLER_83_2258 ();
 b15zdnd11an1n08x5 FILLER_83_2274 ();
 b15zdnd00an1n02x5 FILLER_83_2282 ();
 b15zdnd11an1n64x5 FILLER_84_8 ();
 b15zdnd11an1n64x5 FILLER_84_72 ();
 b15zdnd11an1n64x5 FILLER_84_136 ();
 b15zdnd11an1n64x5 FILLER_84_200 ();
 b15zdnd11an1n64x5 FILLER_84_264 ();
 b15zdnd11an1n64x5 FILLER_84_328 ();
 b15zdnd11an1n64x5 FILLER_84_392 ();
 b15zdnd11an1n04x5 FILLER_84_456 ();
 b15zdnd11an1n64x5 FILLER_84_487 ();
 b15zdnd11an1n64x5 FILLER_84_551 ();
 b15zdnd11an1n64x5 FILLER_84_615 ();
 b15zdnd11an1n32x5 FILLER_84_679 ();
 b15zdnd11an1n04x5 FILLER_84_711 ();
 b15zdnd00an1n02x5 FILLER_84_715 ();
 b15zdnd00an1n01x5 FILLER_84_717 ();
 b15zdnd11an1n04x5 FILLER_84_726 ();
 b15zdnd00an1n01x5 FILLER_84_730 ();
 b15zdnd11an1n08x5 FILLER_84_739 ();
 b15zdnd11an1n04x5 FILLER_84_747 ();
 b15zdnd00an1n02x5 FILLER_84_751 ();
 b15zdnd00an1n01x5 FILLER_84_753 ();
 b15zdnd11an1n64x5 FILLER_84_780 ();
 b15zdnd11an1n64x5 FILLER_84_844 ();
 b15zdnd00an1n02x5 FILLER_84_908 ();
 b15zdnd00an1n01x5 FILLER_84_910 ();
 b15zdnd11an1n04x5 FILLER_84_919 ();
 b15zdnd11an1n64x5 FILLER_84_931 ();
 b15zdnd11an1n64x5 FILLER_84_995 ();
 b15zdnd11an1n64x5 FILLER_84_1059 ();
 b15zdnd11an1n64x5 FILLER_84_1123 ();
 b15zdnd11an1n64x5 FILLER_84_1187 ();
 b15zdnd11an1n64x5 FILLER_84_1251 ();
 b15zdnd11an1n64x5 FILLER_84_1315 ();
 b15zdnd11an1n64x5 FILLER_84_1379 ();
 b15zdnd11an1n64x5 FILLER_84_1443 ();
 b15zdnd11an1n32x5 FILLER_84_1507 ();
 b15zdnd11an1n16x5 FILLER_84_1539 ();
 b15zdnd11an1n08x5 FILLER_84_1555 ();
 b15zdnd11an1n64x5 FILLER_84_1615 ();
 b15zdnd11an1n64x5 FILLER_84_1679 ();
 b15zdnd11an1n64x5 FILLER_84_1743 ();
 b15zdnd11an1n64x5 FILLER_84_1807 ();
 b15zdnd11an1n64x5 FILLER_84_1871 ();
 b15zdnd11an1n32x5 FILLER_84_1935 ();
 b15zdnd11an1n16x5 FILLER_84_1967 ();
 b15zdnd11an1n08x5 FILLER_84_1983 ();
 b15zdnd11an1n04x5 FILLER_84_1991 ();
 b15zdnd00an1n01x5 FILLER_84_1995 ();
 b15zdnd11an1n04x5 FILLER_84_2048 ();
 b15zdnd11an1n32x5 FILLER_84_2094 ();
 b15zdnd11an1n16x5 FILLER_84_2126 ();
 b15zdnd11an1n08x5 FILLER_84_2142 ();
 b15zdnd11an1n04x5 FILLER_84_2150 ();
 b15zdnd11an1n64x5 FILLER_84_2162 ();
 b15zdnd11an1n32x5 FILLER_84_2226 ();
 b15zdnd11an1n16x5 FILLER_84_2258 ();
 b15zdnd00an1n02x5 FILLER_84_2274 ();
 b15zdnd11an1n64x5 FILLER_85_0 ();
 b15zdnd11an1n64x5 FILLER_85_64 ();
 b15zdnd11an1n64x5 FILLER_85_128 ();
 b15zdnd11an1n64x5 FILLER_85_192 ();
 b15zdnd11an1n64x5 FILLER_85_256 ();
 b15zdnd11an1n64x5 FILLER_85_320 ();
 b15zdnd11an1n64x5 FILLER_85_384 ();
 b15zdnd11an1n64x5 FILLER_85_448 ();
 b15zdnd11an1n64x5 FILLER_85_512 ();
 b15zdnd11an1n64x5 FILLER_85_576 ();
 b15zdnd11an1n64x5 FILLER_85_640 ();
 b15zdnd11an1n64x5 FILLER_85_704 ();
 b15zdnd11an1n64x5 FILLER_85_768 ();
 b15zdnd11an1n64x5 FILLER_85_832 ();
 b15zdnd11an1n64x5 FILLER_85_896 ();
 b15zdnd11an1n64x5 FILLER_85_960 ();
 b15zdnd11an1n64x5 FILLER_85_1024 ();
 b15zdnd11an1n64x5 FILLER_85_1088 ();
 b15zdnd11an1n64x5 FILLER_85_1152 ();
 b15zdnd11an1n64x5 FILLER_85_1216 ();
 b15zdnd11an1n64x5 FILLER_85_1280 ();
 b15zdnd11an1n64x5 FILLER_85_1344 ();
 b15zdnd11an1n64x5 FILLER_85_1408 ();
 b15zdnd11an1n64x5 FILLER_85_1472 ();
 b15zdnd11an1n16x5 FILLER_85_1536 ();
 b15zdnd11an1n08x5 FILLER_85_1552 ();
 b15zdnd11an1n64x5 FILLER_85_1602 ();
 b15zdnd11an1n64x5 FILLER_85_1666 ();
 b15zdnd11an1n64x5 FILLER_85_1730 ();
 b15zdnd11an1n64x5 FILLER_85_1794 ();
 b15zdnd11an1n64x5 FILLER_85_1858 ();
 b15zdnd11an1n64x5 FILLER_85_1922 ();
 b15zdnd11an1n32x5 FILLER_85_1986 ();
 b15zdnd00an1n02x5 FILLER_85_2018 ();
 b15zdnd00an1n01x5 FILLER_85_2020 ();
 b15zdnd11an1n64x5 FILLER_85_2024 ();
 b15zdnd11an1n64x5 FILLER_85_2088 ();
 b15zdnd11an1n64x5 FILLER_85_2152 ();
 b15zdnd11an1n64x5 FILLER_85_2216 ();
 b15zdnd11an1n04x5 FILLER_85_2280 ();
 b15zdnd11an1n64x5 FILLER_86_8 ();
 b15zdnd11an1n64x5 FILLER_86_72 ();
 b15zdnd11an1n64x5 FILLER_86_136 ();
 b15zdnd11an1n64x5 FILLER_86_200 ();
 b15zdnd11an1n64x5 FILLER_86_264 ();
 b15zdnd11an1n32x5 FILLER_86_328 ();
 b15zdnd11an1n16x5 FILLER_86_360 ();
 b15zdnd11an1n08x5 FILLER_86_376 ();
 b15zdnd11an1n04x5 FILLER_86_384 ();
 b15zdnd00an1n02x5 FILLER_86_388 ();
 b15zdnd11an1n64x5 FILLER_86_394 ();
 b15zdnd11an1n32x5 FILLER_86_458 ();
 b15zdnd11an1n16x5 FILLER_86_490 ();
 b15zdnd00an1n01x5 FILLER_86_506 ();
 b15zdnd11an1n64x5 FILLER_86_510 ();
 b15zdnd11an1n64x5 FILLER_86_574 ();
 b15zdnd11an1n64x5 FILLER_86_638 ();
 b15zdnd11an1n16x5 FILLER_86_702 ();
 b15zdnd11an1n64x5 FILLER_86_726 ();
 b15zdnd11an1n64x5 FILLER_86_790 ();
 b15zdnd11an1n64x5 FILLER_86_854 ();
 b15zdnd11an1n64x5 FILLER_86_918 ();
 b15zdnd11an1n64x5 FILLER_86_982 ();
 b15zdnd11an1n64x5 FILLER_86_1046 ();
 b15zdnd11an1n64x5 FILLER_86_1110 ();
 b15zdnd11an1n64x5 FILLER_86_1174 ();
 b15zdnd11an1n16x5 FILLER_86_1238 ();
 b15zdnd11an1n04x5 FILLER_86_1254 ();
 b15zdnd00an1n02x5 FILLER_86_1258 ();
 b15zdnd00an1n01x5 FILLER_86_1260 ();
 b15zdnd11an1n64x5 FILLER_86_1279 ();
 b15zdnd11an1n64x5 FILLER_86_1343 ();
 b15zdnd11an1n64x5 FILLER_86_1407 ();
 b15zdnd11an1n64x5 FILLER_86_1471 ();
 b15zdnd11an1n32x5 FILLER_86_1535 ();
 b15zdnd11an1n16x5 FILLER_86_1567 ();
 b15zdnd11an1n04x5 FILLER_86_1583 ();
 b15zdnd00an1n01x5 FILLER_86_1587 ();
 b15zdnd11an1n64x5 FILLER_86_1591 ();
 b15zdnd11an1n64x5 FILLER_86_1655 ();
 b15zdnd11an1n64x5 FILLER_86_1719 ();
 b15zdnd11an1n64x5 FILLER_86_1783 ();
 b15zdnd11an1n32x5 FILLER_86_1847 ();
 b15zdnd11an1n16x5 FILLER_86_1879 ();
 b15zdnd11an1n04x5 FILLER_86_1898 ();
 b15zdnd11an1n64x5 FILLER_86_1905 ();
 b15zdnd11an1n32x5 FILLER_86_1969 ();
 b15zdnd11an1n16x5 FILLER_86_2001 ();
 b15zdnd11an1n04x5 FILLER_86_2017 ();
 b15zdnd11an1n64x5 FILLER_86_2024 ();
 b15zdnd11an1n64x5 FILLER_86_2088 ();
 b15zdnd00an1n02x5 FILLER_86_2152 ();
 b15zdnd11an1n64x5 FILLER_86_2162 ();
 b15zdnd11an1n32x5 FILLER_86_2226 ();
 b15zdnd11an1n16x5 FILLER_86_2258 ();
 b15zdnd00an1n02x5 FILLER_86_2274 ();
 b15zdnd11an1n64x5 FILLER_87_0 ();
 b15zdnd11an1n64x5 FILLER_87_64 ();
 b15zdnd11an1n64x5 FILLER_87_128 ();
 b15zdnd11an1n64x5 FILLER_87_192 ();
 b15zdnd11an1n64x5 FILLER_87_256 ();
 b15zdnd11an1n64x5 FILLER_87_320 ();
 b15zdnd11an1n64x5 FILLER_87_384 ();
 b15zdnd11an1n32x5 FILLER_87_448 ();
 b15zdnd11an1n64x5 FILLER_87_532 ();
 b15zdnd11an1n64x5 FILLER_87_596 ();
 b15zdnd11an1n64x5 FILLER_87_660 ();
 b15zdnd11an1n64x5 FILLER_87_724 ();
 b15zdnd11an1n64x5 FILLER_87_788 ();
 b15zdnd11an1n64x5 FILLER_87_852 ();
 b15zdnd11an1n64x5 FILLER_87_916 ();
 b15zdnd11an1n64x5 FILLER_87_980 ();
 b15zdnd11an1n64x5 FILLER_87_1044 ();
 b15zdnd11an1n64x5 FILLER_87_1108 ();
 b15zdnd11an1n08x5 FILLER_87_1172 ();
 b15zdnd00an1n02x5 FILLER_87_1180 ();
 b15zdnd00an1n01x5 FILLER_87_1182 ();
 b15zdnd11an1n32x5 FILLER_87_1197 ();
 b15zdnd11an1n16x5 FILLER_87_1229 ();
 b15zdnd11an1n08x5 FILLER_87_1245 ();
 b15zdnd11an1n04x5 FILLER_87_1253 ();
 b15zdnd11an1n64x5 FILLER_87_1264 ();
 b15zdnd11an1n64x5 FILLER_87_1328 ();
 b15zdnd11an1n64x5 FILLER_87_1392 ();
 b15zdnd11an1n64x5 FILLER_87_1456 ();
 b15zdnd11an1n64x5 FILLER_87_1520 ();
 b15zdnd11an1n64x5 FILLER_87_1584 ();
 b15zdnd11an1n64x5 FILLER_87_1648 ();
 b15zdnd11an1n64x5 FILLER_87_1712 ();
 b15zdnd11an1n64x5 FILLER_87_1776 ();
 b15zdnd11an1n16x5 FILLER_87_1840 ();
 b15zdnd11an1n08x5 FILLER_87_1856 ();
 b15zdnd11an1n64x5 FILLER_87_1904 ();
 b15zdnd11an1n64x5 FILLER_87_1968 ();
 b15zdnd11an1n64x5 FILLER_87_2032 ();
 b15zdnd11an1n64x5 FILLER_87_2096 ();
 b15zdnd11an1n64x5 FILLER_87_2160 ();
 b15zdnd11an1n32x5 FILLER_87_2224 ();
 b15zdnd11an1n16x5 FILLER_87_2256 ();
 b15zdnd11an1n08x5 FILLER_87_2272 ();
 b15zdnd11an1n04x5 FILLER_87_2280 ();
 b15zdnd11an1n64x5 FILLER_88_8 ();
 b15zdnd11an1n64x5 FILLER_88_72 ();
 b15zdnd11an1n64x5 FILLER_88_136 ();
 b15zdnd11an1n64x5 FILLER_88_200 ();
 b15zdnd11an1n64x5 FILLER_88_264 ();
 b15zdnd11an1n64x5 FILLER_88_328 ();
 b15zdnd11an1n64x5 FILLER_88_392 ();
 b15zdnd11an1n32x5 FILLER_88_456 ();
 b15zdnd11an1n08x5 FILLER_88_488 ();
 b15zdnd00an1n02x5 FILLER_88_496 ();
 b15zdnd11an1n04x5 FILLER_88_501 ();
 b15zdnd11an1n64x5 FILLER_88_508 ();
 b15zdnd11an1n64x5 FILLER_88_572 ();
 b15zdnd11an1n64x5 FILLER_88_636 ();
 b15zdnd11an1n16x5 FILLER_88_700 ();
 b15zdnd00an1n02x5 FILLER_88_716 ();
 b15zdnd11an1n64x5 FILLER_88_726 ();
 b15zdnd11an1n64x5 FILLER_88_790 ();
 b15zdnd11an1n64x5 FILLER_88_854 ();
 b15zdnd11an1n64x5 FILLER_88_918 ();
 b15zdnd11an1n64x5 FILLER_88_982 ();
 b15zdnd11an1n32x5 FILLER_88_1046 ();
 b15zdnd00an1n01x5 FILLER_88_1078 ();
 b15zdnd11an1n64x5 FILLER_88_1083 ();
 b15zdnd11an1n64x5 FILLER_88_1147 ();
 b15zdnd11an1n64x5 FILLER_88_1211 ();
 b15zdnd11an1n64x5 FILLER_88_1275 ();
 b15zdnd11an1n64x5 FILLER_88_1339 ();
 b15zdnd11an1n64x5 FILLER_88_1403 ();
 b15zdnd11an1n64x5 FILLER_88_1467 ();
 b15zdnd11an1n64x5 FILLER_88_1531 ();
 b15zdnd11an1n64x5 FILLER_88_1595 ();
 b15zdnd11an1n64x5 FILLER_88_1659 ();
 b15zdnd11an1n08x5 FILLER_88_1723 ();
 b15zdnd11an1n04x5 FILLER_88_1731 ();
 b15zdnd00an1n01x5 FILLER_88_1735 ();
 b15zdnd11an1n64x5 FILLER_88_1741 ();
 b15zdnd11an1n64x5 FILLER_88_1805 ();
 b15zdnd11an1n64x5 FILLER_88_1869 ();
 b15zdnd11an1n64x5 FILLER_88_1933 ();
 b15zdnd11an1n64x5 FILLER_88_1997 ();
 b15zdnd11an1n64x5 FILLER_88_2061 ();
 b15zdnd11an1n16x5 FILLER_88_2125 ();
 b15zdnd11an1n08x5 FILLER_88_2141 ();
 b15zdnd11an1n04x5 FILLER_88_2149 ();
 b15zdnd00an1n01x5 FILLER_88_2153 ();
 b15zdnd11an1n64x5 FILLER_88_2162 ();
 b15zdnd11an1n32x5 FILLER_88_2226 ();
 b15zdnd11an1n16x5 FILLER_88_2258 ();
 b15zdnd00an1n02x5 FILLER_88_2274 ();
 b15zdnd11an1n64x5 FILLER_89_0 ();
 b15zdnd11an1n64x5 FILLER_89_64 ();
 b15zdnd11an1n64x5 FILLER_89_128 ();
 b15zdnd11an1n64x5 FILLER_89_192 ();
 b15zdnd11an1n64x5 FILLER_89_256 ();
 b15zdnd11an1n64x5 FILLER_89_320 ();
 b15zdnd11an1n64x5 FILLER_89_384 ();
 b15zdnd11an1n64x5 FILLER_89_448 ();
 b15zdnd11an1n64x5 FILLER_89_512 ();
 b15zdnd11an1n64x5 FILLER_89_576 ();
 b15zdnd11an1n64x5 FILLER_89_640 ();
 b15zdnd11an1n64x5 FILLER_89_704 ();
 b15zdnd11an1n08x5 FILLER_89_768 ();
 b15zdnd11an1n04x5 FILLER_89_776 ();
 b15zdnd00an1n02x5 FILLER_89_780 ();
 b15zdnd00an1n01x5 FILLER_89_782 ();
 b15zdnd11an1n64x5 FILLER_89_787 ();
 b15zdnd11an1n64x5 FILLER_89_851 ();
 b15zdnd11an1n64x5 FILLER_89_915 ();
 b15zdnd11an1n64x5 FILLER_89_979 ();
 b15zdnd11an1n64x5 FILLER_89_1043 ();
 b15zdnd11an1n64x5 FILLER_89_1107 ();
 b15zdnd11an1n64x5 FILLER_89_1171 ();
 b15zdnd11an1n64x5 FILLER_89_1235 ();
 b15zdnd11an1n64x5 FILLER_89_1299 ();
 b15zdnd11an1n64x5 FILLER_89_1363 ();
 b15zdnd11an1n64x5 FILLER_89_1427 ();
 b15zdnd11an1n64x5 FILLER_89_1491 ();
 b15zdnd11an1n64x5 FILLER_89_1555 ();
 b15zdnd11an1n64x5 FILLER_89_1619 ();
 b15zdnd11an1n32x5 FILLER_89_1683 ();
 b15zdnd11an1n16x5 FILLER_89_1715 ();
 b15zdnd11an1n04x5 FILLER_89_1731 ();
 b15zdnd11an1n64x5 FILLER_89_1777 ();
 b15zdnd11an1n64x5 FILLER_89_1841 ();
 b15zdnd11an1n64x5 FILLER_89_1905 ();
 b15zdnd11an1n64x5 FILLER_89_1969 ();
 b15zdnd11an1n64x5 FILLER_89_2033 ();
 b15zdnd11an1n64x5 FILLER_89_2097 ();
 b15zdnd11an1n64x5 FILLER_89_2161 ();
 b15zdnd11an1n32x5 FILLER_89_2225 ();
 b15zdnd11an1n16x5 FILLER_89_2257 ();
 b15zdnd11an1n08x5 FILLER_89_2273 ();
 b15zdnd00an1n02x5 FILLER_89_2281 ();
 b15zdnd00an1n01x5 FILLER_89_2283 ();
 b15zdnd11an1n64x5 FILLER_90_8 ();
 b15zdnd11an1n64x5 FILLER_90_72 ();
 b15zdnd11an1n32x5 FILLER_90_136 ();
 b15zdnd11an1n16x5 FILLER_90_168 ();
 b15zdnd11an1n08x5 FILLER_90_184 ();
 b15zdnd11an1n64x5 FILLER_90_195 ();
 b15zdnd11an1n64x5 FILLER_90_259 ();
 b15zdnd11an1n32x5 FILLER_90_323 ();
 b15zdnd11an1n16x5 FILLER_90_355 ();
 b15zdnd11an1n08x5 FILLER_90_371 ();
 b15zdnd11an1n04x5 FILLER_90_379 ();
 b15zdnd11an1n32x5 FILLER_90_425 ();
 b15zdnd11an1n16x5 FILLER_90_457 ();
 b15zdnd11an1n08x5 FILLER_90_473 ();
 b15zdnd00an1n01x5 FILLER_90_481 ();
 b15zdnd11an1n64x5 FILLER_90_524 ();
 b15zdnd11an1n64x5 FILLER_90_588 ();
 b15zdnd11an1n64x5 FILLER_90_652 ();
 b15zdnd00an1n02x5 FILLER_90_716 ();
 b15zdnd11an1n16x5 FILLER_90_726 ();
 b15zdnd11an1n04x5 FILLER_90_742 ();
 b15zdnd00an1n02x5 FILLER_90_746 ();
 b15zdnd11an1n64x5 FILLER_90_754 ();
 b15zdnd11an1n64x5 FILLER_90_818 ();
 b15zdnd11an1n64x5 FILLER_90_882 ();
 b15zdnd11an1n64x5 FILLER_90_946 ();
 b15zdnd11an1n32x5 FILLER_90_1010 ();
 b15zdnd11an1n16x5 FILLER_90_1042 ();
 b15zdnd11an1n08x5 FILLER_90_1058 ();
 b15zdnd11an1n04x5 FILLER_90_1066 ();
 b15zdnd11an1n64x5 FILLER_90_1074 ();
 b15zdnd11an1n32x5 FILLER_90_1138 ();
 b15zdnd11an1n16x5 FILLER_90_1170 ();
 b15zdnd00an1n02x5 FILLER_90_1186 ();
 b15zdnd00an1n01x5 FILLER_90_1188 ();
 b15zdnd11an1n32x5 FILLER_90_1233 ();
 b15zdnd11an1n16x5 FILLER_90_1265 ();
 b15zdnd00an1n02x5 FILLER_90_1281 ();
 b15zdnd00an1n01x5 FILLER_90_1283 ();
 b15zdnd11an1n04x5 FILLER_90_1287 ();
 b15zdnd11an1n64x5 FILLER_90_1294 ();
 b15zdnd11an1n64x5 FILLER_90_1358 ();
 b15zdnd11an1n64x5 FILLER_90_1422 ();
 b15zdnd11an1n64x5 FILLER_90_1486 ();
 b15zdnd11an1n64x5 FILLER_90_1550 ();
 b15zdnd11an1n64x5 FILLER_90_1614 ();
 b15zdnd11an1n64x5 FILLER_90_1678 ();
 b15zdnd11an1n64x5 FILLER_90_1742 ();
 b15zdnd11an1n16x5 FILLER_90_1806 ();
 b15zdnd11an1n08x5 FILLER_90_1822 ();
 b15zdnd11an1n04x5 FILLER_90_1830 ();
 b15zdnd00an1n01x5 FILLER_90_1834 ();
 b15zdnd11an1n64x5 FILLER_90_1887 ();
 b15zdnd11an1n64x5 FILLER_90_1951 ();
 b15zdnd11an1n64x5 FILLER_90_2015 ();
 b15zdnd11an1n64x5 FILLER_90_2079 ();
 b15zdnd11an1n08x5 FILLER_90_2143 ();
 b15zdnd00an1n02x5 FILLER_90_2151 ();
 b15zdnd00an1n01x5 FILLER_90_2153 ();
 b15zdnd11an1n64x5 FILLER_90_2162 ();
 b15zdnd11an1n32x5 FILLER_90_2226 ();
 b15zdnd11an1n16x5 FILLER_90_2258 ();
 b15zdnd00an1n02x5 FILLER_90_2274 ();
 b15zdnd11an1n64x5 FILLER_91_0 ();
 b15zdnd11an1n64x5 FILLER_91_64 ();
 b15zdnd11an1n32x5 FILLER_91_128 ();
 b15zdnd11an1n16x5 FILLER_91_160 ();
 b15zdnd11an1n08x5 FILLER_91_176 ();
 b15zdnd00an1n02x5 FILLER_91_184 ();
 b15zdnd11an1n08x5 FILLER_91_189 ();
 b15zdnd00an1n02x5 FILLER_91_197 ();
 b15zdnd11an1n16x5 FILLER_91_206 ();
 b15zdnd11an1n04x5 FILLER_91_222 ();
 b15zdnd00an1n01x5 FILLER_91_226 ();
 b15zdnd11an1n64x5 FILLER_91_253 ();
 b15zdnd11an1n64x5 FILLER_91_317 ();
 b15zdnd11an1n64x5 FILLER_91_381 ();
 b15zdnd11an1n32x5 FILLER_91_445 ();
 b15zdnd00an1n01x5 FILLER_91_477 ();
 b15zdnd11an1n04x5 FILLER_91_509 ();
 b15zdnd00an1n01x5 FILLER_91_513 ();
 b15zdnd11an1n64x5 FILLER_91_517 ();
 b15zdnd11an1n64x5 FILLER_91_581 ();
 b15zdnd11an1n64x5 FILLER_91_645 ();
 b15zdnd11an1n32x5 FILLER_91_709 ();
 b15zdnd11an1n16x5 FILLER_91_741 ();
 b15zdnd00an1n01x5 FILLER_91_757 ();
 b15zdnd11an1n04x5 FILLER_91_764 ();
 b15zdnd00an1n01x5 FILLER_91_768 ();
 b15zdnd11an1n64x5 FILLER_91_773 ();
 b15zdnd11an1n64x5 FILLER_91_837 ();
 b15zdnd11an1n64x5 FILLER_91_901 ();
 b15zdnd11an1n64x5 FILLER_91_965 ();
 b15zdnd11an1n64x5 FILLER_91_1029 ();
 b15zdnd11an1n64x5 FILLER_91_1093 ();
 b15zdnd11an1n32x5 FILLER_91_1157 ();
 b15zdnd00an1n02x5 FILLER_91_1189 ();
 b15zdnd00an1n01x5 FILLER_91_1191 ();
 b15zdnd11an1n04x5 FILLER_91_1200 ();
 b15zdnd11an1n04x5 FILLER_91_1207 ();
 b15zdnd11an1n04x5 FILLER_91_1214 ();
 b15zdnd11an1n32x5 FILLER_91_1221 ();
 b15zdnd11an1n16x5 FILLER_91_1253 ();
 b15zdnd11an1n64x5 FILLER_91_1313 ();
 b15zdnd11an1n64x5 FILLER_91_1377 ();
 b15zdnd11an1n64x5 FILLER_91_1441 ();
 b15zdnd11an1n64x5 FILLER_91_1505 ();
 b15zdnd11an1n64x5 FILLER_91_1569 ();
 b15zdnd11an1n64x5 FILLER_91_1633 ();
 b15zdnd11an1n64x5 FILLER_91_1697 ();
 b15zdnd11an1n64x5 FILLER_91_1761 ();
 b15zdnd11an1n32x5 FILLER_91_1825 ();
 b15zdnd00an1n02x5 FILLER_91_1857 ();
 b15zdnd00an1n01x5 FILLER_91_1859 ();
 b15zdnd11an1n04x5 FILLER_91_1863 ();
 b15zdnd11an1n64x5 FILLER_91_1870 ();
 b15zdnd11an1n64x5 FILLER_91_1934 ();
 b15zdnd11an1n64x5 FILLER_91_1998 ();
 b15zdnd11an1n32x5 FILLER_91_2062 ();
 b15zdnd11an1n16x5 FILLER_91_2094 ();
 b15zdnd11an1n08x5 FILLER_91_2113 ();
 b15zdnd00an1n01x5 FILLER_91_2121 ();
 b15zdnd11an1n64x5 FILLER_91_2125 ();
 b15zdnd11an1n64x5 FILLER_91_2189 ();
 b15zdnd11an1n16x5 FILLER_91_2253 ();
 b15zdnd11an1n08x5 FILLER_91_2269 ();
 b15zdnd11an1n04x5 FILLER_91_2277 ();
 b15zdnd00an1n02x5 FILLER_91_2281 ();
 b15zdnd00an1n01x5 FILLER_91_2283 ();
 b15zdnd11an1n64x5 FILLER_92_8 ();
 b15zdnd11an1n64x5 FILLER_92_72 ();
 b15zdnd11an1n32x5 FILLER_92_136 ();
 b15zdnd11an1n04x5 FILLER_92_168 ();
 b15zdnd00an1n02x5 FILLER_92_172 ();
 b15zdnd00an1n01x5 FILLER_92_174 ();
 b15zdnd11an1n04x5 FILLER_92_227 ();
 b15zdnd00an1n02x5 FILLER_92_231 ();
 b15zdnd00an1n01x5 FILLER_92_233 ();
 b15zdnd11an1n64x5 FILLER_92_238 ();
 b15zdnd11an1n64x5 FILLER_92_302 ();
 b15zdnd11an1n64x5 FILLER_92_366 ();
 b15zdnd11an1n32x5 FILLER_92_430 ();
 b15zdnd11an1n08x5 FILLER_92_462 ();
 b15zdnd00an1n02x5 FILLER_92_470 ();
 b15zdnd00an1n01x5 FILLER_92_472 ();
 b15zdnd11an1n64x5 FILLER_92_513 ();
 b15zdnd11an1n64x5 FILLER_92_577 ();
 b15zdnd11an1n64x5 FILLER_92_641 ();
 b15zdnd11an1n08x5 FILLER_92_705 ();
 b15zdnd11an1n04x5 FILLER_92_713 ();
 b15zdnd00an1n01x5 FILLER_92_717 ();
 b15zdnd11an1n64x5 FILLER_92_726 ();
 b15zdnd11an1n64x5 FILLER_92_790 ();
 b15zdnd11an1n64x5 FILLER_92_854 ();
 b15zdnd11an1n64x5 FILLER_92_918 ();
 b15zdnd11an1n64x5 FILLER_92_982 ();
 b15zdnd11an1n16x5 FILLER_92_1046 ();
 b15zdnd11an1n04x5 FILLER_92_1062 ();
 b15zdnd00an1n02x5 FILLER_92_1066 ();
 b15zdnd00an1n01x5 FILLER_92_1068 ();
 b15zdnd11an1n64x5 FILLER_92_1073 ();
 b15zdnd11an1n32x5 FILLER_92_1137 ();
 b15zdnd11an1n16x5 FILLER_92_1169 ();
 b15zdnd11an1n04x5 FILLER_92_1185 ();
 b15zdnd00an1n02x5 FILLER_92_1189 ();
 b15zdnd11an1n64x5 FILLER_92_1198 ();
 b15zdnd11an1n16x5 FILLER_92_1262 ();
 b15zdnd11an1n08x5 FILLER_92_1278 ();
 b15zdnd11an1n04x5 FILLER_92_1286 ();
 b15zdnd00an1n02x5 FILLER_92_1290 ();
 b15zdnd11an1n64x5 FILLER_92_1295 ();
 b15zdnd11an1n64x5 FILLER_92_1359 ();
 b15zdnd11an1n64x5 FILLER_92_1423 ();
 b15zdnd11an1n64x5 FILLER_92_1487 ();
 b15zdnd11an1n64x5 FILLER_92_1551 ();
 b15zdnd11an1n64x5 FILLER_92_1615 ();
 b15zdnd11an1n64x5 FILLER_92_1679 ();
 b15zdnd11an1n64x5 FILLER_92_1743 ();
 b15zdnd11an1n32x5 FILLER_92_1807 ();
 b15zdnd11an1n16x5 FILLER_92_1839 ();
 b15zdnd11an1n04x5 FILLER_92_1855 ();
 b15zdnd00an1n02x5 FILLER_92_1859 ();
 b15zdnd11an1n64x5 FILLER_92_1864 ();
 b15zdnd11an1n64x5 FILLER_92_1928 ();
 b15zdnd11an1n64x5 FILLER_92_1992 ();
 b15zdnd11an1n16x5 FILLER_92_2056 ();
 b15zdnd11an1n08x5 FILLER_92_2072 ();
 b15zdnd11an1n04x5 FILLER_92_2080 ();
 b15zdnd00an1n02x5 FILLER_92_2084 ();
 b15zdnd00an1n01x5 FILLER_92_2086 ();
 b15zdnd11an1n08x5 FILLER_92_2139 ();
 b15zdnd11an1n04x5 FILLER_92_2147 ();
 b15zdnd00an1n02x5 FILLER_92_2151 ();
 b15zdnd00an1n01x5 FILLER_92_2153 ();
 b15zdnd11an1n64x5 FILLER_92_2162 ();
 b15zdnd11an1n32x5 FILLER_92_2226 ();
 b15zdnd11an1n16x5 FILLER_92_2258 ();
 b15zdnd00an1n02x5 FILLER_92_2274 ();
 b15zdnd11an1n64x5 FILLER_93_0 ();
 b15zdnd11an1n64x5 FILLER_93_64 ();
 b15zdnd11an1n32x5 FILLER_93_128 ();
 b15zdnd11an1n16x5 FILLER_93_160 ();
 b15zdnd11an1n04x5 FILLER_93_176 ();
 b15zdnd00an1n01x5 FILLER_93_180 ();
 b15zdnd11an1n04x5 FILLER_93_184 ();
 b15zdnd11an1n04x5 FILLER_93_191 ();
 b15zdnd11an1n04x5 FILLER_93_200 ();
 b15zdnd11an1n04x5 FILLER_93_213 ();
 b15zdnd11an1n08x5 FILLER_93_222 ();
 b15zdnd11an1n64x5 FILLER_93_272 ();
 b15zdnd11an1n64x5 FILLER_93_336 ();
 b15zdnd11an1n64x5 FILLER_93_400 ();
 b15zdnd11an1n32x5 FILLER_93_464 ();
 b15zdnd11an1n08x5 FILLER_93_496 ();
 b15zdnd11an1n04x5 FILLER_93_504 ();
 b15zdnd11an1n32x5 FILLER_93_511 ();
 b15zdnd11an1n04x5 FILLER_93_543 ();
 b15zdnd00an1n01x5 FILLER_93_547 ();
 b15zdnd11an1n16x5 FILLER_93_590 ();
 b15zdnd11an1n08x5 FILLER_93_606 ();
 b15zdnd00an1n02x5 FILLER_93_614 ();
 b15zdnd11an1n64x5 FILLER_93_622 ();
 b15zdnd11an1n64x5 FILLER_93_686 ();
 b15zdnd11an1n08x5 FILLER_93_750 ();
 b15zdnd00an1n02x5 FILLER_93_758 ();
 b15zdnd00an1n01x5 FILLER_93_760 ();
 b15zdnd11an1n08x5 FILLER_93_765 ();
 b15zdnd00an1n01x5 FILLER_93_773 ();
 b15zdnd11an1n64x5 FILLER_93_778 ();
 b15zdnd11an1n64x5 FILLER_93_842 ();
 b15zdnd11an1n16x5 FILLER_93_906 ();
 b15zdnd11an1n08x5 FILLER_93_922 ();
 b15zdnd11an1n04x5 FILLER_93_930 ();
 b15zdnd00an1n02x5 FILLER_93_934 ();
 b15zdnd11an1n64x5 FILLER_93_940 ();
 b15zdnd11an1n64x5 FILLER_93_1004 ();
 b15zdnd11an1n08x5 FILLER_93_1068 ();
 b15zdnd11an1n04x5 FILLER_93_1076 ();
 b15zdnd11an1n64x5 FILLER_93_1084 ();
 b15zdnd11an1n32x5 FILLER_93_1148 ();
 b15zdnd11an1n04x5 FILLER_93_1180 ();
 b15zdnd00an1n01x5 FILLER_93_1184 ();
 b15zdnd11an1n64x5 FILLER_93_1216 ();
 b15zdnd11an1n64x5 FILLER_93_1280 ();
 b15zdnd11an1n32x5 FILLER_93_1344 ();
 b15zdnd00an1n02x5 FILLER_93_1376 ();
 b15zdnd00an1n01x5 FILLER_93_1378 ();
 b15zdnd11an1n64x5 FILLER_93_1406 ();
 b15zdnd11an1n64x5 FILLER_93_1470 ();
 b15zdnd11an1n64x5 FILLER_93_1534 ();
 b15zdnd11an1n64x5 FILLER_93_1598 ();
 b15zdnd11an1n64x5 FILLER_93_1662 ();
 b15zdnd11an1n64x5 FILLER_93_1726 ();
 b15zdnd11an1n64x5 FILLER_93_1790 ();
 b15zdnd11an1n64x5 FILLER_93_1854 ();
 b15zdnd11an1n64x5 FILLER_93_1918 ();
 b15zdnd11an1n64x5 FILLER_93_1982 ();
 b15zdnd11an1n32x5 FILLER_93_2046 ();
 b15zdnd11an1n16x5 FILLER_93_2078 ();
 b15zdnd11an1n08x5 FILLER_93_2094 ();
 b15zdnd11an1n04x5 FILLER_93_2102 ();
 b15zdnd00an1n02x5 FILLER_93_2106 ();
 b15zdnd00an1n01x5 FILLER_93_2108 ();
 b15zdnd11an1n64x5 FILLER_93_2112 ();
 b15zdnd11an1n64x5 FILLER_93_2176 ();
 b15zdnd11an1n32x5 FILLER_93_2240 ();
 b15zdnd11an1n08x5 FILLER_93_2272 ();
 b15zdnd11an1n04x5 FILLER_93_2280 ();
 b15zdnd11an1n64x5 FILLER_94_8 ();
 b15zdnd11an1n64x5 FILLER_94_72 ();
 b15zdnd11an1n32x5 FILLER_94_136 ();
 b15zdnd11an1n16x5 FILLER_94_168 ();
 b15zdnd11an1n04x5 FILLER_94_195 ();
 b15zdnd11an1n64x5 FILLER_94_241 ();
 b15zdnd11an1n64x5 FILLER_94_305 ();
 b15zdnd11an1n08x5 FILLER_94_369 ();
 b15zdnd11an1n04x5 FILLER_94_377 ();
 b15zdnd00an1n01x5 FILLER_94_381 ();
 b15zdnd11an1n64x5 FILLER_94_424 ();
 b15zdnd11an1n64x5 FILLER_94_488 ();
 b15zdnd11an1n64x5 FILLER_94_552 ();
 b15zdnd11an1n64x5 FILLER_94_616 ();
 b15zdnd11an1n32x5 FILLER_94_680 ();
 b15zdnd11an1n04x5 FILLER_94_712 ();
 b15zdnd00an1n02x5 FILLER_94_716 ();
 b15zdnd11an1n64x5 FILLER_94_726 ();
 b15zdnd11an1n64x5 FILLER_94_790 ();
 b15zdnd11an1n64x5 FILLER_94_854 ();
 b15zdnd11an1n04x5 FILLER_94_918 ();
 b15zdnd00an1n02x5 FILLER_94_922 ();
 b15zdnd00an1n01x5 FILLER_94_924 ();
 b15zdnd11an1n64x5 FILLER_94_931 ();
 b15zdnd11an1n64x5 FILLER_94_995 ();
 b15zdnd11an1n64x5 FILLER_94_1059 ();
 b15zdnd11an1n64x5 FILLER_94_1123 ();
 b15zdnd11an1n64x5 FILLER_94_1187 ();
 b15zdnd11an1n64x5 FILLER_94_1251 ();
 b15zdnd11an1n64x5 FILLER_94_1315 ();
 b15zdnd11an1n64x5 FILLER_94_1379 ();
 b15zdnd11an1n64x5 FILLER_94_1443 ();
 b15zdnd11an1n64x5 FILLER_94_1507 ();
 b15zdnd11an1n64x5 FILLER_94_1571 ();
 b15zdnd11an1n64x5 FILLER_94_1635 ();
 b15zdnd11an1n64x5 FILLER_94_1699 ();
 b15zdnd11an1n64x5 FILLER_94_1763 ();
 b15zdnd11an1n64x5 FILLER_94_1827 ();
 b15zdnd11an1n64x5 FILLER_94_1891 ();
 b15zdnd11an1n64x5 FILLER_94_1955 ();
 b15zdnd11an1n64x5 FILLER_94_2019 ();
 b15zdnd11an1n08x5 FILLER_94_2083 ();
 b15zdnd11an1n04x5 FILLER_94_2091 ();
 b15zdnd00an1n02x5 FILLER_94_2095 ();
 b15zdnd00an1n01x5 FILLER_94_2097 ();
 b15zdnd11an1n32x5 FILLER_94_2102 ();
 b15zdnd11an1n16x5 FILLER_94_2134 ();
 b15zdnd11an1n04x5 FILLER_94_2150 ();
 b15zdnd11an1n64x5 FILLER_94_2162 ();
 b15zdnd11an1n32x5 FILLER_94_2226 ();
 b15zdnd11an1n16x5 FILLER_94_2258 ();
 b15zdnd00an1n02x5 FILLER_94_2274 ();
 b15zdnd11an1n64x5 FILLER_95_0 ();
 b15zdnd11an1n64x5 FILLER_95_64 ();
 b15zdnd11an1n32x5 FILLER_95_128 ();
 b15zdnd11an1n16x5 FILLER_95_160 ();
 b15zdnd11an1n08x5 FILLER_95_176 ();
 b15zdnd11an1n04x5 FILLER_95_184 ();
 b15zdnd11an1n64x5 FILLER_95_230 ();
 b15zdnd11an1n64x5 FILLER_95_294 ();
 b15zdnd11an1n64x5 FILLER_95_358 ();
 b15zdnd11an1n64x5 FILLER_95_422 ();
 b15zdnd11an1n64x5 FILLER_95_486 ();
 b15zdnd00an1n02x5 FILLER_95_550 ();
 b15zdnd00an1n01x5 FILLER_95_552 ();
 b15zdnd11an1n32x5 FILLER_95_557 ();
 b15zdnd11an1n16x5 FILLER_95_589 ();
 b15zdnd11an1n04x5 FILLER_95_605 ();
 b15zdnd11an1n04x5 FILLER_95_628 ();
 b15zdnd11an1n64x5 FILLER_95_636 ();
 b15zdnd11an1n64x5 FILLER_95_700 ();
 b15zdnd11an1n32x5 FILLER_95_764 ();
 b15zdnd11an1n16x5 FILLER_95_796 ();
 b15zdnd11an1n04x5 FILLER_95_812 ();
 b15zdnd00an1n02x5 FILLER_95_816 ();
 b15zdnd11an1n64x5 FILLER_95_825 ();
 b15zdnd11an1n32x5 FILLER_95_889 ();
 b15zdnd11an1n08x5 FILLER_95_921 ();
 b15zdnd11an1n04x5 FILLER_95_929 ();
 b15zdnd11an1n32x5 FILLER_95_937 ();
 b15zdnd11an1n04x5 FILLER_95_969 ();
 b15zdnd00an1n02x5 FILLER_95_973 ();
 b15zdnd11an1n64x5 FILLER_95_992 ();
 b15zdnd11an1n64x5 FILLER_95_1056 ();
 b15zdnd11an1n32x5 FILLER_95_1120 ();
 b15zdnd11an1n08x5 FILLER_95_1152 ();
 b15zdnd11an1n64x5 FILLER_95_1204 ();
 b15zdnd11an1n64x5 FILLER_95_1268 ();
 b15zdnd11an1n64x5 FILLER_95_1332 ();
 b15zdnd11an1n64x5 FILLER_95_1396 ();
 b15zdnd11an1n64x5 FILLER_95_1460 ();
 b15zdnd11an1n64x5 FILLER_95_1524 ();
 b15zdnd11an1n64x5 FILLER_95_1588 ();
 b15zdnd11an1n64x5 FILLER_95_1652 ();
 b15zdnd11an1n32x5 FILLER_95_1716 ();
 b15zdnd11an1n64x5 FILLER_95_1752 ();
 b15zdnd11an1n64x5 FILLER_95_1816 ();
 b15zdnd11an1n64x5 FILLER_95_1880 ();
 b15zdnd11an1n64x5 FILLER_95_1944 ();
 b15zdnd00an1n02x5 FILLER_95_2008 ();
 b15zdnd11an1n64x5 FILLER_95_2013 ();
 b15zdnd11an1n16x5 FILLER_95_2077 ();
 b15zdnd00an1n02x5 FILLER_95_2093 ();
 b15zdnd11an1n04x5 FILLER_95_2101 ();
 b15zdnd00an1n02x5 FILLER_95_2105 ();
 b15zdnd00an1n01x5 FILLER_95_2107 ();
 b15zdnd11an1n64x5 FILLER_95_2112 ();
 b15zdnd11an1n64x5 FILLER_95_2176 ();
 b15zdnd11an1n32x5 FILLER_95_2240 ();
 b15zdnd11an1n08x5 FILLER_95_2272 ();
 b15zdnd11an1n04x5 FILLER_95_2280 ();
 b15zdnd11an1n64x5 FILLER_96_8 ();
 b15zdnd11an1n64x5 FILLER_96_72 ();
 b15zdnd11an1n32x5 FILLER_96_136 ();
 b15zdnd11an1n16x5 FILLER_96_168 ();
 b15zdnd11an1n04x5 FILLER_96_184 ();
 b15zdnd00an1n02x5 FILLER_96_188 ();
 b15zdnd11an1n08x5 FILLER_96_232 ();
 b15zdnd11an1n04x5 FILLER_96_240 ();
 b15zdnd11an1n64x5 FILLER_96_250 ();
 b15zdnd11an1n64x5 FILLER_96_314 ();
 b15zdnd11an1n64x5 FILLER_96_378 ();
 b15zdnd11an1n64x5 FILLER_96_442 ();
 b15zdnd11an1n32x5 FILLER_96_506 ();
 b15zdnd11an1n16x5 FILLER_96_538 ();
 b15zdnd11an1n04x5 FILLER_96_554 ();
 b15zdnd00an1n02x5 FILLER_96_558 ();
 b15zdnd11an1n08x5 FILLER_96_599 ();
 b15zdnd11an1n04x5 FILLER_96_607 ();
 b15zdnd00an1n02x5 FILLER_96_611 ();
 b15zdnd11an1n08x5 FILLER_96_619 ();
 b15zdnd11an1n04x5 FILLER_96_627 ();
 b15zdnd00an1n02x5 FILLER_96_631 ();
 b15zdnd11an1n08x5 FILLER_96_637 ();
 b15zdnd00an1n01x5 FILLER_96_645 ();
 b15zdnd11an1n64x5 FILLER_96_652 ();
 b15zdnd00an1n02x5 FILLER_96_716 ();
 b15zdnd11an1n32x5 FILLER_96_726 ();
 b15zdnd11an1n08x5 FILLER_96_758 ();
 b15zdnd00an1n02x5 FILLER_96_766 ();
 b15zdnd00an1n01x5 FILLER_96_768 ();
 b15zdnd11an1n64x5 FILLER_96_777 ();
 b15zdnd00an1n02x5 FILLER_96_841 ();
 b15zdnd11an1n64x5 FILLER_96_847 ();
 b15zdnd11an1n16x5 FILLER_96_911 ();
 b15zdnd11an1n64x5 FILLER_96_933 ();
 b15zdnd11an1n32x5 FILLER_96_997 ();
 b15zdnd11an1n16x5 FILLER_96_1029 ();
 b15zdnd11an1n08x5 FILLER_96_1045 ();
 b15zdnd00an1n01x5 FILLER_96_1053 ();
 b15zdnd11an1n08x5 FILLER_96_1057 ();
 b15zdnd11an1n04x5 FILLER_96_1065 ();
 b15zdnd00an1n01x5 FILLER_96_1069 ();
 b15zdnd11an1n64x5 FILLER_96_1074 ();
 b15zdnd11an1n32x5 FILLER_96_1138 ();
 b15zdnd11an1n04x5 FILLER_96_1170 ();
 b15zdnd00an1n01x5 FILLER_96_1174 ();
 b15zdnd11an1n04x5 FILLER_96_1178 ();
 b15zdnd11an1n04x5 FILLER_96_1185 ();
 b15zdnd11an1n64x5 FILLER_96_1192 ();
 b15zdnd11an1n64x5 FILLER_96_1256 ();
 b15zdnd11an1n64x5 FILLER_96_1320 ();
 b15zdnd11an1n64x5 FILLER_96_1384 ();
 b15zdnd11an1n64x5 FILLER_96_1448 ();
 b15zdnd11an1n64x5 FILLER_96_1512 ();
 b15zdnd11an1n64x5 FILLER_96_1576 ();
 b15zdnd11an1n64x5 FILLER_96_1640 ();
 b15zdnd11an1n64x5 FILLER_96_1704 ();
 b15zdnd11an1n64x5 FILLER_96_1768 ();
 b15zdnd11an1n64x5 FILLER_96_1832 ();
 b15zdnd11an1n64x5 FILLER_96_1896 ();
 b15zdnd11an1n32x5 FILLER_96_1960 ();
 b15zdnd11an1n08x5 FILLER_96_1992 ();
 b15zdnd00an1n02x5 FILLER_96_2000 ();
 b15zdnd00an1n01x5 FILLER_96_2002 ();
 b15zdnd11an1n04x5 FILLER_96_2009 ();
 b15zdnd11an1n04x5 FILLER_96_2018 ();
 b15zdnd11an1n32x5 FILLER_96_2026 ();
 b15zdnd11an1n16x5 FILLER_96_2058 ();
 b15zdnd11an1n08x5 FILLER_96_2074 ();
 b15zdnd11an1n04x5 FILLER_96_2082 ();
 b15zdnd00an1n01x5 FILLER_96_2086 ();
 b15zdnd11an1n32x5 FILLER_96_2091 ();
 b15zdnd11an1n16x5 FILLER_96_2123 ();
 b15zdnd11an1n08x5 FILLER_96_2139 ();
 b15zdnd11an1n04x5 FILLER_96_2147 ();
 b15zdnd00an1n02x5 FILLER_96_2151 ();
 b15zdnd00an1n01x5 FILLER_96_2153 ();
 b15zdnd11an1n64x5 FILLER_96_2162 ();
 b15zdnd11an1n32x5 FILLER_96_2226 ();
 b15zdnd11an1n16x5 FILLER_96_2258 ();
 b15zdnd00an1n02x5 FILLER_96_2274 ();
 b15zdnd11an1n64x5 FILLER_97_0 ();
 b15zdnd11an1n64x5 FILLER_97_64 ();
 b15zdnd11an1n64x5 FILLER_97_128 ();
 b15zdnd11an1n04x5 FILLER_97_199 ();
 b15zdnd11an1n04x5 FILLER_97_216 ();
 b15zdnd11an1n64x5 FILLER_97_226 ();
 b15zdnd11an1n32x5 FILLER_97_290 ();
 b15zdnd11an1n08x5 FILLER_97_322 ();
 b15zdnd11an1n64x5 FILLER_97_382 ();
 b15zdnd11an1n64x5 FILLER_97_446 ();
 b15zdnd11an1n64x5 FILLER_97_510 ();
 b15zdnd11an1n08x5 FILLER_97_574 ();
 b15zdnd00an1n02x5 FILLER_97_582 ();
 b15zdnd11an1n32x5 FILLER_97_592 ();
 b15zdnd11an1n16x5 FILLER_97_624 ();
 b15zdnd00an1n02x5 FILLER_97_640 ();
 b15zdnd11an1n64x5 FILLER_97_646 ();
 b15zdnd11an1n64x5 FILLER_97_710 ();
 b15zdnd11an1n32x5 FILLER_97_774 ();
 b15zdnd11an1n16x5 FILLER_97_806 ();
 b15zdnd11an1n04x5 FILLER_97_822 ();
 b15zdnd11an1n32x5 FILLER_97_836 ();
 b15zdnd11an1n08x5 FILLER_97_868 ();
 b15zdnd00an1n02x5 FILLER_97_876 ();
 b15zdnd00an1n01x5 FILLER_97_878 ();
 b15zdnd11an1n04x5 FILLER_97_883 ();
 b15zdnd11an1n32x5 FILLER_97_891 ();
 b15zdnd11an1n04x5 FILLER_97_923 ();
 b15zdnd11an1n04x5 FILLER_97_931 ();
 b15zdnd11an1n04x5 FILLER_97_939 ();
 b15zdnd11an1n64x5 FILLER_97_947 ();
 b15zdnd11an1n16x5 FILLER_97_1011 ();
 b15zdnd00an1n02x5 FILLER_97_1027 ();
 b15zdnd00an1n01x5 FILLER_97_1029 ();
 b15zdnd11an1n64x5 FILLER_97_1082 ();
 b15zdnd11an1n64x5 FILLER_97_1146 ();
 b15zdnd11an1n32x5 FILLER_97_1210 ();
 b15zdnd11an1n16x5 FILLER_97_1242 ();
 b15zdnd11an1n08x5 FILLER_97_1258 ();
 b15zdnd00an1n01x5 FILLER_97_1266 ();
 b15zdnd11an1n64x5 FILLER_97_1270 ();
 b15zdnd11an1n64x5 FILLER_97_1334 ();
 b15zdnd11an1n32x5 FILLER_97_1398 ();
 b15zdnd11an1n04x5 FILLER_97_1430 ();
 b15zdnd00an1n02x5 FILLER_97_1434 ();
 b15zdnd00an1n01x5 FILLER_97_1436 ();
 b15zdnd11an1n64x5 FILLER_97_1455 ();
 b15zdnd11an1n64x5 FILLER_97_1519 ();
 b15zdnd11an1n64x5 FILLER_97_1583 ();
 b15zdnd11an1n64x5 FILLER_97_1647 ();
 b15zdnd11an1n16x5 FILLER_97_1711 ();
 b15zdnd11an1n08x5 FILLER_97_1727 ();
 b15zdnd11an1n04x5 FILLER_97_1735 ();
 b15zdnd11an1n08x5 FILLER_97_1742 ();
 b15zdnd11an1n04x5 FILLER_97_1750 ();
 b15zdnd00an1n02x5 FILLER_97_1754 ();
 b15zdnd00an1n01x5 FILLER_97_1756 ();
 b15zdnd11an1n64x5 FILLER_97_1799 ();
 b15zdnd11an1n04x5 FILLER_97_1863 ();
 b15zdnd00an1n02x5 FILLER_97_1867 ();
 b15zdnd11an1n64x5 FILLER_97_1911 ();
 b15zdnd11an1n16x5 FILLER_97_1975 ();
 b15zdnd00an1n02x5 FILLER_97_1991 ();
 b15zdnd11an1n08x5 FILLER_97_1999 ();
 b15zdnd00an1n02x5 FILLER_97_2007 ();
 b15zdnd00an1n01x5 FILLER_97_2009 ();
 b15zdnd11an1n04x5 FILLER_97_2022 ();
 b15zdnd11an1n64x5 FILLER_97_2029 ();
 b15zdnd11an1n64x5 FILLER_97_2093 ();
 b15zdnd11an1n64x5 FILLER_97_2157 ();
 b15zdnd11an1n32x5 FILLER_97_2221 ();
 b15zdnd11an1n16x5 FILLER_97_2253 ();
 b15zdnd11an1n08x5 FILLER_97_2269 ();
 b15zdnd11an1n04x5 FILLER_97_2277 ();
 b15zdnd00an1n02x5 FILLER_97_2281 ();
 b15zdnd00an1n01x5 FILLER_97_2283 ();
 b15zdnd11an1n64x5 FILLER_98_8 ();
 b15zdnd11an1n64x5 FILLER_98_72 ();
 b15zdnd11an1n32x5 FILLER_98_136 ();
 b15zdnd11an1n16x5 FILLER_98_168 ();
 b15zdnd11an1n08x5 FILLER_98_184 ();
 b15zdnd00an1n02x5 FILLER_98_192 ();
 b15zdnd11an1n16x5 FILLER_98_198 ();
 b15zdnd00an1n01x5 FILLER_98_214 ();
 b15zdnd11an1n64x5 FILLER_98_257 ();
 b15zdnd11an1n16x5 FILLER_98_321 ();
 b15zdnd11an1n08x5 FILLER_98_337 ();
 b15zdnd00an1n01x5 FILLER_98_345 ();
 b15zdnd11an1n64x5 FILLER_98_388 ();
 b15zdnd11an1n64x5 FILLER_98_452 ();
 b15zdnd11an1n64x5 FILLER_98_516 ();
 b15zdnd11an1n32x5 FILLER_98_580 ();
 b15zdnd11an1n16x5 FILLER_98_612 ();
 b15zdnd11an1n08x5 FILLER_98_628 ();
 b15zdnd11an1n04x5 FILLER_98_640 ();
 b15zdnd00an1n02x5 FILLER_98_644 ();
 b15zdnd11an1n64x5 FILLER_98_652 ();
 b15zdnd00an1n02x5 FILLER_98_716 ();
 b15zdnd11an1n16x5 FILLER_98_726 ();
 b15zdnd11an1n08x5 FILLER_98_742 ();
 b15zdnd11an1n04x5 FILLER_98_750 ();
 b15zdnd00an1n02x5 FILLER_98_754 ();
 b15zdnd11an1n64x5 FILLER_98_760 ();
 b15zdnd11an1n64x5 FILLER_98_824 ();
 b15zdnd11an1n08x5 FILLER_98_888 ();
 b15zdnd00an1n02x5 FILLER_98_896 ();
 b15zdnd00an1n01x5 FILLER_98_898 ();
 b15zdnd11an1n32x5 FILLER_98_941 ();
 b15zdnd11an1n04x5 FILLER_98_973 ();
 b15zdnd11an1n64x5 FILLER_98_985 ();
 b15zdnd00an1n02x5 FILLER_98_1049 ();
 b15zdnd11an1n64x5 FILLER_98_1054 ();
 b15zdnd11an1n64x5 FILLER_98_1118 ();
 b15zdnd11an1n64x5 FILLER_98_1182 ();
 b15zdnd11an1n64x5 FILLER_98_1246 ();
 b15zdnd11an1n16x5 FILLER_98_1310 ();
 b15zdnd11an1n08x5 FILLER_98_1326 ();
 b15zdnd11an1n04x5 FILLER_98_1334 ();
 b15zdnd00an1n02x5 FILLER_98_1338 ();
 b15zdnd11an1n64x5 FILLER_98_1348 ();
 b15zdnd11an1n64x5 FILLER_98_1412 ();
 b15zdnd11an1n64x5 FILLER_98_1476 ();
 b15zdnd11an1n32x5 FILLER_98_1540 ();
 b15zdnd00an1n02x5 FILLER_98_1572 ();
 b15zdnd11an1n64x5 FILLER_98_1578 ();
 b15zdnd11an1n64x5 FILLER_98_1642 ();
 b15zdnd11an1n16x5 FILLER_98_1706 ();
 b15zdnd11an1n08x5 FILLER_98_1722 ();
 b15zdnd00an1n02x5 FILLER_98_1730 ();
 b15zdnd00an1n01x5 FILLER_98_1732 ();
 b15zdnd11an1n04x5 FILLER_98_1736 ();
 b15zdnd11an1n64x5 FILLER_98_1743 ();
 b15zdnd11an1n64x5 FILLER_98_1807 ();
 b15zdnd11an1n64x5 FILLER_98_1871 ();
 b15zdnd11an1n32x5 FILLER_98_1935 ();
 b15zdnd11an1n16x5 FILLER_98_1967 ();
 b15zdnd11an1n08x5 FILLER_98_1983 ();
 b15zdnd11an1n04x5 FILLER_98_2004 ();
 b15zdnd11an1n64x5 FILLER_98_2050 ();
 b15zdnd11an1n32x5 FILLER_98_2114 ();
 b15zdnd11an1n08x5 FILLER_98_2146 ();
 b15zdnd11an1n64x5 FILLER_98_2162 ();
 b15zdnd11an1n32x5 FILLER_98_2226 ();
 b15zdnd11an1n16x5 FILLER_98_2258 ();
 b15zdnd00an1n02x5 FILLER_98_2274 ();
 b15zdnd11an1n64x5 FILLER_99_0 ();
 b15zdnd11an1n64x5 FILLER_99_64 ();
 b15zdnd11an1n64x5 FILLER_99_128 ();
 b15zdnd11an1n64x5 FILLER_99_192 ();
 b15zdnd11an1n64x5 FILLER_99_256 ();
 b15zdnd11an1n16x5 FILLER_99_320 ();
 b15zdnd11an1n08x5 FILLER_99_336 ();
 b15zdnd11an1n04x5 FILLER_99_344 ();
 b15zdnd00an1n01x5 FILLER_99_348 ();
 b15zdnd11an1n04x5 FILLER_99_352 ();
 b15zdnd11an1n04x5 FILLER_99_359 ();
 b15zdnd11an1n64x5 FILLER_99_366 ();
 b15zdnd11an1n64x5 FILLER_99_430 ();
 b15zdnd11an1n64x5 FILLER_99_494 ();
 b15zdnd11an1n64x5 FILLER_99_558 ();
 b15zdnd11an1n64x5 FILLER_99_622 ();
 b15zdnd11an1n64x5 FILLER_99_686 ();
 b15zdnd11an1n64x5 FILLER_99_750 ();
 b15zdnd11an1n08x5 FILLER_99_814 ();
 b15zdnd00an1n02x5 FILLER_99_822 ();
 b15zdnd11an1n64x5 FILLER_99_832 ();
 b15zdnd11an1n32x5 FILLER_99_896 ();
 b15zdnd11an1n16x5 FILLER_99_928 ();
 b15zdnd11an1n08x5 FILLER_99_944 ();
 b15zdnd11an1n04x5 FILLER_99_952 ();
 b15zdnd00an1n02x5 FILLER_99_956 ();
 b15zdnd11an1n64x5 FILLER_99_972 ();
 b15zdnd11an1n08x5 FILLER_99_1036 ();
 b15zdnd11an1n04x5 FILLER_99_1044 ();
 b15zdnd00an1n02x5 FILLER_99_1048 ();
 b15zdnd11an1n16x5 FILLER_99_1053 ();
 b15zdnd11an1n04x5 FILLER_99_1069 ();
 b15zdnd00an1n02x5 FILLER_99_1073 ();
 b15zdnd00an1n01x5 FILLER_99_1075 ();
 b15zdnd11an1n64x5 FILLER_99_1082 ();
 b15zdnd11an1n64x5 FILLER_99_1146 ();
 b15zdnd11an1n64x5 FILLER_99_1210 ();
 b15zdnd11an1n64x5 FILLER_99_1274 ();
 b15zdnd11an1n64x5 FILLER_99_1338 ();
 b15zdnd11an1n64x5 FILLER_99_1402 ();
 b15zdnd11an1n64x5 FILLER_99_1466 ();
 b15zdnd11an1n64x5 FILLER_99_1530 ();
 b15zdnd11an1n64x5 FILLER_99_1594 ();
 b15zdnd11an1n32x5 FILLER_99_1658 ();
 b15zdnd11an1n16x5 FILLER_99_1690 ();
 b15zdnd11an1n08x5 FILLER_99_1706 ();
 b15zdnd00an1n01x5 FILLER_99_1714 ();
 b15zdnd11an1n64x5 FILLER_99_1767 ();
 b15zdnd11an1n64x5 FILLER_99_1831 ();
 b15zdnd11an1n64x5 FILLER_99_1895 ();
 b15zdnd11an1n08x5 FILLER_99_1959 ();
 b15zdnd11an1n04x5 FILLER_99_1967 ();
 b15zdnd11an1n04x5 FILLER_99_2023 ();
 b15zdnd11an1n64x5 FILLER_99_2069 ();
 b15zdnd11an1n64x5 FILLER_99_2133 ();
 b15zdnd11an1n64x5 FILLER_99_2197 ();
 b15zdnd11an1n16x5 FILLER_99_2261 ();
 b15zdnd11an1n04x5 FILLER_99_2277 ();
 b15zdnd00an1n02x5 FILLER_99_2281 ();
 b15zdnd00an1n01x5 FILLER_99_2283 ();
 b15zdnd11an1n64x5 FILLER_100_8 ();
 b15zdnd11an1n64x5 FILLER_100_72 ();
 b15zdnd11an1n64x5 FILLER_100_136 ();
 b15zdnd11an1n16x5 FILLER_100_200 ();
 b15zdnd11an1n08x5 FILLER_100_216 ();
 b15zdnd00an1n02x5 FILLER_100_224 ();
 b15zdnd11an1n64x5 FILLER_100_229 ();
 b15zdnd11an1n64x5 FILLER_100_293 ();
 b15zdnd11an1n64x5 FILLER_100_357 ();
 b15zdnd11an1n64x5 FILLER_100_421 ();
 b15zdnd11an1n64x5 FILLER_100_485 ();
 b15zdnd11an1n64x5 FILLER_100_549 ();
 b15zdnd11an1n64x5 FILLER_100_613 ();
 b15zdnd11an1n32x5 FILLER_100_677 ();
 b15zdnd11an1n08x5 FILLER_100_709 ();
 b15zdnd00an1n01x5 FILLER_100_717 ();
 b15zdnd11an1n64x5 FILLER_100_726 ();
 b15zdnd11an1n64x5 FILLER_100_790 ();
 b15zdnd11an1n64x5 FILLER_100_854 ();
 b15zdnd11an1n64x5 FILLER_100_918 ();
 b15zdnd11an1n32x5 FILLER_100_982 ();
 b15zdnd11an1n04x5 FILLER_100_1014 ();
 b15zdnd00an1n01x5 FILLER_100_1018 ();
 b15zdnd11an1n64x5 FILLER_100_1030 ();
 b15zdnd11an1n64x5 FILLER_100_1094 ();
 b15zdnd11an1n64x5 FILLER_100_1158 ();
 b15zdnd11an1n64x5 FILLER_100_1222 ();
 b15zdnd11an1n32x5 FILLER_100_1286 ();
 b15zdnd11an1n08x5 FILLER_100_1318 ();
 b15zdnd00an1n01x5 FILLER_100_1326 ();
 b15zdnd11an1n08x5 FILLER_100_1336 ();
 b15zdnd11an1n04x5 FILLER_100_1344 ();
 b15zdnd00an1n02x5 FILLER_100_1348 ();
 b15zdnd00an1n01x5 FILLER_100_1350 ();
 b15zdnd11an1n04x5 FILLER_100_1355 ();
 b15zdnd11an1n64x5 FILLER_100_1363 ();
 b15zdnd11an1n04x5 FILLER_100_1427 ();
 b15zdnd00an1n02x5 FILLER_100_1431 ();
 b15zdnd00an1n01x5 FILLER_100_1433 ();
 b15zdnd11an1n04x5 FILLER_100_1437 ();
 b15zdnd11an1n64x5 FILLER_100_1444 ();
 b15zdnd11an1n64x5 FILLER_100_1508 ();
 b15zdnd11an1n64x5 FILLER_100_1572 ();
 b15zdnd11an1n64x5 FILLER_100_1636 ();
 b15zdnd11an1n64x5 FILLER_100_1700 ();
 b15zdnd11an1n04x5 FILLER_100_1764 ();
 b15zdnd11an1n64x5 FILLER_100_1788 ();
 b15zdnd11an1n64x5 FILLER_100_1852 ();
 b15zdnd11an1n64x5 FILLER_100_1916 ();
 b15zdnd11an1n04x5 FILLER_100_1980 ();
 b15zdnd11an1n04x5 FILLER_100_1987 ();
 b15zdnd11an1n08x5 FILLER_100_2001 ();
 b15zdnd00an1n02x5 FILLER_100_2009 ();
 b15zdnd11an1n64x5 FILLER_100_2053 ();
 b15zdnd11an1n32x5 FILLER_100_2117 ();
 b15zdnd11an1n04x5 FILLER_100_2149 ();
 b15zdnd00an1n01x5 FILLER_100_2153 ();
 b15zdnd11an1n64x5 FILLER_100_2162 ();
 b15zdnd11an1n32x5 FILLER_100_2226 ();
 b15zdnd11an1n16x5 FILLER_100_2258 ();
 b15zdnd00an1n02x5 FILLER_100_2274 ();
 b15zdnd11an1n64x5 FILLER_101_0 ();
 b15zdnd11an1n64x5 FILLER_101_64 ();
 b15zdnd11an1n64x5 FILLER_101_128 ();
 b15zdnd11an1n04x5 FILLER_101_192 ();
 b15zdnd00an1n02x5 FILLER_101_196 ();
 b15zdnd00an1n01x5 FILLER_101_198 ();
 b15zdnd11an1n64x5 FILLER_101_251 ();
 b15zdnd11an1n64x5 FILLER_101_315 ();
 b15zdnd11an1n64x5 FILLER_101_379 ();
 b15zdnd11an1n64x5 FILLER_101_443 ();
 b15zdnd11an1n64x5 FILLER_101_507 ();
 b15zdnd11an1n64x5 FILLER_101_571 ();
 b15zdnd11an1n32x5 FILLER_101_635 ();
 b15zdnd11an1n16x5 FILLER_101_667 ();
 b15zdnd11an1n04x5 FILLER_101_683 ();
 b15zdnd00an1n02x5 FILLER_101_687 ();
 b15zdnd11an1n64x5 FILLER_101_720 ();
 b15zdnd11an1n64x5 FILLER_101_784 ();
 b15zdnd11an1n64x5 FILLER_101_848 ();
 b15zdnd11an1n64x5 FILLER_101_912 ();
 b15zdnd11an1n32x5 FILLER_101_976 ();
 b15zdnd11an1n08x5 FILLER_101_1008 ();
 b15zdnd11an1n04x5 FILLER_101_1016 ();
 b15zdnd00an1n02x5 FILLER_101_1020 ();
 b15zdnd00an1n01x5 FILLER_101_1022 ();
 b15zdnd11an1n64x5 FILLER_101_1043 ();
 b15zdnd11an1n64x5 FILLER_101_1107 ();
 b15zdnd11an1n64x5 FILLER_101_1171 ();
 b15zdnd11an1n16x5 FILLER_101_1235 ();
 b15zdnd11an1n08x5 FILLER_101_1251 ();
 b15zdnd11an1n04x5 FILLER_101_1259 ();
 b15zdnd00an1n02x5 FILLER_101_1263 ();
 b15zdnd11an1n64x5 FILLER_101_1279 ();
 b15zdnd11an1n64x5 FILLER_101_1343 ();
 b15zdnd11an1n16x5 FILLER_101_1407 ();
 b15zdnd00an1n02x5 FILLER_101_1423 ();
 b15zdnd11an1n04x5 FILLER_101_1428 ();
 b15zdnd11an1n64x5 FILLER_101_1441 ();
 b15zdnd11an1n64x5 FILLER_101_1505 ();
 b15zdnd11an1n64x5 FILLER_101_1569 ();
 b15zdnd11an1n64x5 FILLER_101_1633 ();
 b15zdnd11an1n64x5 FILLER_101_1697 ();
 b15zdnd11an1n64x5 FILLER_101_1761 ();
 b15zdnd11an1n16x5 FILLER_101_1825 ();
 b15zdnd11an1n08x5 FILLER_101_1841 ();
 b15zdnd00an1n02x5 FILLER_101_1849 ();
 b15zdnd00an1n01x5 FILLER_101_1851 ();
 b15zdnd11an1n64x5 FILLER_101_1856 ();
 b15zdnd11an1n64x5 FILLER_101_1920 ();
 b15zdnd00an1n02x5 FILLER_101_1984 ();
 b15zdnd11an1n04x5 FILLER_101_1992 ();
 b15zdnd11an1n04x5 FILLER_101_1999 ();
 b15zdnd00an1n02x5 FILLER_101_2003 ();
 b15zdnd11an1n04x5 FILLER_101_2008 ();
 b15zdnd00an1n01x5 FILLER_101_2012 ();
 b15zdnd11an1n64x5 FILLER_101_2017 ();
 b15zdnd11an1n64x5 FILLER_101_2081 ();
 b15zdnd11an1n64x5 FILLER_101_2145 ();
 b15zdnd11an1n64x5 FILLER_101_2209 ();
 b15zdnd11an1n08x5 FILLER_101_2273 ();
 b15zdnd00an1n02x5 FILLER_101_2281 ();
 b15zdnd00an1n01x5 FILLER_101_2283 ();
 b15zdnd11an1n64x5 FILLER_102_8 ();
 b15zdnd11an1n64x5 FILLER_102_72 ();
 b15zdnd11an1n64x5 FILLER_102_136 ();
 b15zdnd11an1n16x5 FILLER_102_200 ();
 b15zdnd00an1n02x5 FILLER_102_216 ();
 b15zdnd11an1n04x5 FILLER_102_221 ();
 b15zdnd11an1n64x5 FILLER_102_228 ();
 b15zdnd11an1n64x5 FILLER_102_292 ();
 b15zdnd11an1n16x5 FILLER_102_356 ();
 b15zdnd11an1n08x5 FILLER_102_372 ();
 b15zdnd11an1n04x5 FILLER_102_380 ();
 b15zdnd00an1n02x5 FILLER_102_384 ();
 b15zdnd00an1n01x5 FILLER_102_386 ();
 b15zdnd11an1n64x5 FILLER_102_427 ();
 b15zdnd11an1n64x5 FILLER_102_491 ();
 b15zdnd11an1n64x5 FILLER_102_555 ();
 b15zdnd11an1n32x5 FILLER_102_619 ();
 b15zdnd11an1n16x5 FILLER_102_651 ();
 b15zdnd11an1n08x5 FILLER_102_667 ();
 b15zdnd00an1n01x5 FILLER_102_675 ();
 b15zdnd11an1n32x5 FILLER_102_680 ();
 b15zdnd11an1n04x5 FILLER_102_712 ();
 b15zdnd00an1n02x5 FILLER_102_716 ();
 b15zdnd11an1n64x5 FILLER_102_726 ();
 b15zdnd11an1n04x5 FILLER_102_790 ();
 b15zdnd11an1n64x5 FILLER_102_803 ();
 b15zdnd11an1n64x5 FILLER_102_867 ();
 b15zdnd11an1n64x5 FILLER_102_931 ();
 b15zdnd11an1n64x5 FILLER_102_995 ();
 b15zdnd11an1n64x5 FILLER_102_1059 ();
 b15zdnd11an1n08x5 FILLER_102_1137 ();
 b15zdnd00an1n02x5 FILLER_102_1145 ();
 b15zdnd00an1n01x5 FILLER_102_1147 ();
 b15zdnd11an1n64x5 FILLER_102_1159 ();
 b15zdnd11an1n32x5 FILLER_102_1223 ();
 b15zdnd11an1n16x5 FILLER_102_1255 ();
 b15zdnd11an1n08x5 FILLER_102_1271 ();
 b15zdnd11an1n04x5 FILLER_102_1279 ();
 b15zdnd00an1n02x5 FILLER_102_1283 ();
 b15zdnd00an1n01x5 FILLER_102_1285 ();
 b15zdnd11an1n08x5 FILLER_102_1292 ();
 b15zdnd11an1n04x5 FILLER_102_1300 ();
 b15zdnd00an1n02x5 FILLER_102_1304 ();
 b15zdnd00an1n01x5 FILLER_102_1306 ();
 b15zdnd11an1n16x5 FILLER_102_1311 ();
 b15zdnd11an1n04x5 FILLER_102_1327 ();
 b15zdnd00an1n02x5 FILLER_102_1331 ();
 b15zdnd11an1n64x5 FILLER_102_1341 ();
 b15zdnd00an1n02x5 FILLER_102_1405 ();
 b15zdnd00an1n01x5 FILLER_102_1407 ();
 b15zdnd11an1n64x5 FILLER_102_1460 ();
 b15zdnd11an1n64x5 FILLER_102_1524 ();
 b15zdnd11an1n64x5 FILLER_102_1588 ();
 b15zdnd11an1n32x5 FILLER_102_1652 ();
 b15zdnd11an1n16x5 FILLER_102_1684 ();
 b15zdnd11an1n08x5 FILLER_102_1700 ();
 b15zdnd11an1n04x5 FILLER_102_1711 ();
 b15zdnd11an1n64x5 FILLER_102_1718 ();
 b15zdnd11an1n32x5 FILLER_102_1782 ();
 b15zdnd11an1n16x5 FILLER_102_1814 ();
 b15zdnd11an1n04x5 FILLER_102_1830 ();
 b15zdnd00an1n01x5 FILLER_102_1834 ();
 b15zdnd11an1n04x5 FILLER_102_1838 ();
 b15zdnd11an1n04x5 FILLER_102_1845 ();
 b15zdnd11an1n04x5 FILLER_102_1856 ();
 b15zdnd11an1n04x5 FILLER_102_1865 ();
 b15zdnd11an1n64x5 FILLER_102_1874 ();
 b15zdnd11an1n64x5 FILLER_102_1938 ();
 b15zdnd11an1n64x5 FILLER_102_2002 ();
 b15zdnd11an1n64x5 FILLER_102_2066 ();
 b15zdnd11an1n16x5 FILLER_102_2130 ();
 b15zdnd11an1n08x5 FILLER_102_2146 ();
 b15zdnd11an1n64x5 FILLER_102_2162 ();
 b15zdnd11an1n32x5 FILLER_102_2226 ();
 b15zdnd11an1n16x5 FILLER_102_2258 ();
 b15zdnd00an1n02x5 FILLER_102_2274 ();
 b15zdnd11an1n64x5 FILLER_103_0 ();
 b15zdnd11an1n64x5 FILLER_103_64 ();
 b15zdnd11an1n64x5 FILLER_103_128 ();
 b15zdnd11an1n64x5 FILLER_103_192 ();
 b15zdnd11an1n64x5 FILLER_103_256 ();
 b15zdnd11an1n64x5 FILLER_103_320 ();
 b15zdnd11an1n32x5 FILLER_103_384 ();
 b15zdnd00an1n02x5 FILLER_103_416 ();
 b15zdnd11an1n04x5 FILLER_103_421 ();
 b15zdnd11an1n64x5 FILLER_103_428 ();
 b15zdnd11an1n64x5 FILLER_103_492 ();
 b15zdnd11an1n64x5 FILLER_103_556 ();
 b15zdnd11an1n32x5 FILLER_103_620 ();
 b15zdnd11an1n08x5 FILLER_103_652 ();
 b15zdnd11an1n04x5 FILLER_103_660 ();
 b15zdnd00an1n02x5 FILLER_103_664 ();
 b15zdnd11an1n04x5 FILLER_103_670 ();
 b15zdnd11an1n64x5 FILLER_103_678 ();
 b15zdnd11an1n64x5 FILLER_103_742 ();
 b15zdnd11an1n08x5 FILLER_103_806 ();
 b15zdnd11an1n04x5 FILLER_103_814 ();
 b15zdnd00an1n02x5 FILLER_103_818 ();
 b15zdnd11an1n64x5 FILLER_103_862 ();
 b15zdnd11an1n08x5 FILLER_103_926 ();
 b15zdnd11an1n04x5 FILLER_103_934 ();
 b15zdnd00an1n02x5 FILLER_103_938 ();
 b15zdnd11an1n64x5 FILLER_103_954 ();
 b15zdnd11an1n64x5 FILLER_103_1018 ();
 b15zdnd11an1n16x5 FILLER_103_1082 ();
 b15zdnd11an1n08x5 FILLER_103_1098 ();
 b15zdnd11an1n64x5 FILLER_103_1127 ();
 b15zdnd11an1n64x5 FILLER_103_1191 ();
 b15zdnd11an1n16x5 FILLER_103_1255 ();
 b15zdnd11an1n08x5 FILLER_103_1271 ();
 b15zdnd11an1n04x5 FILLER_103_1279 ();
 b15zdnd00an1n02x5 FILLER_103_1283 ();
 b15zdnd11an1n64x5 FILLER_103_1297 ();
 b15zdnd11an1n32x5 FILLER_103_1361 ();
 b15zdnd11an1n16x5 FILLER_103_1393 ();
 b15zdnd00an1n01x5 FILLER_103_1409 ();
 b15zdnd11an1n64x5 FILLER_103_1413 ();
 b15zdnd11an1n64x5 FILLER_103_1477 ();
 b15zdnd11an1n64x5 FILLER_103_1541 ();
 b15zdnd11an1n64x5 FILLER_103_1605 ();
 b15zdnd11an1n04x5 FILLER_103_1669 ();
 b15zdnd00an1n02x5 FILLER_103_1673 ();
 b15zdnd00an1n01x5 FILLER_103_1675 ();
 b15zdnd11an1n64x5 FILLER_103_1716 ();
 b15zdnd11an1n32x5 FILLER_103_1780 ();
 b15zdnd11an1n04x5 FILLER_103_1812 ();
 b15zdnd00an1n02x5 FILLER_103_1816 ();
 b15zdnd11an1n04x5 FILLER_103_1870 ();
 b15zdnd11an1n64x5 FILLER_103_1884 ();
 b15zdnd11an1n64x5 FILLER_103_1948 ();
 b15zdnd11an1n64x5 FILLER_103_2012 ();
 b15zdnd11an1n64x5 FILLER_103_2076 ();
 b15zdnd11an1n64x5 FILLER_103_2140 ();
 b15zdnd11an1n64x5 FILLER_103_2204 ();
 b15zdnd11an1n16x5 FILLER_103_2268 ();
 b15zdnd11an1n64x5 FILLER_104_8 ();
 b15zdnd11an1n64x5 FILLER_104_72 ();
 b15zdnd11an1n64x5 FILLER_104_136 ();
 b15zdnd11an1n64x5 FILLER_104_200 ();
 b15zdnd11an1n64x5 FILLER_104_264 ();
 b15zdnd11an1n32x5 FILLER_104_328 ();
 b15zdnd11an1n04x5 FILLER_104_360 ();
 b15zdnd00an1n01x5 FILLER_104_364 ();
 b15zdnd11an1n64x5 FILLER_104_374 ();
 b15zdnd11an1n64x5 FILLER_104_438 ();
 b15zdnd11an1n64x5 FILLER_104_502 ();
 b15zdnd11an1n32x5 FILLER_104_566 ();
 b15zdnd11an1n16x5 FILLER_104_598 ();
 b15zdnd11an1n08x5 FILLER_104_614 ();
 b15zdnd11an1n04x5 FILLER_104_622 ();
 b15zdnd11an1n64x5 FILLER_104_629 ();
 b15zdnd11an1n16x5 FILLER_104_693 ();
 b15zdnd11an1n08x5 FILLER_104_709 ();
 b15zdnd00an1n01x5 FILLER_104_717 ();
 b15zdnd11an1n64x5 FILLER_104_726 ();
 b15zdnd11an1n64x5 FILLER_104_790 ();
 b15zdnd11an1n16x5 FILLER_104_854 ();
 b15zdnd11an1n04x5 FILLER_104_870 ();
 b15zdnd00an1n01x5 FILLER_104_874 ();
 b15zdnd11an1n04x5 FILLER_104_927 ();
 b15zdnd11an1n64x5 FILLER_104_942 ();
 b15zdnd11an1n32x5 FILLER_104_1006 ();
 b15zdnd11an1n64x5 FILLER_104_1048 ();
 b15zdnd11an1n08x5 FILLER_104_1112 ();
 b15zdnd11an1n04x5 FILLER_104_1120 ();
 b15zdnd11an1n64x5 FILLER_104_1176 ();
 b15zdnd11an1n32x5 FILLER_104_1240 ();
 b15zdnd11an1n16x5 FILLER_104_1272 ();
 b15zdnd11an1n64x5 FILLER_104_1292 ();
 b15zdnd11an1n32x5 FILLER_104_1356 ();
 b15zdnd11an1n16x5 FILLER_104_1388 ();
 b15zdnd11an1n04x5 FILLER_104_1404 ();
 b15zdnd11an1n04x5 FILLER_104_1411 ();
 b15zdnd11an1n08x5 FILLER_104_1418 ();
 b15zdnd00an1n01x5 FILLER_104_1426 ();
 b15zdnd11an1n64x5 FILLER_104_1435 ();
 b15zdnd11an1n32x5 FILLER_104_1499 ();
 b15zdnd11an1n04x5 FILLER_104_1531 ();
 b15zdnd00an1n02x5 FILLER_104_1535 ();
 b15zdnd11an1n04x5 FILLER_104_1540 ();
 b15zdnd11an1n04x5 FILLER_104_1547 ();
 b15zdnd11an1n64x5 FILLER_104_1554 ();
 b15zdnd11an1n64x5 FILLER_104_1618 ();
 b15zdnd11an1n64x5 FILLER_104_1682 ();
 b15zdnd11an1n64x5 FILLER_104_1746 ();
 b15zdnd11an1n16x5 FILLER_104_1810 ();
 b15zdnd11an1n08x5 FILLER_104_1826 ();
 b15zdnd11an1n04x5 FILLER_104_1834 ();
 b15zdnd00an1n01x5 FILLER_104_1838 ();
 b15zdnd11an1n08x5 FILLER_104_1845 ();
 b15zdnd00an1n02x5 FILLER_104_1853 ();
 b15zdnd11an1n64x5 FILLER_104_1897 ();
 b15zdnd11an1n64x5 FILLER_104_1961 ();
 b15zdnd11an1n64x5 FILLER_104_2025 ();
 b15zdnd11an1n64x5 FILLER_104_2089 ();
 b15zdnd00an1n01x5 FILLER_104_2153 ();
 b15zdnd11an1n64x5 FILLER_104_2162 ();
 b15zdnd11an1n32x5 FILLER_104_2226 ();
 b15zdnd11an1n16x5 FILLER_104_2258 ();
 b15zdnd00an1n02x5 FILLER_104_2274 ();
 b15zdnd11an1n64x5 FILLER_105_0 ();
 b15zdnd11an1n64x5 FILLER_105_64 ();
 b15zdnd11an1n64x5 FILLER_105_128 ();
 b15zdnd11an1n64x5 FILLER_105_192 ();
 b15zdnd11an1n64x5 FILLER_105_256 ();
 b15zdnd11an1n64x5 FILLER_105_320 ();
 b15zdnd11an1n64x5 FILLER_105_384 ();
 b15zdnd11an1n64x5 FILLER_105_448 ();
 b15zdnd11an1n64x5 FILLER_105_512 ();
 b15zdnd11an1n32x5 FILLER_105_576 ();
 b15zdnd11an1n16x5 FILLER_105_608 ();
 b15zdnd11an1n08x5 FILLER_105_624 ();
 b15zdnd00an1n01x5 FILLER_105_632 ();
 b15zdnd11an1n64x5 FILLER_105_647 ();
 b15zdnd11an1n64x5 FILLER_105_711 ();
 b15zdnd11an1n64x5 FILLER_105_775 ();
 b15zdnd11an1n64x5 FILLER_105_839 ();
 b15zdnd11an1n16x5 FILLER_105_903 ();
 b15zdnd11an1n08x5 FILLER_105_919 ();
 b15zdnd00an1n02x5 FILLER_105_927 ();
 b15zdnd11an1n64x5 FILLER_105_933 ();
 b15zdnd11an1n32x5 FILLER_105_997 ();
 b15zdnd11an1n08x5 FILLER_105_1029 ();
 b15zdnd11an1n64x5 FILLER_105_1044 ();
 b15zdnd11an1n16x5 FILLER_105_1108 ();
 b15zdnd11an1n04x5 FILLER_105_1124 ();
 b15zdnd00an1n02x5 FILLER_105_1128 ();
 b15zdnd11an1n64x5 FILLER_105_1150 ();
 b15zdnd11an1n16x5 FILLER_105_1214 ();
 b15zdnd11an1n08x5 FILLER_105_1230 ();
 b15zdnd00an1n02x5 FILLER_105_1238 ();
 b15zdnd00an1n01x5 FILLER_105_1240 ();
 b15zdnd11an1n64x5 FILLER_105_1249 ();
 b15zdnd11an1n64x5 FILLER_105_1313 ();
 b15zdnd11an1n04x5 FILLER_105_1377 ();
 b15zdnd00an1n02x5 FILLER_105_1381 ();
 b15zdnd00an1n01x5 FILLER_105_1383 ();
 b15zdnd11an1n64x5 FILLER_105_1436 ();
 b15zdnd11an1n16x5 FILLER_105_1500 ();
 b15zdnd00an1n02x5 FILLER_105_1516 ();
 b15zdnd00an1n01x5 FILLER_105_1518 ();
 b15zdnd11an1n64x5 FILLER_105_1571 ();
 b15zdnd11an1n16x5 FILLER_105_1635 ();
 b15zdnd00an1n01x5 FILLER_105_1651 ();
 b15zdnd11an1n64x5 FILLER_105_1656 ();
 b15zdnd11an1n64x5 FILLER_105_1720 ();
 b15zdnd11an1n32x5 FILLER_105_1784 ();
 b15zdnd11an1n16x5 FILLER_105_1816 ();
 b15zdnd11an1n08x5 FILLER_105_1832 ();
 b15zdnd00an1n02x5 FILLER_105_1840 ();
 b15zdnd11an1n04x5 FILLER_105_1845 ();
 b15zdnd11an1n08x5 FILLER_105_1855 ();
 b15zdnd00an1n02x5 FILLER_105_1863 ();
 b15zdnd11an1n64x5 FILLER_105_1907 ();
 b15zdnd11an1n64x5 FILLER_105_1971 ();
 b15zdnd11an1n64x5 FILLER_105_2035 ();
 b15zdnd11an1n64x5 FILLER_105_2099 ();
 b15zdnd11an1n64x5 FILLER_105_2163 ();
 b15zdnd11an1n32x5 FILLER_105_2227 ();
 b15zdnd11an1n16x5 FILLER_105_2259 ();
 b15zdnd11an1n08x5 FILLER_105_2275 ();
 b15zdnd00an1n01x5 FILLER_105_2283 ();
 b15zdnd11an1n64x5 FILLER_106_8 ();
 b15zdnd11an1n64x5 FILLER_106_72 ();
 b15zdnd11an1n64x5 FILLER_106_136 ();
 b15zdnd11an1n64x5 FILLER_106_200 ();
 b15zdnd11an1n64x5 FILLER_106_264 ();
 b15zdnd11an1n64x5 FILLER_106_328 ();
 b15zdnd11an1n64x5 FILLER_106_392 ();
 b15zdnd11an1n64x5 FILLER_106_456 ();
 b15zdnd11an1n64x5 FILLER_106_520 ();
 b15zdnd11an1n64x5 FILLER_106_584 ();
 b15zdnd11an1n16x5 FILLER_106_648 ();
 b15zdnd00an1n01x5 FILLER_106_664 ();
 b15zdnd11an1n32x5 FILLER_106_671 ();
 b15zdnd11an1n08x5 FILLER_106_703 ();
 b15zdnd11an1n04x5 FILLER_106_711 ();
 b15zdnd00an1n02x5 FILLER_106_715 ();
 b15zdnd00an1n01x5 FILLER_106_717 ();
 b15zdnd11an1n64x5 FILLER_106_726 ();
 b15zdnd11an1n64x5 FILLER_106_790 ();
 b15zdnd11an1n64x5 FILLER_106_854 ();
 b15zdnd11an1n32x5 FILLER_106_918 ();
 b15zdnd11an1n16x5 FILLER_106_950 ();
 b15zdnd11an1n08x5 FILLER_106_966 ();
 b15zdnd11an1n04x5 FILLER_106_974 ();
 b15zdnd11an1n32x5 FILLER_106_989 ();
 b15zdnd11an1n04x5 FILLER_106_1021 ();
 b15zdnd00an1n02x5 FILLER_106_1025 ();
 b15zdnd11an1n64x5 FILLER_106_1047 ();
 b15zdnd11an1n16x5 FILLER_106_1111 ();
 b15zdnd00an1n02x5 FILLER_106_1127 ();
 b15zdnd00an1n01x5 FILLER_106_1129 ();
 b15zdnd11an1n64x5 FILLER_106_1142 ();
 b15zdnd11an1n64x5 FILLER_106_1206 ();
 b15zdnd11an1n32x5 FILLER_106_1270 ();
 b15zdnd11an1n16x5 FILLER_106_1302 ();
 b15zdnd11an1n04x5 FILLER_106_1318 ();
 b15zdnd11an1n64x5 FILLER_106_1326 ();
 b15zdnd11an1n32x5 FILLER_106_1390 ();
 b15zdnd11an1n08x5 FILLER_106_1422 ();
 b15zdnd00an1n02x5 FILLER_106_1430 ();
 b15zdnd00an1n01x5 FILLER_106_1432 ();
 b15zdnd11an1n64x5 FILLER_106_1436 ();
 b15zdnd11an1n32x5 FILLER_106_1500 ();
 b15zdnd11an1n08x5 FILLER_106_1532 ();
 b15zdnd11an1n64x5 FILLER_106_1567 ();
 b15zdnd11an1n64x5 FILLER_106_1631 ();
 b15zdnd11an1n64x5 FILLER_106_1695 ();
 b15zdnd11an1n64x5 FILLER_106_1759 ();
 b15zdnd11an1n16x5 FILLER_106_1823 ();
 b15zdnd11an1n08x5 FILLER_106_1839 ();
 b15zdnd11an1n04x5 FILLER_106_1847 ();
 b15zdnd00an1n01x5 FILLER_106_1851 ();
 b15zdnd11an1n04x5 FILLER_106_1856 ();
 b15zdnd11an1n64x5 FILLER_106_1864 ();
 b15zdnd11an1n64x5 FILLER_106_1928 ();
 b15zdnd11an1n64x5 FILLER_106_1992 ();
 b15zdnd11an1n64x5 FILLER_106_2056 ();
 b15zdnd11an1n32x5 FILLER_106_2120 ();
 b15zdnd00an1n02x5 FILLER_106_2152 ();
 b15zdnd11an1n64x5 FILLER_106_2162 ();
 b15zdnd11an1n32x5 FILLER_106_2226 ();
 b15zdnd11an1n16x5 FILLER_106_2258 ();
 b15zdnd00an1n02x5 FILLER_106_2274 ();
 b15zdnd11an1n64x5 FILLER_107_0 ();
 b15zdnd11an1n64x5 FILLER_107_64 ();
 b15zdnd11an1n64x5 FILLER_107_128 ();
 b15zdnd11an1n64x5 FILLER_107_192 ();
 b15zdnd11an1n64x5 FILLER_107_256 ();
 b15zdnd11an1n64x5 FILLER_107_320 ();
 b15zdnd11an1n64x5 FILLER_107_384 ();
 b15zdnd11an1n64x5 FILLER_107_448 ();
 b15zdnd11an1n64x5 FILLER_107_512 ();
 b15zdnd11an1n64x5 FILLER_107_576 ();
 b15zdnd11an1n16x5 FILLER_107_640 ();
 b15zdnd00an1n01x5 FILLER_107_656 ();
 b15zdnd11an1n64x5 FILLER_107_663 ();
 b15zdnd11an1n64x5 FILLER_107_727 ();
 b15zdnd11an1n64x5 FILLER_107_791 ();
 b15zdnd11an1n64x5 FILLER_107_855 ();
 b15zdnd11an1n64x5 FILLER_107_919 ();
 b15zdnd11an1n64x5 FILLER_107_983 ();
 b15zdnd11an1n64x5 FILLER_107_1047 ();
 b15zdnd11an1n64x5 FILLER_107_1111 ();
 b15zdnd11an1n64x5 FILLER_107_1175 ();
 b15zdnd11an1n16x5 FILLER_107_1239 ();
 b15zdnd11an1n08x5 FILLER_107_1255 ();
 b15zdnd11an1n04x5 FILLER_107_1263 ();
 b15zdnd00an1n02x5 FILLER_107_1267 ();
 b15zdnd11an1n64x5 FILLER_107_1275 ();
 b15zdnd11an1n64x5 FILLER_107_1339 ();
 b15zdnd11an1n04x5 FILLER_107_1403 ();
 b15zdnd00an1n02x5 FILLER_107_1407 ();
 b15zdnd11an1n04x5 FILLER_107_1461 ();
 b15zdnd11an1n32x5 FILLER_107_1474 ();
 b15zdnd11an1n08x5 FILLER_107_1506 ();
 b15zdnd00an1n02x5 FILLER_107_1514 ();
 b15zdnd11an1n16x5 FILLER_107_1525 ();
 b15zdnd11an1n04x5 FILLER_107_1541 ();
 b15zdnd00an1n01x5 FILLER_107_1545 ();
 b15zdnd11an1n32x5 FILLER_107_1598 ();
 b15zdnd11an1n08x5 FILLER_107_1630 ();
 b15zdnd11an1n64x5 FILLER_107_1642 ();
 b15zdnd11an1n32x5 FILLER_107_1706 ();
 b15zdnd11an1n16x5 FILLER_107_1738 ();
 b15zdnd11an1n08x5 FILLER_107_1754 ();
 b15zdnd11an1n64x5 FILLER_107_1804 ();
 b15zdnd11an1n64x5 FILLER_107_1868 ();
 b15zdnd11an1n64x5 FILLER_107_1932 ();
 b15zdnd11an1n64x5 FILLER_107_1996 ();
 b15zdnd11an1n64x5 FILLER_107_2060 ();
 b15zdnd11an1n64x5 FILLER_107_2124 ();
 b15zdnd11an1n64x5 FILLER_107_2188 ();
 b15zdnd11an1n32x5 FILLER_107_2252 ();
 b15zdnd11an1n64x5 FILLER_108_8 ();
 b15zdnd11an1n64x5 FILLER_108_72 ();
 b15zdnd11an1n64x5 FILLER_108_136 ();
 b15zdnd11an1n64x5 FILLER_108_200 ();
 b15zdnd11an1n64x5 FILLER_108_264 ();
 b15zdnd11an1n64x5 FILLER_108_328 ();
 b15zdnd11an1n64x5 FILLER_108_392 ();
 b15zdnd11an1n64x5 FILLER_108_456 ();
 b15zdnd11an1n64x5 FILLER_108_520 ();
 b15zdnd11an1n64x5 FILLER_108_584 ();
 b15zdnd11an1n08x5 FILLER_108_648 ();
 b15zdnd11an1n04x5 FILLER_108_656 ();
 b15zdnd00an1n02x5 FILLER_108_660 ();
 b15zdnd00an1n01x5 FILLER_108_662 ();
 b15zdnd11an1n32x5 FILLER_108_669 ();
 b15zdnd11an1n16x5 FILLER_108_701 ();
 b15zdnd00an1n01x5 FILLER_108_717 ();
 b15zdnd11an1n64x5 FILLER_108_726 ();
 b15zdnd11an1n16x5 FILLER_108_790 ();
 b15zdnd11an1n04x5 FILLER_108_806 ();
 b15zdnd00an1n01x5 FILLER_108_810 ();
 b15zdnd11an1n64x5 FILLER_108_819 ();
 b15zdnd11an1n64x5 FILLER_108_883 ();
 b15zdnd11an1n64x5 FILLER_108_947 ();
 b15zdnd11an1n64x5 FILLER_108_1011 ();
 b15zdnd11an1n64x5 FILLER_108_1075 ();
 b15zdnd11an1n32x5 FILLER_108_1139 ();
 b15zdnd11an1n08x5 FILLER_108_1171 ();
 b15zdnd11an1n04x5 FILLER_108_1179 ();
 b15zdnd11an1n64x5 FILLER_108_1186 ();
 b15zdnd11an1n16x5 FILLER_108_1250 ();
 b15zdnd11an1n08x5 FILLER_108_1266 ();
 b15zdnd11an1n04x5 FILLER_108_1274 ();
 b15zdnd11an1n64x5 FILLER_108_1281 ();
 b15zdnd11an1n32x5 FILLER_108_1345 ();
 b15zdnd11an1n16x5 FILLER_108_1377 ();
 b15zdnd11an1n08x5 FILLER_108_1393 ();
 b15zdnd11an1n04x5 FILLER_108_1401 ();
 b15zdnd00an1n01x5 FILLER_108_1405 ();
 b15zdnd11an1n16x5 FILLER_108_1458 ();
 b15zdnd11an1n04x5 FILLER_108_1474 ();
 b15zdnd00an1n02x5 FILLER_108_1478 ();
 b15zdnd11an1n08x5 FILLER_108_1488 ();
 b15zdnd11an1n04x5 FILLER_108_1496 ();
 b15zdnd00an1n01x5 FILLER_108_1500 ();
 b15zdnd11an1n16x5 FILLER_108_1510 ();
 b15zdnd11an1n08x5 FILLER_108_1526 ();
 b15zdnd00an1n02x5 FILLER_108_1534 ();
 b15zdnd00an1n01x5 FILLER_108_1536 ();
 b15zdnd11an1n08x5 FILLER_108_1540 ();
 b15zdnd11an1n04x5 FILLER_108_1548 ();
 b15zdnd00an1n01x5 FILLER_108_1552 ();
 b15zdnd11an1n64x5 FILLER_108_1605 ();
 b15zdnd11an1n64x5 FILLER_108_1669 ();
 b15zdnd11an1n04x5 FILLER_108_1733 ();
 b15zdnd00an1n01x5 FILLER_108_1737 ();
 b15zdnd11an1n64x5 FILLER_108_1780 ();
 b15zdnd11an1n64x5 FILLER_108_1844 ();
 b15zdnd11an1n64x5 FILLER_108_1908 ();
 b15zdnd11an1n64x5 FILLER_108_1972 ();
 b15zdnd11an1n64x5 FILLER_108_2036 ();
 b15zdnd11an1n32x5 FILLER_108_2100 ();
 b15zdnd11an1n16x5 FILLER_108_2132 ();
 b15zdnd11an1n04x5 FILLER_108_2148 ();
 b15zdnd00an1n02x5 FILLER_108_2152 ();
 b15zdnd11an1n64x5 FILLER_108_2162 ();
 b15zdnd11an1n16x5 FILLER_108_2226 ();
 b15zdnd11an1n08x5 FILLER_108_2242 ();
 b15zdnd00an1n02x5 FILLER_108_2250 ();
 b15zdnd11an1n16x5 FILLER_108_2258 ();
 b15zdnd00an1n02x5 FILLER_108_2274 ();
 b15zdnd11an1n16x5 FILLER_109_0 ();
 b15zdnd11an1n08x5 FILLER_109_16 ();
 b15zdnd00an1n02x5 FILLER_109_24 ();
 b15zdnd00an1n01x5 FILLER_109_26 ();
 b15zdnd11an1n04x5 FILLER_109_31 ();
 b15zdnd11an1n64x5 FILLER_109_40 ();
 b15zdnd11an1n64x5 FILLER_109_104 ();
 b15zdnd11an1n64x5 FILLER_109_168 ();
 b15zdnd11an1n64x5 FILLER_109_232 ();
 b15zdnd11an1n64x5 FILLER_109_296 ();
 b15zdnd11an1n64x5 FILLER_109_360 ();
 b15zdnd11an1n64x5 FILLER_109_424 ();
 b15zdnd11an1n64x5 FILLER_109_488 ();
 b15zdnd11an1n64x5 FILLER_109_552 ();
 b15zdnd11an1n64x5 FILLER_109_616 ();
 b15zdnd11an1n64x5 FILLER_109_680 ();
 b15zdnd11an1n64x5 FILLER_109_744 ();
 b15zdnd11an1n64x5 FILLER_109_808 ();
 b15zdnd11an1n64x5 FILLER_109_872 ();
 b15zdnd11an1n64x5 FILLER_109_936 ();
 b15zdnd11an1n64x5 FILLER_109_1000 ();
 b15zdnd11an1n64x5 FILLER_109_1064 ();
 b15zdnd11an1n64x5 FILLER_109_1128 ();
 b15zdnd11an1n64x5 FILLER_109_1192 ();
 b15zdnd11an1n08x5 FILLER_109_1256 ();
 b15zdnd11an1n04x5 FILLER_109_1264 ();
 b15zdnd00an1n02x5 FILLER_109_1268 ();
 b15zdnd00an1n01x5 FILLER_109_1270 ();
 b15zdnd11an1n04x5 FILLER_109_1284 ();
 b15zdnd00an1n02x5 FILLER_109_1288 ();
 b15zdnd00an1n01x5 FILLER_109_1290 ();
 b15zdnd11an1n64x5 FILLER_109_1297 ();
 b15zdnd11an1n32x5 FILLER_109_1361 ();
 b15zdnd11an1n16x5 FILLER_109_1393 ();
 b15zdnd11an1n08x5 FILLER_109_1409 ();
 b15zdnd11an1n04x5 FILLER_109_1417 ();
 b15zdnd00an1n02x5 FILLER_109_1421 ();
 b15zdnd00an1n01x5 FILLER_109_1423 ();
 b15zdnd11an1n04x5 FILLER_109_1427 ();
 b15zdnd11an1n04x5 FILLER_109_1434 ();
 b15zdnd11an1n04x5 FILLER_109_1441 ();
 b15zdnd11an1n64x5 FILLER_109_1448 ();
 b15zdnd11an1n32x5 FILLER_109_1512 ();
 b15zdnd11an1n16x5 FILLER_109_1544 ();
 b15zdnd00an1n02x5 FILLER_109_1560 ();
 b15zdnd11an1n04x5 FILLER_109_1565 ();
 b15zdnd11an1n04x5 FILLER_109_1572 ();
 b15zdnd11an1n04x5 FILLER_109_1579 ();
 b15zdnd11an1n64x5 FILLER_109_1586 ();
 b15zdnd11an1n64x5 FILLER_109_1650 ();
 b15zdnd11an1n64x5 FILLER_109_1714 ();
 b15zdnd11an1n64x5 FILLER_109_1778 ();
 b15zdnd11an1n64x5 FILLER_109_1842 ();
 b15zdnd11an1n64x5 FILLER_109_1906 ();
 b15zdnd11an1n64x5 FILLER_109_1970 ();
 b15zdnd11an1n64x5 FILLER_109_2034 ();
 b15zdnd11an1n08x5 FILLER_109_2098 ();
 b15zdnd00an1n02x5 FILLER_109_2106 ();
 b15zdnd11an1n64x5 FILLER_109_2160 ();
 b15zdnd11an1n32x5 FILLER_109_2224 ();
 b15zdnd11an1n16x5 FILLER_109_2256 ();
 b15zdnd11an1n08x5 FILLER_109_2272 ();
 b15zdnd11an1n04x5 FILLER_109_2280 ();
 b15zdnd00an1n02x5 FILLER_110_8 ();
 b15zdnd11an1n64x5 FILLER_110_52 ();
 b15zdnd11an1n64x5 FILLER_110_116 ();
 b15zdnd11an1n64x5 FILLER_110_180 ();
 b15zdnd11an1n64x5 FILLER_110_244 ();
 b15zdnd11an1n08x5 FILLER_110_308 ();
 b15zdnd00an1n02x5 FILLER_110_316 ();
 b15zdnd00an1n01x5 FILLER_110_318 ();
 b15zdnd11an1n64x5 FILLER_110_322 ();
 b15zdnd11an1n64x5 FILLER_110_386 ();
 b15zdnd11an1n64x5 FILLER_110_450 ();
 b15zdnd11an1n32x5 FILLER_110_514 ();
 b15zdnd00an1n01x5 FILLER_110_546 ();
 b15zdnd11an1n32x5 FILLER_110_552 ();
 b15zdnd00an1n02x5 FILLER_110_584 ();
 b15zdnd00an1n01x5 FILLER_110_586 ();
 b15zdnd11an1n64x5 FILLER_110_593 ();
 b15zdnd11an1n08x5 FILLER_110_657 ();
 b15zdnd00an1n01x5 FILLER_110_665 ();
 b15zdnd11an1n32x5 FILLER_110_672 ();
 b15zdnd11an1n08x5 FILLER_110_704 ();
 b15zdnd11an1n04x5 FILLER_110_712 ();
 b15zdnd00an1n02x5 FILLER_110_716 ();
 b15zdnd11an1n16x5 FILLER_110_726 ();
 b15zdnd11an1n04x5 FILLER_110_742 ();
 b15zdnd00an1n02x5 FILLER_110_746 ();
 b15zdnd00an1n01x5 FILLER_110_748 ();
 b15zdnd11an1n04x5 FILLER_110_752 ();
 b15zdnd11an1n64x5 FILLER_110_759 ();
 b15zdnd11an1n64x5 FILLER_110_823 ();
 b15zdnd11an1n64x5 FILLER_110_887 ();
 b15zdnd11an1n64x5 FILLER_110_951 ();
 b15zdnd11an1n64x5 FILLER_110_1015 ();
 b15zdnd11an1n64x5 FILLER_110_1079 ();
 b15zdnd11an1n32x5 FILLER_110_1143 ();
 b15zdnd00an1n01x5 FILLER_110_1175 ();
 b15zdnd11an1n04x5 FILLER_110_1179 ();
 b15zdnd11an1n64x5 FILLER_110_1197 ();
 b15zdnd11an1n64x5 FILLER_110_1261 ();
 b15zdnd11an1n64x5 FILLER_110_1325 ();
 b15zdnd11an1n32x5 FILLER_110_1389 ();
 b15zdnd11an1n08x5 FILLER_110_1421 ();
 b15zdnd11an1n04x5 FILLER_110_1429 ();
 b15zdnd00an1n01x5 FILLER_110_1433 ();
 b15zdnd11an1n64x5 FILLER_110_1437 ();
 b15zdnd11an1n64x5 FILLER_110_1501 ();
 b15zdnd11an1n04x5 FILLER_110_1565 ();
 b15zdnd00an1n02x5 FILLER_110_1569 ();
 b15zdnd11an1n04x5 FILLER_110_1574 ();
 b15zdnd11an1n64x5 FILLER_110_1581 ();
 b15zdnd11an1n64x5 FILLER_110_1645 ();
 b15zdnd11an1n64x5 FILLER_110_1709 ();
 b15zdnd11an1n64x5 FILLER_110_1773 ();
 b15zdnd11an1n64x5 FILLER_110_1837 ();
 b15zdnd11an1n64x5 FILLER_110_1901 ();
 b15zdnd11an1n64x5 FILLER_110_1965 ();
 b15zdnd11an1n64x5 FILLER_110_2029 ();
 b15zdnd11an1n32x5 FILLER_110_2093 ();
 b15zdnd00an1n01x5 FILLER_110_2125 ();
 b15zdnd11an1n04x5 FILLER_110_2129 ();
 b15zdnd11an1n16x5 FILLER_110_2136 ();
 b15zdnd00an1n02x5 FILLER_110_2152 ();
 b15zdnd11an1n64x5 FILLER_110_2162 ();
 b15zdnd11an1n32x5 FILLER_110_2226 ();
 b15zdnd11an1n16x5 FILLER_110_2258 ();
 b15zdnd00an1n02x5 FILLER_110_2274 ();
 b15zdnd11an1n64x5 FILLER_111_0 ();
 b15zdnd11an1n32x5 FILLER_111_64 ();
 b15zdnd11an1n16x5 FILLER_111_96 ();
 b15zdnd11an1n08x5 FILLER_111_154 ();
 b15zdnd11an1n32x5 FILLER_111_204 ();
 b15zdnd11an1n08x5 FILLER_111_236 ();
 b15zdnd00an1n02x5 FILLER_111_244 ();
 b15zdnd00an1n01x5 FILLER_111_246 ();
 b15zdnd11an1n32x5 FILLER_111_250 ();
 b15zdnd11an1n08x5 FILLER_111_282 ();
 b15zdnd00an1n02x5 FILLER_111_290 ();
 b15zdnd11an1n64x5 FILLER_111_344 ();
 b15zdnd11an1n32x5 FILLER_111_408 ();
 b15zdnd11an1n08x5 FILLER_111_440 ();
 b15zdnd00an1n02x5 FILLER_111_448 ();
 b15zdnd11an1n64x5 FILLER_111_502 ();
 b15zdnd11an1n32x5 FILLER_111_566 ();
 b15zdnd11an1n16x5 FILLER_111_598 ();
 b15zdnd00an1n01x5 FILLER_111_614 ();
 b15zdnd11an1n64x5 FILLER_111_618 ();
 b15zdnd11an1n32x5 FILLER_111_682 ();
 b15zdnd11an1n08x5 FILLER_111_714 ();
 b15zdnd11an1n04x5 FILLER_111_722 ();
 b15zdnd00an1n02x5 FILLER_111_726 ();
 b15zdnd00an1n01x5 FILLER_111_728 ();
 b15zdnd11an1n64x5 FILLER_111_781 ();
 b15zdnd11an1n64x5 FILLER_111_845 ();
 b15zdnd11an1n64x5 FILLER_111_909 ();
 b15zdnd11an1n64x5 FILLER_111_973 ();
 b15zdnd11an1n64x5 FILLER_111_1037 ();
 b15zdnd11an1n64x5 FILLER_111_1101 ();
 b15zdnd11an1n64x5 FILLER_111_1165 ();
 b15zdnd11an1n64x5 FILLER_111_1229 ();
 b15zdnd11an1n64x5 FILLER_111_1293 ();
 b15zdnd11an1n64x5 FILLER_111_1357 ();
 b15zdnd11an1n64x5 FILLER_111_1421 ();
 b15zdnd11an1n64x5 FILLER_111_1485 ();
 b15zdnd11an1n64x5 FILLER_111_1549 ();
 b15zdnd11an1n64x5 FILLER_111_1613 ();
 b15zdnd11an1n64x5 FILLER_111_1677 ();
 b15zdnd11an1n64x5 FILLER_111_1741 ();
 b15zdnd11an1n32x5 FILLER_111_1805 ();
 b15zdnd11an1n08x5 FILLER_111_1837 ();
 b15zdnd00an1n02x5 FILLER_111_1845 ();
 b15zdnd11an1n64x5 FILLER_111_1889 ();
 b15zdnd11an1n64x5 FILLER_111_1953 ();
 b15zdnd11an1n64x5 FILLER_111_2017 ();
 b15zdnd11an1n04x5 FILLER_111_2081 ();
 b15zdnd00an1n01x5 FILLER_111_2085 ();
 b15zdnd11an1n16x5 FILLER_111_2089 ();
 b15zdnd11an1n04x5 FILLER_111_2105 ();
 b15zdnd00an1n01x5 FILLER_111_2109 ();
 b15zdnd11an1n04x5 FILLER_111_2114 ();
 b15zdnd11an1n64x5 FILLER_111_2160 ();
 b15zdnd11an1n32x5 FILLER_111_2224 ();
 b15zdnd11an1n16x5 FILLER_111_2256 ();
 b15zdnd11an1n08x5 FILLER_111_2272 ();
 b15zdnd11an1n04x5 FILLER_111_2280 ();
 b15zdnd11an1n64x5 FILLER_112_8 ();
 b15zdnd11an1n64x5 FILLER_112_72 ();
 b15zdnd11an1n64x5 FILLER_112_136 ();
 b15zdnd11an1n16x5 FILLER_112_200 ();
 b15zdnd11an1n08x5 FILLER_112_216 ();
 b15zdnd11an1n04x5 FILLER_112_224 ();
 b15zdnd00an1n01x5 FILLER_112_228 ();
 b15zdnd11an1n32x5 FILLER_112_271 ();
 b15zdnd11an1n08x5 FILLER_112_303 ();
 b15zdnd11an1n04x5 FILLER_112_314 ();
 b15zdnd11an1n16x5 FILLER_112_321 ();
 b15zdnd11an1n08x5 FILLER_112_337 ();
 b15zdnd00an1n01x5 FILLER_112_345 ();
 b15zdnd11an1n64x5 FILLER_112_388 ();
 b15zdnd11an1n16x5 FILLER_112_452 ();
 b15zdnd00an1n02x5 FILLER_112_468 ();
 b15zdnd11an1n04x5 FILLER_112_473 ();
 b15zdnd11an1n04x5 FILLER_112_480 ();
 b15zdnd11an1n64x5 FILLER_112_487 ();
 b15zdnd11an1n64x5 FILLER_112_551 ();
 b15zdnd11an1n32x5 FILLER_112_615 ();
 b15zdnd11an1n16x5 FILLER_112_647 ();
 b15zdnd00an1n01x5 FILLER_112_663 ();
 b15zdnd11an1n32x5 FILLER_112_675 ();
 b15zdnd11an1n08x5 FILLER_112_707 ();
 b15zdnd00an1n02x5 FILLER_112_715 ();
 b15zdnd00an1n01x5 FILLER_112_717 ();
 b15zdnd11an1n16x5 FILLER_112_726 ();
 b15zdnd11an1n04x5 FILLER_112_742 ();
 b15zdnd00an1n01x5 FILLER_112_746 ();
 b15zdnd11an1n04x5 FILLER_112_750 ();
 b15zdnd11an1n64x5 FILLER_112_757 ();
 b15zdnd11an1n32x5 FILLER_112_821 ();
 b15zdnd11an1n16x5 FILLER_112_853 ();
 b15zdnd11an1n08x5 FILLER_112_869 ();
 b15zdnd00an1n01x5 FILLER_112_877 ();
 b15zdnd11an1n64x5 FILLER_112_881 ();
 b15zdnd11an1n64x5 FILLER_112_945 ();
 b15zdnd11an1n64x5 FILLER_112_1009 ();
 b15zdnd00an1n02x5 FILLER_112_1073 ();
 b15zdnd11an1n64x5 FILLER_112_1078 ();
 b15zdnd11an1n64x5 FILLER_112_1142 ();
 b15zdnd11an1n64x5 FILLER_112_1206 ();
 b15zdnd11an1n04x5 FILLER_112_1270 ();
 b15zdnd11an1n64x5 FILLER_112_1290 ();
 b15zdnd11an1n32x5 FILLER_112_1354 ();
 b15zdnd11an1n16x5 FILLER_112_1386 ();
 b15zdnd11an1n08x5 FILLER_112_1402 ();
 b15zdnd11an1n04x5 FILLER_112_1410 ();
 b15zdnd00an1n01x5 FILLER_112_1414 ();
 b15zdnd11an1n04x5 FILLER_112_1418 ();
 b15zdnd00an1n02x5 FILLER_112_1422 ();
 b15zdnd11an1n04x5 FILLER_112_1427 ();
 b15zdnd11an1n64x5 FILLER_112_1434 ();
 b15zdnd11an1n64x5 FILLER_112_1498 ();
 b15zdnd11an1n64x5 FILLER_112_1562 ();
 b15zdnd11an1n32x5 FILLER_112_1626 ();
 b15zdnd11an1n16x5 FILLER_112_1658 ();
 b15zdnd00an1n01x5 FILLER_112_1674 ();
 b15zdnd11an1n32x5 FILLER_112_1679 ();
 b15zdnd11an1n16x5 FILLER_112_1711 ();
 b15zdnd11an1n64x5 FILLER_112_1758 ();
 b15zdnd11an1n64x5 FILLER_112_1822 ();
 b15zdnd11an1n64x5 FILLER_112_1886 ();
 b15zdnd11an1n64x5 FILLER_112_1950 ();
 b15zdnd11an1n64x5 FILLER_112_2014 ();
 b15zdnd11an1n04x5 FILLER_112_2078 ();
 b15zdnd00an1n02x5 FILLER_112_2082 ();
 b15zdnd11an1n04x5 FILLER_112_2091 ();
 b15zdnd11an1n32x5 FILLER_112_2100 ();
 b15zdnd11an1n16x5 FILLER_112_2135 ();
 b15zdnd00an1n02x5 FILLER_112_2151 ();
 b15zdnd00an1n01x5 FILLER_112_2153 ();
 b15zdnd11an1n64x5 FILLER_112_2162 ();
 b15zdnd11an1n32x5 FILLER_112_2226 ();
 b15zdnd11an1n16x5 FILLER_112_2258 ();
 b15zdnd00an1n02x5 FILLER_112_2274 ();
 b15zdnd11an1n64x5 FILLER_113_0 ();
 b15zdnd11an1n64x5 FILLER_113_64 ();
 b15zdnd11an1n64x5 FILLER_113_128 ();
 b15zdnd11an1n32x5 FILLER_113_192 ();
 b15zdnd11an1n08x5 FILLER_113_224 ();
 b15zdnd11an1n04x5 FILLER_113_232 ();
 b15zdnd00an1n02x5 FILLER_113_236 ();
 b15zdnd00an1n01x5 FILLER_113_238 ();
 b15zdnd11an1n64x5 FILLER_113_281 ();
 b15zdnd11an1n32x5 FILLER_113_345 ();
 b15zdnd00an1n02x5 FILLER_113_377 ();
 b15zdnd11an1n32x5 FILLER_113_421 ();
 b15zdnd11an1n16x5 FILLER_113_453 ();
 b15zdnd11an1n08x5 FILLER_113_469 ();
 b15zdnd00an1n01x5 FILLER_113_477 ();
 b15zdnd11an1n64x5 FILLER_113_481 ();
 b15zdnd11an1n64x5 FILLER_113_545 ();
 b15zdnd11an1n64x5 FILLER_113_609 ();
 b15zdnd11an1n16x5 FILLER_113_673 ();
 b15zdnd11an1n08x5 FILLER_113_689 ();
 b15zdnd11an1n04x5 FILLER_113_697 ();
 b15zdnd00an1n02x5 FILLER_113_701 ();
 b15zdnd11an1n04x5 FILLER_113_723 ();
 b15zdnd11an1n64x5 FILLER_113_779 ();
 b15zdnd11an1n08x5 FILLER_113_843 ();
 b15zdnd00an1n01x5 FILLER_113_851 ();
 b15zdnd11an1n64x5 FILLER_113_904 ();
 b15zdnd11an1n64x5 FILLER_113_968 ();
 b15zdnd11an1n64x5 FILLER_113_1032 ();
 b15zdnd11an1n16x5 FILLER_113_1096 ();
 b15zdnd11an1n04x5 FILLER_113_1112 ();
 b15zdnd00an1n02x5 FILLER_113_1116 ();
 b15zdnd00an1n01x5 FILLER_113_1118 ();
 b15zdnd11an1n08x5 FILLER_113_1164 ();
 b15zdnd00an1n01x5 FILLER_113_1172 ();
 b15zdnd11an1n64x5 FILLER_113_1193 ();
 b15zdnd11an1n08x5 FILLER_113_1257 ();
 b15zdnd11an1n64x5 FILLER_113_1269 ();
 b15zdnd11an1n64x5 FILLER_113_1333 ();
 b15zdnd11an1n04x5 FILLER_113_1397 ();
 b15zdnd00an1n02x5 FILLER_113_1401 ();
 b15zdnd11an1n64x5 FILLER_113_1455 ();
 b15zdnd11an1n64x5 FILLER_113_1519 ();
 b15zdnd11an1n64x5 FILLER_113_1583 ();
 b15zdnd11an1n64x5 FILLER_113_1647 ();
 b15zdnd00an1n02x5 FILLER_113_1711 ();
 b15zdnd00an1n01x5 FILLER_113_1713 ();
 b15zdnd11an1n64x5 FILLER_113_1718 ();
 b15zdnd11an1n64x5 FILLER_113_1782 ();
 b15zdnd11an1n64x5 FILLER_113_1846 ();
 b15zdnd11an1n64x5 FILLER_113_1910 ();
 b15zdnd11an1n64x5 FILLER_113_1974 ();
 b15zdnd11an1n64x5 FILLER_113_2038 ();
 b15zdnd11an1n32x5 FILLER_113_2102 ();
 b15zdnd00an1n02x5 FILLER_113_2134 ();
 b15zdnd11an1n64x5 FILLER_113_2178 ();
 b15zdnd11an1n32x5 FILLER_113_2242 ();
 b15zdnd11an1n08x5 FILLER_113_2274 ();
 b15zdnd00an1n02x5 FILLER_113_2282 ();
 b15zdnd11an1n64x5 FILLER_114_8 ();
 b15zdnd11an1n64x5 FILLER_114_72 ();
 b15zdnd11an1n64x5 FILLER_114_136 ();
 b15zdnd11an1n08x5 FILLER_114_200 ();
 b15zdnd11an1n04x5 FILLER_114_208 ();
 b15zdnd11an1n04x5 FILLER_114_252 ();
 b15zdnd11an1n64x5 FILLER_114_298 ();
 b15zdnd11an1n64x5 FILLER_114_362 ();
 b15zdnd11an1n64x5 FILLER_114_426 ();
 b15zdnd11an1n16x5 FILLER_114_490 ();
 b15zdnd11an1n08x5 FILLER_114_506 ();
 b15zdnd00an1n02x5 FILLER_114_514 ();
 b15zdnd11an1n32x5 FILLER_114_547 ();
 b15zdnd11an1n04x5 FILLER_114_579 ();
 b15zdnd00an1n02x5 FILLER_114_583 ();
 b15zdnd11an1n08x5 FILLER_114_592 ();
 b15zdnd11an1n04x5 FILLER_114_600 ();
 b15zdnd00an1n02x5 FILLER_114_604 ();
 b15zdnd00an1n01x5 FILLER_114_606 ();
 b15zdnd11an1n64x5 FILLER_114_620 ();
 b15zdnd11an1n32x5 FILLER_114_684 ();
 b15zdnd00an1n02x5 FILLER_114_716 ();
 b15zdnd11an1n16x5 FILLER_114_726 ();
 b15zdnd00an1n02x5 FILLER_114_742 ();
 b15zdnd00an1n01x5 FILLER_114_744 ();
 b15zdnd11an1n04x5 FILLER_114_748 ();
 b15zdnd11an1n64x5 FILLER_114_755 ();
 b15zdnd11an1n32x5 FILLER_114_819 ();
 b15zdnd11an1n08x5 FILLER_114_851 ();
 b15zdnd00an1n02x5 FILLER_114_859 ();
 b15zdnd00an1n01x5 FILLER_114_861 ();
 b15zdnd11an1n64x5 FILLER_114_914 ();
 b15zdnd11an1n08x5 FILLER_114_978 ();
 b15zdnd00an1n01x5 FILLER_114_986 ();
 b15zdnd11an1n64x5 FILLER_114_991 ();
 b15zdnd11an1n64x5 FILLER_114_1055 ();
 b15zdnd11an1n32x5 FILLER_114_1119 ();
 b15zdnd11an1n08x5 FILLER_114_1151 ();
 b15zdnd00an1n02x5 FILLER_114_1159 ();
 b15zdnd00an1n01x5 FILLER_114_1161 ();
 b15zdnd11an1n64x5 FILLER_114_1176 ();
 b15zdnd11an1n16x5 FILLER_114_1240 ();
 b15zdnd11an1n04x5 FILLER_114_1256 ();
 b15zdnd00an1n02x5 FILLER_114_1260 ();
 b15zdnd00an1n01x5 FILLER_114_1262 ();
 b15zdnd11an1n04x5 FILLER_114_1266 ();
 b15zdnd11an1n64x5 FILLER_114_1273 ();
 b15zdnd11an1n64x5 FILLER_114_1337 ();
 b15zdnd11an1n64x5 FILLER_114_1401 ();
 b15zdnd11an1n64x5 FILLER_114_1465 ();
 b15zdnd11an1n64x5 FILLER_114_1529 ();
 b15zdnd11an1n64x5 FILLER_114_1593 ();
 b15zdnd11an1n64x5 FILLER_114_1657 ();
 b15zdnd11an1n64x5 FILLER_114_1721 ();
 b15zdnd11an1n32x5 FILLER_114_1785 ();
 b15zdnd11an1n16x5 FILLER_114_1817 ();
 b15zdnd11an1n08x5 FILLER_114_1833 ();
 b15zdnd11an1n04x5 FILLER_114_1841 ();
 b15zdnd11an1n64x5 FILLER_114_1887 ();
 b15zdnd11an1n64x5 FILLER_114_1951 ();
 b15zdnd11an1n64x5 FILLER_114_2015 ();
 b15zdnd11an1n64x5 FILLER_114_2079 ();
 b15zdnd11an1n08x5 FILLER_114_2143 ();
 b15zdnd00an1n02x5 FILLER_114_2151 ();
 b15zdnd00an1n01x5 FILLER_114_2153 ();
 b15zdnd11an1n64x5 FILLER_114_2162 ();
 b15zdnd11an1n32x5 FILLER_114_2226 ();
 b15zdnd11an1n16x5 FILLER_114_2258 ();
 b15zdnd00an1n02x5 FILLER_114_2274 ();
 b15zdnd11an1n08x5 FILLER_115_0 ();
 b15zdnd00an1n02x5 FILLER_115_8 ();
 b15zdnd11an1n08x5 FILLER_115_14 ();
 b15zdnd00an1n01x5 FILLER_115_22 ();
 b15zdnd11an1n64x5 FILLER_115_27 ();
 b15zdnd11an1n32x5 FILLER_115_91 ();
 b15zdnd11an1n16x5 FILLER_115_123 ();
 b15zdnd11an1n08x5 FILLER_115_139 ();
 b15zdnd00an1n01x5 FILLER_115_147 ();
 b15zdnd11an1n64x5 FILLER_115_190 ();
 b15zdnd00an1n02x5 FILLER_115_254 ();
 b15zdnd00an1n01x5 FILLER_115_256 ();
 b15zdnd11an1n64x5 FILLER_115_260 ();
 b15zdnd11an1n64x5 FILLER_115_324 ();
 b15zdnd11an1n64x5 FILLER_115_388 ();
 b15zdnd00an1n02x5 FILLER_115_452 ();
 b15zdnd11an1n04x5 FILLER_115_506 ();
 b15zdnd00an1n02x5 FILLER_115_510 ();
 b15zdnd11an1n64x5 FILLER_115_554 ();
 b15zdnd11an1n08x5 FILLER_115_618 ();
 b15zdnd11an1n04x5 FILLER_115_626 ();
 b15zdnd00an1n01x5 FILLER_115_630 ();
 b15zdnd11an1n64x5 FILLER_115_647 ();
 b15zdnd11an1n64x5 FILLER_115_711 ();
 b15zdnd11an1n64x5 FILLER_115_775 ();
 b15zdnd11an1n32x5 FILLER_115_839 ();
 b15zdnd11an1n04x5 FILLER_115_871 ();
 b15zdnd11an1n04x5 FILLER_115_878 ();
 b15zdnd11an1n04x5 FILLER_115_885 ();
 b15zdnd11an1n64x5 FILLER_115_892 ();
 b15zdnd11an1n64x5 FILLER_115_956 ();
 b15zdnd11an1n64x5 FILLER_115_1020 ();
 b15zdnd11an1n64x5 FILLER_115_1084 ();
 b15zdnd11an1n64x5 FILLER_115_1148 ();
 b15zdnd11an1n16x5 FILLER_115_1212 ();
 b15zdnd11an1n08x5 FILLER_115_1228 ();
 b15zdnd00an1n02x5 FILLER_115_1236 ();
 b15zdnd11an1n16x5 FILLER_115_1290 ();
 b15zdnd11an1n04x5 FILLER_115_1306 ();
 b15zdnd00an1n02x5 FILLER_115_1310 ();
 b15zdnd00an1n01x5 FILLER_115_1312 ();
 b15zdnd11an1n64x5 FILLER_115_1316 ();
 b15zdnd11an1n64x5 FILLER_115_1380 ();
 b15zdnd11an1n64x5 FILLER_115_1444 ();
 b15zdnd11an1n64x5 FILLER_115_1508 ();
 b15zdnd11an1n64x5 FILLER_115_1572 ();
 b15zdnd11an1n64x5 FILLER_115_1636 ();
 b15zdnd11an1n64x5 FILLER_115_1700 ();
 b15zdnd11an1n64x5 FILLER_115_1764 ();
 b15zdnd11an1n64x5 FILLER_115_1828 ();
 b15zdnd11an1n64x5 FILLER_115_1892 ();
 b15zdnd11an1n64x5 FILLER_115_1956 ();
 b15zdnd11an1n04x5 FILLER_115_2020 ();
 b15zdnd11an1n64x5 FILLER_115_2029 ();
 b15zdnd11an1n64x5 FILLER_115_2093 ();
 b15zdnd11an1n64x5 FILLER_115_2157 ();
 b15zdnd11an1n32x5 FILLER_115_2221 ();
 b15zdnd11an1n16x5 FILLER_115_2253 ();
 b15zdnd11an1n08x5 FILLER_115_2269 ();
 b15zdnd11an1n04x5 FILLER_115_2277 ();
 b15zdnd00an1n02x5 FILLER_115_2281 ();
 b15zdnd00an1n01x5 FILLER_115_2283 ();
 b15zdnd00an1n02x5 FILLER_116_8 ();
 b15zdnd11an1n64x5 FILLER_116_52 ();
 b15zdnd11an1n32x5 FILLER_116_116 ();
 b15zdnd00an1n02x5 FILLER_116_148 ();
 b15zdnd00an1n01x5 FILLER_116_150 ();
 b15zdnd11an1n64x5 FILLER_116_193 ();
 b15zdnd11an1n64x5 FILLER_116_257 ();
 b15zdnd11an1n64x5 FILLER_116_321 ();
 b15zdnd11an1n64x5 FILLER_116_385 ();
 b15zdnd11an1n16x5 FILLER_116_449 ();
 b15zdnd11an1n04x5 FILLER_116_465 ();
 b15zdnd00an1n02x5 FILLER_116_469 ();
 b15zdnd00an1n01x5 FILLER_116_471 ();
 b15zdnd11an1n04x5 FILLER_116_475 ();
 b15zdnd11an1n64x5 FILLER_116_482 ();
 b15zdnd11an1n64x5 FILLER_116_546 ();
 b15zdnd11an1n64x5 FILLER_116_610 ();
 b15zdnd11an1n32x5 FILLER_116_674 ();
 b15zdnd11an1n08x5 FILLER_116_706 ();
 b15zdnd11an1n04x5 FILLER_116_714 ();
 b15zdnd11an1n64x5 FILLER_116_726 ();
 b15zdnd11an1n04x5 FILLER_116_790 ();
 b15zdnd11an1n32x5 FILLER_116_803 ();
 b15zdnd11an1n08x5 FILLER_116_835 ();
 b15zdnd11an1n04x5 FILLER_116_843 ();
 b15zdnd00an1n02x5 FILLER_116_847 ();
 b15zdnd11an1n16x5 FILLER_116_858 ();
 b15zdnd00an1n02x5 FILLER_116_874 ();
 b15zdnd00an1n01x5 FILLER_116_876 ();
 b15zdnd11an1n04x5 FILLER_116_880 ();
 b15zdnd11an1n64x5 FILLER_116_887 ();
 b15zdnd11an1n32x5 FILLER_116_951 ();
 b15zdnd11an1n16x5 FILLER_116_983 ();
 b15zdnd11an1n64x5 FILLER_116_1003 ();
 b15zdnd11an1n64x5 FILLER_116_1067 ();
 b15zdnd11an1n16x5 FILLER_116_1131 ();
 b15zdnd11an1n08x5 FILLER_116_1147 ();
 b15zdnd00an1n02x5 FILLER_116_1155 ();
 b15zdnd11an1n08x5 FILLER_116_1171 ();
 b15zdnd00an1n01x5 FILLER_116_1179 ();
 b15zdnd11an1n04x5 FILLER_116_1196 ();
 b15zdnd11an1n16x5 FILLER_116_1242 ();
 b15zdnd11an1n04x5 FILLER_116_1258 ();
 b15zdnd00an1n02x5 FILLER_116_1262 ();
 b15zdnd11an1n32x5 FILLER_116_1267 ();
 b15zdnd11an1n08x5 FILLER_116_1299 ();
 b15zdnd11an1n04x5 FILLER_116_1307 ();
 b15zdnd00an1n02x5 FILLER_116_1311 ();
 b15zdnd11an1n64x5 FILLER_116_1327 ();
 b15zdnd11an1n32x5 FILLER_116_1391 ();
 b15zdnd11an1n16x5 FILLER_116_1423 ();
 b15zdnd00an1n02x5 FILLER_116_1439 ();
 b15zdnd00an1n01x5 FILLER_116_1441 ();
 b15zdnd11an1n64x5 FILLER_116_1450 ();
 b15zdnd11an1n64x5 FILLER_116_1514 ();
 b15zdnd11an1n64x5 FILLER_116_1578 ();
 b15zdnd11an1n64x5 FILLER_116_1642 ();
 b15zdnd11an1n32x5 FILLER_116_1706 ();
 b15zdnd11an1n16x5 FILLER_116_1738 ();
 b15zdnd11an1n08x5 FILLER_116_1754 ();
 b15zdnd00an1n02x5 FILLER_116_1762 ();
 b15zdnd11an1n64x5 FILLER_116_1767 ();
 b15zdnd11an1n64x5 FILLER_116_1831 ();
 b15zdnd11an1n64x5 FILLER_116_1895 ();
 b15zdnd11an1n32x5 FILLER_116_1959 ();
 b15zdnd11an1n16x5 FILLER_116_1991 ();
 b15zdnd00an1n01x5 FILLER_116_2007 ();
 b15zdnd11an1n04x5 FILLER_116_2017 ();
 b15zdnd11an1n64x5 FILLER_116_2031 ();
 b15zdnd11an1n32x5 FILLER_116_2095 ();
 b15zdnd11an1n16x5 FILLER_116_2127 ();
 b15zdnd11an1n08x5 FILLER_116_2143 ();
 b15zdnd00an1n02x5 FILLER_116_2151 ();
 b15zdnd00an1n01x5 FILLER_116_2153 ();
 b15zdnd11an1n64x5 FILLER_116_2162 ();
 b15zdnd11an1n32x5 FILLER_116_2226 ();
 b15zdnd11an1n16x5 FILLER_116_2258 ();
 b15zdnd00an1n02x5 FILLER_116_2274 ();
 b15zdnd11an1n04x5 FILLER_117_0 ();
 b15zdnd00an1n02x5 FILLER_117_4 ();
 b15zdnd00an1n01x5 FILLER_117_6 ();
 b15zdnd11an1n64x5 FILLER_117_49 ();
 b15zdnd11an1n64x5 FILLER_117_113 ();
 b15zdnd11an1n32x5 FILLER_117_177 ();
 b15zdnd11an1n08x5 FILLER_117_209 ();
 b15zdnd11an1n04x5 FILLER_117_217 ();
 b15zdnd00an1n01x5 FILLER_117_221 ();
 b15zdnd11an1n64x5 FILLER_117_226 ();
 b15zdnd11an1n64x5 FILLER_117_290 ();
 b15zdnd11an1n64x5 FILLER_117_354 ();
 b15zdnd11an1n32x5 FILLER_117_418 ();
 b15zdnd11an1n16x5 FILLER_117_450 ();
 b15zdnd11an1n04x5 FILLER_117_466 ();
 b15zdnd00an1n01x5 FILLER_117_470 ();
 b15zdnd11an1n64x5 FILLER_117_482 ();
 b15zdnd11an1n64x5 FILLER_117_546 ();
 b15zdnd11an1n64x5 FILLER_117_610 ();
 b15zdnd11an1n64x5 FILLER_117_674 ();
 b15zdnd11an1n64x5 FILLER_117_738 ();
 b15zdnd11an1n64x5 FILLER_117_802 ();
 b15zdnd11an1n64x5 FILLER_117_866 ();
 b15zdnd11an1n64x5 FILLER_117_930 ();
 b15zdnd11an1n32x5 FILLER_117_994 ();
 b15zdnd11an1n16x5 FILLER_117_1026 ();
 b15zdnd11an1n04x5 FILLER_117_1042 ();
 b15zdnd11an1n16x5 FILLER_117_1053 ();
 b15zdnd11an1n08x5 FILLER_117_1069 ();
 b15zdnd00an1n01x5 FILLER_117_1077 ();
 b15zdnd11an1n64x5 FILLER_117_1092 ();
 b15zdnd11an1n64x5 FILLER_117_1156 ();
 b15zdnd11an1n64x5 FILLER_117_1220 ();
 b15zdnd11an1n32x5 FILLER_117_1284 ();
 b15zdnd00an1n01x5 FILLER_117_1316 ();
 b15zdnd11an1n64x5 FILLER_117_1320 ();
 b15zdnd11an1n64x5 FILLER_117_1384 ();
 b15zdnd11an1n64x5 FILLER_117_1448 ();
 b15zdnd11an1n64x5 FILLER_117_1512 ();
 b15zdnd11an1n64x5 FILLER_117_1576 ();
 b15zdnd11an1n16x5 FILLER_117_1640 ();
 b15zdnd11an1n08x5 FILLER_117_1656 ();
 b15zdnd11an1n04x5 FILLER_117_1664 ();
 b15zdnd11an1n32x5 FILLER_117_1678 ();
 b15zdnd11an1n16x5 FILLER_117_1710 ();
 b15zdnd11an1n08x5 FILLER_117_1726 ();
 b15zdnd11an1n04x5 FILLER_117_1734 ();
 b15zdnd11an1n64x5 FILLER_117_1790 ();
 b15zdnd11an1n64x5 FILLER_117_1854 ();
 b15zdnd11an1n64x5 FILLER_117_1918 ();
 b15zdnd11an1n16x5 FILLER_117_1982 ();
 b15zdnd11an1n08x5 FILLER_117_1998 ();
 b15zdnd00an1n01x5 FILLER_117_2006 ();
 b15zdnd11an1n04x5 FILLER_117_2020 ();
 b15zdnd00an1n01x5 FILLER_117_2024 ();
 b15zdnd11an1n64x5 FILLER_117_2067 ();
 b15zdnd11an1n64x5 FILLER_117_2131 ();
 b15zdnd11an1n64x5 FILLER_117_2195 ();
 b15zdnd11an1n16x5 FILLER_117_2259 ();
 b15zdnd11an1n08x5 FILLER_117_2275 ();
 b15zdnd00an1n01x5 FILLER_117_2283 ();
 b15zdnd11an1n64x5 FILLER_118_8 ();
 b15zdnd11an1n64x5 FILLER_118_72 ();
 b15zdnd11an1n64x5 FILLER_118_136 ();
 b15zdnd11an1n16x5 FILLER_118_200 ();
 b15zdnd00an1n02x5 FILLER_118_216 ();
 b15zdnd00an1n01x5 FILLER_118_218 ();
 b15zdnd11an1n04x5 FILLER_118_237 ();
 b15zdnd00an1n02x5 FILLER_118_241 ();
 b15zdnd11an1n64x5 FILLER_118_248 ();
 b15zdnd11an1n64x5 FILLER_118_312 ();
 b15zdnd11an1n64x5 FILLER_118_376 ();
 b15zdnd11an1n64x5 FILLER_118_440 ();
 b15zdnd11an1n64x5 FILLER_118_504 ();
 b15zdnd11an1n64x5 FILLER_118_568 ();
 b15zdnd11an1n64x5 FILLER_118_632 ();
 b15zdnd11an1n16x5 FILLER_118_696 ();
 b15zdnd11an1n04x5 FILLER_118_712 ();
 b15zdnd00an1n02x5 FILLER_118_716 ();
 b15zdnd11an1n16x5 FILLER_118_726 ();
 b15zdnd11an1n08x5 FILLER_118_742 ();
 b15zdnd00an1n02x5 FILLER_118_750 ();
 b15zdnd00an1n01x5 FILLER_118_752 ();
 b15zdnd11an1n64x5 FILLER_118_756 ();
 b15zdnd11an1n08x5 FILLER_118_820 ();
 b15zdnd11an1n04x5 FILLER_118_828 ();
 b15zdnd00an1n02x5 FILLER_118_832 ();
 b15zdnd11an1n64x5 FILLER_118_843 ();
 b15zdnd11an1n64x5 FILLER_118_907 ();
 b15zdnd11an1n64x5 FILLER_118_971 ();
 b15zdnd11an1n32x5 FILLER_118_1035 ();
 b15zdnd11an1n04x5 FILLER_118_1067 ();
 b15zdnd00an1n01x5 FILLER_118_1071 ();
 b15zdnd11an1n04x5 FILLER_118_1085 ();
 b15zdnd11an1n64x5 FILLER_118_1092 ();
 b15zdnd11an1n64x5 FILLER_118_1156 ();
 b15zdnd11an1n64x5 FILLER_118_1220 ();
 b15zdnd11an1n16x5 FILLER_118_1284 ();
 b15zdnd00an1n02x5 FILLER_118_1300 ();
 b15zdnd00an1n01x5 FILLER_118_1302 ();
 b15zdnd11an1n64x5 FILLER_118_1317 ();
 b15zdnd11an1n64x5 FILLER_118_1381 ();
 b15zdnd11an1n64x5 FILLER_118_1445 ();
 b15zdnd11an1n64x5 FILLER_118_1509 ();
 b15zdnd11an1n64x5 FILLER_118_1573 ();
 b15zdnd11an1n16x5 FILLER_118_1637 ();
 b15zdnd11an1n08x5 FILLER_118_1653 ();
 b15zdnd00an1n01x5 FILLER_118_1661 ();
 b15zdnd11an1n64x5 FILLER_118_1673 ();
 b15zdnd11an1n16x5 FILLER_118_1737 ();
 b15zdnd00an1n02x5 FILLER_118_1753 ();
 b15zdnd00an1n01x5 FILLER_118_1755 ();
 b15zdnd11an1n04x5 FILLER_118_1759 ();
 b15zdnd11an1n64x5 FILLER_118_1766 ();
 b15zdnd11an1n16x5 FILLER_118_1830 ();
 b15zdnd11an1n04x5 FILLER_118_1846 ();
 b15zdnd00an1n01x5 FILLER_118_1850 ();
 b15zdnd11an1n64x5 FILLER_118_1856 ();
 b15zdnd11an1n64x5 FILLER_118_1920 ();
 b15zdnd11an1n08x5 FILLER_118_1984 ();
 b15zdnd11an1n04x5 FILLER_118_1992 ();
 b15zdnd00an1n02x5 FILLER_118_1996 ();
 b15zdnd00an1n01x5 FILLER_118_1998 ();
 b15zdnd11an1n04x5 FILLER_118_2005 ();
 b15zdnd00an1n02x5 FILLER_118_2009 ();
 b15zdnd11an1n64x5 FILLER_118_2053 ();
 b15zdnd11an1n32x5 FILLER_118_2117 ();
 b15zdnd11an1n04x5 FILLER_118_2149 ();
 b15zdnd00an1n01x5 FILLER_118_2153 ();
 b15zdnd11an1n64x5 FILLER_118_2162 ();
 b15zdnd11an1n32x5 FILLER_118_2226 ();
 b15zdnd11an1n16x5 FILLER_118_2258 ();
 b15zdnd00an1n02x5 FILLER_118_2274 ();
 b15zdnd11an1n64x5 FILLER_119_0 ();
 b15zdnd11an1n64x5 FILLER_119_64 ();
 b15zdnd11an1n64x5 FILLER_119_128 ();
 b15zdnd11an1n32x5 FILLER_119_192 ();
 b15zdnd11an1n04x5 FILLER_119_224 ();
 b15zdnd00an1n02x5 FILLER_119_228 ();
 b15zdnd00an1n01x5 FILLER_119_230 ();
 b15zdnd11an1n64x5 FILLER_119_251 ();
 b15zdnd11an1n64x5 FILLER_119_315 ();
 b15zdnd11an1n64x5 FILLER_119_379 ();
 b15zdnd11an1n64x5 FILLER_119_443 ();
 b15zdnd11an1n64x5 FILLER_119_507 ();
 b15zdnd11an1n64x5 FILLER_119_571 ();
 b15zdnd11an1n64x5 FILLER_119_635 ();
 b15zdnd11an1n16x5 FILLER_119_699 ();
 b15zdnd11an1n08x5 FILLER_119_715 ();
 b15zdnd00an1n02x5 FILLER_119_723 ();
 b15zdnd00an1n01x5 FILLER_119_725 ();
 b15zdnd11an1n64x5 FILLER_119_778 ();
 b15zdnd11an1n16x5 FILLER_119_842 ();
 b15zdnd11an1n08x5 FILLER_119_858 ();
 b15zdnd00an1n02x5 FILLER_119_866 ();
 b15zdnd11an1n64x5 FILLER_119_895 ();
 b15zdnd11an1n64x5 FILLER_119_959 ();
 b15zdnd11an1n64x5 FILLER_119_1023 ();
 b15zdnd11an1n64x5 FILLER_119_1087 ();
 b15zdnd11an1n64x5 FILLER_119_1151 ();
 b15zdnd11an1n64x5 FILLER_119_1215 ();
 b15zdnd11an1n64x5 FILLER_119_1279 ();
 b15zdnd11an1n64x5 FILLER_119_1343 ();
 b15zdnd11an1n64x5 FILLER_119_1407 ();
 b15zdnd11an1n64x5 FILLER_119_1471 ();
 b15zdnd11an1n64x5 FILLER_119_1535 ();
 b15zdnd11an1n64x5 FILLER_119_1599 ();
 b15zdnd11an1n64x5 FILLER_119_1663 ();
 b15zdnd11an1n64x5 FILLER_119_1727 ();
 b15zdnd11an1n32x5 FILLER_119_1791 ();
 b15zdnd11an1n16x5 FILLER_119_1823 ();
 b15zdnd11an1n08x5 FILLER_119_1839 ();
 b15zdnd00an1n02x5 FILLER_119_1847 ();
 b15zdnd00an1n01x5 FILLER_119_1849 ();
 b15zdnd11an1n08x5 FILLER_119_1853 ();
 b15zdnd11an1n04x5 FILLER_119_1861 ();
 b15zdnd00an1n02x5 FILLER_119_1865 ();
 b15zdnd11an1n64x5 FILLER_119_1873 ();
 b15zdnd11an1n64x5 FILLER_119_1937 ();
 b15zdnd00an1n01x5 FILLER_119_2001 ();
 b15zdnd11an1n64x5 FILLER_119_2044 ();
 b15zdnd11an1n64x5 FILLER_119_2108 ();
 b15zdnd11an1n64x5 FILLER_119_2172 ();
 b15zdnd11an1n32x5 FILLER_119_2236 ();
 b15zdnd11an1n16x5 FILLER_119_2268 ();
 b15zdnd11an1n64x5 FILLER_120_8 ();
 b15zdnd11an1n64x5 FILLER_120_72 ();
 b15zdnd11an1n64x5 FILLER_120_136 ();
 b15zdnd11an1n16x5 FILLER_120_200 ();
 b15zdnd00an1n02x5 FILLER_120_216 ();
 b15zdnd11an1n64x5 FILLER_120_260 ();
 b15zdnd11an1n64x5 FILLER_120_324 ();
 b15zdnd11an1n64x5 FILLER_120_388 ();
 b15zdnd11an1n64x5 FILLER_120_452 ();
 b15zdnd11an1n32x5 FILLER_120_516 ();
 b15zdnd11an1n08x5 FILLER_120_548 ();
 b15zdnd11an1n04x5 FILLER_120_556 ();
 b15zdnd00an1n01x5 FILLER_120_560 ();
 b15zdnd11an1n64x5 FILLER_120_565 ();
 b15zdnd11an1n64x5 FILLER_120_629 ();
 b15zdnd11an1n16x5 FILLER_120_693 ();
 b15zdnd11an1n08x5 FILLER_120_709 ();
 b15zdnd00an1n01x5 FILLER_120_717 ();
 b15zdnd00an1n02x5 FILLER_120_726 ();
 b15zdnd11an1n64x5 FILLER_120_780 ();
 b15zdnd11an1n16x5 FILLER_120_844 ();
 b15zdnd11an1n04x5 FILLER_120_860 ();
 b15zdnd00an1n02x5 FILLER_120_864 ();
 b15zdnd00an1n01x5 FILLER_120_866 ();
 b15zdnd11an1n16x5 FILLER_120_870 ();
 b15zdnd11an1n04x5 FILLER_120_886 ();
 b15zdnd00an1n01x5 FILLER_120_890 ();
 b15zdnd11an1n64x5 FILLER_120_894 ();
 b15zdnd11an1n64x5 FILLER_120_958 ();
 b15zdnd11an1n32x5 FILLER_120_1022 ();
 b15zdnd11an1n08x5 FILLER_120_1054 ();
 b15zdnd11an1n04x5 FILLER_120_1062 ();
 b15zdnd00an1n02x5 FILLER_120_1066 ();
 b15zdnd00an1n01x5 FILLER_120_1068 ();
 b15zdnd11an1n64x5 FILLER_120_1083 ();
 b15zdnd00an1n02x5 FILLER_120_1147 ();
 b15zdnd00an1n01x5 FILLER_120_1149 ();
 b15zdnd11an1n64x5 FILLER_120_1192 ();
 b15zdnd11an1n64x5 FILLER_120_1256 ();
 b15zdnd00an1n01x5 FILLER_120_1320 ();
 b15zdnd11an1n64x5 FILLER_120_1337 ();
 b15zdnd11an1n64x5 FILLER_120_1401 ();
 b15zdnd11an1n64x5 FILLER_120_1465 ();
 b15zdnd11an1n64x5 FILLER_120_1529 ();
 b15zdnd11an1n64x5 FILLER_120_1593 ();
 b15zdnd11an1n64x5 FILLER_120_1657 ();
 b15zdnd11an1n64x5 FILLER_120_1721 ();
 b15zdnd11an1n64x5 FILLER_120_1785 ();
 b15zdnd11an1n08x5 FILLER_120_1849 ();
 b15zdnd11an1n04x5 FILLER_120_1857 ();
 b15zdnd11an1n04x5 FILLER_120_1864 ();
 b15zdnd00an1n02x5 FILLER_120_1868 ();
 b15zdnd11an1n08x5 FILLER_120_1910 ();
 b15zdnd00an1n02x5 FILLER_120_1918 ();
 b15zdnd00an1n01x5 FILLER_120_1920 ();
 b15zdnd11an1n32x5 FILLER_120_1930 ();
 b15zdnd11an1n08x5 FILLER_120_1962 ();
 b15zdnd11an1n04x5 FILLER_120_1970 ();
 b15zdnd00an1n01x5 FILLER_120_1974 ();
 b15zdnd11an1n04x5 FILLER_120_2027 ();
 b15zdnd11an1n64x5 FILLER_120_2035 ();
 b15zdnd11an1n32x5 FILLER_120_2099 ();
 b15zdnd11an1n16x5 FILLER_120_2131 ();
 b15zdnd11an1n04x5 FILLER_120_2147 ();
 b15zdnd00an1n02x5 FILLER_120_2151 ();
 b15zdnd00an1n01x5 FILLER_120_2153 ();
 b15zdnd11an1n64x5 FILLER_120_2162 ();
 b15zdnd11an1n32x5 FILLER_120_2226 ();
 b15zdnd11an1n16x5 FILLER_120_2258 ();
 b15zdnd00an1n02x5 FILLER_120_2274 ();
 b15zdnd11an1n64x5 FILLER_121_0 ();
 b15zdnd00an1n01x5 FILLER_121_64 ();
 b15zdnd11an1n64x5 FILLER_121_110 ();
 b15zdnd11an1n32x5 FILLER_121_174 ();
 b15zdnd11an1n04x5 FILLER_121_206 ();
 b15zdnd11an1n04x5 FILLER_121_250 ();
 b15zdnd00an1n01x5 FILLER_121_254 ();
 b15zdnd11an1n64x5 FILLER_121_258 ();
 b15zdnd11an1n64x5 FILLER_121_322 ();
 b15zdnd11an1n64x5 FILLER_121_386 ();
 b15zdnd11an1n64x5 FILLER_121_450 ();
 b15zdnd11an1n64x5 FILLER_121_514 ();
 b15zdnd11an1n16x5 FILLER_121_578 ();
 b15zdnd11an1n08x5 FILLER_121_594 ();
 b15zdnd00an1n02x5 FILLER_121_602 ();
 b15zdnd00an1n01x5 FILLER_121_604 ();
 b15zdnd11an1n64x5 FILLER_121_609 ();
 b15zdnd11an1n32x5 FILLER_121_673 ();
 b15zdnd11an1n16x5 FILLER_121_705 ();
 b15zdnd11an1n04x5 FILLER_121_721 ();
 b15zdnd00an1n02x5 FILLER_121_725 ();
 b15zdnd00an1n01x5 FILLER_121_727 ();
 b15zdnd11an1n08x5 FILLER_121_735 ();
 b15zdnd11an1n04x5 FILLER_121_743 ();
 b15zdnd11an1n04x5 FILLER_121_750 ();
 b15zdnd11an1n04x5 FILLER_121_757 ();
 b15zdnd11an1n64x5 FILLER_121_764 ();
 b15zdnd11an1n32x5 FILLER_121_828 ();
 b15zdnd11an1n16x5 FILLER_121_860 ();
 b15zdnd11an1n08x5 FILLER_121_876 ();
 b15zdnd00an1n02x5 FILLER_121_884 ();
 b15zdnd11an1n64x5 FILLER_121_889 ();
 b15zdnd11an1n32x5 FILLER_121_953 ();
 b15zdnd11an1n16x5 FILLER_121_985 ();
 b15zdnd00an1n02x5 FILLER_121_1001 ();
 b15zdnd00an1n01x5 FILLER_121_1003 ();
 b15zdnd11an1n16x5 FILLER_121_1008 ();
 b15zdnd00an1n02x5 FILLER_121_1024 ();
 b15zdnd00an1n01x5 FILLER_121_1026 ();
 b15zdnd11an1n04x5 FILLER_121_1046 ();
 b15zdnd00an1n02x5 FILLER_121_1050 ();
 b15zdnd11an1n32x5 FILLER_121_1063 ();
 b15zdnd11an1n08x5 FILLER_121_1095 ();
 b15zdnd00an1n01x5 FILLER_121_1103 ();
 b15zdnd11an1n08x5 FILLER_121_1112 ();
 b15zdnd11an1n64x5 FILLER_121_1124 ();
 b15zdnd11an1n64x5 FILLER_121_1188 ();
 b15zdnd11an1n64x5 FILLER_121_1252 ();
 b15zdnd11an1n08x5 FILLER_121_1316 ();
 b15zdnd11an1n64x5 FILLER_121_1340 ();
 b15zdnd11an1n64x5 FILLER_121_1404 ();
 b15zdnd11an1n64x5 FILLER_121_1468 ();
 b15zdnd11an1n64x5 FILLER_121_1532 ();
 b15zdnd11an1n64x5 FILLER_121_1596 ();
 b15zdnd11an1n64x5 FILLER_121_1660 ();
 b15zdnd11an1n64x5 FILLER_121_1724 ();
 b15zdnd11an1n64x5 FILLER_121_1788 ();
 b15zdnd00an1n02x5 FILLER_121_1852 ();
 b15zdnd00an1n01x5 FILLER_121_1854 ();
 b15zdnd11an1n16x5 FILLER_121_1897 ();
 b15zdnd00an1n01x5 FILLER_121_1913 ();
 b15zdnd11an1n64x5 FILLER_121_1917 ();
 b15zdnd11an1n16x5 FILLER_121_1981 ();
 b15zdnd00an1n02x5 FILLER_121_1997 ();
 b15zdnd11an1n04x5 FILLER_121_2002 ();
 b15zdnd00an1n02x5 FILLER_121_2006 ();
 b15zdnd00an1n01x5 FILLER_121_2008 ();
 b15zdnd11an1n04x5 FILLER_121_2016 ();
 b15zdnd11an1n64x5 FILLER_121_2025 ();
 b15zdnd11an1n64x5 FILLER_121_2089 ();
 b15zdnd11an1n64x5 FILLER_121_2153 ();
 b15zdnd11an1n64x5 FILLER_121_2217 ();
 b15zdnd00an1n02x5 FILLER_121_2281 ();
 b15zdnd00an1n01x5 FILLER_121_2283 ();
 b15zdnd11an1n64x5 FILLER_122_8 ();
 b15zdnd11an1n64x5 FILLER_122_72 ();
 b15zdnd11an1n64x5 FILLER_122_136 ();
 b15zdnd11an1n16x5 FILLER_122_200 ();
 b15zdnd11an1n08x5 FILLER_122_216 ();
 b15zdnd00an1n02x5 FILLER_122_224 ();
 b15zdnd00an1n01x5 FILLER_122_226 ();
 b15zdnd11an1n04x5 FILLER_122_240 ();
 b15zdnd00an1n01x5 FILLER_122_244 ();
 b15zdnd11an1n64x5 FILLER_122_248 ();
 b15zdnd11an1n16x5 FILLER_122_312 ();
 b15zdnd11an1n08x5 FILLER_122_328 ();
 b15zdnd00an1n01x5 FILLER_122_336 ();
 b15zdnd11an1n64x5 FILLER_122_340 ();
 b15zdnd11an1n64x5 FILLER_122_404 ();
 b15zdnd11an1n64x5 FILLER_122_468 ();
 b15zdnd11an1n64x5 FILLER_122_532 ();
 b15zdnd11an1n64x5 FILLER_122_596 ();
 b15zdnd11an1n32x5 FILLER_122_660 ();
 b15zdnd11an1n16x5 FILLER_122_692 ();
 b15zdnd11an1n08x5 FILLER_122_708 ();
 b15zdnd00an1n02x5 FILLER_122_716 ();
 b15zdnd11an1n16x5 FILLER_122_726 ();
 b15zdnd11an1n08x5 FILLER_122_742 ();
 b15zdnd00an1n01x5 FILLER_122_750 ();
 b15zdnd11an1n04x5 FILLER_122_754 ();
 b15zdnd11an1n64x5 FILLER_122_761 ();
 b15zdnd11an1n32x5 FILLER_122_825 ();
 b15zdnd11an1n16x5 FILLER_122_857 ();
 b15zdnd11an1n08x5 FILLER_122_873 ();
 b15zdnd00an1n02x5 FILLER_122_881 ();
 b15zdnd11an1n04x5 FILLER_122_886 ();
 b15zdnd11an1n32x5 FILLER_122_942 ();
 b15zdnd11an1n08x5 FILLER_122_974 ();
 b15zdnd11an1n04x5 FILLER_122_982 ();
 b15zdnd11an1n64x5 FILLER_122_992 ();
 b15zdnd11an1n32x5 FILLER_122_1056 ();
 b15zdnd11an1n16x5 FILLER_122_1088 ();
 b15zdnd11an1n04x5 FILLER_122_1104 ();
 b15zdnd00an1n02x5 FILLER_122_1108 ();
 b15zdnd11an1n04x5 FILLER_122_1114 ();
 b15zdnd11an1n64x5 FILLER_122_1124 ();
 b15zdnd11an1n64x5 FILLER_122_1188 ();
 b15zdnd11an1n64x5 FILLER_122_1252 ();
 b15zdnd11an1n64x5 FILLER_122_1316 ();
 b15zdnd11an1n64x5 FILLER_122_1380 ();
 b15zdnd11an1n64x5 FILLER_122_1444 ();
 b15zdnd11an1n32x5 FILLER_122_1508 ();
 b15zdnd11an1n16x5 FILLER_122_1540 ();
 b15zdnd11an1n08x5 FILLER_122_1556 ();
 b15zdnd11an1n64x5 FILLER_122_1568 ();
 b15zdnd11an1n64x5 FILLER_122_1632 ();
 b15zdnd11an1n64x5 FILLER_122_1696 ();
 b15zdnd11an1n64x5 FILLER_122_1760 ();
 b15zdnd11an1n08x5 FILLER_122_1824 ();
 b15zdnd11an1n04x5 FILLER_122_1832 ();
 b15zdnd11an1n16x5 FILLER_122_1888 ();
 b15zdnd00an1n02x5 FILLER_122_1904 ();
 b15zdnd11an1n64x5 FILLER_122_1909 ();
 b15zdnd11an1n16x5 FILLER_122_1973 ();
 b15zdnd11an1n04x5 FILLER_122_1989 ();
 b15zdnd00an1n02x5 FILLER_122_1993 ();
 b15zdnd00an1n01x5 FILLER_122_1995 ();
 b15zdnd11an1n04x5 FILLER_122_1999 ();
 b15zdnd00an1n02x5 FILLER_122_2003 ();
 b15zdnd00an1n01x5 FILLER_122_2005 ();
 b15zdnd11an1n64x5 FILLER_122_2009 ();
 b15zdnd11an1n64x5 FILLER_122_2073 ();
 b15zdnd11an1n16x5 FILLER_122_2137 ();
 b15zdnd00an1n01x5 FILLER_122_2153 ();
 b15zdnd11an1n64x5 FILLER_122_2162 ();
 b15zdnd11an1n32x5 FILLER_122_2226 ();
 b15zdnd11an1n16x5 FILLER_122_2258 ();
 b15zdnd00an1n02x5 FILLER_122_2274 ();
 b15zdnd11an1n64x5 FILLER_123_0 ();
 b15zdnd11an1n64x5 FILLER_123_64 ();
 b15zdnd11an1n64x5 FILLER_123_128 ();
 b15zdnd11an1n16x5 FILLER_123_192 ();
 b15zdnd11an1n08x5 FILLER_123_208 ();
 b15zdnd11an1n04x5 FILLER_123_216 ();
 b15zdnd00an1n02x5 FILLER_123_220 ();
 b15zdnd11an1n64x5 FILLER_123_237 ();
 b15zdnd11an1n08x5 FILLER_123_301 ();
 b15zdnd00an1n01x5 FILLER_123_309 ();
 b15zdnd11an1n04x5 FILLER_123_342 ();
 b15zdnd11an1n64x5 FILLER_123_349 ();
 b15zdnd11an1n64x5 FILLER_123_413 ();
 b15zdnd11an1n64x5 FILLER_123_477 ();
 b15zdnd11an1n64x5 FILLER_123_541 ();
 b15zdnd11an1n64x5 FILLER_123_605 ();
 b15zdnd11an1n64x5 FILLER_123_669 ();
 b15zdnd11an1n64x5 FILLER_123_733 ();
 b15zdnd11an1n16x5 FILLER_123_797 ();
 b15zdnd11an1n08x5 FILLER_123_813 ();
 b15zdnd11an1n04x5 FILLER_123_821 ();
 b15zdnd00an1n01x5 FILLER_123_825 ();
 b15zdnd11an1n32x5 FILLER_123_844 ();
 b15zdnd11an1n08x5 FILLER_123_876 ();
 b15zdnd11an1n32x5 FILLER_123_887 ();
 b15zdnd11an1n16x5 FILLER_123_919 ();
 b15zdnd11an1n08x5 FILLER_123_935 ();
 b15zdnd11an1n64x5 FILLER_123_950 ();
 b15zdnd11an1n64x5 FILLER_123_1014 ();
 b15zdnd11an1n64x5 FILLER_123_1078 ();
 b15zdnd11an1n64x5 FILLER_123_1142 ();
 b15zdnd11an1n64x5 FILLER_123_1206 ();
 b15zdnd11an1n64x5 FILLER_123_1270 ();
 b15zdnd11an1n64x5 FILLER_123_1334 ();
 b15zdnd11an1n64x5 FILLER_123_1398 ();
 b15zdnd11an1n64x5 FILLER_123_1462 ();
 b15zdnd11an1n32x5 FILLER_123_1526 ();
 b15zdnd11an1n08x5 FILLER_123_1558 ();
 b15zdnd11an1n04x5 FILLER_123_1566 ();
 b15zdnd00an1n01x5 FILLER_123_1570 ();
 b15zdnd11an1n64x5 FILLER_123_1575 ();
 b15zdnd11an1n64x5 FILLER_123_1639 ();
 b15zdnd11an1n64x5 FILLER_123_1703 ();
 b15zdnd11an1n64x5 FILLER_123_1767 ();
 b15zdnd11an1n16x5 FILLER_123_1831 ();
 b15zdnd11an1n04x5 FILLER_123_1847 ();
 b15zdnd00an1n02x5 FILLER_123_1851 ();
 b15zdnd00an1n01x5 FILLER_123_1853 ();
 b15zdnd11an1n04x5 FILLER_123_1857 ();
 b15zdnd11an1n16x5 FILLER_123_1864 ();
 b15zdnd00an1n02x5 FILLER_123_1880 ();
 b15zdnd00an1n01x5 FILLER_123_1882 ();
 b15zdnd11an1n64x5 FILLER_123_1925 ();
 b15zdnd11an1n64x5 FILLER_123_1989 ();
 b15zdnd11an1n64x5 FILLER_123_2053 ();
 b15zdnd11an1n64x5 FILLER_123_2117 ();
 b15zdnd11an1n64x5 FILLER_123_2181 ();
 b15zdnd11an1n32x5 FILLER_123_2245 ();
 b15zdnd11an1n04x5 FILLER_123_2277 ();
 b15zdnd00an1n02x5 FILLER_123_2281 ();
 b15zdnd00an1n01x5 FILLER_123_2283 ();
 b15zdnd11an1n64x5 FILLER_124_8 ();
 b15zdnd11an1n64x5 FILLER_124_72 ();
 b15zdnd11an1n64x5 FILLER_124_136 ();
 b15zdnd11an1n16x5 FILLER_124_200 ();
 b15zdnd11an1n08x5 FILLER_124_216 ();
 b15zdnd11an1n04x5 FILLER_124_224 ();
 b15zdnd11an1n64x5 FILLER_124_232 ();
 b15zdnd11an1n64x5 FILLER_124_296 ();
 b15zdnd11an1n64x5 FILLER_124_360 ();
 b15zdnd11an1n64x5 FILLER_124_424 ();
 b15zdnd11an1n64x5 FILLER_124_488 ();
 b15zdnd11an1n64x5 FILLER_124_552 ();
 b15zdnd11an1n64x5 FILLER_124_616 ();
 b15zdnd11an1n32x5 FILLER_124_680 ();
 b15zdnd11an1n04x5 FILLER_124_712 ();
 b15zdnd00an1n02x5 FILLER_124_716 ();
 b15zdnd11an1n64x5 FILLER_124_726 ();
 b15zdnd11an1n64x5 FILLER_124_790 ();
 b15zdnd00an1n02x5 FILLER_124_854 ();
 b15zdnd00an1n01x5 FILLER_124_856 ();
 b15zdnd11an1n32x5 FILLER_124_909 ();
 b15zdnd11an1n08x5 FILLER_124_941 ();
 b15zdnd11an1n32x5 FILLER_124_953 ();
 b15zdnd11an1n16x5 FILLER_124_985 ();
 b15zdnd11an1n08x5 FILLER_124_1001 ();
 b15zdnd11an1n04x5 FILLER_124_1009 ();
 b15zdnd11an1n64x5 FILLER_124_1017 ();
 b15zdnd11an1n64x5 FILLER_124_1081 ();
 b15zdnd11an1n64x5 FILLER_124_1145 ();
 b15zdnd11an1n04x5 FILLER_124_1209 ();
 b15zdnd11an1n64x5 FILLER_124_1216 ();
 b15zdnd11an1n64x5 FILLER_124_1280 ();
 b15zdnd11an1n64x5 FILLER_124_1344 ();
 b15zdnd11an1n64x5 FILLER_124_1408 ();
 b15zdnd11an1n64x5 FILLER_124_1472 ();
 b15zdnd11an1n64x5 FILLER_124_1536 ();
 b15zdnd11an1n64x5 FILLER_124_1600 ();
 b15zdnd11an1n64x5 FILLER_124_1664 ();
 b15zdnd11an1n64x5 FILLER_124_1728 ();
 b15zdnd11an1n64x5 FILLER_124_1792 ();
 b15zdnd11an1n16x5 FILLER_124_1856 ();
 b15zdnd11an1n04x5 FILLER_124_1872 ();
 b15zdnd00an1n01x5 FILLER_124_1876 ();
 b15zdnd11an1n64x5 FILLER_124_1892 ();
 b15zdnd11an1n64x5 FILLER_124_1956 ();
 b15zdnd11an1n64x5 FILLER_124_2020 ();
 b15zdnd11an1n64x5 FILLER_124_2084 ();
 b15zdnd11an1n04x5 FILLER_124_2148 ();
 b15zdnd00an1n02x5 FILLER_124_2152 ();
 b15zdnd11an1n32x5 FILLER_124_2162 ();
 b15zdnd11an1n08x5 FILLER_124_2194 ();
 b15zdnd11an1n04x5 FILLER_124_2202 ();
 b15zdnd00an1n02x5 FILLER_124_2206 ();
 b15zdnd11an1n32x5 FILLER_124_2216 ();
 b15zdnd11an1n16x5 FILLER_124_2248 ();
 b15zdnd11an1n08x5 FILLER_124_2264 ();
 b15zdnd11an1n04x5 FILLER_124_2272 ();
 b15zdnd11an1n64x5 FILLER_125_0 ();
 b15zdnd11an1n64x5 FILLER_125_64 ();
 b15zdnd11an1n64x5 FILLER_125_128 ();
 b15zdnd11an1n16x5 FILLER_125_192 ();
 b15zdnd11an1n08x5 FILLER_125_208 ();
 b15zdnd00an1n02x5 FILLER_125_216 ();
 b15zdnd11an1n08x5 FILLER_125_222 ();
 b15zdnd11an1n04x5 FILLER_125_230 ();
 b15zdnd11an1n64x5 FILLER_125_248 ();
 b15zdnd11an1n64x5 FILLER_125_312 ();
 b15zdnd11an1n64x5 FILLER_125_376 ();
 b15zdnd11an1n64x5 FILLER_125_440 ();
 b15zdnd11an1n64x5 FILLER_125_504 ();
 b15zdnd11an1n64x5 FILLER_125_568 ();
 b15zdnd11an1n64x5 FILLER_125_632 ();
 b15zdnd11an1n64x5 FILLER_125_696 ();
 b15zdnd11an1n64x5 FILLER_125_760 ();
 b15zdnd11an1n32x5 FILLER_125_824 ();
 b15zdnd11an1n16x5 FILLER_125_856 ();
 b15zdnd11an1n08x5 FILLER_125_872 ();
 b15zdnd00an1n02x5 FILLER_125_880 ();
 b15zdnd00an1n01x5 FILLER_125_882 ();
 b15zdnd11an1n04x5 FILLER_125_886 ();
 b15zdnd11an1n64x5 FILLER_125_893 ();
 b15zdnd11an1n16x5 FILLER_125_957 ();
 b15zdnd11an1n08x5 FILLER_125_973 ();
 b15zdnd11an1n04x5 FILLER_125_981 ();
 b15zdnd00an1n02x5 FILLER_125_985 ();
 b15zdnd00an1n01x5 FILLER_125_987 ();
 b15zdnd11an1n04x5 FILLER_125_994 ();
 b15zdnd11an1n64x5 FILLER_125_1002 ();
 b15zdnd11an1n32x5 FILLER_125_1066 ();
 b15zdnd11an1n08x5 FILLER_125_1098 ();
 b15zdnd11an1n04x5 FILLER_125_1106 ();
 b15zdnd00an1n02x5 FILLER_125_1110 ();
 b15zdnd11an1n64x5 FILLER_125_1116 ();
 b15zdnd11an1n32x5 FILLER_125_1180 ();
 b15zdnd11an1n04x5 FILLER_125_1212 ();
 b15zdnd00an1n02x5 FILLER_125_1216 ();
 b15zdnd11an1n16x5 FILLER_125_1221 ();
 b15zdnd11an1n08x5 FILLER_125_1237 ();
 b15zdnd00an1n02x5 FILLER_125_1245 ();
 b15zdnd11an1n64x5 FILLER_125_1257 ();
 b15zdnd11an1n64x5 FILLER_125_1321 ();
 b15zdnd11an1n64x5 FILLER_125_1385 ();
 b15zdnd11an1n64x5 FILLER_125_1449 ();
 b15zdnd11an1n64x5 FILLER_125_1513 ();
 b15zdnd11an1n64x5 FILLER_125_1577 ();
 b15zdnd11an1n64x5 FILLER_125_1641 ();
 b15zdnd11an1n64x5 FILLER_125_1705 ();
 b15zdnd11an1n64x5 FILLER_125_1769 ();
 b15zdnd11an1n64x5 FILLER_125_1833 ();
 b15zdnd11an1n64x5 FILLER_125_1897 ();
 b15zdnd11an1n64x5 FILLER_125_1961 ();
 b15zdnd11an1n32x5 FILLER_125_2025 ();
 b15zdnd11an1n16x5 FILLER_125_2057 ();
 b15zdnd11an1n08x5 FILLER_125_2073 ();
 b15zdnd00an1n02x5 FILLER_125_2081 ();
 b15zdnd11an1n32x5 FILLER_125_2101 ();
 b15zdnd11an1n08x5 FILLER_125_2133 ();
 b15zdnd11an1n04x5 FILLER_125_2141 ();
 b15zdnd00an1n02x5 FILLER_125_2145 ();
 b15zdnd00an1n01x5 FILLER_125_2147 ();
 b15zdnd11an1n64x5 FILLER_125_2200 ();
 b15zdnd11an1n16x5 FILLER_125_2264 ();
 b15zdnd11an1n04x5 FILLER_125_2280 ();
 b15zdnd11an1n64x5 FILLER_126_8 ();
 b15zdnd11an1n64x5 FILLER_126_72 ();
 b15zdnd11an1n64x5 FILLER_126_136 ();
 b15zdnd11an1n16x5 FILLER_126_200 ();
 b15zdnd00an1n02x5 FILLER_126_216 ();
 b15zdnd00an1n01x5 FILLER_126_218 ();
 b15zdnd11an1n64x5 FILLER_126_229 ();
 b15zdnd11an1n64x5 FILLER_126_293 ();
 b15zdnd11an1n64x5 FILLER_126_357 ();
 b15zdnd11an1n64x5 FILLER_126_421 ();
 b15zdnd11an1n64x5 FILLER_126_485 ();
 b15zdnd11an1n64x5 FILLER_126_549 ();
 b15zdnd11an1n64x5 FILLER_126_613 ();
 b15zdnd11an1n32x5 FILLER_126_677 ();
 b15zdnd11an1n08x5 FILLER_126_709 ();
 b15zdnd00an1n01x5 FILLER_126_717 ();
 b15zdnd11an1n64x5 FILLER_126_726 ();
 b15zdnd11an1n64x5 FILLER_126_790 ();
 b15zdnd11an1n64x5 FILLER_126_854 ();
 b15zdnd11an1n32x5 FILLER_126_918 ();
 b15zdnd11an1n08x5 FILLER_126_950 ();
 b15zdnd00an1n01x5 FILLER_126_958 ();
 b15zdnd11an1n08x5 FILLER_126_1001 ();
 b15zdnd00an1n01x5 FILLER_126_1009 ();
 b15zdnd11an1n64x5 FILLER_126_1018 ();
 b15zdnd11an1n64x5 FILLER_126_1082 ();
 b15zdnd11an1n32x5 FILLER_126_1146 ();
 b15zdnd00an1n02x5 FILLER_126_1178 ();
 b15zdnd00an1n01x5 FILLER_126_1180 ();
 b15zdnd11an1n04x5 FILLER_126_1201 ();
 b15zdnd00an1n02x5 FILLER_126_1205 ();
 b15zdnd11an1n64x5 FILLER_126_1221 ();
 b15zdnd11an1n64x5 FILLER_126_1285 ();
 b15zdnd11an1n32x5 FILLER_126_1349 ();
 b15zdnd11an1n08x5 FILLER_126_1381 ();
 b15zdnd00an1n02x5 FILLER_126_1389 ();
 b15zdnd11an1n32x5 FILLER_126_1405 ();
 b15zdnd11an1n16x5 FILLER_126_1437 ();
 b15zdnd11an1n08x5 FILLER_126_1453 ();
 b15zdnd11an1n04x5 FILLER_126_1461 ();
 b15zdnd00an1n02x5 FILLER_126_1465 ();
 b15zdnd11an1n64x5 FILLER_126_1487 ();
 b15zdnd11an1n64x5 FILLER_126_1551 ();
 b15zdnd11an1n64x5 FILLER_126_1615 ();
 b15zdnd11an1n64x5 FILLER_126_1679 ();
 b15zdnd11an1n64x5 FILLER_126_1743 ();
 b15zdnd11an1n64x5 FILLER_126_1807 ();
 b15zdnd11an1n64x5 FILLER_126_1871 ();
 b15zdnd11an1n64x5 FILLER_126_1935 ();
 b15zdnd11an1n64x5 FILLER_126_1999 ();
 b15zdnd11an1n16x5 FILLER_126_2063 ();
 b15zdnd11an1n04x5 FILLER_126_2079 ();
 b15zdnd00an1n01x5 FILLER_126_2083 ();
 b15zdnd11an1n16x5 FILLER_126_2126 ();
 b15zdnd11an1n08x5 FILLER_126_2142 ();
 b15zdnd11an1n04x5 FILLER_126_2150 ();
 b15zdnd11an1n04x5 FILLER_126_2162 ();
 b15zdnd11an1n04x5 FILLER_126_2169 ();
 b15zdnd11an1n04x5 FILLER_126_2176 ();
 b15zdnd11an1n64x5 FILLER_126_2183 ();
 b15zdnd11an1n16x5 FILLER_126_2247 ();
 b15zdnd11an1n08x5 FILLER_126_2263 ();
 b15zdnd11an1n04x5 FILLER_126_2271 ();
 b15zdnd00an1n01x5 FILLER_126_2275 ();
 b15zdnd11an1n64x5 FILLER_127_0 ();
 b15zdnd11an1n64x5 FILLER_127_64 ();
 b15zdnd11an1n64x5 FILLER_127_128 ();
 b15zdnd11an1n16x5 FILLER_127_192 ();
 b15zdnd11an1n08x5 FILLER_127_208 ();
 b15zdnd11an1n04x5 FILLER_127_216 ();
 b15zdnd00an1n01x5 FILLER_127_220 ();
 b15zdnd11an1n64x5 FILLER_127_230 ();
 b15zdnd11an1n32x5 FILLER_127_294 ();
 b15zdnd11an1n16x5 FILLER_127_326 ();
 b15zdnd11an1n04x5 FILLER_127_342 ();
 b15zdnd00an1n02x5 FILLER_127_346 ();
 b15zdnd00an1n01x5 FILLER_127_348 ();
 b15zdnd11an1n16x5 FILLER_127_391 ();
 b15zdnd00an1n02x5 FILLER_127_407 ();
 b15zdnd11an1n64x5 FILLER_127_412 ();
 b15zdnd11an1n32x5 FILLER_127_476 ();
 b15zdnd11an1n08x5 FILLER_127_508 ();
 b15zdnd11an1n04x5 FILLER_127_516 ();
 b15zdnd11an1n64x5 FILLER_127_523 ();
 b15zdnd11an1n08x5 FILLER_127_587 ();
 b15zdnd11an1n04x5 FILLER_127_595 ();
 b15zdnd00an1n02x5 FILLER_127_599 ();
 b15zdnd00an1n01x5 FILLER_127_601 ();
 b15zdnd11an1n64x5 FILLER_127_622 ();
 b15zdnd11an1n64x5 FILLER_127_686 ();
 b15zdnd11an1n64x5 FILLER_127_750 ();
 b15zdnd11an1n64x5 FILLER_127_814 ();
 b15zdnd11an1n64x5 FILLER_127_878 ();
 b15zdnd11an1n16x5 FILLER_127_942 ();
 b15zdnd11an1n08x5 FILLER_127_958 ();
 b15zdnd11an1n64x5 FILLER_127_980 ();
 b15zdnd11an1n64x5 FILLER_127_1044 ();
 b15zdnd11an1n64x5 FILLER_127_1108 ();
 b15zdnd11an1n64x5 FILLER_127_1172 ();
 b15zdnd11an1n64x5 FILLER_127_1236 ();
 b15zdnd11an1n64x5 FILLER_127_1300 ();
 b15zdnd11an1n64x5 FILLER_127_1364 ();
 b15zdnd11an1n64x5 FILLER_127_1428 ();
 b15zdnd11an1n04x5 FILLER_127_1492 ();
 b15zdnd00an1n02x5 FILLER_127_1496 ();
 b15zdnd11an1n64x5 FILLER_127_1512 ();
 b15zdnd11an1n64x5 FILLER_127_1576 ();
 b15zdnd11an1n32x5 FILLER_127_1640 ();
 b15zdnd11an1n08x5 FILLER_127_1672 ();
 b15zdnd11an1n04x5 FILLER_127_1680 ();
 b15zdnd00an1n02x5 FILLER_127_1684 ();
 b15zdnd11an1n08x5 FILLER_127_1689 ();
 b15zdnd11an1n04x5 FILLER_127_1737 ();
 b15zdnd11an1n64x5 FILLER_127_1744 ();
 b15zdnd11an1n64x5 FILLER_127_1808 ();
 b15zdnd11an1n64x5 FILLER_127_1872 ();
 b15zdnd11an1n64x5 FILLER_127_1936 ();
 b15zdnd11an1n64x5 FILLER_127_2000 ();
 b15zdnd11an1n16x5 FILLER_127_2064 ();
 b15zdnd00an1n02x5 FILLER_127_2080 ();
 b15zdnd11an1n16x5 FILLER_127_2134 ();
 b15zdnd11an1n64x5 FILLER_127_2192 ();
 b15zdnd11an1n16x5 FILLER_127_2256 ();
 b15zdnd11an1n08x5 FILLER_127_2272 ();
 b15zdnd11an1n04x5 FILLER_127_2280 ();
 b15zdnd11an1n08x5 FILLER_128_8 ();
 b15zdnd11an1n04x5 FILLER_128_16 ();
 b15zdnd00an1n01x5 FILLER_128_20 ();
 b15zdnd11an1n64x5 FILLER_128_25 ();
 b15zdnd11an1n64x5 FILLER_128_89 ();
 b15zdnd11an1n64x5 FILLER_128_153 ();
 b15zdnd11an1n64x5 FILLER_128_217 ();
 b15zdnd11an1n64x5 FILLER_128_281 ();
 b15zdnd11an1n32x5 FILLER_128_345 ();
 b15zdnd11an1n04x5 FILLER_128_377 ();
 b15zdnd00an1n01x5 FILLER_128_381 ();
 b15zdnd11an1n64x5 FILLER_128_434 ();
 b15zdnd11an1n08x5 FILLER_128_498 ();
 b15zdnd11an1n04x5 FILLER_128_509 ();
 b15zdnd00an1n01x5 FILLER_128_513 ();
 b15zdnd11an1n16x5 FILLER_128_517 ();
 b15zdnd11an1n04x5 FILLER_128_533 ();
 b15zdnd00an1n02x5 FILLER_128_537 ();
 b15zdnd11an1n16x5 FILLER_128_546 ();
 b15zdnd11an1n64x5 FILLER_128_614 ();
 b15zdnd11an1n32x5 FILLER_128_678 ();
 b15zdnd11an1n08x5 FILLER_128_710 ();
 b15zdnd11an1n64x5 FILLER_128_726 ();
 b15zdnd11an1n64x5 FILLER_128_790 ();
 b15zdnd11an1n64x5 FILLER_128_854 ();
 b15zdnd11an1n32x5 FILLER_128_918 ();
 b15zdnd11an1n16x5 FILLER_128_950 ();
 b15zdnd00an1n01x5 FILLER_128_966 ();
 b15zdnd11an1n64x5 FILLER_128_984 ();
 b15zdnd11an1n64x5 FILLER_128_1048 ();
 b15zdnd11an1n64x5 FILLER_128_1112 ();
 b15zdnd11an1n04x5 FILLER_128_1176 ();
 b15zdnd00an1n02x5 FILLER_128_1180 ();
 b15zdnd00an1n01x5 FILLER_128_1182 ();
 b15zdnd11an1n32x5 FILLER_128_1201 ();
 b15zdnd11an1n04x5 FILLER_128_1233 ();
 b15zdnd00an1n02x5 FILLER_128_1237 ();
 b15zdnd00an1n01x5 FILLER_128_1239 ();
 b15zdnd11an1n16x5 FILLER_128_1248 ();
 b15zdnd11an1n16x5 FILLER_128_1280 ();
 b15zdnd11an1n04x5 FILLER_128_1296 ();
 b15zdnd00an1n02x5 FILLER_128_1300 ();
 b15zdnd11an1n04x5 FILLER_128_1326 ();
 b15zdnd00an1n02x5 FILLER_128_1330 ();
 b15zdnd11an1n04x5 FILLER_128_1340 ();
 b15zdnd00an1n02x5 FILLER_128_1344 ();
 b15zdnd00an1n01x5 FILLER_128_1346 ();
 b15zdnd11an1n64x5 FILLER_128_1356 ();
 b15zdnd11an1n64x5 FILLER_128_1420 ();
 b15zdnd11an1n64x5 FILLER_128_1484 ();
 b15zdnd11an1n64x5 FILLER_128_1548 ();
 b15zdnd11an1n32x5 FILLER_128_1612 ();
 b15zdnd11an1n16x5 FILLER_128_1644 ();
 b15zdnd11an1n16x5 FILLER_128_1712 ();
 b15zdnd11an1n04x5 FILLER_128_1728 ();
 b15zdnd00an1n01x5 FILLER_128_1732 ();
 b15zdnd11an1n64x5 FILLER_128_1736 ();
 b15zdnd11an1n64x5 FILLER_128_1800 ();
 b15zdnd11an1n64x5 FILLER_128_1864 ();
 b15zdnd11an1n64x5 FILLER_128_1928 ();
 b15zdnd11an1n64x5 FILLER_128_1992 ();
 b15zdnd11an1n32x5 FILLER_128_2056 ();
 b15zdnd11an1n08x5 FILLER_128_2088 ();
 b15zdnd11an1n04x5 FILLER_128_2096 ();
 b15zdnd00an1n01x5 FILLER_128_2100 ();
 b15zdnd11an1n04x5 FILLER_128_2104 ();
 b15zdnd11an1n32x5 FILLER_128_2111 ();
 b15zdnd11an1n08x5 FILLER_128_2143 ();
 b15zdnd00an1n02x5 FILLER_128_2151 ();
 b15zdnd00an1n01x5 FILLER_128_2153 ();
 b15zdnd11an1n64x5 FILLER_128_2162 ();
 b15zdnd11an1n32x5 FILLER_128_2226 ();
 b15zdnd11an1n16x5 FILLER_128_2258 ();
 b15zdnd00an1n02x5 FILLER_128_2274 ();
 b15zdnd11an1n64x5 FILLER_129_0 ();
 b15zdnd11an1n64x5 FILLER_129_64 ();
 b15zdnd11an1n64x5 FILLER_129_128 ();
 b15zdnd11an1n16x5 FILLER_129_192 ();
 b15zdnd11an1n08x5 FILLER_129_208 ();
 b15zdnd11an1n04x5 FILLER_129_216 ();
 b15zdnd00an1n02x5 FILLER_129_220 ();
 b15zdnd00an1n01x5 FILLER_129_222 ();
 b15zdnd11an1n64x5 FILLER_129_263 ();
 b15zdnd11an1n64x5 FILLER_129_327 ();
 b15zdnd11an1n08x5 FILLER_129_391 ();
 b15zdnd00an1n02x5 FILLER_129_399 ();
 b15zdnd11an1n04x5 FILLER_129_404 ();
 b15zdnd11an1n64x5 FILLER_129_411 ();
 b15zdnd11an1n08x5 FILLER_129_475 ();
 b15zdnd11an1n04x5 FILLER_129_535 ();
 b15zdnd11an1n64x5 FILLER_129_581 ();
 b15zdnd11an1n08x5 FILLER_129_645 ();
 b15zdnd11an1n04x5 FILLER_129_653 ();
 b15zdnd11an1n16x5 FILLER_129_660 ();
 b15zdnd11an1n64x5 FILLER_129_684 ();
 b15zdnd11an1n64x5 FILLER_129_748 ();
 b15zdnd11an1n64x5 FILLER_129_812 ();
 b15zdnd11an1n64x5 FILLER_129_876 ();
 b15zdnd11an1n64x5 FILLER_129_940 ();
 b15zdnd11an1n64x5 FILLER_129_1004 ();
 b15zdnd11an1n64x5 FILLER_129_1068 ();
 b15zdnd11an1n64x5 FILLER_129_1132 ();
 b15zdnd00an1n02x5 FILLER_129_1196 ();
 b15zdnd11an1n64x5 FILLER_129_1219 ();
 b15zdnd11an1n64x5 FILLER_129_1283 ();
 b15zdnd11an1n64x5 FILLER_129_1347 ();
 b15zdnd11an1n64x5 FILLER_129_1411 ();
 b15zdnd11an1n64x5 FILLER_129_1475 ();
 b15zdnd11an1n64x5 FILLER_129_1539 ();
 b15zdnd11an1n16x5 FILLER_129_1603 ();
 b15zdnd11an1n08x5 FILLER_129_1619 ();
 b15zdnd00an1n02x5 FILLER_129_1627 ();
 b15zdnd11an1n16x5 FILLER_129_1649 ();
 b15zdnd11an1n08x5 FILLER_129_1665 ();
 b15zdnd11an1n04x5 FILLER_129_1673 ();
 b15zdnd00an1n01x5 FILLER_129_1677 ();
 b15zdnd11an1n04x5 FILLER_129_1681 ();
 b15zdnd11an1n64x5 FILLER_129_1688 ();
 b15zdnd11an1n64x5 FILLER_129_1752 ();
 b15zdnd11an1n64x5 FILLER_129_1816 ();
 b15zdnd11an1n64x5 FILLER_129_1880 ();
 b15zdnd11an1n64x5 FILLER_129_1944 ();
 b15zdnd11an1n64x5 FILLER_129_2008 ();
 b15zdnd11an1n32x5 FILLER_129_2072 ();
 b15zdnd00an1n02x5 FILLER_129_2104 ();
 b15zdnd11an1n64x5 FILLER_129_2109 ();
 b15zdnd11an1n64x5 FILLER_129_2173 ();
 b15zdnd11an1n32x5 FILLER_129_2237 ();
 b15zdnd11an1n08x5 FILLER_129_2269 ();
 b15zdnd11an1n04x5 FILLER_129_2277 ();
 b15zdnd00an1n02x5 FILLER_129_2281 ();
 b15zdnd00an1n01x5 FILLER_129_2283 ();
 b15zdnd11an1n16x5 FILLER_130_8 ();
 b15zdnd11an1n04x5 FILLER_130_24 ();
 b15zdnd00an1n02x5 FILLER_130_28 ();
 b15zdnd11an1n64x5 FILLER_130_34 ();
 b15zdnd11an1n64x5 FILLER_130_98 ();
 b15zdnd11an1n64x5 FILLER_130_162 ();
 b15zdnd11an1n64x5 FILLER_130_226 ();
 b15zdnd11an1n04x5 FILLER_130_290 ();
 b15zdnd00an1n01x5 FILLER_130_294 ();
 b15zdnd11an1n64x5 FILLER_130_337 ();
 b15zdnd11an1n32x5 FILLER_130_401 ();
 b15zdnd00an1n02x5 FILLER_130_433 ();
 b15zdnd00an1n01x5 FILLER_130_435 ();
 b15zdnd11an1n04x5 FILLER_130_440 ();
 b15zdnd11an1n04x5 FILLER_130_455 ();
 b15zdnd11an1n32x5 FILLER_130_501 ();
 b15zdnd00an1n02x5 FILLER_130_533 ();
 b15zdnd00an1n01x5 FILLER_130_535 ();
 b15zdnd11an1n04x5 FILLER_130_588 ();
 b15zdnd11an1n08x5 FILLER_130_595 ();
 b15zdnd11an1n04x5 FILLER_130_603 ();
 b15zdnd00an1n02x5 FILLER_130_607 ();
 b15zdnd11an1n32x5 FILLER_130_616 ();
 b15zdnd11an1n08x5 FILLER_130_648 ();
 b15zdnd11an1n04x5 FILLER_130_656 ();
 b15zdnd00an1n01x5 FILLER_130_660 ();
 b15zdnd11an1n04x5 FILLER_130_713 ();
 b15zdnd00an1n01x5 FILLER_130_717 ();
 b15zdnd11an1n16x5 FILLER_130_726 ();
 b15zdnd11an1n08x5 FILLER_130_742 ();
 b15zdnd00an1n01x5 FILLER_130_750 ();
 b15zdnd11an1n64x5 FILLER_130_769 ();
 b15zdnd11an1n64x5 FILLER_130_833 ();
 b15zdnd11an1n64x5 FILLER_130_897 ();
 b15zdnd11an1n64x5 FILLER_130_961 ();
 b15zdnd11an1n64x5 FILLER_130_1025 ();
 b15zdnd11an1n64x5 FILLER_130_1089 ();
 b15zdnd11an1n08x5 FILLER_130_1153 ();
 b15zdnd00an1n02x5 FILLER_130_1161 ();
 b15zdnd11an1n32x5 FILLER_130_1167 ();
 b15zdnd11an1n64x5 FILLER_130_1218 ();
 b15zdnd11an1n64x5 FILLER_130_1282 ();
 b15zdnd11an1n64x5 FILLER_130_1346 ();
 b15zdnd11an1n64x5 FILLER_130_1410 ();
 b15zdnd11an1n64x5 FILLER_130_1474 ();
 b15zdnd11an1n64x5 FILLER_130_1538 ();
 b15zdnd11an1n64x5 FILLER_130_1602 ();
 b15zdnd11an1n16x5 FILLER_130_1666 ();
 b15zdnd11an1n08x5 FILLER_130_1682 ();
 b15zdnd11an1n04x5 FILLER_130_1690 ();
 b15zdnd11an1n64x5 FILLER_130_1736 ();
 b15zdnd11an1n64x5 FILLER_130_1800 ();
 b15zdnd11an1n64x5 FILLER_130_1864 ();
 b15zdnd11an1n64x5 FILLER_130_1928 ();
 b15zdnd11an1n64x5 FILLER_130_1992 ();
 b15zdnd11an1n16x5 FILLER_130_2056 ();
 b15zdnd11an1n08x5 FILLER_130_2072 ();
 b15zdnd11an1n04x5 FILLER_130_2080 ();
 b15zdnd00an1n01x5 FILLER_130_2084 ();
 b15zdnd11an1n32x5 FILLER_130_2096 ();
 b15zdnd11an1n16x5 FILLER_130_2128 ();
 b15zdnd11an1n08x5 FILLER_130_2144 ();
 b15zdnd00an1n02x5 FILLER_130_2152 ();
 b15zdnd11an1n32x5 FILLER_130_2162 ();
 b15zdnd11an1n08x5 FILLER_130_2194 ();
 b15zdnd00an1n01x5 FILLER_130_2202 ();
 b15zdnd11an1n32x5 FILLER_130_2213 ();
 b15zdnd11an1n16x5 FILLER_130_2245 ();
 b15zdnd11an1n08x5 FILLER_130_2261 ();
 b15zdnd11an1n04x5 FILLER_130_2269 ();
 b15zdnd00an1n02x5 FILLER_130_2273 ();
 b15zdnd00an1n01x5 FILLER_130_2275 ();
 b15zdnd11an1n16x5 FILLER_131_0 ();
 b15zdnd11an1n04x5 FILLER_131_16 ();
 b15zdnd00an1n01x5 FILLER_131_20 ();
 b15zdnd11an1n16x5 FILLER_131_25 ();
 b15zdnd11an1n08x5 FILLER_131_41 ();
 b15zdnd11an1n04x5 FILLER_131_49 ();
 b15zdnd11an1n64x5 FILLER_131_61 ();
 b15zdnd11an1n64x5 FILLER_131_125 ();
 b15zdnd11an1n08x5 FILLER_131_189 ();
 b15zdnd11an1n04x5 FILLER_131_197 ();
 b15zdnd00an1n02x5 FILLER_131_201 ();
 b15zdnd00an1n01x5 FILLER_131_203 ();
 b15zdnd11an1n64x5 FILLER_131_246 ();
 b15zdnd11an1n64x5 FILLER_131_310 ();
 b15zdnd11an1n64x5 FILLER_131_374 ();
 b15zdnd11an1n32x5 FILLER_131_438 ();
 b15zdnd00an1n01x5 FILLER_131_470 ();
 b15zdnd11an1n64x5 FILLER_131_491 ();
 b15zdnd00an1n01x5 FILLER_131_555 ();
 b15zdnd11an1n04x5 FILLER_131_559 ();
 b15zdnd11an1n04x5 FILLER_131_566 ();
 b15zdnd11an1n08x5 FILLER_131_573 ();
 b15zdnd00an1n02x5 FILLER_131_581 ();
 b15zdnd00an1n01x5 FILLER_131_583 ();
 b15zdnd11an1n64x5 FILLER_131_587 ();
 b15zdnd11an1n08x5 FILLER_131_651 ();
 b15zdnd11an1n04x5 FILLER_131_659 ();
 b15zdnd11an1n64x5 FILLER_131_715 ();
 b15zdnd11an1n64x5 FILLER_131_779 ();
 b15zdnd11an1n64x5 FILLER_131_843 ();
 b15zdnd11an1n64x5 FILLER_131_907 ();
 b15zdnd11an1n64x5 FILLER_131_971 ();
 b15zdnd11an1n64x5 FILLER_131_1035 ();
 b15zdnd11an1n32x5 FILLER_131_1099 ();
 b15zdnd11an1n64x5 FILLER_131_1134 ();
 b15zdnd11an1n32x5 FILLER_131_1198 ();
 b15zdnd11an1n16x5 FILLER_131_1230 ();
 b15zdnd00an1n02x5 FILLER_131_1246 ();
 b15zdnd11an1n16x5 FILLER_131_1256 ();
 b15zdnd11an1n04x5 FILLER_131_1272 ();
 b15zdnd00an1n02x5 FILLER_131_1276 ();
 b15zdnd00an1n01x5 FILLER_131_1278 ();
 b15zdnd11an1n64x5 FILLER_131_1298 ();
 b15zdnd11an1n32x5 FILLER_131_1362 ();
 b15zdnd11an1n16x5 FILLER_131_1394 ();
 b15zdnd11an1n08x5 FILLER_131_1410 ();
 b15zdnd00an1n02x5 FILLER_131_1418 ();
 b15zdnd11an1n32x5 FILLER_131_1424 ();
 b15zdnd11an1n16x5 FILLER_131_1456 ();
 b15zdnd00an1n01x5 FILLER_131_1472 ();
 b15zdnd11an1n64x5 FILLER_131_1484 ();
 b15zdnd11an1n64x5 FILLER_131_1548 ();
 b15zdnd11an1n64x5 FILLER_131_1612 ();
 b15zdnd11an1n32x5 FILLER_131_1676 ();
 b15zdnd11an1n16x5 FILLER_131_1708 ();
 b15zdnd00an1n01x5 FILLER_131_1724 ();
 b15zdnd11an1n32x5 FILLER_131_1733 ();
 b15zdnd11an1n08x5 FILLER_131_1765 ();
 b15zdnd00an1n01x5 FILLER_131_1773 ();
 b15zdnd11an1n64x5 FILLER_131_1786 ();
 b15zdnd11an1n64x5 FILLER_131_1850 ();
 b15zdnd11an1n64x5 FILLER_131_1914 ();
 b15zdnd11an1n64x5 FILLER_131_1978 ();
 b15zdnd11an1n64x5 FILLER_131_2042 ();
 b15zdnd11an1n08x5 FILLER_131_2106 ();
 b15zdnd11an1n64x5 FILLER_131_2156 ();
 b15zdnd11an1n64x5 FILLER_131_2220 ();
 b15zdnd00an1n02x5 FILLER_132_8 ();
 b15zdnd11an1n04x5 FILLER_132_52 ();
 b15zdnd11an1n64x5 FILLER_132_59 ();
 b15zdnd11an1n04x5 FILLER_132_123 ();
 b15zdnd00an1n02x5 FILLER_132_127 ();
 b15zdnd00an1n01x5 FILLER_132_129 ();
 b15zdnd11an1n08x5 FILLER_132_172 ();
 b15zdnd11an1n64x5 FILLER_132_200 ();
 b15zdnd11an1n64x5 FILLER_132_264 ();
 b15zdnd11an1n32x5 FILLER_132_328 ();
 b15zdnd11an1n16x5 FILLER_132_360 ();
 b15zdnd11an1n08x5 FILLER_132_376 ();
 b15zdnd11an1n04x5 FILLER_132_384 ();
 b15zdnd00an1n01x5 FILLER_132_388 ();
 b15zdnd11an1n64x5 FILLER_132_392 ();
 b15zdnd11an1n16x5 FILLER_132_456 ();
 b15zdnd11an1n04x5 FILLER_132_472 ();
 b15zdnd00an1n01x5 FILLER_132_476 ();
 b15zdnd11an1n04x5 FILLER_132_503 ();
 b15zdnd11an1n64x5 FILLER_132_521 ();
 b15zdnd00an1n01x5 FILLER_132_585 ();
 b15zdnd11an1n64x5 FILLER_132_589 ();
 b15zdnd11an1n16x5 FILLER_132_653 ();
 b15zdnd11an1n04x5 FILLER_132_672 ();
 b15zdnd11an1n04x5 FILLER_132_679 ();
 b15zdnd00an1n02x5 FILLER_132_683 ();
 b15zdnd00an1n01x5 FILLER_132_685 ();
 b15zdnd11an1n04x5 FILLER_132_689 ();
 b15zdnd11an1n16x5 FILLER_132_696 ();
 b15zdnd11an1n04x5 FILLER_132_712 ();
 b15zdnd00an1n02x5 FILLER_132_716 ();
 b15zdnd11an1n32x5 FILLER_132_726 ();
 b15zdnd00an1n01x5 FILLER_132_758 ();
 b15zdnd11an1n64x5 FILLER_132_767 ();
 b15zdnd11an1n64x5 FILLER_132_831 ();
 b15zdnd11an1n64x5 FILLER_132_895 ();
 b15zdnd11an1n64x5 FILLER_132_959 ();
 b15zdnd11an1n64x5 FILLER_132_1023 ();
 b15zdnd11an1n32x5 FILLER_132_1087 ();
 b15zdnd11an1n08x5 FILLER_132_1119 ();
 b15zdnd11an1n04x5 FILLER_132_1127 ();
 b15zdnd11an1n64x5 FILLER_132_1158 ();
 b15zdnd11an1n32x5 FILLER_132_1222 ();
 b15zdnd11an1n16x5 FILLER_132_1254 ();
 b15zdnd00an1n02x5 FILLER_132_1270 ();
 b15zdnd00an1n01x5 FILLER_132_1272 ();
 b15zdnd11an1n04x5 FILLER_132_1315 ();
 b15zdnd11an1n64x5 FILLER_132_1332 ();
 b15zdnd11an1n64x5 FILLER_132_1396 ();
 b15zdnd11an1n64x5 FILLER_132_1460 ();
 b15zdnd11an1n64x5 FILLER_132_1524 ();
 b15zdnd11an1n64x5 FILLER_132_1588 ();
 b15zdnd11an1n32x5 FILLER_132_1652 ();
 b15zdnd11an1n16x5 FILLER_132_1684 ();
 b15zdnd11an1n08x5 FILLER_132_1700 ();
 b15zdnd00an1n02x5 FILLER_132_1708 ();
 b15zdnd11an1n64x5 FILLER_132_1752 ();
 b15zdnd11an1n64x5 FILLER_132_1816 ();
 b15zdnd11an1n64x5 FILLER_132_1880 ();
 b15zdnd11an1n64x5 FILLER_132_1944 ();
 b15zdnd11an1n64x5 FILLER_132_2008 ();
 b15zdnd11an1n64x5 FILLER_132_2072 ();
 b15zdnd11an1n16x5 FILLER_132_2136 ();
 b15zdnd00an1n02x5 FILLER_132_2152 ();
 b15zdnd11an1n64x5 FILLER_132_2162 ();
 b15zdnd11an1n32x5 FILLER_132_2226 ();
 b15zdnd11an1n16x5 FILLER_132_2258 ();
 b15zdnd00an1n02x5 FILLER_132_2274 ();
 b15zdnd11an1n16x5 FILLER_133_0 ();
 b15zdnd11an1n08x5 FILLER_133_16 ();
 b15zdnd11an1n64x5 FILLER_133_76 ();
 b15zdnd11an1n64x5 FILLER_133_140 ();
 b15zdnd11an1n64x5 FILLER_133_204 ();
 b15zdnd11an1n64x5 FILLER_133_268 ();
 b15zdnd11an1n16x5 FILLER_133_332 ();
 b15zdnd11an1n08x5 FILLER_133_348 ();
 b15zdnd11an1n04x5 FILLER_133_356 ();
 b15zdnd00an1n01x5 FILLER_133_360 ();
 b15zdnd11an1n64x5 FILLER_133_393 ();
 b15zdnd11an1n64x5 FILLER_133_457 ();
 b15zdnd11an1n64x5 FILLER_133_521 ();
 b15zdnd11an1n64x5 FILLER_133_585 ();
 b15zdnd11an1n16x5 FILLER_133_649 ();
 b15zdnd11an1n08x5 FILLER_133_665 ();
 b15zdnd00an1n02x5 FILLER_133_673 ();
 b15zdnd00an1n01x5 FILLER_133_675 ();
 b15zdnd11an1n64x5 FILLER_133_679 ();
 b15zdnd11an1n64x5 FILLER_133_743 ();
 b15zdnd11an1n64x5 FILLER_133_807 ();
 b15zdnd11an1n64x5 FILLER_133_871 ();
 b15zdnd11an1n64x5 FILLER_133_935 ();
 b15zdnd11an1n64x5 FILLER_133_999 ();
 b15zdnd11an1n04x5 FILLER_133_1063 ();
 b15zdnd11an1n64x5 FILLER_133_1075 ();
 b15zdnd11an1n64x5 FILLER_133_1139 ();
 b15zdnd11an1n64x5 FILLER_133_1203 ();
 b15zdnd11an1n64x5 FILLER_133_1267 ();
 b15zdnd11an1n64x5 FILLER_133_1331 ();
 b15zdnd11an1n64x5 FILLER_133_1395 ();
 b15zdnd11an1n64x5 FILLER_133_1459 ();
 b15zdnd11an1n16x5 FILLER_133_1523 ();
 b15zdnd11an1n04x5 FILLER_133_1548 ();
 b15zdnd11an1n32x5 FILLER_133_1555 ();
 b15zdnd00an1n01x5 FILLER_133_1587 ();
 b15zdnd11an1n04x5 FILLER_133_1591 ();
 b15zdnd11an1n64x5 FILLER_133_1598 ();
 b15zdnd11an1n64x5 FILLER_133_1662 ();
 b15zdnd11an1n64x5 FILLER_133_1726 ();
 b15zdnd11an1n64x5 FILLER_133_1790 ();
 b15zdnd11an1n64x5 FILLER_133_1854 ();
 b15zdnd11an1n64x5 FILLER_133_1918 ();
 b15zdnd11an1n64x5 FILLER_133_1982 ();
 b15zdnd11an1n64x5 FILLER_133_2046 ();
 b15zdnd11an1n64x5 FILLER_133_2110 ();
 b15zdnd11an1n64x5 FILLER_133_2174 ();
 b15zdnd11an1n32x5 FILLER_133_2238 ();
 b15zdnd11an1n08x5 FILLER_133_2270 ();
 b15zdnd11an1n04x5 FILLER_133_2278 ();
 b15zdnd00an1n02x5 FILLER_133_2282 ();
 b15zdnd11an1n32x5 FILLER_134_8 ();
 b15zdnd00an1n02x5 FILLER_134_40 ();
 b15zdnd00an1n01x5 FILLER_134_42 ();
 b15zdnd11an1n04x5 FILLER_134_46 ();
 b15zdnd11an1n64x5 FILLER_134_53 ();
 b15zdnd11an1n64x5 FILLER_134_117 ();
 b15zdnd11an1n64x5 FILLER_134_181 ();
 b15zdnd11an1n64x5 FILLER_134_245 ();
 b15zdnd11an1n64x5 FILLER_134_309 ();
 b15zdnd11an1n16x5 FILLER_134_373 ();
 b15zdnd11an1n64x5 FILLER_134_392 ();
 b15zdnd11an1n64x5 FILLER_134_456 ();
 b15zdnd11an1n64x5 FILLER_134_520 ();
 b15zdnd11an1n64x5 FILLER_134_584 ();
 b15zdnd11an1n64x5 FILLER_134_648 ();
 b15zdnd11an1n04x5 FILLER_134_712 ();
 b15zdnd00an1n02x5 FILLER_134_716 ();
 b15zdnd11an1n64x5 FILLER_134_726 ();
 b15zdnd11an1n64x5 FILLER_134_790 ();
 b15zdnd11an1n64x5 FILLER_134_854 ();
 b15zdnd11an1n64x5 FILLER_134_918 ();
 b15zdnd11an1n64x5 FILLER_134_982 ();
 b15zdnd11an1n16x5 FILLER_134_1046 ();
 b15zdnd00an1n02x5 FILLER_134_1062 ();
 b15zdnd11an1n32x5 FILLER_134_1072 ();
 b15zdnd11an1n16x5 FILLER_134_1104 ();
 b15zdnd11an1n08x5 FILLER_134_1120 ();
 b15zdnd00an1n02x5 FILLER_134_1128 ();
 b15zdnd11an1n64x5 FILLER_134_1140 ();
 b15zdnd11an1n64x5 FILLER_134_1204 ();
 b15zdnd11an1n64x5 FILLER_134_1268 ();
 b15zdnd11an1n64x5 FILLER_134_1332 ();
 b15zdnd11an1n32x5 FILLER_134_1396 ();
 b15zdnd11an1n08x5 FILLER_134_1428 ();
 b15zdnd00an1n01x5 FILLER_134_1436 ();
 b15zdnd11an1n32x5 FILLER_134_1446 ();
 b15zdnd00an1n02x5 FILLER_134_1478 ();
 b15zdnd11an1n16x5 FILLER_134_1501 ();
 b15zdnd11an1n04x5 FILLER_134_1517 ();
 b15zdnd00an1n02x5 FILLER_134_1521 ();
 b15zdnd00an1n01x5 FILLER_134_1523 ();
 b15zdnd11an1n04x5 FILLER_134_1531 ();
 b15zdnd11an1n08x5 FILLER_134_1551 ();
 b15zdnd11an1n04x5 FILLER_134_1559 ();
 b15zdnd00an1n01x5 FILLER_134_1563 ();
 b15zdnd11an1n04x5 FILLER_134_1567 ();
 b15zdnd00an1n02x5 FILLER_134_1571 ();
 b15zdnd11an1n64x5 FILLER_134_1617 ();
 b15zdnd11an1n16x5 FILLER_134_1681 ();
 b15zdnd11an1n08x5 FILLER_134_1697 ();
 b15zdnd00an1n02x5 FILLER_134_1705 ();
 b15zdnd00an1n01x5 FILLER_134_1707 ();
 b15zdnd11an1n64x5 FILLER_134_1722 ();
 b15zdnd11an1n64x5 FILLER_134_1786 ();
 b15zdnd11an1n64x5 FILLER_134_1850 ();
 b15zdnd11an1n64x5 FILLER_134_1914 ();
 b15zdnd11an1n64x5 FILLER_134_1978 ();
 b15zdnd11an1n64x5 FILLER_134_2042 ();
 b15zdnd11an1n32x5 FILLER_134_2106 ();
 b15zdnd11an1n16x5 FILLER_134_2138 ();
 b15zdnd11an1n64x5 FILLER_134_2162 ();
 b15zdnd11an1n32x5 FILLER_134_2226 ();
 b15zdnd11an1n16x5 FILLER_134_2258 ();
 b15zdnd00an1n02x5 FILLER_134_2274 ();
 b15zdnd11an1n64x5 FILLER_135_0 ();
 b15zdnd11an1n08x5 FILLER_135_64 ();
 b15zdnd00an1n02x5 FILLER_135_72 ();
 b15zdnd00an1n01x5 FILLER_135_74 ();
 b15zdnd11an1n64x5 FILLER_135_120 ();
 b15zdnd11an1n64x5 FILLER_135_184 ();
 b15zdnd11an1n64x5 FILLER_135_248 ();
 b15zdnd11an1n64x5 FILLER_135_312 ();
 b15zdnd11an1n64x5 FILLER_135_376 ();
 b15zdnd11an1n64x5 FILLER_135_440 ();
 b15zdnd11an1n64x5 FILLER_135_504 ();
 b15zdnd11an1n32x5 FILLER_135_568 ();
 b15zdnd11an1n16x5 FILLER_135_600 ();
 b15zdnd11an1n08x5 FILLER_135_616 ();
 b15zdnd00an1n02x5 FILLER_135_624 ();
 b15zdnd00an1n01x5 FILLER_135_626 ();
 b15zdnd11an1n64x5 FILLER_135_636 ();
 b15zdnd11an1n64x5 FILLER_135_700 ();
 b15zdnd11an1n64x5 FILLER_135_764 ();
 b15zdnd11an1n08x5 FILLER_135_828 ();
 b15zdnd00an1n02x5 FILLER_135_836 ();
 b15zdnd11an1n64x5 FILLER_135_849 ();
 b15zdnd11an1n64x5 FILLER_135_913 ();
 b15zdnd11an1n64x5 FILLER_135_977 ();
 b15zdnd11an1n64x5 FILLER_135_1041 ();
 b15zdnd11an1n64x5 FILLER_135_1105 ();
 b15zdnd11an1n64x5 FILLER_135_1169 ();
 b15zdnd11an1n64x5 FILLER_135_1233 ();
 b15zdnd11an1n32x5 FILLER_135_1297 ();
 b15zdnd11an1n16x5 FILLER_135_1329 ();
 b15zdnd11an1n64x5 FILLER_135_1354 ();
 b15zdnd11an1n64x5 FILLER_135_1418 ();
 b15zdnd00an1n02x5 FILLER_135_1482 ();
 b15zdnd00an1n01x5 FILLER_135_1484 ();
 b15zdnd11an1n32x5 FILLER_135_1494 ();
 b15zdnd11an1n08x5 FILLER_135_1526 ();
 b15zdnd00an1n02x5 FILLER_135_1534 ();
 b15zdnd11an1n08x5 FILLER_135_1546 ();
 b15zdnd00an1n02x5 FILLER_135_1554 ();
 b15zdnd11an1n04x5 FILLER_135_1598 ();
 b15zdnd11an1n64x5 FILLER_135_1605 ();
 b15zdnd11an1n16x5 FILLER_135_1669 ();
 b15zdnd11an1n08x5 FILLER_135_1685 ();
 b15zdnd00an1n01x5 FILLER_135_1693 ();
 b15zdnd11an1n64x5 FILLER_135_1736 ();
 b15zdnd11an1n64x5 FILLER_135_1800 ();
 b15zdnd11an1n64x5 FILLER_135_1864 ();
 b15zdnd11an1n64x5 FILLER_135_1928 ();
 b15zdnd11an1n64x5 FILLER_135_1992 ();
 b15zdnd11an1n64x5 FILLER_135_2056 ();
 b15zdnd11an1n64x5 FILLER_135_2120 ();
 b15zdnd11an1n64x5 FILLER_135_2184 ();
 b15zdnd11an1n32x5 FILLER_135_2248 ();
 b15zdnd11an1n04x5 FILLER_135_2280 ();
 b15zdnd11an1n64x5 FILLER_136_8 ();
 b15zdnd11an1n64x5 FILLER_136_72 ();
 b15zdnd11an1n64x5 FILLER_136_136 ();
 b15zdnd11an1n64x5 FILLER_136_200 ();
 b15zdnd11an1n64x5 FILLER_136_264 ();
 b15zdnd11an1n64x5 FILLER_136_328 ();
 b15zdnd11an1n64x5 FILLER_136_392 ();
 b15zdnd11an1n64x5 FILLER_136_456 ();
 b15zdnd11an1n64x5 FILLER_136_520 ();
 b15zdnd11an1n64x5 FILLER_136_584 ();
 b15zdnd11an1n64x5 FILLER_136_648 ();
 b15zdnd11an1n04x5 FILLER_136_712 ();
 b15zdnd00an1n02x5 FILLER_136_716 ();
 b15zdnd11an1n16x5 FILLER_136_726 ();
 b15zdnd11an1n08x5 FILLER_136_742 ();
 b15zdnd00an1n02x5 FILLER_136_750 ();
 b15zdnd11an1n64x5 FILLER_136_756 ();
 b15zdnd11an1n64x5 FILLER_136_820 ();
 b15zdnd11an1n64x5 FILLER_136_884 ();
 b15zdnd11an1n64x5 FILLER_136_948 ();
 b15zdnd11an1n64x5 FILLER_136_1012 ();
 b15zdnd11an1n64x5 FILLER_136_1076 ();
 b15zdnd11an1n08x5 FILLER_136_1140 ();
 b15zdnd11an1n64x5 FILLER_136_1156 ();
 b15zdnd11an1n64x5 FILLER_136_1220 ();
 b15zdnd11an1n64x5 FILLER_136_1284 ();
 b15zdnd11an1n64x5 FILLER_136_1348 ();
 b15zdnd11an1n64x5 FILLER_136_1412 ();
 b15zdnd11an1n64x5 FILLER_136_1476 ();
 b15zdnd11an1n04x5 FILLER_136_1540 ();
 b15zdnd11an1n04x5 FILLER_136_1547 ();
 b15zdnd11an1n04x5 FILLER_136_1564 ();
 b15zdnd11an1n08x5 FILLER_136_1571 ();
 b15zdnd11an1n04x5 FILLER_136_1579 ();
 b15zdnd00an1n01x5 FILLER_136_1583 ();
 b15zdnd11an1n64x5 FILLER_136_1626 ();
 b15zdnd11an1n16x5 FILLER_136_1690 ();
 b15zdnd11an1n04x5 FILLER_136_1706 ();
 b15zdnd00an1n02x5 FILLER_136_1710 ();
 b15zdnd00an1n01x5 FILLER_136_1712 ();
 b15zdnd11an1n64x5 FILLER_136_1724 ();
 b15zdnd11an1n64x5 FILLER_136_1788 ();
 b15zdnd11an1n64x5 FILLER_136_1852 ();
 b15zdnd11an1n64x5 FILLER_136_1916 ();
 b15zdnd11an1n32x5 FILLER_136_1980 ();
 b15zdnd11an1n16x5 FILLER_136_2012 ();
 b15zdnd11an1n04x5 FILLER_136_2031 ();
 b15zdnd11an1n64x5 FILLER_136_2038 ();
 b15zdnd11an1n32x5 FILLER_136_2102 ();
 b15zdnd11an1n16x5 FILLER_136_2134 ();
 b15zdnd11an1n04x5 FILLER_136_2150 ();
 b15zdnd11an1n64x5 FILLER_136_2162 ();
 b15zdnd11an1n04x5 FILLER_136_2226 ();
 b15zdnd00an1n02x5 FILLER_136_2230 ();
 b15zdnd00an1n02x5 FILLER_136_2274 ();
 b15zdnd11an1n64x5 FILLER_137_0 ();
 b15zdnd11an1n04x5 FILLER_137_64 ();
 b15zdnd00an1n02x5 FILLER_137_68 ();
 b15zdnd00an1n01x5 FILLER_137_70 ();
 b15zdnd11an1n64x5 FILLER_137_78 ();
 b15zdnd11an1n64x5 FILLER_137_142 ();
 b15zdnd11an1n64x5 FILLER_137_206 ();
 b15zdnd11an1n64x5 FILLER_137_270 ();
 b15zdnd11an1n64x5 FILLER_137_334 ();
 b15zdnd11an1n64x5 FILLER_137_398 ();
 b15zdnd11an1n64x5 FILLER_137_462 ();
 b15zdnd11an1n64x5 FILLER_137_526 ();
 b15zdnd11an1n64x5 FILLER_137_590 ();
 b15zdnd11an1n64x5 FILLER_137_654 ();
 b15zdnd11an1n08x5 FILLER_137_718 ();
 b15zdnd00an1n02x5 FILLER_137_726 ();
 b15zdnd11an1n64x5 FILLER_137_734 ();
 b15zdnd11an1n64x5 FILLER_137_798 ();
 b15zdnd11an1n64x5 FILLER_137_862 ();
 b15zdnd11an1n64x5 FILLER_137_926 ();
 b15zdnd11an1n64x5 FILLER_137_990 ();
 b15zdnd11an1n32x5 FILLER_137_1054 ();
 b15zdnd11an1n16x5 FILLER_137_1086 ();
 b15zdnd11an1n08x5 FILLER_137_1102 ();
 b15zdnd11an1n04x5 FILLER_137_1110 ();
 b15zdnd00an1n02x5 FILLER_137_1114 ();
 b15zdnd11an1n64x5 FILLER_137_1119 ();
 b15zdnd11an1n64x5 FILLER_137_1183 ();
 b15zdnd11an1n64x5 FILLER_137_1247 ();
 b15zdnd11an1n64x5 FILLER_137_1311 ();
 b15zdnd11an1n64x5 FILLER_137_1375 ();
 b15zdnd11an1n64x5 FILLER_137_1439 ();
 b15zdnd11an1n16x5 FILLER_137_1503 ();
 b15zdnd11an1n08x5 FILLER_137_1519 ();
 b15zdnd00an1n02x5 FILLER_137_1527 ();
 b15zdnd00an1n01x5 FILLER_137_1529 ();
 b15zdnd11an1n16x5 FILLER_137_1536 ();
 b15zdnd11an1n08x5 FILLER_137_1552 ();
 b15zdnd11an1n64x5 FILLER_137_1570 ();
 b15zdnd11an1n64x5 FILLER_137_1634 ();
 b15zdnd11an1n64x5 FILLER_137_1698 ();
 b15zdnd11an1n64x5 FILLER_137_1762 ();
 b15zdnd11an1n64x5 FILLER_137_1826 ();
 b15zdnd11an1n64x5 FILLER_137_1890 ();
 b15zdnd11an1n32x5 FILLER_137_1954 ();
 b15zdnd11an1n16x5 FILLER_137_1986 ();
 b15zdnd11an1n08x5 FILLER_137_2002 ();
 b15zdnd11an1n64x5 FILLER_137_2062 ();
 b15zdnd11an1n64x5 FILLER_137_2126 ();
 b15zdnd11an1n32x5 FILLER_137_2190 ();
 b15zdnd11an1n04x5 FILLER_137_2222 ();
 b15zdnd11an1n04x5 FILLER_137_2229 ();
 b15zdnd11an1n04x5 FILLER_137_2236 ();
 b15zdnd00an1n02x5 FILLER_137_2282 ();
 b15zdnd11an1n64x5 FILLER_138_8 ();
 b15zdnd11an1n64x5 FILLER_138_72 ();
 b15zdnd11an1n64x5 FILLER_138_136 ();
 b15zdnd11an1n64x5 FILLER_138_200 ();
 b15zdnd11an1n64x5 FILLER_138_264 ();
 b15zdnd11an1n64x5 FILLER_138_328 ();
 b15zdnd11an1n64x5 FILLER_138_392 ();
 b15zdnd11an1n64x5 FILLER_138_456 ();
 b15zdnd11an1n64x5 FILLER_138_520 ();
 b15zdnd11an1n64x5 FILLER_138_584 ();
 b15zdnd11an1n64x5 FILLER_138_648 ();
 b15zdnd11an1n04x5 FILLER_138_712 ();
 b15zdnd00an1n02x5 FILLER_138_716 ();
 b15zdnd11an1n32x5 FILLER_138_726 ();
 b15zdnd11an1n16x5 FILLER_138_758 ();
 b15zdnd11an1n08x5 FILLER_138_774 ();
 b15zdnd00an1n02x5 FILLER_138_782 ();
 b15zdnd00an1n01x5 FILLER_138_784 ();
 b15zdnd11an1n08x5 FILLER_138_789 ();
 b15zdnd11an1n04x5 FILLER_138_797 ();
 b15zdnd00an1n02x5 FILLER_138_801 ();
 b15zdnd11an1n64x5 FILLER_138_809 ();
 b15zdnd11an1n08x5 FILLER_138_873 ();
 b15zdnd00an1n02x5 FILLER_138_881 ();
 b15zdnd00an1n01x5 FILLER_138_883 ();
 b15zdnd11an1n64x5 FILLER_138_888 ();
 b15zdnd11an1n64x5 FILLER_138_952 ();
 b15zdnd11an1n64x5 FILLER_138_1016 ();
 b15zdnd11an1n08x5 FILLER_138_1080 ();
 b15zdnd11an1n04x5 FILLER_138_1088 ();
 b15zdnd11an1n64x5 FILLER_138_1144 ();
 b15zdnd11an1n64x5 FILLER_138_1208 ();
 b15zdnd00an1n01x5 FILLER_138_1272 ();
 b15zdnd11an1n64x5 FILLER_138_1290 ();
 b15zdnd11an1n64x5 FILLER_138_1354 ();
 b15zdnd11an1n64x5 FILLER_138_1418 ();
 b15zdnd11an1n64x5 FILLER_138_1482 ();
 b15zdnd11an1n08x5 FILLER_138_1546 ();
 b15zdnd11an1n04x5 FILLER_138_1554 ();
 b15zdnd00an1n01x5 FILLER_138_1558 ();
 b15zdnd11an1n64x5 FILLER_138_1580 ();
 b15zdnd11an1n64x5 FILLER_138_1644 ();
 b15zdnd11an1n64x5 FILLER_138_1708 ();
 b15zdnd11an1n64x5 FILLER_138_1772 ();
 b15zdnd11an1n16x5 FILLER_138_1836 ();
 b15zdnd11an1n08x5 FILLER_138_1852 ();
 b15zdnd11an1n04x5 FILLER_138_1860 ();
 b15zdnd00an1n02x5 FILLER_138_1864 ();
 b15zdnd00an1n01x5 FILLER_138_1866 ();
 b15zdnd11an1n04x5 FILLER_138_1870 ();
 b15zdnd11an1n64x5 FILLER_138_1877 ();
 b15zdnd11an1n64x5 FILLER_138_1941 ();
 b15zdnd11an1n16x5 FILLER_138_2005 ();
 b15zdnd11an1n08x5 FILLER_138_2021 ();
 b15zdnd11an1n04x5 FILLER_138_2029 ();
 b15zdnd00an1n02x5 FILLER_138_2033 ();
 b15zdnd11an1n32x5 FILLER_138_2038 ();
 b15zdnd11an1n08x5 FILLER_138_2070 ();
 b15zdnd00an1n02x5 FILLER_138_2078 ();
 b15zdnd00an1n01x5 FILLER_138_2080 ();
 b15zdnd11an1n16x5 FILLER_138_2123 ();
 b15zdnd11an1n08x5 FILLER_138_2139 ();
 b15zdnd11an1n04x5 FILLER_138_2147 ();
 b15zdnd00an1n02x5 FILLER_138_2151 ();
 b15zdnd00an1n01x5 FILLER_138_2153 ();
 b15zdnd11an1n16x5 FILLER_138_2162 ();
 b15zdnd11an1n08x5 FILLER_138_2178 ();
 b15zdnd11an1n04x5 FILLER_138_2186 ();
 b15zdnd00an1n01x5 FILLER_138_2190 ();
 b15zdnd11an1n04x5 FILLER_138_2233 ();
 b15zdnd11an1n08x5 FILLER_138_2240 ();
 b15zdnd00an1n02x5 FILLER_138_2248 ();
 b15zdnd11an1n08x5 FILLER_138_2254 ();
 b15zdnd11an1n04x5 FILLER_138_2262 ();
 b15zdnd00an1n01x5 FILLER_138_2266 ();
 b15zdnd11an1n04x5 FILLER_138_2271 ();
 b15zdnd00an1n01x5 FILLER_138_2275 ();
 b15zdnd11an1n64x5 FILLER_139_0 ();
 b15zdnd11an1n04x5 FILLER_139_64 ();
 b15zdnd00an1n02x5 FILLER_139_68 ();
 b15zdnd00an1n01x5 FILLER_139_70 ();
 b15zdnd11an1n64x5 FILLER_139_98 ();
 b15zdnd11an1n64x5 FILLER_139_162 ();
 b15zdnd11an1n64x5 FILLER_139_226 ();
 b15zdnd11an1n64x5 FILLER_139_290 ();
 b15zdnd11an1n16x5 FILLER_139_354 ();
 b15zdnd11an1n08x5 FILLER_139_370 ();
 b15zdnd11an1n04x5 FILLER_139_378 ();
 b15zdnd00an1n02x5 FILLER_139_382 ();
 b15zdnd00an1n01x5 FILLER_139_384 ();
 b15zdnd11an1n64x5 FILLER_139_427 ();
 b15zdnd11an1n32x5 FILLER_139_491 ();
 b15zdnd11an1n16x5 FILLER_139_523 ();
 b15zdnd11an1n08x5 FILLER_139_539 ();
 b15zdnd00an1n02x5 FILLER_139_547 ();
 b15zdnd00an1n01x5 FILLER_139_549 ();
 b15zdnd11an1n64x5 FILLER_139_553 ();
 b15zdnd11an1n64x5 FILLER_139_617 ();
 b15zdnd11an1n64x5 FILLER_139_681 ();
 b15zdnd11an1n32x5 FILLER_139_745 ();
 b15zdnd11an1n08x5 FILLER_139_777 ();
 b15zdnd00an1n02x5 FILLER_139_785 ();
 b15zdnd11an1n64x5 FILLER_139_798 ();
 b15zdnd11an1n64x5 FILLER_139_862 ();
 b15zdnd11an1n64x5 FILLER_139_926 ();
 b15zdnd11an1n16x5 FILLER_139_990 ();
 b15zdnd11an1n04x5 FILLER_139_1006 ();
 b15zdnd00an1n02x5 FILLER_139_1010 ();
 b15zdnd00an1n01x5 FILLER_139_1012 ();
 b15zdnd11an1n64x5 FILLER_139_1016 ();
 b15zdnd11an1n08x5 FILLER_139_1080 ();
 b15zdnd00an1n01x5 FILLER_139_1088 ();
 b15zdnd11an1n64x5 FILLER_139_1141 ();
 b15zdnd11an1n64x5 FILLER_139_1205 ();
 b15zdnd11an1n64x5 FILLER_139_1269 ();
 b15zdnd11an1n64x5 FILLER_139_1333 ();
 b15zdnd11an1n64x5 FILLER_139_1397 ();
 b15zdnd11an1n64x5 FILLER_139_1461 ();
 b15zdnd11an1n64x5 FILLER_139_1525 ();
 b15zdnd11an1n64x5 FILLER_139_1589 ();
 b15zdnd11an1n64x5 FILLER_139_1653 ();
 b15zdnd11an1n64x5 FILLER_139_1717 ();
 b15zdnd11an1n32x5 FILLER_139_1781 ();
 b15zdnd11an1n16x5 FILLER_139_1813 ();
 b15zdnd11an1n08x5 FILLER_139_1829 ();
 b15zdnd11an1n04x5 FILLER_139_1837 ();
 b15zdnd00an1n01x5 FILLER_139_1841 ();
 b15zdnd11an1n64x5 FILLER_139_1894 ();
 b15zdnd11an1n16x5 FILLER_139_1958 ();
 b15zdnd11an1n08x5 FILLER_139_1974 ();
 b15zdnd11an1n04x5 FILLER_139_1982 ();
 b15zdnd00an1n01x5 FILLER_139_1986 ();
 b15zdnd11an1n16x5 FILLER_139_2029 ();
 b15zdnd00an1n02x5 FILLER_139_2045 ();
 b15zdnd00an1n01x5 FILLER_139_2047 ();
 b15zdnd11an1n64x5 FILLER_139_2090 ();
 b15zdnd11an1n08x5 FILLER_139_2154 ();
 b15zdnd11an1n04x5 FILLER_139_2204 ();
 b15zdnd11an1n16x5 FILLER_139_2260 ();
 b15zdnd11an1n08x5 FILLER_139_2276 ();
 b15zdnd11an1n64x5 FILLER_140_8 ();
 b15zdnd11an1n64x5 FILLER_140_72 ();
 b15zdnd11an1n64x5 FILLER_140_136 ();
 b15zdnd11an1n64x5 FILLER_140_200 ();
 b15zdnd11an1n08x5 FILLER_140_264 ();
 b15zdnd11an1n04x5 FILLER_140_272 ();
 b15zdnd00an1n01x5 FILLER_140_276 ();
 b15zdnd11an1n04x5 FILLER_140_280 ();
 b15zdnd11an1n64x5 FILLER_140_287 ();
 b15zdnd11an1n64x5 FILLER_140_351 ();
 b15zdnd11an1n32x5 FILLER_140_415 ();
 b15zdnd11an1n04x5 FILLER_140_447 ();
 b15zdnd11an1n08x5 FILLER_140_493 ();
 b15zdnd11an1n04x5 FILLER_140_501 ();
 b15zdnd00an1n01x5 FILLER_140_505 ();
 b15zdnd11an1n08x5 FILLER_140_513 ();
 b15zdnd00an1n02x5 FILLER_140_521 ();
 b15zdnd11an1n64x5 FILLER_140_575 ();
 b15zdnd11an1n64x5 FILLER_140_639 ();
 b15zdnd11an1n08x5 FILLER_140_703 ();
 b15zdnd11an1n04x5 FILLER_140_711 ();
 b15zdnd00an1n02x5 FILLER_140_715 ();
 b15zdnd00an1n01x5 FILLER_140_717 ();
 b15zdnd11an1n64x5 FILLER_140_726 ();
 b15zdnd11an1n64x5 FILLER_140_790 ();
 b15zdnd11an1n64x5 FILLER_140_854 ();
 b15zdnd11an1n64x5 FILLER_140_918 ();
 b15zdnd11an1n04x5 FILLER_140_982 ();
 b15zdnd11an1n64x5 FILLER_140_1038 ();
 b15zdnd11an1n04x5 FILLER_140_1102 ();
 b15zdnd00an1n02x5 FILLER_140_1106 ();
 b15zdnd00an1n01x5 FILLER_140_1108 ();
 b15zdnd11an1n04x5 FILLER_140_1112 ();
 b15zdnd11an1n04x5 FILLER_140_1119 ();
 b15zdnd11an1n64x5 FILLER_140_1126 ();
 b15zdnd11an1n64x5 FILLER_140_1190 ();
 b15zdnd11an1n64x5 FILLER_140_1254 ();
 b15zdnd11an1n64x5 FILLER_140_1318 ();
 b15zdnd11an1n64x5 FILLER_140_1382 ();
 b15zdnd11an1n64x5 FILLER_140_1446 ();
 b15zdnd11an1n64x5 FILLER_140_1510 ();
 b15zdnd11an1n64x5 FILLER_140_1574 ();
 b15zdnd11an1n64x5 FILLER_140_1638 ();
 b15zdnd11an1n64x5 FILLER_140_1702 ();
 b15zdnd11an1n64x5 FILLER_140_1766 ();
 b15zdnd11an1n32x5 FILLER_140_1830 ();
 b15zdnd11an1n04x5 FILLER_140_1862 ();
 b15zdnd00an1n01x5 FILLER_140_1866 ();
 b15zdnd11an1n64x5 FILLER_140_1870 ();
 b15zdnd11an1n08x5 FILLER_140_1934 ();
 b15zdnd11an1n04x5 FILLER_140_1942 ();
 b15zdnd00an1n01x5 FILLER_140_1946 ();
 b15zdnd11an1n64x5 FILLER_140_1989 ();
 b15zdnd11an1n64x5 FILLER_140_2053 ();
 b15zdnd11an1n32x5 FILLER_140_2117 ();
 b15zdnd11an1n04x5 FILLER_140_2149 ();
 b15zdnd00an1n01x5 FILLER_140_2153 ();
 b15zdnd11an1n64x5 FILLER_140_2162 ();
 b15zdnd11an1n04x5 FILLER_140_2226 ();
 b15zdnd00an1n01x5 FILLER_140_2230 ();
 b15zdnd11an1n04x5 FILLER_140_2270 ();
 b15zdnd00an1n02x5 FILLER_140_2274 ();
 b15zdnd11an1n64x5 FILLER_141_0 ();
 b15zdnd11an1n64x5 FILLER_141_64 ();
 b15zdnd11an1n64x5 FILLER_141_128 ();
 b15zdnd11an1n16x5 FILLER_141_192 ();
 b15zdnd00an1n02x5 FILLER_141_208 ();
 b15zdnd00an1n01x5 FILLER_141_210 ();
 b15zdnd11an1n08x5 FILLER_141_227 ();
 b15zdnd00an1n02x5 FILLER_141_235 ();
 b15zdnd00an1n01x5 FILLER_141_237 ();
 b15zdnd11an1n04x5 FILLER_141_246 ();
 b15zdnd11an1n08x5 FILLER_141_253 ();
 b15zdnd11an1n04x5 FILLER_141_261 ();
 b15zdnd11an1n64x5 FILLER_141_307 ();
 b15zdnd11an1n64x5 FILLER_141_371 ();
 b15zdnd11an1n64x5 FILLER_141_435 ();
 b15zdnd11an1n16x5 FILLER_141_499 ();
 b15zdnd00an1n01x5 FILLER_141_515 ();
 b15zdnd11an1n64x5 FILLER_141_558 ();
 b15zdnd11an1n64x5 FILLER_141_622 ();
 b15zdnd11an1n64x5 FILLER_141_686 ();
 b15zdnd11an1n04x5 FILLER_141_750 ();
 b15zdnd00an1n01x5 FILLER_141_754 ();
 b15zdnd11an1n64x5 FILLER_141_799 ();
 b15zdnd11an1n64x5 FILLER_141_863 ();
 b15zdnd11an1n64x5 FILLER_141_927 ();
 b15zdnd11an1n08x5 FILLER_141_991 ();
 b15zdnd11an1n04x5 FILLER_141_999 ();
 b15zdnd00an1n01x5 FILLER_141_1003 ();
 b15zdnd11an1n04x5 FILLER_141_1007 ();
 b15zdnd00an1n01x5 FILLER_141_1011 ();
 b15zdnd11an1n64x5 FILLER_141_1015 ();
 b15zdnd11an1n32x5 FILLER_141_1079 ();
 b15zdnd11an1n04x5 FILLER_141_1111 ();
 b15zdnd11an1n04x5 FILLER_141_1118 ();
 b15zdnd11an1n64x5 FILLER_141_1125 ();
 b15zdnd11an1n64x5 FILLER_141_1189 ();
 b15zdnd11an1n08x5 FILLER_141_1253 ();
 b15zdnd11an1n04x5 FILLER_141_1261 ();
 b15zdnd00an1n02x5 FILLER_141_1265 ();
 b15zdnd11an1n32x5 FILLER_141_1275 ();
 b15zdnd11an1n08x5 FILLER_141_1307 ();
 b15zdnd11an1n04x5 FILLER_141_1315 ();
 b15zdnd00an1n02x5 FILLER_141_1319 ();
 b15zdnd00an1n01x5 FILLER_141_1321 ();
 b15zdnd11an1n08x5 FILLER_141_1329 ();
 b15zdnd00an1n01x5 FILLER_141_1337 ();
 b15zdnd11an1n64x5 FILLER_141_1347 ();
 b15zdnd11an1n64x5 FILLER_141_1411 ();
 b15zdnd11an1n64x5 FILLER_141_1475 ();
 b15zdnd11an1n64x5 FILLER_141_1539 ();
 b15zdnd11an1n64x5 FILLER_141_1603 ();
 b15zdnd11an1n04x5 FILLER_141_1667 ();
 b15zdnd11an1n08x5 FILLER_141_1674 ();
 b15zdnd00an1n02x5 FILLER_141_1682 ();
 b15zdnd00an1n01x5 FILLER_141_1684 ();
 b15zdnd11an1n64x5 FILLER_141_1689 ();
 b15zdnd11an1n64x5 FILLER_141_1753 ();
 b15zdnd11an1n64x5 FILLER_141_1817 ();
 b15zdnd11an1n64x5 FILLER_141_1881 ();
 b15zdnd11an1n64x5 FILLER_141_1945 ();
 b15zdnd11an1n64x5 FILLER_141_2009 ();
 b15zdnd11an1n64x5 FILLER_141_2073 ();
 b15zdnd11an1n64x5 FILLER_141_2137 ();
 b15zdnd11an1n64x5 FILLER_141_2201 ();
 b15zdnd11an1n16x5 FILLER_141_2265 ();
 b15zdnd00an1n02x5 FILLER_141_2281 ();
 b15zdnd00an1n01x5 FILLER_141_2283 ();
 b15zdnd11an1n64x5 FILLER_142_8 ();
 b15zdnd11an1n64x5 FILLER_142_72 ();
 b15zdnd11an1n64x5 FILLER_142_136 ();
 b15zdnd11an1n32x5 FILLER_142_200 ();
 b15zdnd11an1n16x5 FILLER_142_232 ();
 b15zdnd00an1n02x5 FILLER_142_248 ();
 b15zdnd11an1n04x5 FILLER_142_253 ();
 b15zdnd11an1n64x5 FILLER_142_309 ();
 b15zdnd11an1n08x5 FILLER_142_373 ();
 b15zdnd00an1n02x5 FILLER_142_381 ();
 b15zdnd00an1n01x5 FILLER_142_383 ();
 b15zdnd11an1n64x5 FILLER_142_426 ();
 b15zdnd11an1n32x5 FILLER_142_490 ();
 b15zdnd11an1n16x5 FILLER_142_522 ();
 b15zdnd11an1n04x5 FILLER_142_538 ();
 b15zdnd11an1n04x5 FILLER_142_545 ();
 b15zdnd11an1n64x5 FILLER_142_552 ();
 b15zdnd11an1n64x5 FILLER_142_616 ();
 b15zdnd11an1n32x5 FILLER_142_680 ();
 b15zdnd11an1n04x5 FILLER_142_712 ();
 b15zdnd00an1n02x5 FILLER_142_716 ();
 b15zdnd11an1n08x5 FILLER_142_726 ();
 b15zdnd11an1n04x5 FILLER_142_734 ();
 b15zdnd11an1n16x5 FILLER_142_749 ();
 b15zdnd11an1n04x5 FILLER_142_765 ();
 b15zdnd00an1n02x5 FILLER_142_769 ();
 b15zdnd00an1n01x5 FILLER_142_771 ();
 b15zdnd11an1n04x5 FILLER_142_775 ();
 b15zdnd11an1n64x5 FILLER_142_782 ();
 b15zdnd11an1n64x5 FILLER_142_846 ();
 b15zdnd11an1n64x5 FILLER_142_910 ();
 b15zdnd11an1n64x5 FILLER_142_974 ();
 b15zdnd11an1n64x5 FILLER_142_1038 ();
 b15zdnd11an1n64x5 FILLER_142_1102 ();
 b15zdnd11an1n64x5 FILLER_142_1166 ();
 b15zdnd11an1n64x5 FILLER_142_1230 ();
 b15zdnd11an1n64x5 FILLER_142_1294 ();
 b15zdnd11an1n64x5 FILLER_142_1358 ();
 b15zdnd11an1n64x5 FILLER_142_1422 ();
 b15zdnd11an1n64x5 FILLER_142_1486 ();
 b15zdnd11an1n08x5 FILLER_142_1550 ();
 b15zdnd11an1n64x5 FILLER_142_1568 ();
 b15zdnd11an1n64x5 FILLER_142_1632 ();
 b15zdnd11an1n64x5 FILLER_142_1696 ();
 b15zdnd11an1n08x5 FILLER_142_1760 ();
 b15zdnd11an1n04x5 FILLER_142_1768 ();
 b15zdnd00an1n02x5 FILLER_142_1772 ();
 b15zdnd11an1n64x5 FILLER_142_1785 ();
 b15zdnd11an1n64x5 FILLER_142_1849 ();
 b15zdnd11an1n64x5 FILLER_142_1913 ();
 b15zdnd11an1n64x5 FILLER_142_1977 ();
 b15zdnd11an1n08x5 FILLER_142_2041 ();
 b15zdnd11an1n32x5 FILLER_142_2091 ();
 b15zdnd11an1n16x5 FILLER_142_2123 ();
 b15zdnd11an1n08x5 FILLER_142_2139 ();
 b15zdnd11an1n04x5 FILLER_142_2147 ();
 b15zdnd00an1n02x5 FILLER_142_2151 ();
 b15zdnd00an1n01x5 FILLER_142_2153 ();
 b15zdnd11an1n64x5 FILLER_142_2162 ();
 b15zdnd00an1n02x5 FILLER_142_2226 ();
 b15zdnd11an1n16x5 FILLER_142_2259 ();
 b15zdnd00an1n01x5 FILLER_142_2275 ();
 b15zdnd11an1n64x5 FILLER_143_0 ();
 b15zdnd11an1n64x5 FILLER_143_64 ();
 b15zdnd11an1n64x5 FILLER_143_128 ();
 b15zdnd11an1n32x5 FILLER_143_192 ();
 b15zdnd11an1n04x5 FILLER_143_224 ();
 b15zdnd11an1n04x5 FILLER_143_280 ();
 b15zdnd11an1n64x5 FILLER_143_326 ();
 b15zdnd11an1n64x5 FILLER_143_390 ();
 b15zdnd11an1n64x5 FILLER_143_454 ();
 b15zdnd11an1n64x5 FILLER_143_518 ();
 b15zdnd11an1n64x5 FILLER_143_582 ();
 b15zdnd11an1n64x5 FILLER_143_646 ();
 b15zdnd11an1n64x5 FILLER_143_710 ();
 b15zdnd00an1n02x5 FILLER_143_774 ();
 b15zdnd00an1n01x5 FILLER_143_776 ();
 b15zdnd11an1n64x5 FILLER_143_780 ();
 b15zdnd11an1n64x5 FILLER_143_844 ();
 b15zdnd11an1n32x5 FILLER_143_908 ();
 b15zdnd11an1n16x5 FILLER_143_940 ();
 b15zdnd11an1n08x5 FILLER_143_956 ();
 b15zdnd11an1n64x5 FILLER_143_1016 ();
 b15zdnd11an1n64x5 FILLER_143_1080 ();
 b15zdnd11an1n32x5 FILLER_143_1144 ();
 b15zdnd11an1n16x5 FILLER_143_1176 ();
 b15zdnd11an1n04x5 FILLER_143_1192 ();
 b15zdnd00an1n01x5 FILLER_143_1196 ();
 b15zdnd11an1n64x5 FILLER_143_1223 ();
 b15zdnd11an1n64x5 FILLER_143_1287 ();
 b15zdnd11an1n64x5 FILLER_143_1351 ();
 b15zdnd11an1n64x5 FILLER_143_1415 ();
 b15zdnd11an1n64x5 FILLER_143_1479 ();
 b15zdnd11an1n64x5 FILLER_143_1543 ();
 b15zdnd11an1n64x5 FILLER_143_1607 ();
 b15zdnd11an1n64x5 FILLER_143_1671 ();
 b15zdnd11an1n64x5 FILLER_143_1735 ();
 b15zdnd11an1n32x5 FILLER_143_1799 ();
 b15zdnd11an1n08x5 FILLER_143_1831 ();
 b15zdnd11an1n32x5 FILLER_143_1843 ();
 b15zdnd11an1n08x5 FILLER_143_1875 ();
 b15zdnd11an1n64x5 FILLER_143_1907 ();
 b15zdnd11an1n64x5 FILLER_143_1971 ();
 b15zdnd11an1n04x5 FILLER_143_2035 ();
 b15zdnd00an1n02x5 FILLER_143_2039 ();
 b15zdnd11an1n64x5 FILLER_143_2083 ();
 b15zdnd11an1n64x5 FILLER_143_2147 ();
 b15zdnd11an1n16x5 FILLER_143_2211 ();
 b15zdnd11an1n04x5 FILLER_143_2227 ();
 b15zdnd11an1n04x5 FILLER_143_2268 ();
 b15zdnd11an1n08x5 FILLER_143_2276 ();
 b15zdnd11an1n64x5 FILLER_144_8 ();
 b15zdnd11an1n64x5 FILLER_144_72 ();
 b15zdnd11an1n64x5 FILLER_144_136 ();
 b15zdnd11an1n32x5 FILLER_144_200 ();
 b15zdnd11an1n08x5 FILLER_144_232 ();
 b15zdnd11an1n04x5 FILLER_144_240 ();
 b15zdnd00an1n02x5 FILLER_144_244 ();
 b15zdnd00an1n01x5 FILLER_144_246 ();
 b15zdnd11an1n04x5 FILLER_144_250 ();
 b15zdnd11an1n64x5 FILLER_144_296 ();
 b15zdnd11an1n16x5 FILLER_144_360 ();
 b15zdnd11an1n04x5 FILLER_144_376 ();
 b15zdnd00an1n01x5 FILLER_144_380 ();
 b15zdnd11an1n04x5 FILLER_144_413 ();
 b15zdnd11an1n64x5 FILLER_144_420 ();
 b15zdnd11an1n64x5 FILLER_144_484 ();
 b15zdnd11an1n64x5 FILLER_144_548 ();
 b15zdnd11an1n16x5 FILLER_144_612 ();
 b15zdnd00an1n02x5 FILLER_144_628 ();
 b15zdnd11an1n64x5 FILLER_144_639 ();
 b15zdnd11an1n08x5 FILLER_144_703 ();
 b15zdnd11an1n04x5 FILLER_144_711 ();
 b15zdnd00an1n02x5 FILLER_144_715 ();
 b15zdnd00an1n01x5 FILLER_144_717 ();
 b15zdnd11an1n64x5 FILLER_144_726 ();
 b15zdnd11an1n64x5 FILLER_144_790 ();
 b15zdnd11an1n64x5 FILLER_144_854 ();
 b15zdnd11an1n64x5 FILLER_144_918 ();
 b15zdnd00an1n01x5 FILLER_144_982 ();
 b15zdnd11an1n04x5 FILLER_144_986 ();
 b15zdnd11an1n04x5 FILLER_144_993 ();
 b15zdnd11an1n64x5 FILLER_144_1000 ();
 b15zdnd11an1n64x5 FILLER_144_1064 ();
 b15zdnd11an1n32x5 FILLER_144_1128 ();
 b15zdnd11an1n08x5 FILLER_144_1160 ();
 b15zdnd11an1n64x5 FILLER_144_1171 ();
 b15zdnd11an1n64x5 FILLER_144_1235 ();
 b15zdnd11an1n64x5 FILLER_144_1299 ();
 b15zdnd11an1n64x5 FILLER_144_1363 ();
 b15zdnd11an1n64x5 FILLER_144_1427 ();
 b15zdnd11an1n64x5 FILLER_144_1491 ();
 b15zdnd11an1n64x5 FILLER_144_1555 ();
 b15zdnd11an1n32x5 FILLER_144_1619 ();
 b15zdnd11an1n16x5 FILLER_144_1651 ();
 b15zdnd11an1n32x5 FILLER_144_1688 ();
 b15zdnd11an1n16x5 FILLER_144_1720 ();
 b15zdnd11an1n08x5 FILLER_144_1736 ();
 b15zdnd00an1n01x5 FILLER_144_1744 ();
 b15zdnd11an1n04x5 FILLER_144_1765 ();
 b15zdnd00an1n02x5 FILLER_144_1769 ();
 b15zdnd00an1n01x5 FILLER_144_1771 ();
 b15zdnd11an1n64x5 FILLER_144_1787 ();
 b15zdnd11an1n32x5 FILLER_144_1851 ();
 b15zdnd11an1n16x5 FILLER_144_1883 ();
 b15zdnd11an1n04x5 FILLER_144_1899 ();
 b15zdnd11an1n04x5 FILLER_144_1906 ();
 b15zdnd11an1n08x5 FILLER_144_1913 ();
 b15zdnd00an1n01x5 FILLER_144_1921 ();
 b15zdnd11an1n64x5 FILLER_144_1925 ();
 b15zdnd11an1n32x5 FILLER_144_1989 ();
 b15zdnd11an1n08x5 FILLER_144_2021 ();
 b15zdnd11an1n04x5 FILLER_144_2029 ();
 b15zdnd00an1n01x5 FILLER_144_2033 ();
 b15zdnd11an1n64x5 FILLER_144_2037 ();
 b15zdnd11an1n32x5 FILLER_144_2101 ();
 b15zdnd11an1n16x5 FILLER_144_2133 ();
 b15zdnd11an1n04x5 FILLER_144_2149 ();
 b15zdnd00an1n01x5 FILLER_144_2153 ();
 b15zdnd11an1n64x5 FILLER_144_2162 ();
 b15zdnd11an1n32x5 FILLER_144_2226 ();
 b15zdnd11an1n16x5 FILLER_144_2258 ();
 b15zdnd00an1n02x5 FILLER_144_2274 ();
 b15zdnd11an1n64x5 FILLER_145_0 ();
 b15zdnd11an1n64x5 FILLER_145_64 ();
 b15zdnd11an1n64x5 FILLER_145_128 ();
 b15zdnd11an1n32x5 FILLER_145_192 ();
 b15zdnd11an1n16x5 FILLER_145_224 ();
 b15zdnd11an1n08x5 FILLER_145_240 ();
 b15zdnd11an1n04x5 FILLER_145_248 ();
 b15zdnd00an1n02x5 FILLER_145_252 ();
 b15zdnd00an1n01x5 FILLER_145_254 ();
 b15zdnd11an1n16x5 FILLER_145_258 ();
 b15zdnd11an1n08x5 FILLER_145_274 ();
 b15zdnd00an1n02x5 FILLER_145_282 ();
 b15zdnd11an1n64x5 FILLER_145_287 ();
 b15zdnd11an1n32x5 FILLER_145_351 ();
 b15zdnd11an1n16x5 FILLER_145_383 ();
 b15zdnd11an1n04x5 FILLER_145_399 ();
 b15zdnd00an1n01x5 FILLER_145_403 ();
 b15zdnd11an1n64x5 FILLER_145_407 ();
 b15zdnd11an1n64x5 FILLER_145_471 ();
 b15zdnd11an1n64x5 FILLER_145_535 ();
 b15zdnd11an1n16x5 FILLER_145_599 ();
 b15zdnd11an1n08x5 FILLER_145_615 ();
 b15zdnd11an1n04x5 FILLER_145_623 ();
 b15zdnd11an1n64x5 FILLER_145_636 ();
 b15zdnd11an1n64x5 FILLER_145_700 ();
 b15zdnd11an1n64x5 FILLER_145_764 ();
 b15zdnd11an1n64x5 FILLER_145_828 ();
 b15zdnd11an1n64x5 FILLER_145_892 ();
 b15zdnd11an1n16x5 FILLER_145_956 ();
 b15zdnd11an1n08x5 FILLER_145_972 ();
 b15zdnd00an1n01x5 FILLER_145_980 ();
 b15zdnd11an1n04x5 FILLER_145_984 ();
 b15zdnd11an1n04x5 FILLER_145_1015 ();
 b15zdnd11an1n16x5 FILLER_145_1028 ();
 b15zdnd11an1n08x5 FILLER_145_1044 ();
 b15zdnd11an1n04x5 FILLER_145_1052 ();
 b15zdnd00an1n02x5 FILLER_145_1056 ();
 b15zdnd11an1n04x5 FILLER_145_1067 ();
 b15zdnd11an1n32x5 FILLER_145_1080 ();
 b15zdnd11an1n16x5 FILLER_145_1112 ();
 b15zdnd11an1n08x5 FILLER_145_1128 ();
 b15zdnd11an1n04x5 FILLER_145_1136 ();
 b15zdnd00an1n02x5 FILLER_145_1140 ();
 b15zdnd11an1n64x5 FILLER_145_1194 ();
 b15zdnd11an1n64x5 FILLER_145_1258 ();
 b15zdnd11an1n16x5 FILLER_145_1330 ();
 b15zdnd11an1n04x5 FILLER_145_1346 ();
 b15zdnd00an1n02x5 FILLER_145_1350 ();
 b15zdnd00an1n01x5 FILLER_145_1352 ();
 b15zdnd11an1n16x5 FILLER_145_1356 ();
 b15zdnd00an1n02x5 FILLER_145_1372 ();
 b15zdnd11an1n32x5 FILLER_145_1377 ();
 b15zdnd11an1n04x5 FILLER_145_1409 ();
 b15zdnd11an1n64x5 FILLER_145_1455 ();
 b15zdnd11an1n64x5 FILLER_145_1519 ();
 b15zdnd11an1n64x5 FILLER_145_1583 ();
 b15zdnd11an1n64x5 FILLER_145_1647 ();
 b15zdnd11an1n64x5 FILLER_145_1711 ();
 b15zdnd11an1n64x5 FILLER_145_1775 ();
 b15zdnd11an1n32x5 FILLER_145_1839 ();
 b15zdnd11an1n08x5 FILLER_145_1871 ();
 b15zdnd00an1n01x5 FILLER_145_1879 ();
 b15zdnd11an1n64x5 FILLER_145_1932 ();
 b15zdnd11an1n16x5 FILLER_145_1996 ();
 b15zdnd11an1n08x5 FILLER_145_2012 ();
 b15zdnd00an1n02x5 FILLER_145_2020 ();
 b15zdnd00an1n01x5 FILLER_145_2022 ();
 b15zdnd11an1n04x5 FILLER_145_2026 ();
 b15zdnd11an1n04x5 FILLER_145_2039 ();
 b15zdnd11an1n04x5 FILLER_145_2052 ();
 b15zdnd11an1n64x5 FILLER_145_2063 ();
 b15zdnd11an1n64x5 FILLER_145_2127 ();
 b15zdnd11an1n64x5 FILLER_145_2191 ();
 b15zdnd00an1n02x5 FILLER_145_2255 ();
 b15zdnd00an1n01x5 FILLER_145_2257 ();
 b15zdnd11an1n16x5 FILLER_145_2262 ();
 b15zdnd11an1n04x5 FILLER_145_2278 ();
 b15zdnd00an1n02x5 FILLER_145_2282 ();
 b15zdnd11an1n08x5 FILLER_146_8 ();
 b15zdnd11an1n04x5 FILLER_146_16 ();
 b15zdnd00an1n02x5 FILLER_146_20 ();
 b15zdnd00an1n01x5 FILLER_146_22 ();
 b15zdnd11an1n04x5 FILLER_146_27 ();
 b15zdnd11an1n64x5 FILLER_146_35 ();
 b15zdnd11an1n64x5 FILLER_146_99 ();
 b15zdnd11an1n64x5 FILLER_146_163 ();
 b15zdnd11an1n64x5 FILLER_146_227 ();
 b15zdnd11an1n64x5 FILLER_146_291 ();
 b15zdnd11an1n64x5 FILLER_146_355 ();
 b15zdnd11an1n64x5 FILLER_146_419 ();
 b15zdnd11an1n64x5 FILLER_146_483 ();
 b15zdnd11an1n64x5 FILLER_146_547 ();
 b15zdnd11an1n64x5 FILLER_146_611 ();
 b15zdnd11an1n32x5 FILLER_146_675 ();
 b15zdnd11an1n08x5 FILLER_146_707 ();
 b15zdnd00an1n02x5 FILLER_146_715 ();
 b15zdnd00an1n01x5 FILLER_146_717 ();
 b15zdnd11an1n64x5 FILLER_146_726 ();
 b15zdnd11an1n64x5 FILLER_146_790 ();
 b15zdnd11an1n64x5 FILLER_146_854 ();
 b15zdnd11an1n32x5 FILLER_146_918 ();
 b15zdnd11an1n08x5 FILLER_146_950 ();
 b15zdnd11an1n04x5 FILLER_146_958 ();
 b15zdnd00an1n02x5 FILLER_146_962 ();
 b15zdnd00an1n01x5 FILLER_146_964 ();
 b15zdnd11an1n64x5 FILLER_146_1017 ();
 b15zdnd11an1n64x5 FILLER_146_1081 ();
 b15zdnd11an1n16x5 FILLER_146_1145 ();
 b15zdnd11an1n04x5 FILLER_146_1161 ();
 b15zdnd11an1n04x5 FILLER_146_1168 ();
 b15zdnd11an1n64x5 FILLER_146_1175 ();
 b15zdnd11an1n16x5 FILLER_146_1239 ();
 b15zdnd00an1n02x5 FILLER_146_1255 ();
 b15zdnd00an1n01x5 FILLER_146_1257 ();
 b15zdnd11an1n16x5 FILLER_146_1300 ();
 b15zdnd00an1n01x5 FILLER_146_1316 ();
 b15zdnd11an1n04x5 FILLER_146_1359 ();
 b15zdnd00an1n02x5 FILLER_146_1363 ();
 b15zdnd11an1n04x5 FILLER_146_1368 ();
 b15zdnd11an1n64x5 FILLER_146_1375 ();
 b15zdnd11an1n16x5 FILLER_146_1439 ();
 b15zdnd11an1n64x5 FILLER_146_1458 ();
 b15zdnd11an1n64x5 FILLER_146_1522 ();
 b15zdnd11an1n64x5 FILLER_146_1586 ();
 b15zdnd11an1n64x5 FILLER_146_1650 ();
 b15zdnd11an1n64x5 FILLER_146_1714 ();
 b15zdnd11an1n32x5 FILLER_146_1778 ();
 b15zdnd11an1n04x5 FILLER_146_1810 ();
 b15zdnd00an1n02x5 FILLER_146_1814 ();
 b15zdnd00an1n01x5 FILLER_146_1816 ();
 b15zdnd11an1n64x5 FILLER_146_1822 ();
 b15zdnd11an1n64x5 FILLER_146_1886 ();
 b15zdnd11an1n32x5 FILLER_146_1950 ();
 b15zdnd11an1n16x5 FILLER_146_1982 ();
 b15zdnd11an1n08x5 FILLER_146_1998 ();
 b15zdnd11an1n64x5 FILLER_146_2058 ();
 b15zdnd11an1n32x5 FILLER_146_2122 ();
 b15zdnd11an1n32x5 FILLER_146_2162 ();
 b15zdnd11an1n16x5 FILLER_146_2194 ();
 b15zdnd00an1n01x5 FILLER_146_2210 ();
 b15zdnd11an1n32x5 FILLER_146_2242 ();
 b15zdnd00an1n02x5 FILLER_146_2274 ();
 b15zdnd00an1n02x5 FILLER_147_0 ();
 b15zdnd11an1n64x5 FILLER_147_7 ();
 b15zdnd11an1n64x5 FILLER_147_71 ();
 b15zdnd11an1n64x5 FILLER_147_135 ();
 b15zdnd11an1n64x5 FILLER_147_199 ();
 b15zdnd11an1n64x5 FILLER_147_263 ();
 b15zdnd11an1n64x5 FILLER_147_327 ();
 b15zdnd11an1n64x5 FILLER_147_391 ();
 b15zdnd11an1n64x5 FILLER_147_455 ();
 b15zdnd11an1n64x5 FILLER_147_519 ();
 b15zdnd11an1n64x5 FILLER_147_583 ();
 b15zdnd11an1n64x5 FILLER_147_647 ();
 b15zdnd11an1n64x5 FILLER_147_711 ();
 b15zdnd11an1n64x5 FILLER_147_775 ();
 b15zdnd11an1n32x5 FILLER_147_839 ();
 b15zdnd11an1n08x5 FILLER_147_871 ();
 b15zdnd11an1n04x5 FILLER_147_879 ();
 b15zdnd00an1n02x5 FILLER_147_883 ();
 b15zdnd00an1n01x5 FILLER_147_885 ();
 b15zdnd11an1n64x5 FILLER_147_905 ();
 b15zdnd11an1n16x5 FILLER_147_969 ();
 b15zdnd11an1n04x5 FILLER_147_988 ();
 b15zdnd11an1n64x5 FILLER_147_995 ();
 b15zdnd11an1n64x5 FILLER_147_1059 ();
 b15zdnd11an1n32x5 FILLER_147_1123 ();
 b15zdnd11an1n08x5 FILLER_147_1155 ();
 b15zdnd11an1n04x5 FILLER_147_1163 ();
 b15zdnd00an1n02x5 FILLER_147_1167 ();
 b15zdnd11an1n64x5 FILLER_147_1189 ();
 b15zdnd11an1n16x5 FILLER_147_1253 ();
 b15zdnd00an1n02x5 FILLER_147_1269 ();
 b15zdnd00an1n01x5 FILLER_147_1271 ();
 b15zdnd11an1n64x5 FILLER_147_1281 ();
 b15zdnd11an1n04x5 FILLER_147_1345 ();
 b15zdnd11an1n32x5 FILLER_147_1401 ();
 b15zdnd11an1n16x5 FILLER_147_1433 ();
 b15zdnd11an1n04x5 FILLER_147_1452 ();
 b15zdnd11an1n04x5 FILLER_147_1459 ();
 b15zdnd11an1n16x5 FILLER_147_1466 ();
 b15zdnd11an1n04x5 FILLER_147_1482 ();
 b15zdnd00an1n02x5 FILLER_147_1486 ();
 b15zdnd00an1n01x5 FILLER_147_1488 ();
 b15zdnd11an1n32x5 FILLER_147_1497 ();
 b15zdnd11an1n16x5 FILLER_147_1529 ();
 b15zdnd11an1n04x5 FILLER_147_1545 ();
 b15zdnd11an1n64x5 FILLER_147_1565 ();
 b15zdnd11an1n64x5 FILLER_147_1629 ();
 b15zdnd11an1n64x5 FILLER_147_1693 ();
 b15zdnd11an1n64x5 FILLER_147_1757 ();
 b15zdnd11an1n64x5 FILLER_147_1821 ();
 b15zdnd11an1n64x5 FILLER_147_1885 ();
 b15zdnd11an1n64x5 FILLER_147_1949 ();
 b15zdnd11an1n08x5 FILLER_147_2013 ();
 b15zdnd11an1n04x5 FILLER_147_2063 ();
 b15zdnd11an1n64x5 FILLER_147_2109 ();
 b15zdnd11an1n08x5 FILLER_147_2173 ();
 b15zdnd00an1n02x5 FILLER_147_2181 ();
 b15zdnd00an1n01x5 FILLER_147_2183 ();
 b15zdnd11an1n04x5 FILLER_147_2229 ();
 b15zdnd11an1n32x5 FILLER_147_2236 ();
 b15zdnd11an1n16x5 FILLER_147_2268 ();
 b15zdnd11an1n64x5 FILLER_148_8 ();
 b15zdnd11an1n64x5 FILLER_148_72 ();
 b15zdnd11an1n64x5 FILLER_148_136 ();
 b15zdnd11an1n32x5 FILLER_148_200 ();
 b15zdnd11an1n16x5 FILLER_148_232 ();
 b15zdnd11an1n08x5 FILLER_148_248 ();
 b15zdnd00an1n02x5 FILLER_148_256 ();
 b15zdnd00an1n01x5 FILLER_148_258 ();
 b15zdnd11an1n64x5 FILLER_148_301 ();
 b15zdnd11an1n64x5 FILLER_148_365 ();
 b15zdnd11an1n64x5 FILLER_148_429 ();
 b15zdnd11an1n08x5 FILLER_148_493 ();
 b15zdnd11an1n04x5 FILLER_148_501 ();
 b15zdnd00an1n01x5 FILLER_148_505 ();
 b15zdnd11an1n04x5 FILLER_148_509 ();
 b15zdnd00an1n01x5 FILLER_148_513 ();
 b15zdnd11an1n64x5 FILLER_148_517 ();
 b15zdnd11an1n64x5 FILLER_148_581 ();
 b15zdnd11an1n64x5 FILLER_148_645 ();
 b15zdnd11an1n08x5 FILLER_148_709 ();
 b15zdnd00an1n01x5 FILLER_148_717 ();
 b15zdnd11an1n64x5 FILLER_148_726 ();
 b15zdnd11an1n32x5 FILLER_148_790 ();
 b15zdnd11an1n04x5 FILLER_148_822 ();
 b15zdnd00an1n02x5 FILLER_148_826 ();
 b15zdnd00an1n01x5 FILLER_148_828 ();
 b15zdnd11an1n04x5 FILLER_148_842 ();
 b15zdnd11an1n04x5 FILLER_148_849 ();
 b15zdnd11an1n64x5 FILLER_148_863 ();
 b15zdnd11an1n64x5 FILLER_148_927 ();
 b15zdnd00an1n02x5 FILLER_148_991 ();
 b15zdnd11an1n64x5 FILLER_148_996 ();
 b15zdnd11an1n64x5 FILLER_148_1060 ();
 b15zdnd11an1n64x5 FILLER_148_1124 ();
 b15zdnd11an1n64x5 FILLER_148_1188 ();
 b15zdnd11an1n64x5 FILLER_148_1252 ();
 b15zdnd11an1n32x5 FILLER_148_1316 ();
 b15zdnd11an1n04x5 FILLER_148_1348 ();
 b15zdnd11an1n04x5 FILLER_148_1355 ();
 b15zdnd00an1n01x5 FILLER_148_1359 ();
 b15zdnd11an1n64x5 FILLER_148_1363 ();
 b15zdnd00an1n02x5 FILLER_148_1427 ();
 b15zdnd00an1n01x5 FILLER_148_1429 ();
 b15zdnd11an1n64x5 FILLER_148_1482 ();
 b15zdnd11an1n64x5 FILLER_148_1546 ();
 b15zdnd11an1n64x5 FILLER_148_1610 ();
 b15zdnd11an1n64x5 FILLER_148_1674 ();
 b15zdnd11an1n64x5 FILLER_148_1738 ();
 b15zdnd11an1n16x5 FILLER_148_1802 ();
 b15zdnd00an1n02x5 FILLER_148_1818 ();
 b15zdnd11an1n64x5 FILLER_148_1827 ();
 b15zdnd11an1n64x5 FILLER_148_1891 ();
 b15zdnd11an1n64x5 FILLER_148_1955 ();
 b15zdnd11an1n04x5 FILLER_148_2019 ();
 b15zdnd11an1n04x5 FILLER_148_2026 ();
 b15zdnd00an1n01x5 FILLER_148_2030 ();
 b15zdnd11an1n64x5 FILLER_148_2073 ();
 b15zdnd11an1n08x5 FILLER_148_2137 ();
 b15zdnd00an1n02x5 FILLER_148_2151 ();
 b15zdnd00an1n01x5 FILLER_148_2153 ();
 b15zdnd11an1n32x5 FILLER_148_2162 ();
 b15zdnd11an1n16x5 FILLER_148_2194 ();
 b15zdnd11an1n04x5 FILLER_148_2217 ();
 b15zdnd00an1n01x5 FILLER_148_2221 ();
 b15zdnd11an1n04x5 FILLER_148_2225 ();
 b15zdnd00an1n02x5 FILLER_148_2274 ();
 b15zdnd11an1n64x5 FILLER_149_0 ();
 b15zdnd11an1n04x5 FILLER_149_64 ();
 b15zdnd00an1n01x5 FILLER_149_68 ();
 b15zdnd11an1n64x5 FILLER_149_108 ();
 b15zdnd11an1n64x5 FILLER_149_172 ();
 b15zdnd11an1n32x5 FILLER_149_236 ();
 b15zdnd11an1n08x5 FILLER_149_268 ();
 b15zdnd11an1n04x5 FILLER_149_276 ();
 b15zdnd11an1n64x5 FILLER_149_322 ();
 b15zdnd11an1n32x5 FILLER_149_386 ();
 b15zdnd11an1n16x5 FILLER_149_418 ();
 b15zdnd11an1n08x5 FILLER_149_434 ();
 b15zdnd00an1n02x5 FILLER_149_442 ();
 b15zdnd00an1n01x5 FILLER_149_444 ();
 b15zdnd11an1n32x5 FILLER_149_451 ();
 b15zdnd11an1n64x5 FILLER_149_535 ();
 b15zdnd11an1n64x5 FILLER_149_608 ();
 b15zdnd11an1n64x5 FILLER_149_672 ();
 b15zdnd11an1n08x5 FILLER_149_736 ();
 b15zdnd11an1n04x5 FILLER_149_744 ();
 b15zdnd00an1n02x5 FILLER_149_748 ();
 b15zdnd00an1n01x5 FILLER_149_750 ();
 b15zdnd11an1n32x5 FILLER_149_757 ();
 b15zdnd11an1n16x5 FILLER_149_789 ();
 b15zdnd11an1n04x5 FILLER_149_805 ();
 b15zdnd00an1n01x5 FILLER_149_809 ();
 b15zdnd11an1n32x5 FILLER_149_834 ();
 b15zdnd11an1n16x5 FILLER_149_866 ();
 b15zdnd11an1n04x5 FILLER_149_882 ();
 b15zdnd00an1n02x5 FILLER_149_886 ();
 b15zdnd00an1n01x5 FILLER_149_888 ();
 b15zdnd11an1n04x5 FILLER_149_909 ();
 b15zdnd11an1n64x5 FILLER_149_923 ();
 b15zdnd11an1n64x5 FILLER_149_987 ();
 b15zdnd11an1n64x5 FILLER_149_1051 ();
 b15zdnd00an1n02x5 FILLER_149_1115 ();
 b15zdnd11an1n64x5 FILLER_149_1120 ();
 b15zdnd11an1n64x5 FILLER_149_1184 ();
 b15zdnd11an1n64x5 FILLER_149_1248 ();
 b15zdnd11an1n16x5 FILLER_149_1312 ();
 b15zdnd00an1n01x5 FILLER_149_1328 ();
 b15zdnd11an1n04x5 FILLER_149_1381 ();
 b15zdnd11an1n32x5 FILLER_149_1392 ();
 b15zdnd11an1n08x5 FILLER_149_1424 ();
 b15zdnd11an1n04x5 FILLER_149_1432 ();
 b15zdnd11an1n32x5 FILLER_149_1488 ();
 b15zdnd11an1n04x5 FILLER_149_1520 ();
 b15zdnd11an1n64x5 FILLER_149_1566 ();
 b15zdnd11an1n64x5 FILLER_149_1630 ();
 b15zdnd11an1n08x5 FILLER_149_1694 ();
 b15zdnd00an1n02x5 FILLER_149_1702 ();
 b15zdnd11an1n64x5 FILLER_149_1735 ();
 b15zdnd11an1n16x5 FILLER_149_1799 ();
 b15zdnd11an1n08x5 FILLER_149_1815 ();
 b15zdnd11an1n04x5 FILLER_149_1823 ();
 b15zdnd00an1n01x5 FILLER_149_1827 ();
 b15zdnd11an1n64x5 FILLER_149_1831 ();
 b15zdnd11an1n32x5 FILLER_149_1895 ();
 b15zdnd11an1n16x5 FILLER_149_1927 ();
 b15zdnd11an1n04x5 FILLER_149_1943 ();
 b15zdnd11an1n32x5 FILLER_149_1966 ();
 b15zdnd11an1n16x5 FILLER_149_1998 ();
 b15zdnd11an1n08x5 FILLER_149_2014 ();
 b15zdnd11an1n04x5 FILLER_149_2022 ();
 b15zdnd00an1n01x5 FILLER_149_2026 ();
 b15zdnd11an1n04x5 FILLER_149_2037 ();
 b15zdnd11an1n64x5 FILLER_149_2083 ();
 b15zdnd11an1n16x5 FILLER_149_2147 ();
 b15zdnd11an1n04x5 FILLER_149_2163 ();
 b15zdnd11an1n16x5 FILLER_149_2180 ();
 b15zdnd11an1n08x5 FILLER_149_2196 ();
 b15zdnd11an1n04x5 FILLER_149_2204 ();
 b15zdnd11an1n08x5 FILLER_149_2260 ();
 b15zdnd00an1n01x5 FILLER_149_2268 ();
 b15zdnd11an1n04x5 FILLER_149_2273 ();
 b15zdnd00an1n01x5 FILLER_149_2277 ();
 b15zdnd00an1n02x5 FILLER_149_2282 ();
 b15zdnd11an1n64x5 FILLER_150_8 ();
 b15zdnd11an1n64x5 FILLER_150_72 ();
 b15zdnd11an1n64x5 FILLER_150_136 ();
 b15zdnd11an1n64x5 FILLER_150_200 ();
 b15zdnd11an1n64x5 FILLER_150_264 ();
 b15zdnd11an1n64x5 FILLER_150_328 ();
 b15zdnd11an1n64x5 FILLER_150_392 ();
 b15zdnd11an1n32x5 FILLER_150_456 ();
 b15zdnd11an1n16x5 FILLER_150_488 ();
 b15zdnd11an1n08x5 FILLER_150_504 ();
 b15zdnd11an1n04x5 FILLER_150_512 ();
 b15zdnd00an1n01x5 FILLER_150_516 ();
 b15zdnd11an1n08x5 FILLER_150_520 ();
 b15zdnd11an1n04x5 FILLER_150_528 ();
 b15zdnd11an1n04x5 FILLER_150_574 ();
 b15zdnd11an1n08x5 FILLER_150_581 ();
 b15zdnd00an1n01x5 FILLER_150_589 ();
 b15zdnd11an1n32x5 FILLER_150_617 ();
 b15zdnd11an1n08x5 FILLER_150_649 ();
 b15zdnd11an1n04x5 FILLER_150_657 ();
 b15zdnd00an1n02x5 FILLER_150_661 ();
 b15zdnd00an1n01x5 FILLER_150_663 ();
 b15zdnd11an1n32x5 FILLER_150_674 ();
 b15zdnd11an1n08x5 FILLER_150_706 ();
 b15zdnd11an1n04x5 FILLER_150_714 ();
 b15zdnd11an1n64x5 FILLER_150_726 ();
 b15zdnd11an1n16x5 FILLER_150_790 ();
 b15zdnd11an1n08x5 FILLER_150_806 ();
 b15zdnd00an1n02x5 FILLER_150_814 ();
 b15zdnd11an1n32x5 FILLER_150_837 ();
 b15zdnd11an1n08x5 FILLER_150_869 ();
 b15zdnd11an1n04x5 FILLER_150_877 ();
 b15zdnd00an1n01x5 FILLER_150_881 ();
 b15zdnd11an1n64x5 FILLER_150_902 ();
 b15zdnd11an1n64x5 FILLER_150_966 ();
 b15zdnd11an1n32x5 FILLER_150_1030 ();
 b15zdnd11an1n16x5 FILLER_150_1062 ();
 b15zdnd11an1n08x5 FILLER_150_1078 ();
 b15zdnd11an1n04x5 FILLER_150_1086 ();
 b15zdnd00an1n02x5 FILLER_150_1090 ();
 b15zdnd11an1n04x5 FILLER_150_1144 ();
 b15zdnd11an1n64x5 FILLER_150_1157 ();
 b15zdnd11an1n64x5 FILLER_150_1221 ();
 b15zdnd11an1n64x5 FILLER_150_1285 ();
 b15zdnd11an1n64x5 FILLER_150_1349 ();
 b15zdnd11an1n32x5 FILLER_150_1413 ();
 b15zdnd11an1n08x5 FILLER_150_1445 ();
 b15zdnd00an1n01x5 FILLER_150_1453 ();
 b15zdnd11an1n04x5 FILLER_150_1457 ();
 b15zdnd11an1n64x5 FILLER_150_1464 ();
 b15zdnd11an1n64x5 FILLER_150_1528 ();
 b15zdnd11an1n64x5 FILLER_150_1592 ();
 b15zdnd11an1n64x5 FILLER_150_1656 ();
 b15zdnd11an1n32x5 FILLER_150_1727 ();
 b15zdnd11an1n16x5 FILLER_150_1759 ();
 b15zdnd11an1n04x5 FILLER_150_1775 ();
 b15zdnd00an1n02x5 FILLER_150_1779 ();
 b15zdnd00an1n01x5 FILLER_150_1781 ();
 b15zdnd11an1n04x5 FILLER_150_1794 ();
 b15zdnd11an1n04x5 FILLER_150_1840 ();
 b15zdnd11an1n64x5 FILLER_150_1847 ();
 b15zdnd11an1n64x5 FILLER_150_1911 ();
 b15zdnd11an1n32x5 FILLER_150_1975 ();
 b15zdnd11an1n16x5 FILLER_150_2007 ();
 b15zdnd11an1n04x5 FILLER_150_2023 ();
 b15zdnd00an1n02x5 FILLER_150_2027 ();
 b15zdnd00an1n01x5 FILLER_150_2029 ();
 b15zdnd11an1n04x5 FILLER_150_2050 ();
 b15zdnd11an1n64x5 FILLER_150_2059 ();
 b15zdnd11an1n16x5 FILLER_150_2123 ();
 b15zdnd11an1n08x5 FILLER_150_2139 ();
 b15zdnd11an1n04x5 FILLER_150_2147 ();
 b15zdnd00an1n02x5 FILLER_150_2151 ();
 b15zdnd00an1n01x5 FILLER_150_2153 ();
 b15zdnd11an1n32x5 FILLER_150_2162 ();
 b15zdnd11an1n16x5 FILLER_150_2194 ();
 b15zdnd11an1n04x5 FILLER_150_2210 ();
 b15zdnd00an1n01x5 FILLER_150_2214 ();
 b15zdnd11an1n04x5 FILLER_150_2246 ();
 b15zdnd00an1n02x5 FILLER_150_2250 ();
 b15zdnd00an1n01x5 FILLER_150_2252 ();
 b15zdnd11an1n04x5 FILLER_150_2257 ();
 b15zdnd00an1n01x5 FILLER_150_2261 ();
 b15zdnd11an1n04x5 FILLER_150_2266 ();
 b15zdnd00an1n02x5 FILLER_150_2274 ();
 b15zdnd11an1n64x5 FILLER_151_0 ();
 b15zdnd11an1n64x5 FILLER_151_64 ();
 b15zdnd11an1n64x5 FILLER_151_128 ();
 b15zdnd11an1n64x5 FILLER_151_192 ();
 b15zdnd11an1n64x5 FILLER_151_256 ();
 b15zdnd11an1n64x5 FILLER_151_320 ();
 b15zdnd11an1n32x5 FILLER_151_384 ();
 b15zdnd11an1n64x5 FILLER_151_424 ();
 b15zdnd11an1n32x5 FILLER_151_488 ();
 b15zdnd11an1n08x5 FILLER_151_520 ();
 b15zdnd00an1n02x5 FILLER_151_528 ();
 b15zdnd11an1n64x5 FILLER_151_538 ();
 b15zdnd11an1n64x5 FILLER_151_602 ();
 b15zdnd11an1n64x5 FILLER_151_666 ();
 b15zdnd11an1n64x5 FILLER_151_730 ();
 b15zdnd11an1n16x5 FILLER_151_794 ();
 b15zdnd00an1n02x5 FILLER_151_810 ();
 b15zdnd00an1n01x5 FILLER_151_812 ();
 b15zdnd11an1n08x5 FILLER_151_824 ();
 b15zdnd11an1n04x5 FILLER_151_832 ();
 b15zdnd00an1n02x5 FILLER_151_836 ();
 b15zdnd00an1n01x5 FILLER_151_838 ();
 b15zdnd11an1n04x5 FILLER_151_842 ();
 b15zdnd00an1n01x5 FILLER_151_846 ();
 b15zdnd11an1n64x5 FILLER_151_863 ();
 b15zdnd11an1n64x5 FILLER_151_927 ();
 b15zdnd11an1n64x5 FILLER_151_994 ();
 b15zdnd11an1n16x5 FILLER_151_1058 ();
 b15zdnd11an1n08x5 FILLER_151_1074 ();
 b15zdnd00an1n02x5 FILLER_151_1082 ();
 b15zdnd00an1n01x5 FILLER_151_1084 ();
 b15zdnd11an1n64x5 FILLER_151_1137 ();
 b15zdnd11an1n64x5 FILLER_151_1201 ();
 b15zdnd11an1n64x5 FILLER_151_1265 ();
 b15zdnd11an1n64x5 FILLER_151_1329 ();
 b15zdnd11an1n64x5 FILLER_151_1393 ();
 b15zdnd11an1n64x5 FILLER_151_1457 ();
 b15zdnd11an1n64x5 FILLER_151_1521 ();
 b15zdnd11an1n64x5 FILLER_151_1585 ();
 b15zdnd11an1n64x5 FILLER_151_1649 ();
 b15zdnd11an1n64x5 FILLER_151_1713 ();
 b15zdnd11an1n32x5 FILLER_151_1777 ();
 b15zdnd00an1n01x5 FILLER_151_1809 ();
 b15zdnd11an1n64x5 FILLER_151_1862 ();
 b15zdnd11an1n64x5 FILLER_151_1926 ();
 b15zdnd11an1n32x5 FILLER_151_1990 ();
 b15zdnd11an1n16x5 FILLER_151_2022 ();
 b15zdnd00an1n02x5 FILLER_151_2038 ();
 b15zdnd11an1n04x5 FILLER_151_2047 ();
 b15zdnd11an1n64x5 FILLER_151_2057 ();
 b15zdnd11an1n32x5 FILLER_151_2121 ();
 b15zdnd11an1n16x5 FILLER_151_2153 ();
 b15zdnd00an1n01x5 FILLER_151_2169 ();
 b15zdnd11an1n08x5 FILLER_151_2215 ();
 b15zdnd11an1n08x5 FILLER_151_2230 ();
 b15zdnd00an1n02x5 FILLER_151_2238 ();
 b15zdnd00an1n02x5 FILLER_151_2282 ();
 b15zdnd11an1n64x5 FILLER_152_8 ();
 b15zdnd11an1n64x5 FILLER_152_72 ();
 b15zdnd11an1n64x5 FILLER_152_136 ();
 b15zdnd11an1n64x5 FILLER_152_200 ();
 b15zdnd11an1n64x5 FILLER_152_264 ();
 b15zdnd11an1n64x5 FILLER_152_328 ();
 b15zdnd11an1n64x5 FILLER_152_392 ();
 b15zdnd11an1n64x5 FILLER_152_456 ();
 b15zdnd11an1n64x5 FILLER_152_520 ();
 b15zdnd11an1n64x5 FILLER_152_584 ();
 b15zdnd11an1n64x5 FILLER_152_648 ();
 b15zdnd11an1n04x5 FILLER_152_712 ();
 b15zdnd00an1n02x5 FILLER_152_716 ();
 b15zdnd11an1n64x5 FILLER_152_726 ();
 b15zdnd11an1n64x5 FILLER_152_790 ();
 b15zdnd11an1n64x5 FILLER_152_854 ();
 b15zdnd11an1n32x5 FILLER_152_918 ();
 b15zdnd11an1n08x5 FILLER_152_950 ();
 b15zdnd11an1n04x5 FILLER_152_958 ();
 b15zdnd00an1n02x5 FILLER_152_962 ();
 b15zdnd11an1n64x5 FILLER_152_1016 ();
 b15zdnd11an1n16x5 FILLER_152_1080 ();
 b15zdnd11an1n08x5 FILLER_152_1096 ();
 b15zdnd00an1n01x5 FILLER_152_1104 ();
 b15zdnd11an1n04x5 FILLER_152_1108 ();
 b15zdnd11an1n04x5 FILLER_152_1115 ();
 b15zdnd11an1n04x5 FILLER_152_1122 ();
 b15zdnd11an1n16x5 FILLER_152_1129 ();
 b15zdnd11an1n04x5 FILLER_152_1145 ();
 b15zdnd00an1n02x5 FILLER_152_1149 ();
 b15zdnd00an1n01x5 FILLER_152_1151 ();
 b15zdnd11an1n32x5 FILLER_152_1159 ();
 b15zdnd11an1n16x5 FILLER_152_1191 ();
 b15zdnd00an1n02x5 FILLER_152_1207 ();
 b15zdnd00an1n01x5 FILLER_152_1209 ();
 b15zdnd11an1n64x5 FILLER_152_1230 ();
 b15zdnd00an1n02x5 FILLER_152_1294 ();
 b15zdnd00an1n01x5 FILLER_152_1296 ();
 b15zdnd11an1n64x5 FILLER_152_1306 ();
 b15zdnd11an1n64x5 FILLER_152_1370 ();
 b15zdnd11an1n64x5 FILLER_152_1434 ();
 b15zdnd11an1n16x5 FILLER_152_1498 ();
 b15zdnd11an1n08x5 FILLER_152_1514 ();
 b15zdnd00an1n01x5 FILLER_152_1522 ();
 b15zdnd11an1n32x5 FILLER_152_1532 ();
 b15zdnd11an1n08x5 FILLER_152_1564 ();
 b15zdnd00an1n02x5 FILLER_152_1572 ();
 b15zdnd11an1n64x5 FILLER_152_1591 ();
 b15zdnd11an1n16x5 FILLER_152_1655 ();
 b15zdnd11an1n04x5 FILLER_152_1671 ();
 b15zdnd00an1n02x5 FILLER_152_1675 ();
 b15zdnd11an1n64x5 FILLER_152_1687 ();
 b15zdnd11an1n16x5 FILLER_152_1751 ();
 b15zdnd11an1n08x5 FILLER_152_1772 ();
 b15zdnd11an1n04x5 FILLER_152_1780 ();
 b15zdnd00an1n02x5 FILLER_152_1784 ();
 b15zdnd11an1n08x5 FILLER_152_1793 ();
 b15zdnd11an1n04x5 FILLER_152_1801 ();
 b15zdnd00an1n01x5 FILLER_152_1805 ();
 b15zdnd11an1n16x5 FILLER_152_1810 ();
 b15zdnd11an1n08x5 FILLER_152_1826 ();
 b15zdnd00an1n01x5 FILLER_152_1834 ();
 b15zdnd11an1n32x5 FILLER_152_1838 ();
 b15zdnd11an1n64x5 FILLER_152_1912 ();
 b15zdnd11an1n64x5 FILLER_152_1976 ();
 b15zdnd11an1n64x5 FILLER_152_2040 ();
 b15zdnd11an1n32x5 FILLER_152_2104 ();
 b15zdnd11an1n16x5 FILLER_152_2136 ();
 b15zdnd00an1n02x5 FILLER_152_2152 ();
 b15zdnd11an1n16x5 FILLER_152_2162 ();
 b15zdnd11an1n04x5 FILLER_152_2178 ();
 b15zdnd00an1n02x5 FILLER_152_2182 ();
 b15zdnd00an1n01x5 FILLER_152_2184 ();
 b15zdnd11an1n04x5 FILLER_152_2199 ();
 b15zdnd11an1n08x5 FILLER_152_2234 ();
 b15zdnd11an1n04x5 FILLER_152_2242 ();
 b15zdnd11an1n08x5 FILLER_152_2249 ();
 b15zdnd11an1n04x5 FILLER_152_2257 ();
 b15zdnd00an1n02x5 FILLER_152_2261 ();
 b15zdnd00an1n01x5 FILLER_152_2263 ();
 b15zdnd11an1n08x5 FILLER_152_2268 ();
 b15zdnd11an1n64x5 FILLER_153_0 ();
 b15zdnd11an1n64x5 FILLER_153_64 ();
 b15zdnd11an1n64x5 FILLER_153_128 ();
 b15zdnd11an1n64x5 FILLER_153_192 ();
 b15zdnd11an1n64x5 FILLER_153_256 ();
 b15zdnd11an1n64x5 FILLER_153_320 ();
 b15zdnd11an1n64x5 FILLER_153_384 ();
 b15zdnd11an1n64x5 FILLER_153_448 ();
 b15zdnd11an1n64x5 FILLER_153_512 ();
 b15zdnd11an1n64x5 FILLER_153_576 ();
 b15zdnd11an1n32x5 FILLER_153_640 ();
 b15zdnd11an1n16x5 FILLER_153_672 ();
 b15zdnd00an1n02x5 FILLER_153_688 ();
 b15zdnd11an1n64x5 FILLER_153_693 ();
 b15zdnd11an1n64x5 FILLER_153_757 ();
 b15zdnd11an1n64x5 FILLER_153_821 ();
 b15zdnd11an1n64x5 FILLER_153_885 ();
 b15zdnd11an1n32x5 FILLER_153_949 ();
 b15zdnd00an1n02x5 FILLER_153_981 ();
 b15zdnd11an1n04x5 FILLER_153_986 ();
 b15zdnd11an1n64x5 FILLER_153_993 ();
 b15zdnd11an1n32x5 FILLER_153_1057 ();
 b15zdnd11an1n16x5 FILLER_153_1089 ();
 b15zdnd11an1n04x5 FILLER_153_1105 ();
 b15zdnd00an1n02x5 FILLER_153_1109 ();
 b15zdnd11an1n64x5 FILLER_153_1114 ();
 b15zdnd11an1n64x5 FILLER_153_1178 ();
 b15zdnd11an1n64x5 FILLER_153_1242 ();
 b15zdnd11an1n64x5 FILLER_153_1306 ();
 b15zdnd11an1n64x5 FILLER_153_1370 ();
 b15zdnd11an1n64x5 FILLER_153_1434 ();
 b15zdnd11an1n32x5 FILLER_153_1498 ();
 b15zdnd11an1n16x5 FILLER_153_1530 ();
 b15zdnd11an1n04x5 FILLER_153_1546 ();
 b15zdnd00an1n02x5 FILLER_153_1550 ();
 b15zdnd11an1n08x5 FILLER_153_1558 ();
 b15zdnd11an1n04x5 FILLER_153_1566 ();
 b15zdnd11an1n32x5 FILLER_153_1587 ();
 b15zdnd11an1n04x5 FILLER_153_1619 ();
 b15zdnd00an1n01x5 FILLER_153_1623 ();
 b15zdnd11an1n08x5 FILLER_153_1645 ();
 b15zdnd11an1n04x5 FILLER_153_1653 ();
 b15zdnd00an1n02x5 FILLER_153_1657 ();
 b15zdnd00an1n01x5 FILLER_153_1659 ();
 b15zdnd11an1n08x5 FILLER_153_1663 ();
 b15zdnd00an1n02x5 FILLER_153_1671 ();
 b15zdnd00an1n01x5 FILLER_153_1673 ();
 b15zdnd11an1n04x5 FILLER_153_1677 ();
 b15zdnd11an1n32x5 FILLER_153_1684 ();
 b15zdnd11an1n08x5 FILLER_153_1716 ();
 b15zdnd00an1n01x5 FILLER_153_1724 ();
 b15zdnd11an1n32x5 FILLER_153_1749 ();
 b15zdnd11an1n04x5 FILLER_153_1781 ();
 b15zdnd00an1n02x5 FILLER_153_1785 ();
 b15zdnd11an1n32x5 FILLER_153_1829 ();
 b15zdnd11an1n04x5 FILLER_153_1861 ();
 b15zdnd00an1n02x5 FILLER_153_1865 ();
 b15zdnd11an1n64x5 FILLER_153_1870 ();
 b15zdnd11an1n64x5 FILLER_153_1934 ();
 b15zdnd11an1n64x5 FILLER_153_1998 ();
 b15zdnd11an1n32x5 FILLER_153_2062 ();
 b15zdnd11an1n16x5 FILLER_153_2094 ();
 b15zdnd00an1n02x5 FILLER_153_2110 ();
 b15zdnd00an1n01x5 FILLER_153_2112 ();
 b15zdnd11an1n64x5 FILLER_153_2125 ();
 b15zdnd11an1n04x5 FILLER_153_2189 ();
 b15zdnd00an1n02x5 FILLER_153_2193 ();
 b15zdnd11an1n32x5 FILLER_153_2237 ();
 b15zdnd11an1n08x5 FILLER_153_2269 ();
 b15zdnd11an1n04x5 FILLER_153_2277 ();
 b15zdnd00an1n02x5 FILLER_153_2281 ();
 b15zdnd00an1n01x5 FILLER_153_2283 ();
 b15zdnd11an1n64x5 FILLER_154_8 ();
 b15zdnd11an1n64x5 FILLER_154_72 ();
 b15zdnd11an1n64x5 FILLER_154_136 ();
 b15zdnd11an1n64x5 FILLER_154_200 ();
 b15zdnd11an1n64x5 FILLER_154_264 ();
 b15zdnd11an1n64x5 FILLER_154_328 ();
 b15zdnd11an1n32x5 FILLER_154_392 ();
 b15zdnd11an1n08x5 FILLER_154_424 ();
 b15zdnd11an1n04x5 FILLER_154_432 ();
 b15zdnd00an1n02x5 FILLER_154_436 ();
 b15zdnd11an1n16x5 FILLER_154_450 ();
 b15zdnd11an1n08x5 FILLER_154_466 ();
 b15zdnd00an1n01x5 FILLER_154_474 ();
 b15zdnd11an1n64x5 FILLER_154_489 ();
 b15zdnd11an1n32x5 FILLER_154_553 ();
 b15zdnd11an1n16x5 FILLER_154_585 ();
 b15zdnd11an1n04x5 FILLER_154_601 ();
 b15zdnd00an1n01x5 FILLER_154_605 ();
 b15zdnd11an1n32x5 FILLER_154_624 ();
 b15zdnd11an1n08x5 FILLER_154_656 ();
 b15zdnd00an1n02x5 FILLER_154_716 ();
 b15zdnd11an1n32x5 FILLER_154_726 ();
 b15zdnd11an1n08x5 FILLER_154_758 ();
 b15zdnd00an1n01x5 FILLER_154_766 ();
 b15zdnd11an1n64x5 FILLER_154_771 ();
 b15zdnd11an1n32x5 FILLER_154_835 ();
 b15zdnd11an1n16x5 FILLER_154_867 ();
 b15zdnd11an1n08x5 FILLER_154_883 ();
 b15zdnd00an1n02x5 FILLER_154_891 ();
 b15zdnd00an1n01x5 FILLER_154_893 ();
 b15zdnd11an1n64x5 FILLER_154_908 ();
 b15zdnd11an1n64x5 FILLER_154_972 ();
 b15zdnd11an1n64x5 FILLER_154_1036 ();
 b15zdnd11an1n64x5 FILLER_154_1100 ();
 b15zdnd11an1n64x5 FILLER_154_1164 ();
 b15zdnd11an1n64x5 FILLER_154_1228 ();
 b15zdnd11an1n64x5 FILLER_154_1292 ();
 b15zdnd11an1n32x5 FILLER_154_1356 ();
 b15zdnd11an1n16x5 FILLER_154_1388 ();
 b15zdnd00an1n01x5 FILLER_154_1404 ();
 b15zdnd11an1n64x5 FILLER_154_1414 ();
 b15zdnd11an1n64x5 FILLER_154_1478 ();
 b15zdnd11an1n16x5 FILLER_154_1542 ();
 b15zdnd11an1n08x5 FILLER_154_1558 ();
 b15zdnd11an1n04x5 FILLER_154_1566 ();
 b15zdnd11an1n04x5 FILLER_154_1583 ();
 b15zdnd11an1n04x5 FILLER_154_1605 ();
 b15zdnd11an1n16x5 FILLER_154_1620 ();
 b15zdnd00an1n01x5 FILLER_154_1636 ();
 b15zdnd11an1n04x5 FILLER_154_1647 ();
 b15zdnd11an1n04x5 FILLER_154_1654 ();
 b15zdnd11an1n04x5 FILLER_154_1702 ();
 b15zdnd11an1n64x5 FILLER_154_1713 ();
 b15zdnd11an1n16x5 FILLER_154_1777 ();
 b15zdnd00an1n01x5 FILLER_154_1793 ();
 b15zdnd11an1n64x5 FILLER_154_1809 ();
 b15zdnd11an1n64x5 FILLER_154_1873 ();
 b15zdnd11an1n64x5 FILLER_154_1937 ();
 b15zdnd11an1n64x5 FILLER_154_2001 ();
 b15zdnd11an1n64x5 FILLER_154_2065 ();
 b15zdnd11an1n16x5 FILLER_154_2129 ();
 b15zdnd11an1n08x5 FILLER_154_2145 ();
 b15zdnd00an1n01x5 FILLER_154_2153 ();
 b15zdnd11an1n16x5 FILLER_154_2162 ();
 b15zdnd11an1n08x5 FILLER_154_2178 ();
 b15zdnd00an1n02x5 FILLER_154_2186 ();
 b15zdnd00an1n01x5 FILLER_154_2188 ();
 b15zdnd11an1n32x5 FILLER_154_2192 ();
 b15zdnd11an1n08x5 FILLER_154_2224 ();
 b15zdnd00an1n02x5 FILLER_154_2274 ();
 b15zdnd11an1n64x5 FILLER_155_0 ();
 b15zdnd11an1n64x5 FILLER_155_64 ();
 b15zdnd11an1n64x5 FILLER_155_128 ();
 b15zdnd11an1n64x5 FILLER_155_192 ();
 b15zdnd11an1n64x5 FILLER_155_256 ();
 b15zdnd11an1n64x5 FILLER_155_320 ();
 b15zdnd00an1n02x5 FILLER_155_384 ();
 b15zdnd00an1n01x5 FILLER_155_386 ();
 b15zdnd11an1n32x5 FILLER_155_429 ();
 b15zdnd11an1n16x5 FILLER_155_461 ();
 b15zdnd00an1n02x5 FILLER_155_477 ();
 b15zdnd11an1n64x5 FILLER_155_521 ();
 b15zdnd11an1n64x5 FILLER_155_585 ();
 b15zdnd11an1n32x5 FILLER_155_649 ();
 b15zdnd00an1n01x5 FILLER_155_681 ();
 b15zdnd11an1n04x5 FILLER_155_685 ();
 b15zdnd11an1n08x5 FILLER_155_692 ();
 b15zdnd11an1n64x5 FILLER_155_708 ();
 b15zdnd11an1n64x5 FILLER_155_772 ();
 b15zdnd11an1n64x5 FILLER_155_836 ();
 b15zdnd11an1n64x5 FILLER_155_900 ();
 b15zdnd11an1n16x5 FILLER_155_964 ();
 b15zdnd00an1n02x5 FILLER_155_980 ();
 b15zdnd00an1n01x5 FILLER_155_982 ();
 b15zdnd11an1n64x5 FILLER_155_987 ();
 b15zdnd11an1n64x5 FILLER_155_1051 ();
 b15zdnd11an1n64x5 FILLER_155_1115 ();
 b15zdnd11an1n64x5 FILLER_155_1179 ();
 b15zdnd11an1n64x5 FILLER_155_1243 ();
 b15zdnd11an1n64x5 FILLER_155_1307 ();
 b15zdnd11an1n64x5 FILLER_155_1371 ();
 b15zdnd11an1n64x5 FILLER_155_1435 ();
 b15zdnd11an1n32x5 FILLER_155_1499 ();
 b15zdnd11an1n16x5 FILLER_155_1531 ();
 b15zdnd11an1n08x5 FILLER_155_1547 ();
 b15zdnd00an1n02x5 FILLER_155_1555 ();
 b15zdnd00an1n01x5 FILLER_155_1557 ();
 b15zdnd11an1n04x5 FILLER_155_1564 ();
 b15zdnd11an1n04x5 FILLER_155_1571 ();
 b15zdnd11an1n16x5 FILLER_155_1578 ();
 b15zdnd11an1n08x5 FILLER_155_1594 ();
 b15zdnd11an1n32x5 FILLER_155_1616 ();
 b15zdnd11an1n08x5 FILLER_155_1662 ();
 b15zdnd11an1n64x5 FILLER_155_1712 ();
 b15zdnd00an1n02x5 FILLER_155_1776 ();
 b15zdnd00an1n01x5 FILLER_155_1778 ();
 b15zdnd11an1n64x5 FILLER_155_1793 ();
 b15zdnd11an1n64x5 FILLER_155_1857 ();
 b15zdnd11an1n16x5 FILLER_155_1921 ();
 b15zdnd11an1n04x5 FILLER_155_1937 ();
 b15zdnd00an1n02x5 FILLER_155_1941 ();
 b15zdnd00an1n01x5 FILLER_155_1943 ();
 b15zdnd11an1n64x5 FILLER_155_1964 ();
 b15zdnd11an1n64x5 FILLER_155_2028 ();
 b15zdnd11an1n64x5 FILLER_155_2092 ();
 b15zdnd11an1n08x5 FILLER_155_2156 ();
 b15zdnd11an1n04x5 FILLER_155_2216 ();
 b15zdnd11an1n32x5 FILLER_155_2244 ();
 b15zdnd11an1n08x5 FILLER_155_2276 ();
 b15zdnd11an1n64x5 FILLER_156_8 ();
 b15zdnd11an1n64x5 FILLER_156_72 ();
 b15zdnd11an1n64x5 FILLER_156_136 ();
 b15zdnd11an1n64x5 FILLER_156_200 ();
 b15zdnd11an1n64x5 FILLER_156_264 ();
 b15zdnd11an1n64x5 FILLER_156_328 ();
 b15zdnd11an1n16x5 FILLER_156_392 ();
 b15zdnd11an1n04x5 FILLER_156_408 ();
 b15zdnd11an1n32x5 FILLER_156_417 ();
 b15zdnd11an1n08x5 FILLER_156_449 ();
 b15zdnd00an1n02x5 FILLER_156_457 ();
 b15zdnd00an1n01x5 FILLER_156_459 ();
 b15zdnd11an1n04x5 FILLER_156_466 ();
 b15zdnd11an1n04x5 FILLER_156_476 ();
 b15zdnd00an1n01x5 FILLER_156_480 ();
 b15zdnd11an1n64x5 FILLER_156_501 ();
 b15zdnd11an1n64x5 FILLER_156_565 ();
 b15zdnd11an1n32x5 FILLER_156_629 ();
 b15zdnd11an1n08x5 FILLER_156_661 ();
 b15zdnd11an1n04x5 FILLER_156_669 ();
 b15zdnd11an1n04x5 FILLER_156_676 ();
 b15zdnd00an1n02x5 FILLER_156_680 ();
 b15zdnd11an1n04x5 FILLER_156_685 ();
 b15zdnd11an1n16x5 FILLER_156_692 ();
 b15zdnd11an1n08x5 FILLER_156_708 ();
 b15zdnd00an1n02x5 FILLER_156_716 ();
 b15zdnd11an1n32x5 FILLER_156_726 ();
 b15zdnd11an1n16x5 FILLER_156_758 ();
 b15zdnd11an1n04x5 FILLER_156_774 ();
 b15zdnd00an1n02x5 FILLER_156_778 ();
 b15zdnd11an1n64x5 FILLER_156_788 ();
 b15zdnd11an1n64x5 FILLER_156_852 ();
 b15zdnd11an1n64x5 FILLER_156_916 ();
 b15zdnd00an1n02x5 FILLER_156_980 ();
 b15zdnd11an1n08x5 FILLER_156_986 ();
 b15zdnd00an1n02x5 FILLER_156_994 ();
 b15zdnd11an1n64x5 FILLER_156_1004 ();
 b15zdnd11an1n64x5 FILLER_156_1068 ();
 b15zdnd11an1n64x5 FILLER_156_1132 ();
 b15zdnd11an1n64x5 FILLER_156_1196 ();
 b15zdnd11an1n64x5 FILLER_156_1260 ();
 b15zdnd11an1n64x5 FILLER_156_1324 ();
 b15zdnd11an1n64x5 FILLER_156_1388 ();
 b15zdnd11an1n64x5 FILLER_156_1452 ();
 b15zdnd11an1n32x5 FILLER_156_1516 ();
 b15zdnd11an1n16x5 FILLER_156_1548 ();
 b15zdnd11an1n04x5 FILLER_156_1564 ();
 b15zdnd11an1n32x5 FILLER_156_1578 ();
 b15zdnd11an1n04x5 FILLER_156_1610 ();
 b15zdnd11an1n08x5 FILLER_156_1656 ();
 b15zdnd00an1n02x5 FILLER_156_1664 ();
 b15zdnd11an1n04x5 FILLER_156_1673 ();
 b15zdnd11an1n64x5 FILLER_156_1680 ();
 b15zdnd11an1n64x5 FILLER_156_1744 ();
 b15zdnd11an1n64x5 FILLER_156_1808 ();
 b15zdnd11an1n64x5 FILLER_156_1872 ();
 b15zdnd11an1n64x5 FILLER_156_1936 ();
 b15zdnd11an1n32x5 FILLER_156_2000 ();
 b15zdnd11an1n16x5 FILLER_156_2032 ();
 b15zdnd11an1n64x5 FILLER_156_2051 ();
 b15zdnd11an1n32x5 FILLER_156_2115 ();
 b15zdnd11an1n04x5 FILLER_156_2147 ();
 b15zdnd00an1n02x5 FILLER_156_2151 ();
 b15zdnd00an1n01x5 FILLER_156_2153 ();
 b15zdnd11an1n16x5 FILLER_156_2162 ();
 b15zdnd00an1n02x5 FILLER_156_2178 ();
 b15zdnd00an1n01x5 FILLER_156_2180 ();
 b15zdnd11an1n04x5 FILLER_156_2233 ();
 b15zdnd11an1n32x5 FILLER_156_2244 ();
 b15zdnd11an1n64x5 FILLER_157_0 ();
 b15zdnd11an1n64x5 FILLER_157_64 ();
 b15zdnd11an1n64x5 FILLER_157_128 ();
 b15zdnd11an1n64x5 FILLER_157_192 ();
 b15zdnd11an1n64x5 FILLER_157_256 ();
 b15zdnd11an1n64x5 FILLER_157_320 ();
 b15zdnd11an1n16x5 FILLER_157_384 ();
 b15zdnd00an1n02x5 FILLER_157_400 ();
 b15zdnd00an1n01x5 FILLER_157_402 ();
 b15zdnd11an1n64x5 FILLER_157_410 ();
 b15zdnd11an1n64x5 FILLER_157_474 ();
 b15zdnd11an1n64x5 FILLER_157_538 ();
 b15zdnd11an1n32x5 FILLER_157_602 ();
 b15zdnd11an1n16x5 FILLER_157_634 ();
 b15zdnd11an1n08x5 FILLER_157_650 ();
 b15zdnd11an1n04x5 FILLER_157_658 ();
 b15zdnd00an1n02x5 FILLER_157_662 ();
 b15zdnd00an1n01x5 FILLER_157_664 ();
 b15zdnd11an1n32x5 FILLER_157_717 ();
 b15zdnd11an1n16x5 FILLER_157_749 ();
 b15zdnd11an1n08x5 FILLER_157_765 ();
 b15zdnd00an1n02x5 FILLER_157_773 ();
 b15zdnd00an1n01x5 FILLER_157_775 ();
 b15zdnd11an1n64x5 FILLER_157_784 ();
 b15zdnd11an1n16x5 FILLER_157_848 ();
 b15zdnd11an1n04x5 FILLER_157_864 ();
 b15zdnd00an1n02x5 FILLER_157_868 ();
 b15zdnd00an1n01x5 FILLER_157_870 ();
 b15zdnd11an1n64x5 FILLER_157_885 ();
 b15zdnd11an1n64x5 FILLER_157_949 ();
 b15zdnd11an1n64x5 FILLER_157_1013 ();
 b15zdnd11an1n64x5 FILLER_157_1077 ();
 b15zdnd11an1n64x5 FILLER_157_1141 ();
 b15zdnd11an1n64x5 FILLER_157_1205 ();
 b15zdnd11an1n64x5 FILLER_157_1269 ();
 b15zdnd11an1n64x5 FILLER_157_1333 ();
 b15zdnd11an1n64x5 FILLER_157_1397 ();
 b15zdnd11an1n64x5 FILLER_157_1461 ();
 b15zdnd11an1n64x5 FILLER_157_1525 ();
 b15zdnd11an1n64x5 FILLER_157_1589 ();
 b15zdnd11an1n64x5 FILLER_157_1653 ();
 b15zdnd11an1n64x5 FILLER_157_1717 ();
 b15zdnd11an1n64x5 FILLER_157_1781 ();
 b15zdnd11an1n64x5 FILLER_157_1845 ();
 b15zdnd11an1n64x5 FILLER_157_1909 ();
 b15zdnd11an1n64x5 FILLER_157_1973 ();
 b15zdnd11an1n08x5 FILLER_157_2037 ();
 b15zdnd11an1n64x5 FILLER_157_2051 ();
 b15zdnd11an1n64x5 FILLER_157_2115 ();
 b15zdnd00an1n02x5 FILLER_157_2179 ();
 b15zdnd11an1n08x5 FILLER_157_2184 ();
 b15zdnd00an1n01x5 FILLER_157_2192 ();
 b15zdnd11an1n08x5 FILLER_157_2196 ();
 b15zdnd11an1n04x5 FILLER_157_2207 ();
 b15zdnd11an1n16x5 FILLER_157_2218 ();
 b15zdnd11an1n08x5 FILLER_157_2234 ();
 b15zdnd00an1n02x5 FILLER_157_2242 ();
 b15zdnd11an1n32x5 FILLER_157_2248 ();
 b15zdnd11an1n04x5 FILLER_157_2280 ();
 b15zdnd11an1n64x5 FILLER_158_8 ();
 b15zdnd11an1n64x5 FILLER_158_72 ();
 b15zdnd11an1n64x5 FILLER_158_136 ();
 b15zdnd11an1n64x5 FILLER_158_200 ();
 b15zdnd11an1n08x5 FILLER_158_264 ();
 b15zdnd11an1n04x5 FILLER_158_272 ();
 b15zdnd00an1n02x5 FILLER_158_276 ();
 b15zdnd00an1n01x5 FILLER_158_278 ();
 b15zdnd11an1n04x5 FILLER_158_282 ();
 b15zdnd11an1n64x5 FILLER_158_289 ();
 b15zdnd11an1n64x5 FILLER_158_353 ();
 b15zdnd11an1n64x5 FILLER_158_417 ();
 b15zdnd11an1n64x5 FILLER_158_481 ();
 b15zdnd11an1n08x5 FILLER_158_545 ();
 b15zdnd00an1n02x5 FILLER_158_553 ();
 b15zdnd00an1n01x5 FILLER_158_555 ();
 b15zdnd11an1n64x5 FILLER_158_559 ();
 b15zdnd11an1n64x5 FILLER_158_623 ();
 b15zdnd11an1n08x5 FILLER_158_687 ();
 b15zdnd00an1n02x5 FILLER_158_715 ();
 b15zdnd00an1n01x5 FILLER_158_717 ();
 b15zdnd11an1n64x5 FILLER_158_726 ();
 b15zdnd11an1n64x5 FILLER_158_790 ();
 b15zdnd11an1n16x5 FILLER_158_854 ();
 b15zdnd11an1n08x5 FILLER_158_870 ();
 b15zdnd00an1n02x5 FILLER_158_878 ();
 b15zdnd00an1n01x5 FILLER_158_880 ();
 b15zdnd11an1n16x5 FILLER_158_887 ();
 b15zdnd11an1n08x5 FILLER_158_903 ();
 b15zdnd11an1n04x5 FILLER_158_911 ();
 b15zdnd00an1n01x5 FILLER_158_915 ();
 b15zdnd11an1n64x5 FILLER_158_937 ();
 b15zdnd11an1n64x5 FILLER_158_1001 ();
 b15zdnd11an1n64x5 FILLER_158_1065 ();
 b15zdnd11an1n32x5 FILLER_158_1129 ();
 b15zdnd11an1n08x5 FILLER_158_1161 ();
 b15zdnd11an1n04x5 FILLER_158_1169 ();
 b15zdnd00an1n01x5 FILLER_158_1173 ();
 b15zdnd11an1n64x5 FILLER_158_1193 ();
 b15zdnd11an1n64x5 FILLER_158_1257 ();
 b15zdnd11an1n64x5 FILLER_158_1321 ();
 b15zdnd11an1n64x5 FILLER_158_1385 ();
 b15zdnd11an1n64x5 FILLER_158_1449 ();
 b15zdnd11an1n64x5 FILLER_158_1513 ();
 b15zdnd11an1n32x5 FILLER_158_1577 ();
 b15zdnd11an1n08x5 FILLER_158_1609 ();
 b15zdnd11an1n04x5 FILLER_158_1617 ();
 b15zdnd11an1n04x5 FILLER_158_1635 ();
 b15zdnd11an1n16x5 FILLER_158_1653 ();
 b15zdnd11an1n08x5 FILLER_158_1669 ();
 b15zdnd00an1n02x5 FILLER_158_1677 ();
 b15zdnd00an1n01x5 FILLER_158_1679 ();
 b15zdnd11an1n08x5 FILLER_158_1711 ();
 b15zdnd00an1n01x5 FILLER_158_1719 ();
 b15zdnd11an1n64x5 FILLER_158_1739 ();
 b15zdnd11an1n64x5 FILLER_158_1803 ();
 b15zdnd11an1n64x5 FILLER_158_1867 ();
 b15zdnd11an1n64x5 FILLER_158_1931 ();
 b15zdnd11an1n64x5 FILLER_158_1995 ();
 b15zdnd11an1n64x5 FILLER_158_2059 ();
 b15zdnd11an1n16x5 FILLER_158_2123 ();
 b15zdnd11an1n08x5 FILLER_158_2139 ();
 b15zdnd11an1n04x5 FILLER_158_2147 ();
 b15zdnd00an1n02x5 FILLER_158_2151 ();
 b15zdnd00an1n01x5 FILLER_158_2153 ();
 b15zdnd11an1n16x5 FILLER_158_2162 ();
 b15zdnd11an1n08x5 FILLER_158_2178 ();
 b15zdnd11an1n04x5 FILLER_158_2186 ();
 b15zdnd00an1n02x5 FILLER_158_2190 ();
 b15zdnd11an1n08x5 FILLER_158_2195 ();
 b15zdnd00an1n01x5 FILLER_158_2203 ();
 b15zdnd11an1n64x5 FILLER_158_2207 ();
 b15zdnd11an1n04x5 FILLER_158_2271 ();
 b15zdnd00an1n01x5 FILLER_158_2275 ();
 b15zdnd11an1n64x5 FILLER_159_0 ();
 b15zdnd11an1n64x5 FILLER_159_64 ();
 b15zdnd11an1n64x5 FILLER_159_128 ();
 b15zdnd11an1n32x5 FILLER_159_192 ();
 b15zdnd11an1n16x5 FILLER_159_224 ();
 b15zdnd11an1n08x5 FILLER_159_240 ();
 b15zdnd11an1n04x5 FILLER_159_248 ();
 b15zdnd00an1n02x5 FILLER_159_252 ();
 b15zdnd11an1n64x5 FILLER_159_306 ();
 b15zdnd11an1n64x5 FILLER_159_370 ();
 b15zdnd11an1n64x5 FILLER_159_434 ();
 b15zdnd11an1n32x5 FILLER_159_498 ();
 b15zdnd00an1n01x5 FILLER_159_530 ();
 b15zdnd11an1n64x5 FILLER_159_583 ();
 b15zdnd11an1n64x5 FILLER_159_647 ();
 b15zdnd11an1n32x5 FILLER_159_711 ();
 b15zdnd11an1n16x5 FILLER_159_743 ();
 b15zdnd00an1n02x5 FILLER_159_759 ();
 b15zdnd11an1n64x5 FILLER_159_765 ();
 b15zdnd11an1n32x5 FILLER_159_829 ();
 b15zdnd11an1n08x5 FILLER_159_861 ();
 b15zdnd11an1n04x5 FILLER_159_869 ();
 b15zdnd00an1n02x5 FILLER_159_873 ();
 b15zdnd00an1n01x5 FILLER_159_875 ();
 b15zdnd11an1n04x5 FILLER_159_892 ();
 b15zdnd11an1n64x5 FILLER_159_903 ();
 b15zdnd11an1n64x5 FILLER_159_967 ();
 b15zdnd11an1n64x5 FILLER_159_1031 ();
 b15zdnd11an1n64x5 FILLER_159_1095 ();
 b15zdnd11an1n32x5 FILLER_159_1159 ();
 b15zdnd11an1n16x5 FILLER_159_1191 ();
 b15zdnd11an1n08x5 FILLER_159_1207 ();
 b15zdnd11an1n04x5 FILLER_159_1215 ();
 b15zdnd00an1n01x5 FILLER_159_1219 ();
 b15zdnd11an1n64x5 FILLER_159_1234 ();
 b15zdnd11an1n64x5 FILLER_159_1298 ();
 b15zdnd11an1n64x5 FILLER_159_1362 ();
 b15zdnd11an1n64x5 FILLER_159_1426 ();
 b15zdnd11an1n64x5 FILLER_159_1490 ();
 b15zdnd11an1n64x5 FILLER_159_1554 ();
 b15zdnd11an1n64x5 FILLER_159_1618 ();
 b15zdnd11an1n64x5 FILLER_159_1682 ();
 b15zdnd11an1n64x5 FILLER_159_1746 ();
 b15zdnd11an1n64x5 FILLER_159_1810 ();
 b15zdnd11an1n64x5 FILLER_159_1874 ();
 b15zdnd11an1n64x5 FILLER_159_1938 ();
 b15zdnd11an1n32x5 FILLER_159_2002 ();
 b15zdnd11an1n08x5 FILLER_159_2034 ();
 b15zdnd11an1n04x5 FILLER_159_2042 ();
 b15zdnd00an1n01x5 FILLER_159_2046 ();
 b15zdnd11an1n64x5 FILLER_159_2053 ();
 b15zdnd11an1n64x5 FILLER_159_2117 ();
 b15zdnd11an1n32x5 FILLER_159_2181 ();
 b15zdnd11an1n16x5 FILLER_159_2213 ();
 b15zdnd11an1n04x5 FILLER_159_2229 ();
 b15zdnd00an1n02x5 FILLER_159_2233 ();
 b15zdnd00an1n01x5 FILLER_159_2235 ();
 b15zdnd11an1n04x5 FILLER_159_2278 ();
 b15zdnd00an1n02x5 FILLER_159_2282 ();
 b15zdnd11an1n64x5 FILLER_160_8 ();
 b15zdnd11an1n64x5 FILLER_160_72 ();
 b15zdnd11an1n32x5 FILLER_160_136 ();
 b15zdnd11an1n16x5 FILLER_160_168 ();
 b15zdnd00an1n02x5 FILLER_160_184 ();
 b15zdnd11an1n04x5 FILLER_160_190 ();
 b15zdnd11an1n32x5 FILLER_160_200 ();
 b15zdnd11an1n04x5 FILLER_160_232 ();
 b15zdnd00an1n02x5 FILLER_160_236 ();
 b15zdnd11an1n32x5 FILLER_160_242 ();
 b15zdnd00an1n02x5 FILLER_160_274 ();
 b15zdnd00an1n01x5 FILLER_160_276 ();
 b15zdnd11an1n64x5 FILLER_160_280 ();
 b15zdnd11an1n64x5 FILLER_160_344 ();
 b15zdnd11an1n32x5 FILLER_160_408 ();
 b15zdnd11an1n04x5 FILLER_160_440 ();
 b15zdnd11an1n64x5 FILLER_160_450 ();
 b15zdnd11an1n16x5 FILLER_160_514 ();
 b15zdnd11an1n08x5 FILLER_160_530 ();
 b15zdnd11an1n04x5 FILLER_160_538 ();
 b15zdnd00an1n02x5 FILLER_160_542 ();
 b15zdnd11an1n64x5 FILLER_160_596 ();
 b15zdnd11an1n08x5 FILLER_160_660 ();
 b15zdnd11an1n04x5 FILLER_160_668 ();
 b15zdnd00an1n02x5 FILLER_160_672 ();
 b15zdnd00an1n02x5 FILLER_160_716 ();
 b15zdnd11an1n64x5 FILLER_160_726 ();
 b15zdnd11an1n64x5 FILLER_160_790 ();
 b15zdnd11an1n64x5 FILLER_160_854 ();
 b15zdnd11an1n04x5 FILLER_160_918 ();
 b15zdnd00an1n01x5 FILLER_160_922 ();
 b15zdnd11an1n16x5 FILLER_160_937 ();
 b15zdnd11an1n04x5 FILLER_160_953 ();
 b15zdnd00an1n02x5 FILLER_160_957 ();
 b15zdnd11an1n64x5 FILLER_160_982 ();
 b15zdnd11an1n64x5 FILLER_160_1046 ();
 b15zdnd11an1n64x5 FILLER_160_1110 ();
 b15zdnd11an1n32x5 FILLER_160_1174 ();
 b15zdnd11an1n08x5 FILLER_160_1206 ();
 b15zdnd00an1n02x5 FILLER_160_1214 ();
 b15zdnd00an1n01x5 FILLER_160_1216 ();
 b15zdnd11an1n64x5 FILLER_160_1220 ();
 b15zdnd11an1n64x5 FILLER_160_1284 ();
 b15zdnd11an1n64x5 FILLER_160_1348 ();
 b15zdnd11an1n64x5 FILLER_160_1412 ();
 b15zdnd11an1n64x5 FILLER_160_1476 ();
 b15zdnd11an1n64x5 FILLER_160_1540 ();
 b15zdnd11an1n64x5 FILLER_160_1604 ();
 b15zdnd11an1n32x5 FILLER_160_1668 ();
 b15zdnd11an1n08x5 FILLER_160_1700 ();
 b15zdnd11an1n04x5 FILLER_160_1708 ();
 b15zdnd00an1n01x5 FILLER_160_1712 ();
 b15zdnd11an1n64x5 FILLER_160_1734 ();
 b15zdnd11an1n64x5 FILLER_160_1798 ();
 b15zdnd11an1n64x5 FILLER_160_1862 ();
 b15zdnd11an1n64x5 FILLER_160_1926 ();
 b15zdnd11an1n64x5 FILLER_160_1990 ();
 b15zdnd11an1n64x5 FILLER_160_2054 ();
 b15zdnd11an1n32x5 FILLER_160_2118 ();
 b15zdnd11an1n04x5 FILLER_160_2150 ();
 b15zdnd11an1n64x5 FILLER_160_2162 ();
 b15zdnd11an1n32x5 FILLER_160_2226 ();
 b15zdnd11an1n16x5 FILLER_160_2258 ();
 b15zdnd00an1n02x5 FILLER_160_2274 ();
 b15zdnd11an1n64x5 FILLER_161_0 ();
 b15zdnd11an1n64x5 FILLER_161_64 ();
 b15zdnd11an1n32x5 FILLER_161_128 ();
 b15zdnd11an1n08x5 FILLER_161_160 ();
 b15zdnd00an1n02x5 FILLER_161_168 ();
 b15zdnd11an1n04x5 FILLER_161_173 ();
 b15zdnd11an1n04x5 FILLER_161_189 ();
 b15zdnd11an1n64x5 FILLER_161_211 ();
 b15zdnd11an1n64x5 FILLER_161_275 ();
 b15zdnd11an1n64x5 FILLER_161_339 ();
 b15zdnd11an1n64x5 FILLER_161_403 ();
 b15zdnd11an1n64x5 FILLER_161_467 ();
 b15zdnd11an1n16x5 FILLER_161_531 ();
 b15zdnd11an1n08x5 FILLER_161_547 ();
 b15zdnd00an1n02x5 FILLER_161_555 ();
 b15zdnd11an1n04x5 FILLER_161_560 ();
 b15zdnd11an1n04x5 FILLER_161_567 ();
 b15zdnd11an1n04x5 FILLER_161_574 ();
 b15zdnd11an1n64x5 FILLER_161_581 ();
 b15zdnd11an1n64x5 FILLER_161_645 ();
 b15zdnd11an1n08x5 FILLER_161_709 ();
 b15zdnd00an1n02x5 FILLER_161_717 ();
 b15zdnd00an1n01x5 FILLER_161_719 ();
 b15zdnd11an1n64x5 FILLER_161_724 ();
 b15zdnd11an1n32x5 FILLER_161_788 ();
 b15zdnd11an1n08x5 FILLER_161_820 ();
 b15zdnd11an1n04x5 FILLER_161_828 ();
 b15zdnd00an1n02x5 FILLER_161_832 ();
 b15zdnd11an1n16x5 FILLER_161_854 ();
 b15zdnd11an1n08x5 FILLER_161_870 ();
 b15zdnd11an1n04x5 FILLER_161_878 ();
 b15zdnd00an1n01x5 FILLER_161_882 ();
 b15zdnd11an1n64x5 FILLER_161_903 ();
 b15zdnd11an1n64x5 FILLER_161_967 ();
 b15zdnd11an1n64x5 FILLER_161_1031 ();
 b15zdnd11an1n64x5 FILLER_161_1095 ();
 b15zdnd11an1n08x5 FILLER_161_1159 ();
 b15zdnd11an1n32x5 FILLER_161_1179 ();
 b15zdnd11an1n16x5 FILLER_161_1211 ();
 b15zdnd11an1n08x5 FILLER_161_1227 ();
 b15zdnd11an1n64x5 FILLER_161_1255 ();
 b15zdnd11an1n64x5 FILLER_161_1319 ();
 b15zdnd11an1n16x5 FILLER_161_1383 ();
 b15zdnd11an1n08x5 FILLER_161_1399 ();
 b15zdnd11an1n64x5 FILLER_161_1416 ();
 b15zdnd11an1n64x5 FILLER_161_1480 ();
 b15zdnd11an1n64x5 FILLER_161_1544 ();
 b15zdnd11an1n64x5 FILLER_161_1608 ();
 b15zdnd11an1n64x5 FILLER_161_1672 ();
 b15zdnd11an1n64x5 FILLER_161_1736 ();
 b15zdnd11an1n64x5 FILLER_161_1800 ();
 b15zdnd00an1n01x5 FILLER_161_1864 ();
 b15zdnd11an1n64x5 FILLER_161_1874 ();
 b15zdnd11an1n64x5 FILLER_161_1938 ();
 b15zdnd00an1n02x5 FILLER_161_2002 ();
 b15zdnd00an1n01x5 FILLER_161_2004 ();
 b15zdnd11an1n64x5 FILLER_161_2019 ();
 b15zdnd11an1n64x5 FILLER_161_2083 ();
 b15zdnd11an1n32x5 FILLER_161_2147 ();
 b15zdnd11an1n16x5 FILLER_161_2179 ();
 b15zdnd11an1n08x5 FILLER_161_2195 ();
 b15zdnd00an1n01x5 FILLER_161_2203 ();
 b15zdnd11an1n32x5 FILLER_161_2228 ();
 b15zdnd11an1n16x5 FILLER_161_2260 ();
 b15zdnd11an1n08x5 FILLER_161_2276 ();
 b15zdnd11an1n64x5 FILLER_162_8 ();
 b15zdnd11an1n64x5 FILLER_162_72 ();
 b15zdnd11an1n32x5 FILLER_162_136 ();
 b15zdnd11an1n08x5 FILLER_162_168 ();
 b15zdnd00an1n01x5 FILLER_162_176 ();
 b15zdnd11an1n04x5 FILLER_162_181 ();
 b15zdnd00an1n02x5 FILLER_162_185 ();
 b15zdnd11an1n16x5 FILLER_162_205 ();
 b15zdnd11an1n08x5 FILLER_162_221 ();
 b15zdnd00an1n02x5 FILLER_162_229 ();
 b15zdnd11an1n64x5 FILLER_162_235 ();
 b15zdnd11an1n64x5 FILLER_162_299 ();
 b15zdnd11an1n64x5 FILLER_162_363 ();
 b15zdnd11an1n64x5 FILLER_162_427 ();
 b15zdnd11an1n64x5 FILLER_162_491 ();
 b15zdnd00an1n01x5 FILLER_162_555 ();
 b15zdnd11an1n64x5 FILLER_162_559 ();
 b15zdnd11an1n64x5 FILLER_162_623 ();
 b15zdnd11an1n16x5 FILLER_162_687 ();
 b15zdnd11an1n08x5 FILLER_162_703 ();
 b15zdnd11an1n04x5 FILLER_162_711 ();
 b15zdnd00an1n02x5 FILLER_162_715 ();
 b15zdnd00an1n01x5 FILLER_162_717 ();
 b15zdnd11an1n16x5 FILLER_162_726 ();
 b15zdnd11an1n64x5 FILLER_162_753 ();
 b15zdnd11an1n64x5 FILLER_162_817 ();
 b15zdnd11an1n64x5 FILLER_162_881 ();
 b15zdnd11an1n16x5 FILLER_162_945 ();
 b15zdnd11an1n04x5 FILLER_162_961 ();
 b15zdnd00an1n02x5 FILLER_162_965 ();
 b15zdnd11an1n64x5 FILLER_162_983 ();
 b15zdnd11an1n32x5 FILLER_162_1047 ();
 b15zdnd11an1n08x5 FILLER_162_1079 ();
 b15zdnd11an1n04x5 FILLER_162_1087 ();
 b15zdnd11an1n32x5 FILLER_162_1105 ();
 b15zdnd11an1n16x5 FILLER_162_1137 ();
 b15zdnd11an1n08x5 FILLER_162_1153 ();
 b15zdnd11an1n04x5 FILLER_162_1161 ();
 b15zdnd00an1n01x5 FILLER_162_1165 ();
 b15zdnd11an1n16x5 FILLER_162_1186 ();
 b15zdnd11an1n08x5 FILLER_162_1202 ();
 b15zdnd00an1n01x5 FILLER_162_1210 ();
 b15zdnd11an1n64x5 FILLER_162_1227 ();
 b15zdnd11an1n64x5 FILLER_162_1291 ();
 b15zdnd11an1n64x5 FILLER_162_1355 ();
 b15zdnd11an1n64x5 FILLER_162_1419 ();
 b15zdnd11an1n64x5 FILLER_162_1483 ();
 b15zdnd11an1n64x5 FILLER_162_1547 ();
 b15zdnd11an1n64x5 FILLER_162_1611 ();
 b15zdnd11an1n64x5 FILLER_162_1675 ();
 b15zdnd11an1n64x5 FILLER_162_1739 ();
 b15zdnd11an1n64x5 FILLER_162_1803 ();
 b15zdnd11an1n64x5 FILLER_162_1867 ();
 b15zdnd11an1n64x5 FILLER_162_1931 ();
 b15zdnd11an1n64x5 FILLER_162_1995 ();
 b15zdnd11an1n32x5 FILLER_162_2059 ();
 b15zdnd11an1n16x5 FILLER_162_2091 ();
 b15zdnd11an1n04x5 FILLER_162_2107 ();
 b15zdnd11an1n32x5 FILLER_162_2121 ();
 b15zdnd00an1n01x5 FILLER_162_2153 ();
 b15zdnd11an1n64x5 FILLER_162_2162 ();
 b15zdnd11an1n32x5 FILLER_162_2226 ();
 b15zdnd11an1n16x5 FILLER_162_2258 ();
 b15zdnd00an1n02x5 FILLER_162_2274 ();
 b15zdnd11an1n16x5 FILLER_163_0 ();
 b15zdnd00an1n02x5 FILLER_163_16 ();
 b15zdnd11an1n64x5 FILLER_163_22 ();
 b15zdnd11an1n64x5 FILLER_163_86 ();
 b15zdnd11an1n16x5 FILLER_163_150 ();
 b15zdnd11an1n04x5 FILLER_163_166 ();
 b15zdnd00an1n01x5 FILLER_163_170 ();
 b15zdnd11an1n04x5 FILLER_163_177 ();
 b15zdnd11an1n08x5 FILLER_163_187 ();
 b15zdnd11an1n04x5 FILLER_163_195 ();
 b15zdnd00an1n01x5 FILLER_163_199 ();
 b15zdnd11an1n16x5 FILLER_163_203 ();
 b15zdnd11an1n08x5 FILLER_163_219 ();
 b15zdnd11an1n04x5 FILLER_163_231 ();
 b15zdnd11an1n04x5 FILLER_163_248 ();
 b15zdnd11an1n64x5 FILLER_163_262 ();
 b15zdnd11an1n64x5 FILLER_163_326 ();
 b15zdnd11an1n64x5 FILLER_163_390 ();
 b15zdnd11an1n64x5 FILLER_163_454 ();
 b15zdnd11an1n64x5 FILLER_163_518 ();
 b15zdnd11an1n64x5 FILLER_163_582 ();
 b15zdnd11an1n64x5 FILLER_163_646 ();
 b15zdnd11an1n16x5 FILLER_163_710 ();
 b15zdnd11an1n64x5 FILLER_163_730 ();
 b15zdnd11an1n32x5 FILLER_163_794 ();
 b15zdnd11an1n16x5 FILLER_163_826 ();
 b15zdnd11an1n08x5 FILLER_163_842 ();
 b15zdnd11an1n04x5 FILLER_163_850 ();
 b15zdnd00an1n02x5 FILLER_163_854 ();
 b15zdnd11an1n64x5 FILLER_163_879 ();
 b15zdnd11an1n64x5 FILLER_163_943 ();
 b15zdnd11an1n64x5 FILLER_163_1007 ();
 b15zdnd11an1n64x5 FILLER_163_1071 ();
 b15zdnd11an1n64x5 FILLER_163_1135 ();
 b15zdnd11an1n64x5 FILLER_163_1199 ();
 b15zdnd11an1n64x5 FILLER_163_1263 ();
 b15zdnd11an1n64x5 FILLER_163_1327 ();
 b15zdnd11an1n64x5 FILLER_163_1391 ();
 b15zdnd11an1n64x5 FILLER_163_1455 ();
 b15zdnd11an1n64x5 FILLER_163_1519 ();
 b15zdnd11an1n64x5 FILLER_163_1583 ();
 b15zdnd11an1n64x5 FILLER_163_1647 ();
 b15zdnd11an1n32x5 FILLER_163_1711 ();
 b15zdnd11an1n16x5 FILLER_163_1743 ();
 b15zdnd11an1n04x5 FILLER_163_1770 ();
 b15zdnd11an1n64x5 FILLER_163_1788 ();
 b15zdnd11an1n16x5 FILLER_163_1852 ();
 b15zdnd00an1n01x5 FILLER_163_1868 ();
 b15zdnd11an1n64x5 FILLER_163_1873 ();
 b15zdnd11an1n64x5 FILLER_163_1937 ();
 b15zdnd11an1n64x5 FILLER_163_2001 ();
 b15zdnd11an1n64x5 FILLER_163_2065 ();
 b15zdnd11an1n64x5 FILLER_163_2129 ();
 b15zdnd11an1n32x5 FILLER_163_2193 ();
 b15zdnd11an1n16x5 FILLER_163_2225 ();
 b15zdnd11an1n08x5 FILLER_163_2241 ();
 b15zdnd11an1n04x5 FILLER_163_2249 ();
 b15zdnd00an1n02x5 FILLER_163_2253 ();
 b15zdnd00an1n01x5 FILLER_163_2255 ();
 b15zdnd11an1n16x5 FILLER_163_2260 ();
 b15zdnd11an1n08x5 FILLER_163_2276 ();
 b15zdnd11an1n64x5 FILLER_164_8 ();
 b15zdnd11an1n64x5 FILLER_164_72 ();
 b15zdnd11an1n32x5 FILLER_164_136 ();
 b15zdnd11an1n04x5 FILLER_164_168 ();
 b15zdnd00an1n01x5 FILLER_164_172 ();
 b15zdnd11an1n64x5 FILLER_164_189 ();
 b15zdnd11an1n32x5 FILLER_164_253 ();
 b15zdnd11an1n16x5 FILLER_164_285 ();
 b15zdnd11an1n32x5 FILLER_164_343 ();
 b15zdnd11an1n16x5 FILLER_164_375 ();
 b15zdnd11an1n04x5 FILLER_164_391 ();
 b15zdnd00an1n02x5 FILLER_164_395 ();
 b15zdnd00an1n01x5 FILLER_164_397 ();
 b15zdnd11an1n64x5 FILLER_164_401 ();
 b15zdnd11an1n64x5 FILLER_164_465 ();
 b15zdnd11an1n64x5 FILLER_164_529 ();
 b15zdnd11an1n64x5 FILLER_164_593 ();
 b15zdnd11an1n32x5 FILLER_164_657 ();
 b15zdnd11an1n16x5 FILLER_164_689 ();
 b15zdnd11an1n08x5 FILLER_164_705 ();
 b15zdnd11an1n04x5 FILLER_164_713 ();
 b15zdnd00an1n01x5 FILLER_164_717 ();
 b15zdnd11an1n64x5 FILLER_164_726 ();
 b15zdnd11an1n64x5 FILLER_164_790 ();
 b15zdnd11an1n64x5 FILLER_164_854 ();
 b15zdnd11an1n64x5 FILLER_164_918 ();
 b15zdnd11an1n64x5 FILLER_164_982 ();
 b15zdnd11an1n32x5 FILLER_164_1046 ();
 b15zdnd11an1n16x5 FILLER_164_1078 ();
 b15zdnd11an1n08x5 FILLER_164_1094 ();
 b15zdnd11an1n64x5 FILLER_164_1106 ();
 b15zdnd11an1n64x5 FILLER_164_1170 ();
 b15zdnd11an1n64x5 FILLER_164_1234 ();
 b15zdnd11an1n64x5 FILLER_164_1298 ();
 b15zdnd11an1n04x5 FILLER_164_1377 ();
 b15zdnd11an1n64x5 FILLER_164_1390 ();
 b15zdnd11an1n64x5 FILLER_164_1454 ();
 b15zdnd11an1n32x5 FILLER_164_1518 ();
 b15zdnd11an1n16x5 FILLER_164_1550 ();
 b15zdnd11an1n08x5 FILLER_164_1566 ();
 b15zdnd11an1n04x5 FILLER_164_1574 ();
 b15zdnd00an1n02x5 FILLER_164_1578 ();
 b15zdnd00an1n01x5 FILLER_164_1580 ();
 b15zdnd11an1n32x5 FILLER_164_1589 ();
 b15zdnd11an1n16x5 FILLER_164_1621 ();
 b15zdnd11an1n04x5 FILLER_164_1637 ();
 b15zdnd00an1n02x5 FILLER_164_1641 ();
 b15zdnd11an1n64x5 FILLER_164_1664 ();
 b15zdnd11an1n64x5 FILLER_164_1728 ();
 b15zdnd11an1n64x5 FILLER_164_1792 ();
 b15zdnd00an1n02x5 FILLER_164_1856 ();
 b15zdnd00an1n01x5 FILLER_164_1858 ();
 b15zdnd11an1n04x5 FILLER_164_1863 ();
 b15zdnd11an1n64x5 FILLER_164_1883 ();
 b15zdnd11an1n64x5 FILLER_164_1947 ();
 b15zdnd11an1n08x5 FILLER_164_2011 ();
 b15zdnd11an1n04x5 FILLER_164_2026 ();
 b15zdnd00an1n02x5 FILLER_164_2030 ();
 b15zdnd11an1n64x5 FILLER_164_2044 ();
 b15zdnd11an1n32x5 FILLER_164_2108 ();
 b15zdnd11an1n08x5 FILLER_164_2140 ();
 b15zdnd11an1n04x5 FILLER_164_2148 ();
 b15zdnd00an1n02x5 FILLER_164_2152 ();
 b15zdnd11an1n32x5 FILLER_164_2162 ();
 b15zdnd11an1n08x5 FILLER_164_2194 ();
 b15zdnd11an1n04x5 FILLER_164_2202 ();
 b15zdnd00an1n02x5 FILLER_164_2206 ();
 b15zdnd00an1n01x5 FILLER_164_2208 ();
 b15zdnd11an1n32x5 FILLER_164_2222 ();
 b15zdnd11an1n16x5 FILLER_164_2254 ();
 b15zdnd11an1n04x5 FILLER_164_2270 ();
 b15zdnd00an1n02x5 FILLER_164_2274 ();
 b15zdnd11an1n64x5 FILLER_165_0 ();
 b15zdnd11an1n64x5 FILLER_165_64 ();
 b15zdnd11an1n16x5 FILLER_165_128 ();
 b15zdnd11an1n04x5 FILLER_165_144 ();
 b15zdnd11an1n32x5 FILLER_165_162 ();
 b15zdnd11an1n16x5 FILLER_165_194 ();
 b15zdnd11an1n08x5 FILLER_165_210 ();
 b15zdnd00an1n02x5 FILLER_165_218 ();
 b15zdnd00an1n01x5 FILLER_165_220 ();
 b15zdnd11an1n64x5 FILLER_165_232 ();
 b15zdnd11an1n64x5 FILLER_165_296 ();
 b15zdnd11an1n08x5 FILLER_165_360 ();
 b15zdnd00an1n02x5 FILLER_165_368 ();
 b15zdnd00an1n01x5 FILLER_165_370 ();
 b15zdnd11an1n64x5 FILLER_165_423 ();
 b15zdnd11an1n64x5 FILLER_165_487 ();
 b15zdnd11an1n64x5 FILLER_165_551 ();
 b15zdnd11an1n16x5 FILLER_165_615 ();
 b15zdnd11an1n08x5 FILLER_165_631 ();
 b15zdnd11an1n04x5 FILLER_165_639 ();
 b15zdnd11an1n64x5 FILLER_165_657 ();
 b15zdnd11an1n64x5 FILLER_165_721 ();
 b15zdnd11an1n64x5 FILLER_165_785 ();
 b15zdnd11an1n64x5 FILLER_165_849 ();
 b15zdnd11an1n32x5 FILLER_165_913 ();
 b15zdnd11an1n16x5 FILLER_165_945 ();
 b15zdnd00an1n02x5 FILLER_165_961 ();
 b15zdnd00an1n01x5 FILLER_165_963 ();
 b15zdnd11an1n64x5 FILLER_165_967 ();
 b15zdnd11an1n32x5 FILLER_165_1031 ();
 b15zdnd11an1n16x5 FILLER_165_1063 ();
 b15zdnd11an1n04x5 FILLER_165_1079 ();
 b15zdnd00an1n01x5 FILLER_165_1083 ();
 b15zdnd11an1n32x5 FILLER_165_1087 ();
 b15zdnd11an1n64x5 FILLER_165_1123 ();
 b15zdnd11an1n64x5 FILLER_165_1187 ();
 b15zdnd11an1n64x5 FILLER_165_1251 ();
 b15zdnd11an1n64x5 FILLER_165_1315 ();
 b15zdnd11an1n64x5 FILLER_165_1379 ();
 b15zdnd11an1n64x5 FILLER_165_1443 ();
 b15zdnd11an1n64x5 FILLER_165_1507 ();
 b15zdnd11an1n32x5 FILLER_165_1571 ();
 b15zdnd11an1n04x5 FILLER_165_1603 ();
 b15zdnd00an1n01x5 FILLER_165_1607 ();
 b15zdnd11an1n64x5 FILLER_165_1618 ();
 b15zdnd11an1n64x5 FILLER_165_1682 ();
 b15zdnd11an1n16x5 FILLER_165_1746 ();
 b15zdnd11an1n04x5 FILLER_165_1762 ();
 b15zdnd00an1n02x5 FILLER_165_1766 ();
 b15zdnd11an1n64x5 FILLER_165_1784 ();
 b15zdnd00an1n02x5 FILLER_165_1848 ();
 b15zdnd00an1n01x5 FILLER_165_1850 ();
 b15zdnd11an1n64x5 FILLER_165_1872 ();
 b15zdnd11an1n64x5 FILLER_165_1936 ();
 b15zdnd11an1n64x5 FILLER_165_2000 ();
 b15zdnd11an1n64x5 FILLER_165_2064 ();
 b15zdnd11an1n64x5 FILLER_165_2128 ();
 b15zdnd11an1n64x5 FILLER_165_2192 ();
 b15zdnd11an1n16x5 FILLER_165_2256 ();
 b15zdnd11an1n08x5 FILLER_165_2272 ();
 b15zdnd11an1n04x5 FILLER_165_2280 ();
 b15zdnd11an1n64x5 FILLER_166_8 ();
 b15zdnd11an1n64x5 FILLER_166_72 ();
 b15zdnd11an1n08x5 FILLER_166_136 ();
 b15zdnd11an1n64x5 FILLER_166_149 ();
 b15zdnd11an1n64x5 FILLER_166_213 ();
 b15zdnd11an1n64x5 FILLER_166_277 ();
 b15zdnd11an1n32x5 FILLER_166_341 ();
 b15zdnd11an1n16x5 FILLER_166_373 ();
 b15zdnd11an1n04x5 FILLER_166_392 ();
 b15zdnd11an1n32x5 FILLER_166_399 ();
 b15zdnd00an1n01x5 FILLER_166_431 ();
 b15zdnd11an1n64x5 FILLER_166_441 ();
 b15zdnd11an1n64x5 FILLER_166_505 ();
 b15zdnd11an1n32x5 FILLER_166_569 ();
 b15zdnd11an1n04x5 FILLER_166_601 ();
 b15zdnd00an1n01x5 FILLER_166_605 ();
 b15zdnd11an1n64x5 FILLER_166_616 ();
 b15zdnd11an1n32x5 FILLER_166_680 ();
 b15zdnd11an1n04x5 FILLER_166_712 ();
 b15zdnd00an1n02x5 FILLER_166_716 ();
 b15zdnd00an1n02x5 FILLER_166_726 ();
 b15zdnd11an1n64x5 FILLER_166_749 ();
 b15zdnd11an1n64x5 FILLER_166_813 ();
 b15zdnd11an1n32x5 FILLER_166_877 ();
 b15zdnd11an1n08x5 FILLER_166_909 ();
 b15zdnd11an1n04x5 FILLER_166_917 ();
 b15zdnd11an1n32x5 FILLER_166_934 ();
 b15zdnd11an1n16x5 FILLER_166_966 ();
 b15zdnd11an1n08x5 FILLER_166_982 ();
 b15zdnd00an1n01x5 FILLER_166_990 ();
 b15zdnd11an1n64x5 FILLER_166_995 ();
 b15zdnd11an1n32x5 FILLER_166_1059 ();
 b15zdnd11an1n08x5 FILLER_166_1091 ();
 b15zdnd00an1n02x5 FILLER_166_1099 ();
 b15zdnd00an1n01x5 FILLER_166_1101 ();
 b15zdnd11an1n64x5 FILLER_166_1116 ();
 b15zdnd11an1n08x5 FILLER_166_1180 ();
 b15zdnd11an1n04x5 FILLER_166_1188 ();
 b15zdnd00an1n02x5 FILLER_166_1192 ();
 b15zdnd11an1n64x5 FILLER_166_1208 ();
 b15zdnd11an1n64x5 FILLER_166_1272 ();
 b15zdnd11an1n64x5 FILLER_166_1336 ();
 b15zdnd11an1n64x5 FILLER_166_1400 ();
 b15zdnd11an1n64x5 FILLER_166_1464 ();
 b15zdnd11an1n64x5 FILLER_166_1528 ();
 b15zdnd11an1n16x5 FILLER_166_1592 ();
 b15zdnd11an1n04x5 FILLER_166_1608 ();
 b15zdnd00an1n02x5 FILLER_166_1612 ();
 b15zdnd00an1n01x5 FILLER_166_1614 ();
 b15zdnd11an1n16x5 FILLER_166_1618 ();
 b15zdnd11an1n04x5 FILLER_166_1634 ();
 b15zdnd11an1n64x5 FILLER_166_1652 ();
 b15zdnd11an1n64x5 FILLER_166_1716 ();
 b15zdnd11an1n64x5 FILLER_166_1780 ();
 b15zdnd11an1n64x5 FILLER_166_1844 ();
 b15zdnd11an1n64x5 FILLER_166_1908 ();
 b15zdnd11an1n08x5 FILLER_166_1972 ();
 b15zdnd11an1n04x5 FILLER_166_1980 ();
 b15zdnd00an1n02x5 FILLER_166_1984 ();
 b15zdnd00an1n01x5 FILLER_166_1986 ();
 b15zdnd11an1n64x5 FILLER_166_1996 ();
 b15zdnd11an1n08x5 FILLER_166_2060 ();
 b15zdnd11an1n04x5 FILLER_166_2068 ();
 b15zdnd00an1n02x5 FILLER_166_2072 ();
 b15zdnd11an1n64x5 FILLER_166_2078 ();
 b15zdnd11an1n08x5 FILLER_166_2142 ();
 b15zdnd11an1n04x5 FILLER_166_2150 ();
 b15zdnd11an1n32x5 FILLER_166_2162 ();
 b15zdnd11an1n16x5 FILLER_166_2194 ();
 b15zdnd11an1n08x5 FILLER_166_2210 ();
 b15zdnd00an1n02x5 FILLER_166_2218 ();
 b15zdnd11an1n08x5 FILLER_166_2262 ();
 b15zdnd11an1n04x5 FILLER_166_2270 ();
 b15zdnd00an1n02x5 FILLER_166_2274 ();
 b15zdnd11an1n32x5 FILLER_167_0 ();
 b15zdnd11an1n04x5 FILLER_167_32 ();
 b15zdnd00an1n02x5 FILLER_167_36 ();
 b15zdnd00an1n01x5 FILLER_167_38 ();
 b15zdnd11an1n64x5 FILLER_167_44 ();
 b15zdnd11an1n64x5 FILLER_167_108 ();
 b15zdnd11an1n16x5 FILLER_167_172 ();
 b15zdnd11an1n08x5 FILLER_167_188 ();
 b15zdnd11an1n04x5 FILLER_167_196 ();
 b15zdnd00an1n02x5 FILLER_167_200 ();
 b15zdnd11an1n64x5 FILLER_167_205 ();
 b15zdnd11an1n64x5 FILLER_167_269 ();
 b15zdnd11an1n64x5 FILLER_167_333 ();
 b15zdnd11an1n64x5 FILLER_167_397 ();
 b15zdnd11an1n64x5 FILLER_167_461 ();
 b15zdnd11an1n64x5 FILLER_167_525 ();
 b15zdnd11an1n16x5 FILLER_167_589 ();
 b15zdnd11an1n04x5 FILLER_167_605 ();
 b15zdnd00an1n01x5 FILLER_167_609 ();
 b15zdnd11an1n64x5 FILLER_167_617 ();
 b15zdnd11an1n64x5 FILLER_167_681 ();
 b15zdnd11an1n64x5 FILLER_167_745 ();
 b15zdnd11an1n32x5 FILLER_167_809 ();
 b15zdnd00an1n01x5 FILLER_167_841 ();
 b15zdnd11an1n64x5 FILLER_167_846 ();
 b15zdnd11an1n32x5 FILLER_167_910 ();
 b15zdnd11an1n04x5 FILLER_167_942 ();
 b15zdnd00an1n01x5 FILLER_167_946 ();
 b15zdnd11an1n08x5 FILLER_167_967 ();
 b15zdnd11an1n64x5 FILLER_167_994 ();
 b15zdnd11an1n64x5 FILLER_167_1058 ();
 b15zdnd11an1n32x5 FILLER_167_1122 ();
 b15zdnd11an1n16x5 FILLER_167_1154 ();
 b15zdnd11an1n08x5 FILLER_167_1170 ();
 b15zdnd11an1n04x5 FILLER_167_1178 ();
 b15zdnd00an1n01x5 FILLER_167_1182 ();
 b15zdnd11an1n64x5 FILLER_167_1196 ();
 b15zdnd11an1n08x5 FILLER_167_1260 ();
 b15zdnd11an1n32x5 FILLER_167_1277 ();
 b15zdnd11an1n16x5 FILLER_167_1309 ();
 b15zdnd11an1n08x5 FILLER_167_1325 ();
 b15zdnd11an1n04x5 FILLER_167_1333 ();
 b15zdnd11an1n64x5 FILLER_167_1340 ();
 b15zdnd11an1n64x5 FILLER_167_1404 ();
 b15zdnd11an1n32x5 FILLER_167_1468 ();
 b15zdnd00an1n02x5 FILLER_167_1500 ();
 b15zdnd00an1n01x5 FILLER_167_1502 ();
 b15zdnd11an1n64x5 FILLER_167_1512 ();
 b15zdnd11an1n08x5 FILLER_167_1576 ();
 b15zdnd00an1n02x5 FILLER_167_1584 ();
 b15zdnd11an1n64x5 FILLER_167_1628 ();
 b15zdnd11an1n64x5 FILLER_167_1692 ();
 b15zdnd11an1n08x5 FILLER_167_1756 ();
 b15zdnd11an1n04x5 FILLER_167_1764 ();
 b15zdnd00an1n01x5 FILLER_167_1768 ();
 b15zdnd11an1n64x5 FILLER_167_1780 ();
 b15zdnd11an1n32x5 FILLER_167_1844 ();
 b15zdnd00an1n02x5 FILLER_167_1876 ();
 b15zdnd11an1n64x5 FILLER_167_1930 ();
 b15zdnd11an1n64x5 FILLER_167_1994 ();
 b15zdnd11an1n64x5 FILLER_167_2058 ();
 b15zdnd11an1n64x5 FILLER_167_2122 ();
 b15zdnd11an1n32x5 FILLER_167_2186 ();
 b15zdnd11an1n16x5 FILLER_167_2218 ();
 b15zdnd11an1n08x5 FILLER_167_2234 ();
 b15zdnd11an1n04x5 FILLER_167_2242 ();
 b15zdnd00an1n02x5 FILLER_167_2246 ();
 b15zdnd11an1n16x5 FILLER_167_2259 ();
 b15zdnd11an1n08x5 FILLER_167_2275 ();
 b15zdnd00an1n01x5 FILLER_167_2283 ();
 b15zdnd11an1n64x5 FILLER_168_8 ();
 b15zdnd11an1n64x5 FILLER_168_72 ();
 b15zdnd11an1n64x5 FILLER_168_136 ();
 b15zdnd11an1n32x5 FILLER_168_200 ();
 b15zdnd11an1n08x5 FILLER_168_232 ();
 b15zdnd11an1n64x5 FILLER_168_245 ();
 b15zdnd11an1n64x5 FILLER_168_309 ();
 b15zdnd11an1n32x5 FILLER_168_373 ();
 b15zdnd11an1n16x5 FILLER_168_405 ();
 b15zdnd11an1n04x5 FILLER_168_421 ();
 b15zdnd00an1n02x5 FILLER_168_425 ();
 b15zdnd11an1n64x5 FILLER_168_430 ();
 b15zdnd11an1n64x5 FILLER_168_494 ();
 b15zdnd11an1n32x5 FILLER_168_558 ();
 b15zdnd11an1n16x5 FILLER_168_590 ();
 b15zdnd00an1n02x5 FILLER_168_606 ();
 b15zdnd11an1n64x5 FILLER_168_619 ();
 b15zdnd11an1n32x5 FILLER_168_683 ();
 b15zdnd00an1n02x5 FILLER_168_715 ();
 b15zdnd00an1n01x5 FILLER_168_717 ();
 b15zdnd11an1n64x5 FILLER_168_726 ();
 b15zdnd11an1n32x5 FILLER_168_790 ();
 b15zdnd11an1n16x5 FILLER_168_822 ();
 b15zdnd11an1n04x5 FILLER_168_838 ();
 b15zdnd11an1n64x5 FILLER_168_853 ();
 b15zdnd11an1n32x5 FILLER_168_917 ();
 b15zdnd11an1n16x5 FILLER_168_949 ();
 b15zdnd11an1n04x5 FILLER_168_965 ();
 b15zdnd00an1n02x5 FILLER_168_969 ();
 b15zdnd11an1n64x5 FILLER_168_991 ();
 b15zdnd11an1n16x5 FILLER_168_1055 ();
 b15zdnd11an1n08x5 FILLER_168_1071 ();
 b15zdnd11an1n04x5 FILLER_168_1079 ();
 b15zdnd00an1n02x5 FILLER_168_1083 ();
 b15zdnd11an1n16x5 FILLER_168_1093 ();
 b15zdnd11an1n08x5 FILLER_168_1109 ();
 b15zdnd00an1n01x5 FILLER_168_1117 ();
 b15zdnd11an1n16x5 FILLER_168_1155 ();
 b15zdnd11an1n08x5 FILLER_168_1171 ();
 b15zdnd11an1n04x5 FILLER_168_1179 ();
 b15zdnd00an1n01x5 FILLER_168_1183 ();
 b15zdnd11an1n64x5 FILLER_168_1196 ();
 b15zdnd11an1n16x5 FILLER_168_1260 ();
 b15zdnd11an1n08x5 FILLER_168_1276 ();
 b15zdnd11an1n04x5 FILLER_168_1284 ();
 b15zdnd00an1n01x5 FILLER_168_1288 ();
 b15zdnd11an1n16x5 FILLER_168_1303 ();
 b15zdnd11an1n04x5 FILLER_168_1319 ();
 b15zdnd00an1n01x5 FILLER_168_1323 ();
 b15zdnd11an1n04x5 FILLER_168_1335 ();
 b15zdnd11an1n04x5 FILLER_168_1342 ();
 b15zdnd11an1n64x5 FILLER_168_1349 ();
 b15zdnd11an1n32x5 FILLER_168_1413 ();
 b15zdnd11an1n16x5 FILLER_168_1445 ();
 b15zdnd11an1n04x5 FILLER_168_1461 ();
 b15zdnd00an1n01x5 FILLER_168_1465 ();
 b15zdnd11an1n32x5 FILLER_168_1469 ();
 b15zdnd11an1n08x5 FILLER_168_1501 ();
 b15zdnd11an1n04x5 FILLER_168_1509 ();
 b15zdnd11an1n32x5 FILLER_168_1531 ();
 b15zdnd11an1n08x5 FILLER_168_1563 ();
 b15zdnd00an1n02x5 FILLER_168_1571 ();
 b15zdnd00an1n01x5 FILLER_168_1573 ();
 b15zdnd11an1n04x5 FILLER_168_1616 ();
 b15zdnd11an1n64x5 FILLER_168_1636 ();
 b15zdnd11an1n64x5 FILLER_168_1700 ();
 b15zdnd11an1n64x5 FILLER_168_1764 ();
 b15zdnd11an1n64x5 FILLER_168_1828 ();
 b15zdnd11an1n04x5 FILLER_168_1892 ();
 b15zdnd11an1n04x5 FILLER_168_1899 ();
 b15zdnd11an1n04x5 FILLER_168_1906 ();
 b15zdnd11an1n64x5 FILLER_168_1913 ();
 b15zdnd11an1n64x5 FILLER_168_1977 ();
 b15zdnd11an1n64x5 FILLER_168_2041 ();
 b15zdnd11an1n32x5 FILLER_168_2105 ();
 b15zdnd11an1n16x5 FILLER_168_2137 ();
 b15zdnd00an1n01x5 FILLER_168_2153 ();
 b15zdnd11an1n64x5 FILLER_168_2162 ();
 b15zdnd11an1n08x5 FILLER_168_2226 ();
 b15zdnd11an1n04x5 FILLER_168_2234 ();
 b15zdnd11an1n04x5 FILLER_168_2258 ();
 b15zdnd11an1n08x5 FILLER_168_2267 ();
 b15zdnd00an1n01x5 FILLER_168_2275 ();
 b15zdnd11an1n64x5 FILLER_169_0 ();
 b15zdnd11an1n64x5 FILLER_169_64 ();
 b15zdnd11an1n64x5 FILLER_169_128 ();
 b15zdnd11an1n16x5 FILLER_169_192 ();
 b15zdnd11an1n04x5 FILLER_169_208 ();
 b15zdnd00an1n01x5 FILLER_169_212 ();
 b15zdnd11an1n32x5 FILLER_169_228 ();
 b15zdnd11an1n16x5 FILLER_169_260 ();
 b15zdnd11an1n04x5 FILLER_169_276 ();
 b15zdnd11an1n04x5 FILLER_169_322 ();
 b15zdnd11an1n32x5 FILLER_169_368 ();
 b15zdnd11an1n16x5 FILLER_169_400 ();
 b15zdnd11an1n64x5 FILLER_169_458 ();
 b15zdnd11an1n64x5 FILLER_169_522 ();
 b15zdnd11an1n32x5 FILLER_169_586 ();
 b15zdnd11an1n16x5 FILLER_169_618 ();
 b15zdnd11an1n08x5 FILLER_169_634 ();
 b15zdnd00an1n02x5 FILLER_169_642 ();
 b15zdnd11an1n04x5 FILLER_169_651 ();
 b15zdnd11an1n32x5 FILLER_169_665 ();
 b15zdnd11an1n04x5 FILLER_169_697 ();
 b15zdnd00an1n02x5 FILLER_169_701 ();
 b15zdnd00an1n01x5 FILLER_169_703 ();
 b15zdnd11an1n64x5 FILLER_169_714 ();
 b15zdnd11an1n64x5 FILLER_169_778 ();
 b15zdnd11an1n64x5 FILLER_169_842 ();
 b15zdnd11an1n64x5 FILLER_169_906 ();
 b15zdnd11an1n16x5 FILLER_169_970 ();
 b15zdnd11an1n04x5 FILLER_169_986 ();
 b15zdnd00an1n02x5 FILLER_169_990 ();
 b15zdnd00an1n01x5 FILLER_169_992 ();
 b15zdnd11an1n64x5 FILLER_169_1004 ();
 b15zdnd11an1n64x5 FILLER_169_1068 ();
 b15zdnd11an1n64x5 FILLER_169_1132 ();
 b15zdnd11an1n32x5 FILLER_169_1196 ();
 b15zdnd11an1n16x5 FILLER_169_1228 ();
 b15zdnd11an1n08x5 FILLER_169_1244 ();
 b15zdnd11an1n04x5 FILLER_169_1252 ();
 b15zdnd11an1n16x5 FILLER_169_1276 ();
 b15zdnd00an1n01x5 FILLER_169_1292 ();
 b15zdnd11an1n08x5 FILLER_169_1302 ();
 b15zdnd11an1n04x5 FILLER_169_1310 ();
 b15zdnd11an1n64x5 FILLER_169_1366 ();
 b15zdnd11an1n08x5 FILLER_169_1430 ();
 b15zdnd00an1n02x5 FILLER_169_1438 ();
 b15zdnd11an1n04x5 FILLER_169_1492 ();
 b15zdnd11an1n64x5 FILLER_169_1505 ();
 b15zdnd11an1n04x5 FILLER_169_1583 ();
 b15zdnd11an1n64x5 FILLER_169_1639 ();
 b15zdnd11an1n64x5 FILLER_169_1703 ();
 b15zdnd11an1n32x5 FILLER_169_1767 ();
 b15zdnd11an1n16x5 FILLER_169_1799 ();
 b15zdnd11an1n04x5 FILLER_169_1815 ();
 b15zdnd00an1n02x5 FILLER_169_1819 ();
 b15zdnd11an1n64x5 FILLER_169_1833 ();
 b15zdnd00an1n02x5 FILLER_169_1897 ();
 b15zdnd11an1n64x5 FILLER_169_1915 ();
 b15zdnd11an1n32x5 FILLER_169_1979 ();
 b15zdnd11an1n04x5 FILLER_169_2011 ();
 b15zdnd11an1n32x5 FILLER_169_2057 ();
 b15zdnd11an1n08x5 FILLER_169_2089 ();
 b15zdnd00an1n02x5 FILLER_169_2097 ();
 b15zdnd00an1n01x5 FILLER_169_2099 ();
 b15zdnd11an1n64x5 FILLER_169_2142 ();
 b15zdnd11an1n16x5 FILLER_169_2206 ();
 b15zdnd11an1n08x5 FILLER_169_2222 ();
 b15zdnd11an1n04x5 FILLER_169_2250 ();
 b15zdnd11an1n08x5 FILLER_169_2274 ();
 b15zdnd00an1n02x5 FILLER_169_2282 ();
 b15zdnd11an1n08x5 FILLER_170_8 ();
 b15zdnd00an1n02x5 FILLER_170_16 ();
 b15zdnd11an1n04x5 FILLER_170_22 ();
 b15zdnd00an1n01x5 FILLER_170_26 ();
 b15zdnd11an1n64x5 FILLER_170_32 ();
 b15zdnd11an1n64x5 FILLER_170_96 ();
 b15zdnd11an1n64x5 FILLER_170_160 ();
 b15zdnd11an1n64x5 FILLER_170_224 ();
 b15zdnd11an1n64x5 FILLER_170_288 ();
 b15zdnd11an1n32x5 FILLER_170_352 ();
 b15zdnd11an1n16x5 FILLER_170_384 ();
 b15zdnd11an1n16x5 FILLER_170_452 ();
 b15zdnd11an1n08x5 FILLER_170_468 ();
 b15zdnd00an1n02x5 FILLER_170_476 ();
 b15zdnd11an1n64x5 FILLER_170_486 ();
 b15zdnd11an1n64x5 FILLER_170_550 ();
 b15zdnd11an1n64x5 FILLER_170_614 ();
 b15zdnd11an1n32x5 FILLER_170_678 ();
 b15zdnd11an1n08x5 FILLER_170_710 ();
 b15zdnd11an1n64x5 FILLER_170_726 ();
 b15zdnd11an1n64x5 FILLER_170_790 ();
 b15zdnd11an1n64x5 FILLER_170_854 ();
 b15zdnd11an1n64x5 FILLER_170_918 ();
 b15zdnd11an1n16x5 FILLER_170_982 ();
 b15zdnd11an1n08x5 FILLER_170_998 ();
 b15zdnd11an1n64x5 FILLER_170_1017 ();
 b15zdnd11an1n64x5 FILLER_170_1081 ();
 b15zdnd11an1n64x5 FILLER_170_1145 ();
 b15zdnd11an1n64x5 FILLER_170_1209 ();
 b15zdnd11an1n32x5 FILLER_170_1273 ();
 b15zdnd00an1n02x5 FILLER_170_1305 ();
 b15zdnd00an1n01x5 FILLER_170_1307 ();
 b15zdnd11an1n16x5 FILLER_170_1350 ();
 b15zdnd11an1n04x5 FILLER_170_1366 ();
 b15zdnd00an1n02x5 FILLER_170_1370 ();
 b15zdnd11an1n04x5 FILLER_170_1399 ();
 b15zdnd00an1n02x5 FILLER_170_1403 ();
 b15zdnd00an1n01x5 FILLER_170_1405 ();
 b15zdnd11an1n04x5 FILLER_170_1409 ();
 b15zdnd00an1n02x5 FILLER_170_1413 ();
 b15zdnd11an1n32x5 FILLER_170_1418 ();
 b15zdnd11an1n08x5 FILLER_170_1450 ();
 b15zdnd11an1n04x5 FILLER_170_1458 ();
 b15zdnd00an1n02x5 FILLER_170_1462 ();
 b15zdnd00an1n01x5 FILLER_170_1464 ();
 b15zdnd11an1n16x5 FILLER_170_1468 ();
 b15zdnd11an1n08x5 FILLER_170_1484 ();
 b15zdnd11an1n64x5 FILLER_170_1501 ();
 b15zdnd11an1n32x5 FILLER_170_1565 ();
 b15zdnd11an1n08x5 FILLER_170_1597 ();
 b15zdnd11an1n04x5 FILLER_170_1605 ();
 b15zdnd00an1n02x5 FILLER_170_1609 ();
 b15zdnd00an1n01x5 FILLER_170_1611 ();
 b15zdnd11an1n16x5 FILLER_170_1615 ();
 b15zdnd11an1n32x5 FILLER_170_1654 ();
 b15zdnd11an1n16x5 FILLER_170_1686 ();
 b15zdnd11an1n08x5 FILLER_170_1702 ();
 b15zdnd11an1n04x5 FILLER_170_1710 ();
 b15zdnd00an1n02x5 FILLER_170_1714 ();
 b15zdnd11an1n64x5 FILLER_170_1735 ();
 b15zdnd11an1n32x5 FILLER_170_1799 ();
 b15zdnd00an1n01x5 FILLER_170_1831 ();
 b15zdnd11an1n32x5 FILLER_170_1839 ();
 b15zdnd11an1n16x5 FILLER_170_1871 ();
 b15zdnd11an1n04x5 FILLER_170_1887 ();
 b15zdnd00an1n02x5 FILLER_170_1891 ();
 b15zdnd00an1n01x5 FILLER_170_1893 ();
 b15zdnd11an1n64x5 FILLER_170_1901 ();
 b15zdnd11an1n08x5 FILLER_170_1965 ();
 b15zdnd11an1n32x5 FILLER_170_2015 ();
 b15zdnd11an1n16x5 FILLER_170_2047 ();
 b15zdnd11an1n32x5 FILLER_170_2105 ();
 b15zdnd11an1n16x5 FILLER_170_2137 ();
 b15zdnd00an1n01x5 FILLER_170_2153 ();
 b15zdnd11an1n16x5 FILLER_170_2162 ();
 b15zdnd11an1n08x5 FILLER_170_2178 ();
 b15zdnd11an1n04x5 FILLER_170_2186 ();
 b15zdnd11an1n16x5 FILLER_170_2207 ();
 b15zdnd11an1n08x5 FILLER_170_2223 ();
 b15zdnd00an1n01x5 FILLER_170_2231 ();
 b15zdnd00an1n02x5 FILLER_170_2274 ();
 b15zdnd11an1n64x5 FILLER_171_0 ();
 b15zdnd11an1n64x5 FILLER_171_64 ();
 b15zdnd11an1n64x5 FILLER_171_128 ();
 b15zdnd00an1n01x5 FILLER_171_192 ();
 b15zdnd11an1n16x5 FILLER_171_235 ();
 b15zdnd11an1n04x5 FILLER_171_251 ();
 b15zdnd00an1n01x5 FILLER_171_255 ();
 b15zdnd11an1n04x5 FILLER_171_288 ();
 b15zdnd11an1n64x5 FILLER_171_295 ();
 b15zdnd11an1n32x5 FILLER_171_359 ();
 b15zdnd11an1n16x5 FILLER_171_391 ();
 b15zdnd11an1n08x5 FILLER_171_407 ();
 b15zdnd00an1n02x5 FILLER_171_415 ();
 b15zdnd00an1n01x5 FILLER_171_417 ();
 b15zdnd11an1n04x5 FILLER_171_421 ();
 b15zdnd11an1n32x5 FILLER_171_428 ();
 b15zdnd11an1n04x5 FILLER_171_460 ();
 b15zdnd00an1n01x5 FILLER_171_464 ();
 b15zdnd11an1n04x5 FILLER_171_507 ();
 b15zdnd11an1n64x5 FILLER_171_526 ();
 b15zdnd11an1n64x5 FILLER_171_590 ();
 b15zdnd11an1n64x5 FILLER_171_654 ();
 b15zdnd11an1n16x5 FILLER_171_718 ();
 b15zdnd11an1n04x5 FILLER_171_734 ();
 b15zdnd11an1n64x5 FILLER_171_755 ();
 b15zdnd11an1n64x5 FILLER_171_819 ();
 b15zdnd00an1n01x5 FILLER_171_883 ();
 b15zdnd11an1n32x5 FILLER_171_896 ();
 b15zdnd11an1n16x5 FILLER_171_928 ();
 b15zdnd11an1n04x5 FILLER_171_944 ();
 b15zdnd11an1n64x5 FILLER_171_962 ();
 b15zdnd11an1n64x5 FILLER_171_1026 ();
 b15zdnd11an1n64x5 FILLER_171_1090 ();
 b15zdnd11an1n32x5 FILLER_171_1154 ();
 b15zdnd11an1n16x5 FILLER_171_1186 ();
 b15zdnd11an1n04x5 FILLER_171_1202 ();
 b15zdnd11an1n64x5 FILLER_171_1220 ();
 b15zdnd11an1n32x5 FILLER_171_1284 ();
 b15zdnd11an1n16x5 FILLER_171_1316 ();
 b15zdnd11an1n04x5 FILLER_171_1332 ();
 b15zdnd00an1n02x5 FILLER_171_1336 ();
 b15zdnd11an1n16x5 FILLER_171_1341 ();
 b15zdnd11an1n08x5 FILLER_171_1357 ();
 b15zdnd11an1n04x5 FILLER_171_1365 ();
 b15zdnd00an1n02x5 FILLER_171_1369 ();
 b15zdnd00an1n01x5 FILLER_171_1371 ();
 b15zdnd11an1n08x5 FILLER_171_1375 ();
 b15zdnd00an1n01x5 FILLER_171_1383 ();
 b15zdnd11an1n16x5 FILLER_171_1436 ();
 b15zdnd11an1n08x5 FILLER_171_1452 ();
 b15zdnd11an1n04x5 FILLER_171_1460 ();
 b15zdnd11an1n64x5 FILLER_171_1467 ();
 b15zdnd11an1n64x5 FILLER_171_1531 ();
 b15zdnd11an1n16x5 FILLER_171_1595 ();
 b15zdnd11an1n64x5 FILLER_171_1614 ();
 b15zdnd11an1n64x5 FILLER_171_1678 ();
 b15zdnd11an1n64x5 FILLER_171_1742 ();
 b15zdnd11an1n16x5 FILLER_171_1806 ();
 b15zdnd11an1n08x5 FILLER_171_1822 ();
 b15zdnd11an1n64x5 FILLER_171_1841 ();
 b15zdnd11an1n32x5 FILLER_171_1905 ();
 b15zdnd11an1n16x5 FILLER_171_1937 ();
 b15zdnd11an1n64x5 FILLER_171_1960 ();
 b15zdnd11an1n32x5 FILLER_171_2024 ();
 b15zdnd00an1n01x5 FILLER_171_2056 ();
 b15zdnd11an1n64x5 FILLER_171_2099 ();
 b15zdnd11an1n32x5 FILLER_171_2163 ();
 b15zdnd11an1n08x5 FILLER_171_2195 ();
 b15zdnd11an1n04x5 FILLER_171_2245 ();
 b15zdnd11an1n04x5 FILLER_171_2269 ();
 b15zdnd11an1n04x5 FILLER_171_2277 ();
 b15zdnd00an1n02x5 FILLER_171_2281 ();
 b15zdnd00an1n01x5 FILLER_171_2283 ();
 b15zdnd11an1n64x5 FILLER_172_8 ();
 b15zdnd11an1n64x5 FILLER_172_72 ();
 b15zdnd11an1n64x5 FILLER_172_136 ();
 b15zdnd11an1n16x5 FILLER_172_200 ();
 b15zdnd11an1n08x5 FILLER_172_216 ();
 b15zdnd11an1n04x5 FILLER_172_224 ();
 b15zdnd00an1n01x5 FILLER_172_228 ();
 b15zdnd11an1n64x5 FILLER_172_271 ();
 b15zdnd11an1n64x5 FILLER_172_335 ();
 b15zdnd11an1n64x5 FILLER_172_399 ();
 b15zdnd11an1n64x5 FILLER_172_463 ();
 b15zdnd11an1n64x5 FILLER_172_527 ();
 b15zdnd11an1n64x5 FILLER_172_591 ();
 b15zdnd11an1n32x5 FILLER_172_655 ();
 b15zdnd11an1n16x5 FILLER_172_687 ();
 b15zdnd11an1n08x5 FILLER_172_703 ();
 b15zdnd11an1n04x5 FILLER_172_711 ();
 b15zdnd00an1n02x5 FILLER_172_715 ();
 b15zdnd00an1n01x5 FILLER_172_717 ();
 b15zdnd11an1n32x5 FILLER_172_726 ();
 b15zdnd11an1n08x5 FILLER_172_758 ();
 b15zdnd11an1n04x5 FILLER_172_766 ();
 b15zdnd00an1n02x5 FILLER_172_770 ();
 b15zdnd11an1n64x5 FILLER_172_775 ();
 b15zdnd11an1n64x5 FILLER_172_839 ();
 b15zdnd11an1n64x5 FILLER_172_903 ();
 b15zdnd11an1n64x5 FILLER_172_967 ();
 b15zdnd11an1n64x5 FILLER_172_1031 ();
 b15zdnd11an1n64x5 FILLER_172_1095 ();
 b15zdnd11an1n64x5 FILLER_172_1159 ();
 b15zdnd11an1n64x5 FILLER_172_1223 ();
 b15zdnd11an1n32x5 FILLER_172_1287 ();
 b15zdnd11an1n16x5 FILLER_172_1319 ();
 b15zdnd00an1n02x5 FILLER_172_1335 ();
 b15zdnd00an1n01x5 FILLER_172_1337 ();
 b15zdnd11an1n04x5 FILLER_172_1341 ();
 b15zdnd11an1n32x5 FILLER_172_1348 ();
 b15zdnd11an1n16x5 FILLER_172_1380 ();
 b15zdnd11an1n08x5 FILLER_172_1396 ();
 b15zdnd11an1n64x5 FILLER_172_1407 ();
 b15zdnd11an1n32x5 FILLER_172_1471 ();
 b15zdnd11an1n08x5 FILLER_172_1503 ();
 b15zdnd11an1n04x5 FILLER_172_1511 ();
 b15zdnd11an1n64x5 FILLER_172_1529 ();
 b15zdnd11an1n64x5 FILLER_172_1593 ();
 b15zdnd11an1n64x5 FILLER_172_1657 ();
 b15zdnd11an1n64x5 FILLER_172_1721 ();
 b15zdnd11an1n64x5 FILLER_172_1785 ();
 b15zdnd11an1n64x5 FILLER_172_1849 ();
 b15zdnd11an1n64x5 FILLER_172_1913 ();
 b15zdnd11an1n64x5 FILLER_172_1977 ();
 b15zdnd11an1n16x5 FILLER_172_2041 ();
 b15zdnd11an1n08x5 FILLER_172_2057 ();
 b15zdnd00an1n02x5 FILLER_172_2065 ();
 b15zdnd00an1n01x5 FILLER_172_2067 ();
 b15zdnd11an1n32x5 FILLER_172_2110 ();
 b15zdnd11an1n08x5 FILLER_172_2142 ();
 b15zdnd11an1n04x5 FILLER_172_2150 ();
 b15zdnd11an1n64x5 FILLER_172_2162 ();
 b15zdnd11an1n04x5 FILLER_172_2226 ();
 b15zdnd00an1n02x5 FILLER_172_2230 ();
 b15zdnd00an1n02x5 FILLER_172_2274 ();
 b15zdnd11an1n08x5 FILLER_173_0 ();
 b15zdnd11an1n04x5 FILLER_173_8 ();
 b15zdnd00an1n02x5 FILLER_173_12 ();
 b15zdnd11an1n32x5 FILLER_173_28 ();
 b15zdnd11an1n16x5 FILLER_173_60 ();
 b15zdnd11an1n64x5 FILLER_173_88 ();
 b15zdnd11an1n16x5 FILLER_173_152 ();
 b15zdnd11an1n08x5 FILLER_173_168 ();
 b15zdnd00an1n01x5 FILLER_173_176 ();
 b15zdnd11an1n64x5 FILLER_173_184 ();
 b15zdnd11an1n32x5 FILLER_173_248 ();
 b15zdnd11an1n04x5 FILLER_173_280 ();
 b15zdnd11an1n64x5 FILLER_173_287 ();
 b15zdnd11an1n64x5 FILLER_173_351 ();
 b15zdnd11an1n64x5 FILLER_173_415 ();
 b15zdnd11an1n64x5 FILLER_173_479 ();
 b15zdnd11an1n64x5 FILLER_173_543 ();
 b15zdnd11an1n64x5 FILLER_173_607 ();
 b15zdnd11an1n64x5 FILLER_173_671 ();
 b15zdnd11an1n64x5 FILLER_173_735 ();
 b15zdnd11an1n64x5 FILLER_173_799 ();
 b15zdnd11an1n64x5 FILLER_173_863 ();
 b15zdnd11an1n64x5 FILLER_173_927 ();
 b15zdnd11an1n64x5 FILLER_173_991 ();
 b15zdnd11an1n64x5 FILLER_173_1055 ();
 b15zdnd11an1n08x5 FILLER_173_1119 ();
 b15zdnd11an1n04x5 FILLER_173_1127 ();
 b15zdnd11an1n64x5 FILLER_173_1143 ();
 b15zdnd11an1n08x5 FILLER_173_1207 ();
 b15zdnd11an1n04x5 FILLER_173_1215 ();
 b15zdnd11an1n64x5 FILLER_173_1237 ();
 b15zdnd11an1n08x5 FILLER_173_1301 ();
 b15zdnd11an1n04x5 FILLER_173_1309 ();
 b15zdnd00an1n02x5 FILLER_173_1313 ();
 b15zdnd11an1n64x5 FILLER_173_1367 ();
 b15zdnd11an1n64x5 FILLER_173_1431 ();
 b15zdnd11an1n64x5 FILLER_173_1495 ();
 b15zdnd11an1n32x5 FILLER_173_1559 ();
 b15zdnd00an1n02x5 FILLER_173_1591 ();
 b15zdnd11an1n16x5 FILLER_173_1604 ();
 b15zdnd11an1n08x5 FILLER_173_1620 ();
 b15zdnd00an1n02x5 FILLER_173_1628 ();
 b15zdnd11an1n64x5 FILLER_173_1646 ();
 b15zdnd11an1n64x5 FILLER_173_1710 ();
 b15zdnd11an1n64x5 FILLER_173_1774 ();
 b15zdnd11an1n64x5 FILLER_173_1838 ();
 b15zdnd11an1n64x5 FILLER_173_1902 ();
 b15zdnd11an1n64x5 FILLER_173_1966 ();
 b15zdnd11an1n64x5 FILLER_173_2030 ();
 b15zdnd11an1n64x5 FILLER_173_2094 ();
 b15zdnd11an1n32x5 FILLER_173_2158 ();
 b15zdnd11an1n08x5 FILLER_173_2190 ();
 b15zdnd00an1n02x5 FILLER_173_2198 ();
 b15zdnd00an1n01x5 FILLER_173_2200 ();
 b15zdnd11an1n16x5 FILLER_173_2204 ();
 b15zdnd11an1n08x5 FILLER_173_2220 ();
 b15zdnd11an1n04x5 FILLER_173_2228 ();
 b15zdnd11an1n04x5 FILLER_173_2236 ();
 b15zdnd00an1n02x5 FILLER_173_2282 ();
 b15zdnd11an1n64x5 FILLER_174_8 ();
 b15zdnd11an1n64x5 FILLER_174_72 ();
 b15zdnd11an1n64x5 FILLER_174_136 ();
 b15zdnd00an1n01x5 FILLER_174_200 ();
 b15zdnd11an1n64x5 FILLER_174_243 ();
 b15zdnd11an1n64x5 FILLER_174_307 ();
 b15zdnd11an1n64x5 FILLER_174_371 ();
 b15zdnd11an1n64x5 FILLER_174_435 ();
 b15zdnd11an1n16x5 FILLER_174_499 ();
 b15zdnd11an1n08x5 FILLER_174_515 ();
 b15zdnd00an1n02x5 FILLER_174_523 ();
 b15zdnd11an1n64x5 FILLER_174_542 ();
 b15zdnd11an1n16x5 FILLER_174_606 ();
 b15zdnd00an1n01x5 FILLER_174_622 ();
 b15zdnd11an1n32x5 FILLER_174_636 ();
 b15zdnd11an1n16x5 FILLER_174_668 ();
 b15zdnd11an1n08x5 FILLER_174_684 ();
 b15zdnd11an1n04x5 FILLER_174_692 ();
 b15zdnd00an1n02x5 FILLER_174_696 ();
 b15zdnd00an1n01x5 FILLER_174_698 ();
 b15zdnd00an1n02x5 FILLER_174_716 ();
 b15zdnd11an1n32x5 FILLER_174_726 ();
 b15zdnd00an1n02x5 FILLER_174_758 ();
 b15zdnd00an1n01x5 FILLER_174_760 ();
 b15zdnd11an1n16x5 FILLER_174_775 ();
 b15zdnd11an1n08x5 FILLER_174_791 ();
 b15zdnd00an1n02x5 FILLER_174_799 ();
 b15zdnd00an1n01x5 FILLER_174_801 ();
 b15zdnd11an1n32x5 FILLER_174_805 ();
 b15zdnd11an1n04x5 FILLER_174_837 ();
 b15zdnd11an1n08x5 FILLER_174_854 ();
 b15zdnd11an1n04x5 FILLER_174_862 ();
 b15zdnd00an1n02x5 FILLER_174_866 ();
 b15zdnd11an1n04x5 FILLER_174_880 ();
 b15zdnd11an1n16x5 FILLER_174_894 ();
 b15zdnd00an1n01x5 FILLER_174_910 ();
 b15zdnd11an1n08x5 FILLER_174_925 ();
 b15zdnd11an1n04x5 FILLER_174_933 ();
 b15zdnd00an1n01x5 FILLER_174_937 ();
 b15zdnd11an1n64x5 FILLER_174_946 ();
 b15zdnd11an1n16x5 FILLER_174_1010 ();
 b15zdnd11an1n08x5 FILLER_174_1026 ();
 b15zdnd11an1n04x5 FILLER_174_1034 ();
 b15zdnd00an1n02x5 FILLER_174_1038 ();
 b15zdnd11an1n32x5 FILLER_174_1056 ();
 b15zdnd11an1n16x5 FILLER_174_1088 ();
 b15zdnd11an1n08x5 FILLER_174_1104 ();
 b15zdnd11an1n64x5 FILLER_174_1116 ();
 b15zdnd11an1n64x5 FILLER_174_1180 ();
 b15zdnd11an1n64x5 FILLER_174_1244 ();
 b15zdnd11an1n64x5 FILLER_174_1308 ();
 b15zdnd11an1n64x5 FILLER_174_1372 ();
 b15zdnd11an1n64x5 FILLER_174_1436 ();
 b15zdnd11an1n64x5 FILLER_174_1500 ();
 b15zdnd11an1n64x5 FILLER_174_1564 ();
 b15zdnd11an1n16x5 FILLER_174_1628 ();
 b15zdnd11an1n04x5 FILLER_174_1644 ();
 b15zdnd00an1n02x5 FILLER_174_1648 ();
 b15zdnd11an1n08x5 FILLER_174_1692 ();
 b15zdnd11an1n04x5 FILLER_174_1700 ();
 b15zdnd00an1n02x5 FILLER_174_1704 ();
 b15zdnd00an1n01x5 FILLER_174_1706 ();
 b15zdnd11an1n64x5 FILLER_174_1721 ();
 b15zdnd11an1n64x5 FILLER_174_1785 ();
 b15zdnd11an1n32x5 FILLER_174_1849 ();
 b15zdnd11an1n08x5 FILLER_174_1881 ();
 b15zdnd11an1n04x5 FILLER_174_1889 ();
 b15zdnd00an1n02x5 FILLER_174_1893 ();
 b15zdnd11an1n04x5 FILLER_174_1898 ();
 b15zdnd11an1n64x5 FILLER_174_1905 ();
 b15zdnd11an1n64x5 FILLER_174_1969 ();
 b15zdnd11an1n32x5 FILLER_174_2033 ();
 b15zdnd11an1n16x5 FILLER_174_2065 ();
 b15zdnd11an1n04x5 FILLER_174_2081 ();
 b15zdnd00an1n02x5 FILLER_174_2085 ();
 b15zdnd11an1n32x5 FILLER_174_2101 ();
 b15zdnd11an1n16x5 FILLER_174_2133 ();
 b15zdnd11an1n04x5 FILLER_174_2149 ();
 b15zdnd00an1n01x5 FILLER_174_2153 ();
 b15zdnd11an1n08x5 FILLER_174_2162 ();
 b15zdnd00an1n01x5 FILLER_174_2170 ();
 b15zdnd11an1n08x5 FILLER_174_2213 ();
 b15zdnd00an1n02x5 FILLER_174_2221 ();
 b15zdnd00an1n01x5 FILLER_174_2223 ();
 b15zdnd11an1n04x5 FILLER_174_2228 ();
 b15zdnd00an1n02x5 FILLER_174_2274 ();
 b15zdnd11an1n64x5 FILLER_175_0 ();
 b15zdnd11an1n64x5 FILLER_175_64 ();
 b15zdnd11an1n08x5 FILLER_175_128 ();
 b15zdnd11an1n04x5 FILLER_175_136 ();
 b15zdnd00an1n02x5 FILLER_175_140 ();
 b15zdnd00an1n01x5 FILLER_175_142 ();
 b15zdnd11an1n64x5 FILLER_175_185 ();
 b15zdnd11an1n64x5 FILLER_175_249 ();
 b15zdnd11an1n64x5 FILLER_175_313 ();
 b15zdnd11an1n64x5 FILLER_175_377 ();
 b15zdnd11an1n64x5 FILLER_175_441 ();
 b15zdnd11an1n32x5 FILLER_175_505 ();
 b15zdnd11an1n08x5 FILLER_175_537 ();
 b15zdnd00an1n02x5 FILLER_175_545 ();
 b15zdnd00an1n01x5 FILLER_175_547 ();
 b15zdnd11an1n64x5 FILLER_175_551 ();
 b15zdnd11an1n64x5 FILLER_175_615 ();
 b15zdnd11an1n16x5 FILLER_175_679 ();
 b15zdnd11an1n08x5 FILLER_175_695 ();
 b15zdnd11an1n04x5 FILLER_175_703 ();
 b15zdnd00an1n01x5 FILLER_175_707 ();
 b15zdnd11an1n64x5 FILLER_175_715 ();
 b15zdnd11an1n64x5 FILLER_175_779 ();
 b15zdnd11an1n64x5 FILLER_175_843 ();
 b15zdnd11an1n64x5 FILLER_175_907 ();
 b15zdnd11an1n64x5 FILLER_175_971 ();
 b15zdnd11an1n64x5 FILLER_175_1035 ();
 b15zdnd11an1n64x5 FILLER_175_1099 ();
 b15zdnd11an1n64x5 FILLER_175_1163 ();
 b15zdnd11an1n64x5 FILLER_175_1227 ();
 b15zdnd11an1n64x5 FILLER_175_1291 ();
 b15zdnd11an1n64x5 FILLER_175_1355 ();
 b15zdnd11an1n64x5 FILLER_175_1419 ();
 b15zdnd11an1n64x5 FILLER_175_1483 ();
 b15zdnd11an1n64x5 FILLER_175_1547 ();
 b15zdnd11an1n64x5 FILLER_175_1611 ();
 b15zdnd11an1n64x5 FILLER_175_1675 ();
 b15zdnd11an1n64x5 FILLER_175_1739 ();
 b15zdnd11an1n64x5 FILLER_175_1803 ();
 b15zdnd11an1n08x5 FILLER_175_1867 ();
 b15zdnd00an1n01x5 FILLER_175_1875 ();
 b15zdnd11an1n64x5 FILLER_175_1928 ();
 b15zdnd11an1n64x5 FILLER_175_1992 ();
 b15zdnd11an1n64x5 FILLER_175_2056 ();
 b15zdnd11an1n32x5 FILLER_175_2120 ();
 b15zdnd11an1n32x5 FILLER_175_2159 ();
 b15zdnd11an1n08x5 FILLER_175_2191 ();
 b15zdnd00an1n02x5 FILLER_175_2199 ();
 b15zdnd11an1n16x5 FILLER_175_2204 ();
 b15zdnd11an1n04x5 FILLER_175_2220 ();
 b15zdnd11an1n04x5 FILLER_175_2228 ();
 b15zdnd11an1n04x5 FILLER_175_2236 ();
 b15zdnd00an1n02x5 FILLER_175_2282 ();
 b15zdnd11an1n64x5 FILLER_176_8 ();
 b15zdnd11an1n16x5 FILLER_176_72 ();
 b15zdnd11an1n08x5 FILLER_176_88 ();
 b15zdnd11an1n04x5 FILLER_176_96 ();
 b15zdnd00an1n02x5 FILLER_176_100 ();
 b15zdnd00an1n01x5 FILLER_176_102 ();
 b15zdnd11an1n04x5 FILLER_176_145 ();
 b15zdnd11an1n64x5 FILLER_176_191 ();
 b15zdnd11an1n64x5 FILLER_176_255 ();
 b15zdnd11an1n64x5 FILLER_176_319 ();
 b15zdnd11an1n64x5 FILLER_176_383 ();
 b15zdnd11an1n64x5 FILLER_176_447 ();
 b15zdnd11an1n04x5 FILLER_176_511 ();
 b15zdnd11an1n08x5 FILLER_176_518 ();
 b15zdnd00an1n01x5 FILLER_176_526 ();
 b15zdnd11an1n04x5 FILLER_176_534 ();
 b15zdnd11an1n64x5 FILLER_176_552 ();
 b15zdnd00an1n02x5 FILLER_176_616 ();
 b15zdnd00an1n01x5 FILLER_176_618 ();
 b15zdnd11an1n64x5 FILLER_176_635 ();
 b15zdnd11an1n16x5 FILLER_176_699 ();
 b15zdnd00an1n02x5 FILLER_176_715 ();
 b15zdnd00an1n01x5 FILLER_176_717 ();
 b15zdnd11an1n64x5 FILLER_176_726 ();
 b15zdnd11an1n32x5 FILLER_176_790 ();
 b15zdnd11an1n08x5 FILLER_176_822 ();
 b15zdnd11an1n04x5 FILLER_176_830 ();
 b15zdnd00an1n01x5 FILLER_176_834 ();
 b15zdnd11an1n64x5 FILLER_176_851 ();
 b15zdnd11an1n64x5 FILLER_176_915 ();
 b15zdnd11an1n16x5 FILLER_176_979 ();
 b15zdnd11an1n04x5 FILLER_176_995 ();
 b15zdnd00an1n02x5 FILLER_176_999 ();
 b15zdnd00an1n01x5 FILLER_176_1001 ();
 b15zdnd11an1n04x5 FILLER_176_1022 ();
 b15zdnd00an1n02x5 FILLER_176_1026 ();
 b15zdnd00an1n01x5 FILLER_176_1028 ();
 b15zdnd11an1n64x5 FILLER_176_1043 ();
 b15zdnd11an1n64x5 FILLER_176_1107 ();
 b15zdnd11an1n64x5 FILLER_176_1171 ();
 b15zdnd11an1n32x5 FILLER_176_1235 ();
 b15zdnd00an1n01x5 FILLER_176_1267 ();
 b15zdnd11an1n64x5 FILLER_176_1280 ();
 b15zdnd11an1n32x5 FILLER_176_1344 ();
 b15zdnd00an1n02x5 FILLER_176_1376 ();
 b15zdnd00an1n01x5 FILLER_176_1378 ();
 b15zdnd11an1n64x5 FILLER_176_1395 ();
 b15zdnd11an1n64x5 FILLER_176_1459 ();
 b15zdnd11an1n64x5 FILLER_176_1523 ();
 b15zdnd11an1n64x5 FILLER_176_1587 ();
 b15zdnd11an1n64x5 FILLER_176_1651 ();
 b15zdnd00an1n02x5 FILLER_176_1715 ();
 b15zdnd00an1n01x5 FILLER_176_1717 ();
 b15zdnd11an1n04x5 FILLER_176_1732 ();
 b15zdnd00an1n01x5 FILLER_176_1736 ();
 b15zdnd11an1n32x5 FILLER_176_1740 ();
 b15zdnd11an1n08x5 FILLER_176_1772 ();
 b15zdnd11an1n04x5 FILLER_176_1780 ();
 b15zdnd00an1n01x5 FILLER_176_1784 ();
 b15zdnd11an1n64x5 FILLER_176_1798 ();
 b15zdnd00an1n01x5 FILLER_176_1862 ();
 b15zdnd11an1n04x5 FILLER_176_1870 ();
 b15zdnd11an1n04x5 FILLER_176_1894 ();
 b15zdnd11an1n08x5 FILLER_176_1901 ();
 b15zdnd11an1n64x5 FILLER_176_1915 ();
 b15zdnd11an1n64x5 FILLER_176_1979 ();
 b15zdnd11an1n32x5 FILLER_176_2043 ();
 b15zdnd11an1n16x5 FILLER_176_2075 ();
 b15zdnd11an1n08x5 FILLER_176_2091 ();
 b15zdnd11an1n04x5 FILLER_176_2099 ();
 b15zdnd00an1n01x5 FILLER_176_2103 ();
 b15zdnd11an1n16x5 FILLER_176_2124 ();
 b15zdnd11an1n08x5 FILLER_176_2140 ();
 b15zdnd11an1n04x5 FILLER_176_2148 ();
 b15zdnd00an1n02x5 FILLER_176_2152 ();
 b15zdnd11an1n08x5 FILLER_176_2162 ();
 b15zdnd11an1n04x5 FILLER_176_2170 ();
 b15zdnd00an1n02x5 FILLER_176_2174 ();
 b15zdnd11an1n04x5 FILLER_176_2228 ();
 b15zdnd00an1n02x5 FILLER_176_2274 ();
 b15zdnd11an1n08x5 FILLER_177_0 ();
 b15zdnd00an1n02x5 FILLER_177_8 ();
 b15zdnd11an1n08x5 FILLER_177_14 ();
 b15zdnd11an1n04x5 FILLER_177_22 ();
 b15zdnd11an1n04x5 FILLER_177_30 ();
 b15zdnd11an1n64x5 FILLER_177_38 ();
 b15zdnd11an1n16x5 FILLER_177_102 ();
 b15zdnd00an1n01x5 FILLER_177_118 ();
 b15zdnd11an1n32x5 FILLER_177_161 ();
 b15zdnd11an1n04x5 FILLER_177_193 ();
 b15zdnd00an1n02x5 FILLER_177_197 ();
 b15zdnd00an1n01x5 FILLER_177_199 ();
 b15zdnd11an1n64x5 FILLER_177_217 ();
 b15zdnd11an1n64x5 FILLER_177_281 ();
 b15zdnd11an1n64x5 FILLER_177_345 ();
 b15zdnd11an1n32x5 FILLER_177_409 ();
 b15zdnd11an1n16x5 FILLER_177_441 ();
 b15zdnd11an1n08x5 FILLER_177_457 ();
 b15zdnd00an1n01x5 FILLER_177_465 ();
 b15zdnd11an1n64x5 FILLER_177_481 ();
 b15zdnd11an1n64x5 FILLER_177_545 ();
 b15zdnd11an1n64x5 FILLER_177_609 ();
 b15zdnd11an1n64x5 FILLER_177_673 ();
 b15zdnd11an1n64x5 FILLER_177_737 ();
 b15zdnd11an1n64x5 FILLER_177_801 ();
 b15zdnd11an1n64x5 FILLER_177_865 ();
 b15zdnd11an1n08x5 FILLER_177_929 ();
 b15zdnd11an1n04x5 FILLER_177_937 ();
 b15zdnd11an1n64x5 FILLER_177_955 ();
 b15zdnd11an1n64x5 FILLER_177_1019 ();
 b15zdnd11an1n64x5 FILLER_177_1083 ();
 b15zdnd11an1n64x5 FILLER_177_1147 ();
 b15zdnd11an1n32x5 FILLER_177_1211 ();
 b15zdnd11an1n32x5 FILLER_177_1259 ();
 b15zdnd11an1n16x5 FILLER_177_1333 ();
 b15zdnd11an1n04x5 FILLER_177_1349 ();
 b15zdnd00an1n02x5 FILLER_177_1353 ();
 b15zdnd11an1n64x5 FILLER_177_1397 ();
 b15zdnd11an1n64x5 FILLER_177_1461 ();
 b15zdnd11an1n16x5 FILLER_177_1525 ();
 b15zdnd11an1n08x5 FILLER_177_1541 ();
 b15zdnd11an1n04x5 FILLER_177_1549 ();
 b15zdnd00an1n02x5 FILLER_177_1553 ();
 b15zdnd11an1n04x5 FILLER_177_1569 ();
 b15zdnd11an1n64x5 FILLER_177_1587 ();
 b15zdnd11an1n64x5 FILLER_177_1651 ();
 b15zdnd11an1n04x5 FILLER_177_1715 ();
 b15zdnd00an1n02x5 FILLER_177_1719 ();
 b15zdnd00an1n01x5 FILLER_177_1721 ();
 b15zdnd11an1n04x5 FILLER_177_1735 ();
 b15zdnd00an1n02x5 FILLER_177_1739 ();
 b15zdnd00an1n01x5 FILLER_177_1741 ();
 b15zdnd11an1n08x5 FILLER_177_1745 ();
 b15zdnd11an1n04x5 FILLER_177_1753 ();
 b15zdnd00an1n02x5 FILLER_177_1757 ();
 b15zdnd00an1n01x5 FILLER_177_1759 ();
 b15zdnd11an1n64x5 FILLER_177_1766 ();
 b15zdnd11an1n64x5 FILLER_177_1830 ();
 b15zdnd11an1n04x5 FILLER_177_1894 ();
 b15zdnd11an1n04x5 FILLER_177_1918 ();
 b15zdnd11an1n04x5 FILLER_177_1934 ();
 b15zdnd00an1n01x5 FILLER_177_1938 ();
 b15zdnd11an1n64x5 FILLER_177_1951 ();
 b15zdnd11an1n64x5 FILLER_177_2015 ();
 b15zdnd11an1n64x5 FILLER_177_2079 ();
 b15zdnd11an1n32x5 FILLER_177_2143 ();
 b15zdnd11an1n16x5 FILLER_177_2175 ();
 b15zdnd11an1n08x5 FILLER_177_2191 ();
 b15zdnd00an1n02x5 FILLER_177_2199 ();
 b15zdnd00an1n01x5 FILLER_177_2201 ();
 b15zdnd11an1n32x5 FILLER_177_2205 ();
 b15zdnd00an1n02x5 FILLER_177_2237 ();
 b15zdnd00an1n01x5 FILLER_177_2239 ();
 b15zdnd00an1n02x5 FILLER_177_2282 ();
 b15zdnd00an1n02x5 FILLER_178_8 ();
 b15zdnd11an1n64x5 FILLER_178_52 ();
 b15zdnd11an1n16x5 FILLER_178_116 ();
 b15zdnd11an1n08x5 FILLER_178_132 ();
 b15zdnd11an1n04x5 FILLER_178_140 ();
 b15zdnd11an1n32x5 FILLER_178_148 ();
 b15zdnd11an1n16x5 FILLER_178_180 ();
 b15zdnd11an1n08x5 FILLER_178_196 ();
 b15zdnd00an1n02x5 FILLER_178_204 ();
 b15zdnd11an1n08x5 FILLER_178_225 ();
 b15zdnd11an1n04x5 FILLER_178_233 ();
 b15zdnd00an1n02x5 FILLER_178_237 ();
 b15zdnd00an1n01x5 FILLER_178_239 ();
 b15zdnd11an1n64x5 FILLER_178_245 ();
 b15zdnd11an1n64x5 FILLER_178_309 ();
 b15zdnd11an1n64x5 FILLER_178_373 ();
 b15zdnd11an1n64x5 FILLER_178_437 ();
 b15zdnd11an1n64x5 FILLER_178_501 ();
 b15zdnd11an1n64x5 FILLER_178_565 ();
 b15zdnd11an1n64x5 FILLER_178_629 ();
 b15zdnd11an1n16x5 FILLER_178_693 ();
 b15zdnd11an1n08x5 FILLER_178_709 ();
 b15zdnd00an1n01x5 FILLER_178_717 ();
 b15zdnd11an1n64x5 FILLER_178_726 ();
 b15zdnd11an1n64x5 FILLER_178_790 ();
 b15zdnd11an1n08x5 FILLER_178_854 ();
 b15zdnd11an1n04x5 FILLER_178_874 ();
 b15zdnd00an1n01x5 FILLER_178_878 ();
 b15zdnd11an1n64x5 FILLER_178_887 ();
 b15zdnd11an1n08x5 FILLER_178_951 ();
 b15zdnd00an1n01x5 FILLER_178_959 ();
 b15zdnd11an1n64x5 FILLER_178_981 ();
 b15zdnd11an1n64x5 FILLER_178_1045 ();
 b15zdnd11an1n64x5 FILLER_178_1109 ();
 b15zdnd11an1n64x5 FILLER_178_1173 ();
 b15zdnd11an1n64x5 FILLER_178_1237 ();
 b15zdnd11an1n64x5 FILLER_178_1301 ();
 b15zdnd11an1n64x5 FILLER_178_1365 ();
 b15zdnd11an1n64x5 FILLER_178_1429 ();
 b15zdnd11an1n64x5 FILLER_178_1493 ();
 b15zdnd11an1n64x5 FILLER_178_1557 ();
 b15zdnd11an1n32x5 FILLER_178_1621 ();
 b15zdnd11an1n08x5 FILLER_178_1653 ();
 b15zdnd00an1n01x5 FILLER_178_1661 ();
 b15zdnd11an1n16x5 FILLER_178_1674 ();
 b15zdnd11an1n08x5 FILLER_178_1690 ();
 b15zdnd00an1n02x5 FILLER_178_1698 ();
 b15zdnd11an1n64x5 FILLER_178_1744 ();
 b15zdnd11an1n64x5 FILLER_178_1808 ();
 b15zdnd11an1n32x5 FILLER_178_1872 ();
 b15zdnd11an1n08x5 FILLER_178_1904 ();
 b15zdnd00an1n02x5 FILLER_178_1912 ();
 b15zdnd11an1n64x5 FILLER_178_1921 ();
 b15zdnd11an1n64x5 FILLER_178_1985 ();
 b15zdnd11an1n64x5 FILLER_178_2049 ();
 b15zdnd11an1n32x5 FILLER_178_2113 ();
 b15zdnd11an1n08x5 FILLER_178_2145 ();
 b15zdnd00an1n01x5 FILLER_178_2153 ();
 b15zdnd11an1n64x5 FILLER_178_2162 ();
 b15zdnd11an1n08x5 FILLER_178_2226 ();
 b15zdnd11an1n04x5 FILLER_178_2234 ();
 b15zdnd11an1n04x5 FILLER_178_2246 ();
 b15zdnd11an1n04x5 FILLER_178_2264 ();
 b15zdnd00an1n02x5 FILLER_178_2273 ();
 b15zdnd00an1n01x5 FILLER_178_2275 ();
 b15zdnd11an1n08x5 FILLER_179_0 ();
 b15zdnd11an1n04x5 FILLER_179_8 ();
 b15zdnd00an1n01x5 FILLER_179_12 ();
 b15zdnd11an1n64x5 FILLER_179_55 ();
 b15zdnd11an1n32x5 FILLER_179_119 ();
 b15zdnd11an1n16x5 FILLER_179_151 ();
 b15zdnd00an1n02x5 FILLER_179_167 ();
 b15zdnd00an1n01x5 FILLER_179_169 ();
 b15zdnd11an1n64x5 FILLER_179_174 ();
 b15zdnd11an1n08x5 FILLER_179_238 ();
 b15zdnd11an1n04x5 FILLER_179_246 ();
 b15zdnd00an1n01x5 FILLER_179_250 ();
 b15zdnd11an1n64x5 FILLER_179_258 ();
 b15zdnd11an1n64x5 FILLER_179_322 ();
 b15zdnd11an1n64x5 FILLER_179_386 ();
 b15zdnd11an1n64x5 FILLER_179_450 ();
 b15zdnd11an1n64x5 FILLER_179_514 ();
 b15zdnd11an1n64x5 FILLER_179_578 ();
 b15zdnd11an1n16x5 FILLER_179_642 ();
 b15zdnd11an1n04x5 FILLER_179_658 ();
 b15zdnd00an1n02x5 FILLER_179_662 ();
 b15zdnd11an1n64x5 FILLER_179_690 ();
 b15zdnd11an1n08x5 FILLER_179_754 ();
 b15zdnd11an1n64x5 FILLER_179_782 ();
 b15zdnd11an1n16x5 FILLER_179_846 ();
 b15zdnd11an1n08x5 FILLER_179_862 ();
 b15zdnd11an1n04x5 FILLER_179_870 ();
 b15zdnd00an1n01x5 FILLER_179_874 ();
 b15zdnd11an1n64x5 FILLER_179_895 ();
 b15zdnd11an1n32x5 FILLER_179_959 ();
 b15zdnd11an1n08x5 FILLER_179_991 ();
 b15zdnd11an1n04x5 FILLER_179_999 ();
 b15zdnd00an1n02x5 FILLER_179_1003 ();
 b15zdnd00an1n01x5 FILLER_179_1005 ();
 b15zdnd11an1n04x5 FILLER_179_1020 ();
 b15zdnd00an1n02x5 FILLER_179_1024 ();
 b15zdnd00an1n01x5 FILLER_179_1026 ();
 b15zdnd11an1n64x5 FILLER_179_1040 ();
 b15zdnd11an1n64x5 FILLER_179_1104 ();
 b15zdnd11an1n64x5 FILLER_179_1168 ();
 b15zdnd11an1n64x5 FILLER_179_1232 ();
 b15zdnd11an1n16x5 FILLER_179_1296 ();
 b15zdnd11an1n08x5 FILLER_179_1312 ();
 b15zdnd00an1n01x5 FILLER_179_1320 ();
 b15zdnd11an1n64x5 FILLER_179_1363 ();
 b15zdnd11an1n64x5 FILLER_179_1427 ();
 b15zdnd11an1n08x5 FILLER_179_1491 ();
 b15zdnd00an1n02x5 FILLER_179_1499 ();
 b15zdnd00an1n01x5 FILLER_179_1501 ();
 b15zdnd11an1n64x5 FILLER_179_1515 ();
 b15zdnd11an1n08x5 FILLER_179_1579 ();
 b15zdnd11an1n04x5 FILLER_179_1587 ();
 b15zdnd11an1n64x5 FILLER_179_1611 ();
 b15zdnd11an1n32x5 FILLER_179_1675 ();
 b15zdnd11an1n64x5 FILLER_179_1749 ();
 b15zdnd11an1n64x5 FILLER_179_1813 ();
 b15zdnd11an1n64x5 FILLER_179_1877 ();
 b15zdnd11an1n64x5 FILLER_179_1941 ();
 b15zdnd11an1n32x5 FILLER_179_2005 ();
 b15zdnd11an1n16x5 FILLER_179_2037 ();
 b15zdnd11an1n04x5 FILLER_179_2053 ();
 b15zdnd00an1n01x5 FILLER_179_2057 ();
 b15zdnd11an1n04x5 FILLER_179_2100 ();
 b15zdnd11an1n64x5 FILLER_179_2124 ();
 b15zdnd11an1n16x5 FILLER_179_2188 ();
 b15zdnd11an1n08x5 FILLER_179_2204 ();
 b15zdnd11an1n04x5 FILLER_179_2212 ();
 b15zdnd00an1n02x5 FILLER_179_2216 ();
 b15zdnd00an1n01x5 FILLER_179_2218 ();
 b15zdnd11an1n04x5 FILLER_179_2261 ();
 b15zdnd11an1n04x5 FILLER_179_2277 ();
 b15zdnd00an1n02x5 FILLER_179_2281 ();
 b15zdnd00an1n01x5 FILLER_179_2283 ();
 b15zdnd00an1n02x5 FILLER_180_8 ();
 b15zdnd11an1n64x5 FILLER_180_52 ();
 b15zdnd11an1n64x5 FILLER_180_116 ();
 b15zdnd11an1n16x5 FILLER_180_180 ();
 b15zdnd11an1n08x5 FILLER_180_196 ();
 b15zdnd00an1n02x5 FILLER_180_204 ();
 b15zdnd11an1n08x5 FILLER_180_216 ();
 b15zdnd11an1n04x5 FILLER_180_224 ();
 b15zdnd11an1n64x5 FILLER_180_234 ();
 b15zdnd11an1n64x5 FILLER_180_298 ();
 b15zdnd11an1n64x5 FILLER_180_362 ();
 b15zdnd11an1n64x5 FILLER_180_426 ();
 b15zdnd11an1n64x5 FILLER_180_490 ();
 b15zdnd00an1n01x5 FILLER_180_554 ();
 b15zdnd11an1n64x5 FILLER_180_558 ();
 b15zdnd11an1n64x5 FILLER_180_622 ();
 b15zdnd11an1n32x5 FILLER_180_686 ();
 b15zdnd11an1n64x5 FILLER_180_726 ();
 b15zdnd11an1n64x5 FILLER_180_790 ();
 b15zdnd11an1n04x5 FILLER_180_854 ();
 b15zdnd11an1n08x5 FILLER_180_865 ();
 b15zdnd00an1n01x5 FILLER_180_873 ();
 b15zdnd11an1n32x5 FILLER_180_888 ();
 b15zdnd11an1n16x5 FILLER_180_920 ();
 b15zdnd00an1n02x5 FILLER_180_936 ();
 b15zdnd00an1n01x5 FILLER_180_938 ();
 b15zdnd11an1n64x5 FILLER_180_956 ();
 b15zdnd00an1n01x5 FILLER_180_1020 ();
 b15zdnd11an1n04x5 FILLER_180_1024 ();
 b15zdnd11an1n04x5 FILLER_180_1042 ();
 b15zdnd11an1n08x5 FILLER_180_1063 ();
 b15zdnd11an1n04x5 FILLER_180_1071 ();
 b15zdnd00an1n02x5 FILLER_180_1075 ();
 b15zdnd00an1n01x5 FILLER_180_1077 ();
 b15zdnd11an1n32x5 FILLER_180_1102 ();
 b15zdnd11an1n08x5 FILLER_180_1134 ();
 b15zdnd00an1n02x5 FILLER_180_1142 ();
 b15zdnd00an1n01x5 FILLER_180_1144 ();
 b15zdnd11an1n64x5 FILLER_180_1159 ();
 b15zdnd11an1n32x5 FILLER_180_1223 ();
 b15zdnd11an1n64x5 FILLER_180_1269 ();
 b15zdnd00an1n01x5 FILLER_180_1333 ();
 b15zdnd11an1n64x5 FILLER_180_1345 ();
 b15zdnd11an1n32x5 FILLER_180_1409 ();
 b15zdnd11an1n16x5 FILLER_180_1441 ();
 b15zdnd11an1n08x5 FILLER_180_1457 ();
 b15zdnd00an1n02x5 FILLER_180_1465 ();
 b15zdnd11an1n64x5 FILLER_180_1481 ();
 b15zdnd11an1n64x5 FILLER_180_1545 ();
 b15zdnd11an1n64x5 FILLER_180_1609 ();
 b15zdnd11an1n16x5 FILLER_180_1673 ();
 b15zdnd11an1n08x5 FILLER_180_1689 ();
 b15zdnd00an1n01x5 FILLER_180_1697 ();
 b15zdnd11an1n04x5 FILLER_180_1714 ();
 b15zdnd11an1n04x5 FILLER_180_1721 ();
 b15zdnd00an1n01x5 FILLER_180_1725 ();
 b15zdnd11an1n04x5 FILLER_180_1736 ();
 b15zdnd11an1n64x5 FILLER_180_1752 ();
 b15zdnd11an1n64x5 FILLER_180_1816 ();
 b15zdnd11an1n64x5 FILLER_180_1880 ();
 b15zdnd11an1n64x5 FILLER_180_1944 ();
 b15zdnd11an1n64x5 FILLER_180_2008 ();
 b15zdnd11an1n16x5 FILLER_180_2072 ();
 b15zdnd11an1n04x5 FILLER_180_2088 ();
 b15zdnd11an1n16x5 FILLER_180_2134 ();
 b15zdnd11an1n04x5 FILLER_180_2150 ();
 b15zdnd11an1n64x5 FILLER_180_2162 ();
 b15zdnd11an1n04x5 FILLER_180_2226 ();
 b15zdnd00an1n02x5 FILLER_180_2230 ();
 b15zdnd00an1n02x5 FILLER_180_2274 ();
 b15zdnd11an1n64x5 FILLER_181_0 ();
 b15zdnd11an1n08x5 FILLER_181_64 ();
 b15zdnd00an1n02x5 FILLER_181_72 ();
 b15zdnd00an1n01x5 FILLER_181_74 ();
 b15zdnd11an1n64x5 FILLER_181_114 ();
 b15zdnd11an1n16x5 FILLER_181_178 ();
 b15zdnd11an1n08x5 FILLER_181_194 ();
 b15zdnd11an1n04x5 FILLER_181_202 ();
 b15zdnd11an1n32x5 FILLER_181_225 ();
 b15zdnd11an1n08x5 FILLER_181_257 ();
 b15zdnd11an1n64x5 FILLER_181_268 ();
 b15zdnd11an1n64x5 FILLER_181_332 ();
 b15zdnd11an1n64x5 FILLER_181_396 ();
 b15zdnd11an1n64x5 FILLER_181_460 ();
 b15zdnd11an1n04x5 FILLER_181_524 ();
 b15zdnd00an1n02x5 FILLER_181_528 ();
 b15zdnd00an1n01x5 FILLER_181_530 ();
 b15zdnd11an1n64x5 FILLER_181_575 ();
 b15zdnd11an1n32x5 FILLER_181_639 ();
 b15zdnd11an1n16x5 FILLER_181_671 ();
 b15zdnd11an1n04x5 FILLER_181_687 ();
 b15zdnd00an1n01x5 FILLER_181_691 ();
 b15zdnd11an1n16x5 FILLER_181_706 ();
 b15zdnd11an1n08x5 FILLER_181_722 ();
 b15zdnd00an1n01x5 FILLER_181_730 ();
 b15zdnd11an1n16x5 FILLER_181_747 ();
 b15zdnd11an1n04x5 FILLER_181_763 ();
 b15zdnd00an1n02x5 FILLER_181_767 ();
 b15zdnd11an1n64x5 FILLER_181_790 ();
 b15zdnd11an1n16x5 FILLER_181_854 ();
 b15zdnd11an1n08x5 FILLER_181_870 ();
 b15zdnd11an1n04x5 FILLER_181_878 ();
 b15zdnd00an1n02x5 FILLER_181_882 ();
 b15zdnd00an1n01x5 FILLER_181_884 ();
 b15zdnd11an1n64x5 FILLER_181_888 ();
 b15zdnd11an1n32x5 FILLER_181_952 ();
 b15zdnd11an1n04x5 FILLER_181_984 ();
 b15zdnd11an1n16x5 FILLER_181_1006 ();
 b15zdnd00an1n01x5 FILLER_181_1022 ();
 b15zdnd11an1n04x5 FILLER_181_1065 ();
 b15zdnd11an1n64x5 FILLER_181_1085 ();
 b15zdnd11an1n32x5 FILLER_181_1149 ();
 b15zdnd11an1n08x5 FILLER_181_1181 ();
 b15zdnd11an1n04x5 FILLER_181_1189 ();
 b15zdnd11an1n08x5 FILLER_181_1207 ();
 b15zdnd00an1n02x5 FILLER_181_1215 ();
 b15zdnd11an1n08x5 FILLER_181_1225 ();
 b15zdnd11an1n04x5 FILLER_181_1233 ();
 b15zdnd00an1n02x5 FILLER_181_1237 ();
 b15zdnd00an1n01x5 FILLER_181_1239 ();
 b15zdnd11an1n08x5 FILLER_181_1247 ();
 b15zdnd00an1n02x5 FILLER_181_1255 ();
 b15zdnd00an1n01x5 FILLER_181_1257 ();
 b15zdnd11an1n64x5 FILLER_181_1267 ();
 b15zdnd11an1n64x5 FILLER_181_1331 ();
 b15zdnd11an1n64x5 FILLER_181_1395 ();
 b15zdnd11an1n64x5 FILLER_181_1459 ();
 b15zdnd11an1n64x5 FILLER_181_1523 ();
 b15zdnd11an1n64x5 FILLER_181_1587 ();
 b15zdnd11an1n64x5 FILLER_181_1651 ();
 b15zdnd11an1n04x5 FILLER_181_1715 ();
 b15zdnd00an1n02x5 FILLER_181_1719 ();
 b15zdnd00an1n01x5 FILLER_181_1721 ();
 b15zdnd11an1n04x5 FILLER_181_1725 ();
 b15zdnd11an1n64x5 FILLER_181_1732 ();
 b15zdnd11an1n64x5 FILLER_181_1796 ();
 b15zdnd11an1n64x5 FILLER_181_1860 ();
 b15zdnd11an1n64x5 FILLER_181_1924 ();
 b15zdnd11an1n64x5 FILLER_181_1988 ();
 b15zdnd11an1n32x5 FILLER_181_2052 ();
 b15zdnd11an1n04x5 FILLER_181_2084 ();
 b15zdnd00an1n02x5 FILLER_181_2088 ();
 b15zdnd11an1n64x5 FILLER_181_2093 ();
 b15zdnd11an1n08x5 FILLER_181_2157 ();
 b15zdnd11an1n64x5 FILLER_181_2173 ();
 b15zdnd00an1n02x5 FILLER_181_2237 ();
 b15zdnd00an1n01x5 FILLER_181_2239 ();
 b15zdnd00an1n02x5 FILLER_181_2282 ();
 b15zdnd11an1n08x5 FILLER_182_8 ();
 b15zdnd11an1n04x5 FILLER_182_16 ();
 b15zdnd00an1n01x5 FILLER_182_20 ();
 b15zdnd11an1n16x5 FILLER_182_38 ();
 b15zdnd11an1n08x5 FILLER_182_54 ();
 b15zdnd11an1n04x5 FILLER_182_62 ();
 b15zdnd11an1n64x5 FILLER_182_103 ();
 b15zdnd11an1n16x5 FILLER_182_167 ();
 b15zdnd11an1n08x5 FILLER_182_183 ();
 b15zdnd00an1n02x5 FILLER_182_191 ();
 b15zdnd00an1n01x5 FILLER_182_193 ();
 b15zdnd11an1n04x5 FILLER_182_214 ();
 b15zdnd11an1n16x5 FILLER_182_237 ();
 b15zdnd11an1n08x5 FILLER_182_253 ();
 b15zdnd00an1n02x5 FILLER_182_261 ();
 b15zdnd11an1n08x5 FILLER_182_266 ();
 b15zdnd00an1n01x5 FILLER_182_274 ();
 b15zdnd11an1n64x5 FILLER_182_278 ();
 b15zdnd11an1n04x5 FILLER_182_342 ();
 b15zdnd00an1n01x5 FILLER_182_346 ();
 b15zdnd11an1n64x5 FILLER_182_359 ();
 b15zdnd11an1n64x5 FILLER_182_423 ();
 b15zdnd11an1n64x5 FILLER_182_487 ();
 b15zdnd00an1n02x5 FILLER_182_551 ();
 b15zdnd00an1n01x5 FILLER_182_553 ();
 b15zdnd11an1n32x5 FILLER_182_557 ();
 b15zdnd11an1n16x5 FILLER_182_589 ();
 b15zdnd11an1n08x5 FILLER_182_605 ();
 b15zdnd11an1n04x5 FILLER_182_613 ();
 b15zdnd00an1n02x5 FILLER_182_617 ();
 b15zdnd00an1n01x5 FILLER_182_619 ();
 b15zdnd11an1n04x5 FILLER_182_664 ();
 b15zdnd11an1n04x5 FILLER_182_699 ();
 b15zdnd11an1n04x5 FILLER_182_706 ();
 b15zdnd11an1n04x5 FILLER_182_713 ();
 b15zdnd00an1n01x5 FILLER_182_717 ();
 b15zdnd11an1n04x5 FILLER_182_726 ();
 b15zdnd00an1n02x5 FILLER_182_730 ();
 b15zdnd00an1n01x5 FILLER_182_732 ();
 b15zdnd11an1n64x5 FILLER_182_746 ();
 b15zdnd11an1n64x5 FILLER_182_810 ();
 b15zdnd11an1n64x5 FILLER_182_874 ();
 b15zdnd11an1n64x5 FILLER_182_938 ();
 b15zdnd11an1n64x5 FILLER_182_1002 ();
 b15zdnd11an1n16x5 FILLER_182_1066 ();
 b15zdnd11an1n08x5 FILLER_182_1082 ();
 b15zdnd11an1n64x5 FILLER_182_1110 ();
 b15zdnd11an1n64x5 FILLER_182_1174 ();
 b15zdnd11an1n08x5 FILLER_182_1238 ();
 b15zdnd11an1n04x5 FILLER_182_1246 ();
 b15zdnd00an1n01x5 FILLER_182_1250 ();
 b15zdnd11an1n64x5 FILLER_182_1273 ();
 b15zdnd11an1n64x5 FILLER_182_1337 ();
 b15zdnd11an1n64x5 FILLER_182_1401 ();
 b15zdnd11an1n64x5 FILLER_182_1465 ();
 b15zdnd11an1n64x5 FILLER_182_1529 ();
 b15zdnd11an1n64x5 FILLER_182_1593 ();
 b15zdnd11an1n64x5 FILLER_182_1657 ();
 b15zdnd11an1n64x5 FILLER_182_1721 ();
 b15zdnd11an1n64x5 FILLER_182_1785 ();
 b15zdnd11an1n64x5 FILLER_182_1849 ();
 b15zdnd11an1n64x5 FILLER_182_1913 ();
 b15zdnd11an1n08x5 FILLER_182_1977 ();
 b15zdnd11an1n04x5 FILLER_182_1985 ();
 b15zdnd00an1n02x5 FILLER_182_1989 ();
 b15zdnd00an1n01x5 FILLER_182_1991 ();
 b15zdnd11an1n32x5 FILLER_182_2008 ();
 b15zdnd11an1n16x5 FILLER_182_2040 ();
 b15zdnd11an1n08x5 FILLER_182_2056 ();
 b15zdnd11an1n32x5 FILLER_182_2116 ();
 b15zdnd11an1n04x5 FILLER_182_2148 ();
 b15zdnd00an1n02x5 FILLER_182_2152 ();
 b15zdnd00an1n02x5 FILLER_182_2162 ();
 b15zdnd00an1n01x5 FILLER_182_2164 ();
 b15zdnd11an1n32x5 FILLER_182_2172 ();
 b15zdnd11an1n04x5 FILLER_182_2204 ();
 b15zdnd00an1n02x5 FILLER_182_2208 ();
 b15zdnd00an1n01x5 FILLER_182_2210 ();
 b15zdnd11an1n08x5 FILLER_182_2223 ();
 b15zdnd11an1n04x5 FILLER_182_2235 ();
 b15zdnd11an1n04x5 FILLER_182_2244 ();
 b15zdnd00an1n02x5 FILLER_182_2248 ();
 b15zdnd00an1n01x5 FILLER_182_2250 ();
 b15zdnd11an1n04x5 FILLER_182_2255 ();
 b15zdnd11an1n08x5 FILLER_182_2266 ();
 b15zdnd00an1n02x5 FILLER_182_2274 ();
 b15zdnd11an1n64x5 FILLER_183_0 ();
 b15zdnd11an1n64x5 FILLER_183_64 ();
 b15zdnd11an1n32x5 FILLER_183_128 ();
 b15zdnd11an1n16x5 FILLER_183_160 ();
 b15zdnd11an1n08x5 FILLER_183_176 ();
 b15zdnd11an1n04x5 FILLER_183_184 ();
 b15zdnd00an1n02x5 FILLER_183_188 ();
 b15zdnd00an1n01x5 FILLER_183_190 ();
 b15zdnd11an1n04x5 FILLER_183_201 ();
 b15zdnd11an1n16x5 FILLER_183_221 ();
 b15zdnd00an1n02x5 FILLER_183_237 ();
 b15zdnd00an1n01x5 FILLER_183_239 ();
 b15zdnd11an1n64x5 FILLER_183_292 ();
 b15zdnd11an1n64x5 FILLER_183_356 ();
 b15zdnd11an1n64x5 FILLER_183_420 ();
 b15zdnd11an1n64x5 FILLER_183_484 ();
 b15zdnd11an1n04x5 FILLER_183_548 ();
 b15zdnd11an1n64x5 FILLER_183_555 ();
 b15zdnd11an1n16x5 FILLER_183_619 ();
 b15zdnd00an1n02x5 FILLER_183_635 ();
 b15zdnd00an1n01x5 FILLER_183_637 ();
 b15zdnd11an1n04x5 FILLER_183_641 ();
 b15zdnd11an1n16x5 FILLER_183_648 ();
 b15zdnd00an1n02x5 FILLER_183_664 ();
 b15zdnd00an1n01x5 FILLER_183_666 ();
 b15zdnd11an1n04x5 FILLER_183_681 ();
 b15zdnd00an1n02x5 FILLER_183_685 ();
 b15zdnd00an1n01x5 FILLER_183_687 ();
 b15zdnd11an1n64x5 FILLER_183_730 ();
 b15zdnd11an1n64x5 FILLER_183_803 ();
 b15zdnd11an1n08x5 FILLER_183_867 ();
 b15zdnd11an1n64x5 FILLER_183_887 ();
 b15zdnd11an1n64x5 FILLER_183_951 ();
 b15zdnd11an1n64x5 FILLER_183_1015 ();
 b15zdnd11an1n32x5 FILLER_183_1079 ();
 b15zdnd11an1n04x5 FILLER_183_1111 ();
 b15zdnd11an1n64x5 FILLER_183_1132 ();
 b15zdnd11an1n64x5 FILLER_183_1196 ();
 b15zdnd11an1n08x5 FILLER_183_1260 ();
 b15zdnd11an1n32x5 FILLER_183_1277 ();
 b15zdnd11an1n16x5 FILLER_183_1309 ();
 b15zdnd11an1n04x5 FILLER_183_1325 ();
 b15zdnd00an1n02x5 FILLER_183_1329 ();
 b15zdnd11an1n64x5 FILLER_183_1349 ();
 b15zdnd11an1n16x5 FILLER_183_1413 ();
 b15zdnd11an1n08x5 FILLER_183_1429 ();
 b15zdnd11an1n04x5 FILLER_183_1437 ();
 b15zdnd00an1n02x5 FILLER_183_1441 ();
 b15zdnd00an1n01x5 FILLER_183_1443 ();
 b15zdnd11an1n32x5 FILLER_183_1468 ();
 b15zdnd00an1n01x5 FILLER_183_1500 ();
 b15zdnd11an1n64x5 FILLER_183_1513 ();
 b15zdnd11an1n64x5 FILLER_183_1577 ();
 b15zdnd11an1n64x5 FILLER_183_1641 ();
 b15zdnd11an1n64x5 FILLER_183_1705 ();
 b15zdnd11an1n64x5 FILLER_183_1769 ();
 b15zdnd11an1n64x5 FILLER_183_1833 ();
 b15zdnd11an1n64x5 FILLER_183_1897 ();
 b15zdnd11an1n64x5 FILLER_183_1961 ();
 b15zdnd11an1n32x5 FILLER_183_2025 ();
 b15zdnd11an1n08x5 FILLER_183_2057 ();
 b15zdnd00an1n02x5 FILLER_183_2065 ();
 b15zdnd11an1n04x5 FILLER_183_2085 ();
 b15zdnd11an1n64x5 FILLER_183_2092 ();
 b15zdnd11an1n64x5 FILLER_183_2156 ();
 b15zdnd11an1n04x5 FILLER_183_2242 ();
 b15zdnd11an1n08x5 FILLER_183_2266 ();
 b15zdnd00an1n02x5 FILLER_183_2282 ();
 b15zdnd00an1n02x5 FILLER_184_8 ();
 b15zdnd11an1n64x5 FILLER_184_24 ();
 b15zdnd11an1n64x5 FILLER_184_88 ();
 b15zdnd11an1n16x5 FILLER_184_152 ();
 b15zdnd00an1n02x5 FILLER_184_168 ();
 b15zdnd00an1n01x5 FILLER_184_170 ();
 b15zdnd11an1n04x5 FILLER_184_191 ();
 b15zdnd11an1n64x5 FILLER_184_205 ();
 b15zdnd11an1n32x5 FILLER_184_269 ();
 b15zdnd11an1n04x5 FILLER_184_301 ();
 b15zdnd00an1n02x5 FILLER_184_305 ();
 b15zdnd00an1n01x5 FILLER_184_307 ();
 b15zdnd11an1n64x5 FILLER_184_317 ();
 b15zdnd11an1n64x5 FILLER_184_381 ();
 b15zdnd11an1n64x5 FILLER_184_445 ();
 b15zdnd11an1n64x5 FILLER_184_509 ();
 b15zdnd11an1n16x5 FILLER_184_573 ();
 b15zdnd00an1n02x5 FILLER_184_589 ();
 b15zdnd11an1n32x5 FILLER_184_602 ();
 b15zdnd11an1n04x5 FILLER_184_634 ();
 b15zdnd00an1n01x5 FILLER_184_638 ();
 b15zdnd11an1n64x5 FILLER_184_642 ();
 b15zdnd11an1n08x5 FILLER_184_706 ();
 b15zdnd11an1n04x5 FILLER_184_714 ();
 b15zdnd11an1n08x5 FILLER_184_726 ();
 b15zdnd11an1n04x5 FILLER_184_734 ();
 b15zdnd00an1n02x5 FILLER_184_738 ();
 b15zdnd00an1n01x5 FILLER_184_740 ();
 b15zdnd11an1n32x5 FILLER_184_746 ();
 b15zdnd11an1n08x5 FILLER_184_778 ();
 b15zdnd11an1n64x5 FILLER_184_798 ();
 b15zdnd11an1n64x5 FILLER_184_862 ();
 b15zdnd11an1n32x5 FILLER_184_926 ();
 b15zdnd11an1n16x5 FILLER_184_958 ();
 b15zdnd11an1n08x5 FILLER_184_974 ();
 b15zdnd11an1n32x5 FILLER_184_994 ();
 b15zdnd11an1n08x5 FILLER_184_1026 ();
 b15zdnd11an1n64x5 FILLER_184_1051 ();
 b15zdnd11an1n32x5 FILLER_184_1115 ();
 b15zdnd11an1n16x5 FILLER_184_1147 ();
 b15zdnd11an1n08x5 FILLER_184_1163 ();
 b15zdnd11an1n04x5 FILLER_184_1171 ();
 b15zdnd00an1n01x5 FILLER_184_1175 ();
 b15zdnd11an1n32x5 FILLER_184_1189 ();
 b15zdnd11an1n16x5 FILLER_184_1221 ();
 b15zdnd00an1n02x5 FILLER_184_1237 ();
 b15zdnd00an1n01x5 FILLER_184_1239 ();
 b15zdnd11an1n16x5 FILLER_184_1251 ();
 b15zdnd11an1n04x5 FILLER_184_1267 ();
 b15zdnd00an1n02x5 FILLER_184_1271 ();
 b15zdnd11an1n32x5 FILLER_184_1289 ();
 b15zdnd11an1n04x5 FILLER_184_1321 ();
 b15zdnd00an1n02x5 FILLER_184_1325 ();
 b15zdnd11an1n64x5 FILLER_184_1341 ();
 b15zdnd11an1n32x5 FILLER_184_1405 ();
 b15zdnd11an1n08x5 FILLER_184_1437 ();
 b15zdnd00an1n02x5 FILLER_184_1445 ();
 b15zdnd00an1n01x5 FILLER_184_1447 ();
 b15zdnd11an1n16x5 FILLER_184_1458 ();
 b15zdnd11an1n08x5 FILLER_184_1474 ();
 b15zdnd11an1n04x5 FILLER_184_1482 ();
 b15zdnd00an1n01x5 FILLER_184_1486 ();
 b15zdnd11an1n16x5 FILLER_184_1499 ();
 b15zdnd11an1n04x5 FILLER_184_1515 ();
 b15zdnd00an1n02x5 FILLER_184_1519 ();
 b15zdnd11an1n32x5 FILLER_184_1530 ();
 b15zdnd11an1n16x5 FILLER_184_1562 ();
 b15zdnd00an1n02x5 FILLER_184_1578 ();
 b15zdnd11an1n64x5 FILLER_184_1594 ();
 b15zdnd11an1n64x5 FILLER_184_1658 ();
 b15zdnd11an1n64x5 FILLER_184_1722 ();
 b15zdnd11an1n64x5 FILLER_184_1786 ();
 b15zdnd11an1n64x5 FILLER_184_1850 ();
 b15zdnd11an1n64x5 FILLER_184_1914 ();
 b15zdnd11an1n64x5 FILLER_184_1978 ();
 b15zdnd11an1n32x5 FILLER_184_2042 ();
 b15zdnd11an1n16x5 FILLER_184_2074 ();
 b15zdnd11an1n32x5 FILLER_184_2093 ();
 b15zdnd11an1n16x5 FILLER_184_2125 ();
 b15zdnd11an1n08x5 FILLER_184_2141 ();
 b15zdnd11an1n04x5 FILLER_184_2149 ();
 b15zdnd00an1n01x5 FILLER_184_2153 ();
 b15zdnd11an1n64x5 FILLER_184_2162 ();
 b15zdnd11an1n04x5 FILLER_184_2226 ();
 b15zdnd00an1n02x5 FILLER_184_2230 ();
 b15zdnd00an1n02x5 FILLER_184_2274 ();
 b15zdnd11an1n64x5 FILLER_185_0 ();
 b15zdnd11an1n64x5 FILLER_185_64 ();
 b15zdnd11an1n64x5 FILLER_185_128 ();
 b15zdnd11an1n16x5 FILLER_185_192 ();
 b15zdnd11an1n08x5 FILLER_185_208 ();
 b15zdnd11an1n04x5 FILLER_185_216 ();
 b15zdnd00an1n01x5 FILLER_185_220 ();
 b15zdnd11an1n64x5 FILLER_185_234 ();
 b15zdnd11an1n64x5 FILLER_185_298 ();
 b15zdnd11an1n64x5 FILLER_185_362 ();
 b15zdnd00an1n01x5 FILLER_185_426 ();
 b15zdnd11an1n64x5 FILLER_185_447 ();
 b15zdnd11an1n64x5 FILLER_185_511 ();
 b15zdnd11an1n64x5 FILLER_185_575 ();
 b15zdnd11an1n64x5 FILLER_185_639 ();
 b15zdnd11an1n64x5 FILLER_185_703 ();
 b15zdnd11an1n16x5 FILLER_185_767 ();
 b15zdnd11an1n04x5 FILLER_185_783 ();
 b15zdnd00an1n02x5 FILLER_185_787 ();
 b15zdnd11an1n32x5 FILLER_185_807 ();
 b15zdnd00an1n02x5 FILLER_185_839 ();
 b15zdnd00an1n01x5 FILLER_185_841 ();
 b15zdnd11an1n04x5 FILLER_185_860 ();
 b15zdnd11an1n64x5 FILLER_185_879 ();
 b15zdnd11an1n04x5 FILLER_185_943 ();
 b15zdnd00an1n01x5 FILLER_185_947 ();
 b15zdnd11an1n16x5 FILLER_185_960 ();
 b15zdnd11an1n04x5 FILLER_185_976 ();
 b15zdnd11an1n64x5 FILLER_185_994 ();
 b15zdnd11an1n64x5 FILLER_185_1058 ();
 b15zdnd11an1n16x5 FILLER_185_1122 ();
 b15zdnd11an1n04x5 FILLER_185_1138 ();
 b15zdnd11an1n08x5 FILLER_185_1162 ();
 b15zdnd11an1n04x5 FILLER_185_1170 ();
 b15zdnd11an1n64x5 FILLER_185_1219 ();
 b15zdnd11an1n08x5 FILLER_185_1283 ();
 b15zdnd00an1n01x5 FILLER_185_1291 ();
 b15zdnd11an1n64x5 FILLER_185_1311 ();
 b15zdnd11an1n64x5 FILLER_185_1375 ();
 b15zdnd11an1n32x5 FILLER_185_1439 ();
 b15zdnd11an1n16x5 FILLER_185_1471 ();
 b15zdnd11an1n04x5 FILLER_185_1487 ();
 b15zdnd00an1n02x5 FILLER_185_1491 ();
 b15zdnd00an1n01x5 FILLER_185_1493 ();
 b15zdnd11an1n64x5 FILLER_185_1501 ();
 b15zdnd11an1n64x5 FILLER_185_1565 ();
 b15zdnd11an1n32x5 FILLER_185_1629 ();
 b15zdnd11an1n08x5 FILLER_185_1661 ();
 b15zdnd11an1n04x5 FILLER_185_1669 ();
 b15zdnd00an1n01x5 FILLER_185_1673 ();
 b15zdnd11an1n32x5 FILLER_185_1716 ();
 b15zdnd11an1n08x5 FILLER_185_1748 ();
 b15zdnd00an1n02x5 FILLER_185_1756 ();
 b15zdnd11an1n64x5 FILLER_185_1764 ();
 b15zdnd11an1n64x5 FILLER_185_1828 ();
 b15zdnd11an1n64x5 FILLER_185_1892 ();
 b15zdnd11an1n32x5 FILLER_185_1956 ();
 b15zdnd11an1n04x5 FILLER_185_1988 ();
 b15zdnd00an1n02x5 FILLER_185_1992 ();
 b15zdnd11an1n64x5 FILLER_185_2008 ();
 b15zdnd11an1n64x5 FILLER_185_2072 ();
 b15zdnd11an1n64x5 FILLER_185_2136 ();
 b15zdnd11an1n08x5 FILLER_185_2200 ();
 b15zdnd11an1n04x5 FILLER_185_2208 ();
 b15zdnd11an1n04x5 FILLER_185_2222 ();
 b15zdnd00an1n02x5 FILLER_185_2226 ();
 b15zdnd11an1n08x5 FILLER_185_2270 ();
 b15zdnd11an1n04x5 FILLER_185_2278 ();
 b15zdnd00an1n02x5 FILLER_185_2282 ();
 b15zdnd00an1n02x5 FILLER_186_8 ();
 b15zdnd11an1n08x5 FILLER_186_14 ();
 b15zdnd11an1n04x5 FILLER_186_22 ();
 b15zdnd00an1n01x5 FILLER_186_26 ();
 b15zdnd11an1n64x5 FILLER_186_31 ();
 b15zdnd11an1n64x5 FILLER_186_95 ();
 b15zdnd11an1n64x5 FILLER_186_159 ();
 b15zdnd11an1n64x5 FILLER_186_223 ();
 b15zdnd11an1n64x5 FILLER_186_287 ();
 b15zdnd11an1n32x5 FILLER_186_351 ();
 b15zdnd11an1n16x5 FILLER_186_383 ();
 b15zdnd11an1n08x5 FILLER_186_399 ();
 b15zdnd00an1n02x5 FILLER_186_407 ();
 b15zdnd11an1n64x5 FILLER_186_412 ();
 b15zdnd11an1n64x5 FILLER_186_476 ();
 b15zdnd11an1n32x5 FILLER_186_540 ();
 b15zdnd11an1n08x5 FILLER_186_572 ();
 b15zdnd11an1n04x5 FILLER_186_580 ();
 b15zdnd00an1n02x5 FILLER_186_584 ();
 b15zdnd11an1n64x5 FILLER_186_602 ();
 b15zdnd11an1n32x5 FILLER_186_666 ();
 b15zdnd11an1n16x5 FILLER_186_698 ();
 b15zdnd11an1n04x5 FILLER_186_714 ();
 b15zdnd11an1n64x5 FILLER_186_726 ();
 b15zdnd11an1n64x5 FILLER_186_790 ();
 b15zdnd11an1n04x5 FILLER_186_854 ();
 b15zdnd00an1n01x5 FILLER_186_858 ();
 b15zdnd11an1n64x5 FILLER_186_895 ();
 b15zdnd11an1n32x5 FILLER_186_959 ();
 b15zdnd11an1n08x5 FILLER_186_991 ();
 b15zdnd11an1n64x5 FILLER_186_1009 ();
 b15zdnd11an1n32x5 FILLER_186_1073 ();
 b15zdnd11an1n16x5 FILLER_186_1105 ();
 b15zdnd00an1n01x5 FILLER_186_1121 ();
 b15zdnd11an1n08x5 FILLER_186_1142 ();
 b15zdnd11an1n04x5 FILLER_186_1150 ();
 b15zdnd00an1n02x5 FILLER_186_1154 ();
 b15zdnd11an1n64x5 FILLER_186_1175 ();
 b15zdnd11an1n08x5 FILLER_186_1239 ();
 b15zdnd11an1n04x5 FILLER_186_1247 ();
 b15zdnd00an1n02x5 FILLER_186_1251 ();
 b15zdnd11an1n16x5 FILLER_186_1260 ();
 b15zdnd00an1n02x5 FILLER_186_1276 ();
 b15zdnd00an1n01x5 FILLER_186_1278 ();
 b15zdnd11an1n32x5 FILLER_186_1289 ();
 b15zdnd11an1n16x5 FILLER_186_1321 ();
 b15zdnd11an1n64x5 FILLER_186_1346 ();
 b15zdnd11an1n64x5 FILLER_186_1410 ();
 b15zdnd11an1n64x5 FILLER_186_1474 ();
 b15zdnd11an1n64x5 FILLER_186_1538 ();
 b15zdnd11an1n16x5 FILLER_186_1602 ();
 b15zdnd11an1n08x5 FILLER_186_1618 ();
 b15zdnd00an1n01x5 FILLER_186_1626 ();
 b15zdnd11an1n32x5 FILLER_186_1636 ();
 b15zdnd11an1n04x5 FILLER_186_1668 ();
 b15zdnd00an1n02x5 FILLER_186_1672 ();
 b15zdnd00an1n01x5 FILLER_186_1674 ();
 b15zdnd11an1n64x5 FILLER_186_1693 ();
 b15zdnd11an1n64x5 FILLER_186_1757 ();
 b15zdnd11an1n64x5 FILLER_186_1821 ();
 b15zdnd11an1n64x5 FILLER_186_1885 ();
 b15zdnd11an1n64x5 FILLER_186_1949 ();
 b15zdnd11an1n64x5 FILLER_186_2013 ();
 b15zdnd11an1n64x5 FILLER_186_2077 ();
 b15zdnd11an1n08x5 FILLER_186_2141 ();
 b15zdnd11an1n04x5 FILLER_186_2149 ();
 b15zdnd00an1n01x5 FILLER_186_2153 ();
 b15zdnd11an1n32x5 FILLER_186_2162 ();
 b15zdnd11an1n08x5 FILLER_186_2194 ();
 b15zdnd11an1n04x5 FILLER_186_2202 ();
 b15zdnd00an1n02x5 FILLER_186_2206 ();
 b15zdnd11an1n04x5 FILLER_186_2250 ();
 b15zdnd00an1n02x5 FILLER_186_2254 ();
 b15zdnd11an1n16x5 FILLER_186_2260 ();
 b15zdnd11an1n08x5 FILLER_187_0 ();
 b15zdnd00an1n02x5 FILLER_187_8 ();
 b15zdnd00an1n01x5 FILLER_187_10 ();
 b15zdnd11an1n64x5 FILLER_187_15 ();
 b15zdnd11an1n64x5 FILLER_187_79 ();
 b15zdnd11an1n64x5 FILLER_187_143 ();
 b15zdnd11an1n04x5 FILLER_187_207 ();
 b15zdnd00an1n02x5 FILLER_187_211 ();
 b15zdnd11an1n04x5 FILLER_187_226 ();
 b15zdnd00an1n02x5 FILLER_187_230 ();
 b15zdnd00an1n01x5 FILLER_187_232 ();
 b15zdnd11an1n64x5 FILLER_187_252 ();
 b15zdnd11an1n64x5 FILLER_187_316 ();
 b15zdnd11an1n16x5 FILLER_187_380 ();
 b15zdnd11an1n08x5 FILLER_187_396 ();
 b15zdnd11an1n04x5 FILLER_187_407 ();
 b15zdnd11an1n64x5 FILLER_187_414 ();
 b15zdnd11an1n32x5 FILLER_187_478 ();
 b15zdnd11an1n08x5 FILLER_187_510 ();
 b15zdnd00an1n01x5 FILLER_187_518 ();
 b15zdnd11an1n64x5 FILLER_187_535 ();
 b15zdnd11an1n64x5 FILLER_187_599 ();
 b15zdnd11an1n64x5 FILLER_187_663 ();
 b15zdnd11an1n64x5 FILLER_187_727 ();
 b15zdnd11an1n32x5 FILLER_187_791 ();
 b15zdnd11an1n16x5 FILLER_187_823 ();
 b15zdnd00an1n01x5 FILLER_187_839 ();
 b15zdnd11an1n64x5 FILLER_187_855 ();
 b15zdnd11an1n64x5 FILLER_187_919 ();
 b15zdnd11an1n64x5 FILLER_187_983 ();
 b15zdnd11an1n04x5 FILLER_187_1047 ();
 b15zdnd00an1n02x5 FILLER_187_1051 ();
 b15zdnd11an1n64x5 FILLER_187_1064 ();
 b15zdnd11an1n64x5 FILLER_187_1128 ();
 b15zdnd11an1n64x5 FILLER_187_1192 ();
 b15zdnd11an1n64x5 FILLER_187_1256 ();
 b15zdnd11an1n64x5 FILLER_187_1320 ();
 b15zdnd11an1n64x5 FILLER_187_1384 ();
 b15zdnd11an1n64x5 FILLER_187_1448 ();
 b15zdnd11an1n64x5 FILLER_187_1512 ();
 b15zdnd11an1n32x5 FILLER_187_1576 ();
 b15zdnd11an1n16x5 FILLER_187_1608 ();
 b15zdnd11an1n08x5 FILLER_187_1624 ();
 b15zdnd11an1n16x5 FILLER_187_1648 ();
 b15zdnd11an1n08x5 FILLER_187_1664 ();
 b15zdnd00an1n02x5 FILLER_187_1672 ();
 b15zdnd11an1n04x5 FILLER_187_1694 ();
 b15zdnd11an1n04x5 FILLER_187_1709 ();
 b15zdnd11an1n32x5 FILLER_187_1721 ();
 b15zdnd11an1n64x5 FILLER_187_1774 ();
 b15zdnd11an1n64x5 FILLER_187_1838 ();
 b15zdnd11an1n32x5 FILLER_187_1902 ();
 b15zdnd11an1n08x5 FILLER_187_1934 ();
 b15zdnd11an1n04x5 FILLER_187_1942 ();
 b15zdnd00an1n02x5 FILLER_187_1946 ();
 b15zdnd11an1n16x5 FILLER_187_1967 ();
 b15zdnd11an1n04x5 FILLER_187_1983 ();
 b15zdnd11an1n64x5 FILLER_187_1999 ();
 b15zdnd11an1n64x5 FILLER_187_2063 ();
 b15zdnd11an1n64x5 FILLER_187_2127 ();
 b15zdnd11an1n32x5 FILLER_187_2191 ();
 b15zdnd00an1n01x5 FILLER_187_2223 ();
 b15zdnd11an1n08x5 FILLER_187_2269 ();
 b15zdnd11an1n04x5 FILLER_187_2277 ();
 b15zdnd00an1n02x5 FILLER_187_2281 ();
 b15zdnd00an1n01x5 FILLER_187_2283 ();
 b15zdnd11an1n04x5 FILLER_188_8 ();
 b15zdnd00an1n02x5 FILLER_188_12 ();
 b15zdnd00an1n01x5 FILLER_188_14 ();
 b15zdnd11an1n64x5 FILLER_188_19 ();
 b15zdnd11an1n64x5 FILLER_188_83 ();
 b15zdnd11an1n64x5 FILLER_188_147 ();
 b15zdnd11an1n08x5 FILLER_188_211 ();
 b15zdnd11an1n04x5 FILLER_188_219 ();
 b15zdnd00an1n01x5 FILLER_188_223 ();
 b15zdnd11an1n64x5 FILLER_188_266 ();
 b15zdnd11an1n32x5 FILLER_188_330 ();
 b15zdnd11an1n08x5 FILLER_188_362 ();
 b15zdnd11an1n04x5 FILLER_188_370 ();
 b15zdnd00an1n01x5 FILLER_188_374 ();
 b15zdnd11an1n04x5 FILLER_188_380 ();
 b15zdnd11an1n08x5 FILLER_188_436 ();
 b15zdnd00an1n02x5 FILLER_188_444 ();
 b15zdnd00an1n01x5 FILLER_188_446 ();
 b15zdnd11an1n64x5 FILLER_188_462 ();
 b15zdnd11an1n64x5 FILLER_188_526 ();
 b15zdnd11an1n64x5 FILLER_188_590 ();
 b15zdnd11an1n64x5 FILLER_188_654 ();
 b15zdnd11an1n64x5 FILLER_188_726 ();
 b15zdnd11an1n64x5 FILLER_188_790 ();
 b15zdnd11an1n32x5 FILLER_188_854 ();
 b15zdnd11an1n08x5 FILLER_188_886 ();
 b15zdnd11an1n04x5 FILLER_188_894 ();
 b15zdnd11an1n64x5 FILLER_188_912 ();
 b15zdnd11an1n64x5 FILLER_188_976 ();
 b15zdnd11an1n64x5 FILLER_188_1040 ();
 b15zdnd11an1n64x5 FILLER_188_1104 ();
 b15zdnd11an1n32x5 FILLER_188_1168 ();
 b15zdnd11an1n16x5 FILLER_188_1200 ();
 b15zdnd11an1n08x5 FILLER_188_1216 ();
 b15zdnd00an1n02x5 FILLER_188_1224 ();
 b15zdnd11an1n16x5 FILLER_188_1235 ();
 b15zdnd00an1n02x5 FILLER_188_1251 ();
 b15zdnd11an1n64x5 FILLER_188_1260 ();
 b15zdnd11an1n16x5 FILLER_188_1324 ();
 b15zdnd11an1n08x5 FILLER_188_1340 ();
 b15zdnd00an1n01x5 FILLER_188_1348 ();
 b15zdnd11an1n64x5 FILLER_188_1365 ();
 b15zdnd11an1n64x5 FILLER_188_1429 ();
 b15zdnd11an1n64x5 FILLER_188_1493 ();
 b15zdnd11an1n64x5 FILLER_188_1557 ();
 b15zdnd11an1n08x5 FILLER_188_1621 ();
 b15zdnd11an1n04x5 FILLER_188_1629 ();
 b15zdnd11an1n64x5 FILLER_188_1644 ();
 b15zdnd11an1n64x5 FILLER_188_1708 ();
 b15zdnd11an1n64x5 FILLER_188_1772 ();
 b15zdnd11an1n32x5 FILLER_188_1836 ();
 b15zdnd11an1n04x5 FILLER_188_1868 ();
 b15zdnd11an1n64x5 FILLER_188_1886 ();
 b15zdnd11an1n64x5 FILLER_188_1950 ();
 b15zdnd11an1n64x5 FILLER_188_2014 ();
 b15zdnd11an1n64x5 FILLER_188_2078 ();
 b15zdnd11an1n08x5 FILLER_188_2142 ();
 b15zdnd11an1n04x5 FILLER_188_2150 ();
 b15zdnd11an1n64x5 FILLER_188_2162 ();
 b15zdnd11an1n04x5 FILLER_188_2226 ();
 b15zdnd00an1n02x5 FILLER_188_2230 ();
 b15zdnd11an1n16x5 FILLER_188_2252 ();
 b15zdnd11an1n08x5 FILLER_188_2268 ();
 b15zdnd11an1n64x5 FILLER_189_0 ();
 b15zdnd11an1n08x5 FILLER_189_64 ();
 b15zdnd11an1n04x5 FILLER_189_72 ();
 b15zdnd00an1n02x5 FILLER_189_76 ();
 b15zdnd11an1n64x5 FILLER_189_98 ();
 b15zdnd11an1n64x5 FILLER_189_162 ();
 b15zdnd11an1n32x5 FILLER_189_226 ();
 b15zdnd11an1n16x5 FILLER_189_258 ();
 b15zdnd11an1n04x5 FILLER_189_274 ();
 b15zdnd11an1n32x5 FILLER_189_320 ();
 b15zdnd11an1n16x5 FILLER_189_352 ();
 b15zdnd11an1n08x5 FILLER_189_368 ();
 b15zdnd11an1n04x5 FILLER_189_376 ();
 b15zdnd00an1n01x5 FILLER_189_380 ();
 b15zdnd11an1n16x5 FILLER_189_423 ();
 b15zdnd00an1n02x5 FILLER_189_439 ();
 b15zdnd11an1n08x5 FILLER_189_483 ();
 b15zdnd00an1n02x5 FILLER_189_491 ();
 b15zdnd11an1n64x5 FILLER_189_496 ();
 b15zdnd11an1n64x5 FILLER_189_560 ();
 b15zdnd11an1n64x5 FILLER_189_624 ();
 b15zdnd11an1n64x5 FILLER_189_688 ();
 b15zdnd11an1n64x5 FILLER_189_752 ();
 b15zdnd11an1n64x5 FILLER_189_816 ();
 b15zdnd11an1n64x5 FILLER_189_880 ();
 b15zdnd11an1n64x5 FILLER_189_944 ();
 b15zdnd11an1n64x5 FILLER_189_1008 ();
 b15zdnd11an1n64x5 FILLER_189_1072 ();
 b15zdnd11an1n64x5 FILLER_189_1136 ();
 b15zdnd11an1n64x5 FILLER_189_1200 ();
 b15zdnd11an1n64x5 FILLER_189_1264 ();
 b15zdnd11an1n16x5 FILLER_189_1328 ();
 b15zdnd11an1n04x5 FILLER_189_1355 ();
 b15zdnd00an1n02x5 FILLER_189_1359 ();
 b15zdnd11an1n64x5 FILLER_189_1374 ();
 b15zdnd11an1n64x5 FILLER_189_1438 ();
 b15zdnd11an1n04x5 FILLER_189_1502 ();
 b15zdnd00an1n02x5 FILLER_189_1506 ();
 b15zdnd00an1n01x5 FILLER_189_1508 ();
 b15zdnd11an1n04x5 FILLER_189_1518 ();
 b15zdnd11an1n64x5 FILLER_189_1534 ();
 b15zdnd11an1n32x5 FILLER_189_1598 ();
 b15zdnd00an1n02x5 FILLER_189_1630 ();
 b15zdnd00an1n01x5 FILLER_189_1632 ();
 b15zdnd11an1n64x5 FILLER_189_1641 ();
 b15zdnd11an1n64x5 FILLER_189_1705 ();
 b15zdnd11an1n64x5 FILLER_189_1769 ();
 b15zdnd11an1n32x5 FILLER_189_1833 ();
 b15zdnd11an1n08x5 FILLER_189_1865 ();
 b15zdnd11an1n04x5 FILLER_189_1873 ();
 b15zdnd00an1n02x5 FILLER_189_1877 ();
 b15zdnd00an1n01x5 FILLER_189_1879 ();
 b15zdnd11an1n04x5 FILLER_189_1885 ();
 b15zdnd11an1n64x5 FILLER_189_1909 ();
 b15zdnd11an1n64x5 FILLER_189_1973 ();
 b15zdnd11an1n64x5 FILLER_189_2037 ();
 b15zdnd11an1n64x5 FILLER_189_2101 ();
 b15zdnd11an1n64x5 FILLER_189_2165 ();
 b15zdnd11an1n32x5 FILLER_189_2229 ();
 b15zdnd11an1n16x5 FILLER_189_2261 ();
 b15zdnd11an1n04x5 FILLER_189_2277 ();
 b15zdnd00an1n02x5 FILLER_189_2281 ();
 b15zdnd00an1n01x5 FILLER_189_2283 ();
 b15zdnd11an1n32x5 FILLER_190_8 ();
 b15zdnd00an1n02x5 FILLER_190_40 ();
 b15zdnd00an1n01x5 FILLER_190_42 ();
 b15zdnd11an1n04x5 FILLER_190_46 ();
 b15zdnd11an1n16x5 FILLER_190_53 ();
 b15zdnd11an1n64x5 FILLER_190_77 ();
 b15zdnd11an1n64x5 FILLER_190_141 ();
 b15zdnd11an1n64x5 FILLER_190_205 ();
 b15zdnd11an1n64x5 FILLER_190_269 ();
 b15zdnd11an1n64x5 FILLER_190_333 ();
 b15zdnd11an1n64x5 FILLER_190_417 ();
 b15zdnd11an1n04x5 FILLER_190_481 ();
 b15zdnd11an1n64x5 FILLER_190_537 ();
 b15zdnd11an1n64x5 FILLER_190_601 ();
 b15zdnd11an1n32x5 FILLER_190_665 ();
 b15zdnd11an1n16x5 FILLER_190_697 ();
 b15zdnd11an1n04x5 FILLER_190_713 ();
 b15zdnd00an1n01x5 FILLER_190_717 ();
 b15zdnd11an1n64x5 FILLER_190_726 ();
 b15zdnd11an1n64x5 FILLER_190_790 ();
 b15zdnd00an1n02x5 FILLER_190_854 ();
 b15zdnd00an1n01x5 FILLER_190_856 ();
 b15zdnd11an1n64x5 FILLER_190_888 ();
 b15zdnd11an1n64x5 FILLER_190_952 ();
 b15zdnd11an1n64x5 FILLER_190_1016 ();
 b15zdnd11an1n64x5 FILLER_190_1080 ();
 b15zdnd11an1n64x5 FILLER_190_1144 ();
 b15zdnd11an1n64x5 FILLER_190_1208 ();
 b15zdnd11an1n64x5 FILLER_190_1272 ();
 b15zdnd11an1n64x5 FILLER_190_1336 ();
 b15zdnd11an1n64x5 FILLER_190_1400 ();
 b15zdnd11an1n64x5 FILLER_190_1464 ();
 b15zdnd11an1n64x5 FILLER_190_1528 ();
 b15zdnd11an1n32x5 FILLER_190_1592 ();
 b15zdnd11an1n08x5 FILLER_190_1624 ();
 b15zdnd11an1n04x5 FILLER_190_1632 ();
 b15zdnd00an1n02x5 FILLER_190_1636 ();
 b15zdnd00an1n01x5 FILLER_190_1638 ();
 b15zdnd11an1n04x5 FILLER_190_1651 ();
 b15zdnd00an1n01x5 FILLER_190_1655 ();
 b15zdnd11an1n16x5 FILLER_190_1659 ();
 b15zdnd11an1n08x5 FILLER_190_1675 ();
 b15zdnd11an1n04x5 FILLER_190_1683 ();
 b15zdnd11an1n64x5 FILLER_190_1729 ();
 b15zdnd11an1n32x5 FILLER_190_1793 ();
 b15zdnd11an1n08x5 FILLER_190_1825 ();
 b15zdnd00an1n01x5 FILLER_190_1833 ();
 b15zdnd11an1n16x5 FILLER_190_1848 ();
 b15zdnd11an1n64x5 FILLER_190_1884 ();
 b15zdnd11an1n64x5 FILLER_190_1948 ();
 b15zdnd11an1n64x5 FILLER_190_2012 ();
 b15zdnd11an1n64x5 FILLER_190_2076 ();
 b15zdnd11an1n08x5 FILLER_190_2140 ();
 b15zdnd11an1n04x5 FILLER_190_2148 ();
 b15zdnd00an1n02x5 FILLER_190_2152 ();
 b15zdnd11an1n64x5 FILLER_190_2162 ();
 b15zdnd11an1n16x5 FILLER_190_2226 ();
 b15zdnd00an1n02x5 FILLER_190_2242 ();
 b15zdnd11an1n16x5 FILLER_190_2248 ();
 b15zdnd11an1n08x5 FILLER_190_2264 ();
 b15zdnd11an1n04x5 FILLER_190_2272 ();
 b15zdnd11an1n16x5 FILLER_191_0 ();
 b15zdnd11an1n08x5 FILLER_191_16 ();
 b15zdnd11an1n64x5 FILLER_191_76 ();
 b15zdnd11an1n64x5 FILLER_191_140 ();
 b15zdnd11an1n64x5 FILLER_191_204 ();
 b15zdnd11an1n64x5 FILLER_191_268 ();
 b15zdnd11an1n64x5 FILLER_191_332 ();
 b15zdnd11an1n64x5 FILLER_191_396 ();
 b15zdnd11an1n32x5 FILLER_191_460 ();
 b15zdnd11an1n04x5 FILLER_191_492 ();
 b15zdnd00an1n02x5 FILLER_191_496 ();
 b15zdnd11an1n08x5 FILLER_191_501 ();
 b15zdnd00an1n01x5 FILLER_191_509 ();
 b15zdnd11an1n64x5 FILLER_191_513 ();
 b15zdnd11an1n64x5 FILLER_191_577 ();
 b15zdnd11an1n64x5 FILLER_191_641 ();
 b15zdnd11an1n64x5 FILLER_191_705 ();
 b15zdnd11an1n64x5 FILLER_191_769 ();
 b15zdnd11an1n64x5 FILLER_191_833 ();
 b15zdnd11an1n64x5 FILLER_191_897 ();
 b15zdnd11an1n64x5 FILLER_191_961 ();
 b15zdnd11an1n64x5 FILLER_191_1025 ();
 b15zdnd11an1n64x5 FILLER_191_1089 ();
 b15zdnd11an1n64x5 FILLER_191_1153 ();
 b15zdnd11an1n64x5 FILLER_191_1217 ();
 b15zdnd11an1n64x5 FILLER_191_1281 ();
 b15zdnd11an1n64x5 FILLER_191_1345 ();
 b15zdnd11an1n64x5 FILLER_191_1409 ();
 b15zdnd11an1n64x5 FILLER_191_1473 ();
 b15zdnd11an1n64x5 FILLER_191_1537 ();
 b15zdnd11an1n32x5 FILLER_191_1601 ();
 b15zdnd11an1n08x5 FILLER_191_1633 ();
 b15zdnd11an1n04x5 FILLER_191_1641 ();
 b15zdnd00an1n01x5 FILLER_191_1645 ();
 b15zdnd11an1n04x5 FILLER_191_1656 ();
 b15zdnd11an1n64x5 FILLER_191_1663 ();
 b15zdnd11an1n64x5 FILLER_191_1727 ();
 b15zdnd11an1n32x5 FILLER_191_1791 ();
 b15zdnd11an1n16x5 FILLER_191_1823 ();
 b15zdnd11an1n04x5 FILLER_191_1844 ();
 b15zdnd00an1n01x5 FILLER_191_1848 ();
 b15zdnd11an1n64x5 FILLER_191_1865 ();
 b15zdnd11an1n64x5 FILLER_191_1929 ();
 b15zdnd11an1n16x5 FILLER_191_1993 ();
 b15zdnd11an1n04x5 FILLER_191_2009 ();
 b15zdnd11an1n64x5 FILLER_191_2020 ();
 b15zdnd11an1n64x5 FILLER_191_2084 ();
 b15zdnd11an1n64x5 FILLER_191_2148 ();
 b15zdnd00an1n02x5 FILLER_191_2212 ();
 b15zdnd11an1n16x5 FILLER_191_2256 ();
 b15zdnd11an1n08x5 FILLER_191_2272 ();
 b15zdnd11an1n04x5 FILLER_191_2280 ();
 b15zdnd11an1n04x5 FILLER_192_8 ();
 b15zdnd11an1n04x5 FILLER_192_19 ();
 b15zdnd00an1n02x5 FILLER_192_23 ();
 b15zdnd00an1n01x5 FILLER_192_25 ();
 b15zdnd11an1n08x5 FILLER_192_34 ();
 b15zdnd11an1n04x5 FILLER_192_42 ();
 b15zdnd00an1n01x5 FILLER_192_46 ();
 b15zdnd11an1n16x5 FILLER_192_92 ();
 b15zdnd00an1n02x5 FILLER_192_108 ();
 b15zdnd11an1n64x5 FILLER_192_124 ();
 b15zdnd11an1n64x5 FILLER_192_188 ();
 b15zdnd11an1n64x5 FILLER_192_252 ();
 b15zdnd11an1n64x5 FILLER_192_316 ();
 b15zdnd11an1n64x5 FILLER_192_380 ();
 b15zdnd11an1n64x5 FILLER_192_444 ();
 b15zdnd11an1n64x5 FILLER_192_508 ();
 b15zdnd11an1n64x5 FILLER_192_572 ();
 b15zdnd11an1n64x5 FILLER_192_636 ();
 b15zdnd11an1n16x5 FILLER_192_700 ();
 b15zdnd00an1n02x5 FILLER_192_716 ();
 b15zdnd11an1n64x5 FILLER_192_726 ();
 b15zdnd11an1n64x5 FILLER_192_790 ();
 b15zdnd11an1n64x5 FILLER_192_854 ();
 b15zdnd11an1n64x5 FILLER_192_918 ();
 b15zdnd11an1n08x5 FILLER_192_982 ();
 b15zdnd11an1n04x5 FILLER_192_990 ();
 b15zdnd00an1n02x5 FILLER_192_994 ();
 b15zdnd11an1n64x5 FILLER_192_1011 ();
 b15zdnd11an1n64x5 FILLER_192_1075 ();
 b15zdnd11an1n64x5 FILLER_192_1139 ();
 b15zdnd11an1n64x5 FILLER_192_1203 ();
 b15zdnd11an1n64x5 FILLER_192_1267 ();
 b15zdnd11an1n16x5 FILLER_192_1331 ();
 b15zdnd00an1n02x5 FILLER_192_1347 ();
 b15zdnd00an1n01x5 FILLER_192_1349 ();
 b15zdnd11an1n64x5 FILLER_192_1363 ();
 b15zdnd11an1n64x5 FILLER_192_1427 ();
 b15zdnd11an1n64x5 FILLER_192_1491 ();
 b15zdnd11an1n64x5 FILLER_192_1555 ();
 b15zdnd11an1n08x5 FILLER_192_1619 ();
 b15zdnd11an1n04x5 FILLER_192_1627 ();
 b15zdnd00an1n02x5 FILLER_192_1631 ();
 b15zdnd00an1n01x5 FILLER_192_1633 ();
 b15zdnd11an1n04x5 FILLER_192_1642 ();
 b15zdnd11an1n04x5 FILLER_192_1652 ();
 b15zdnd11an1n64x5 FILLER_192_1669 ();
 b15zdnd11an1n04x5 FILLER_192_1733 ();
 b15zdnd00an1n01x5 FILLER_192_1737 ();
 b15zdnd11an1n64x5 FILLER_192_1747 ();
 b15zdnd11an1n16x5 FILLER_192_1811 ();
 b15zdnd11an1n08x5 FILLER_192_1827 ();
 b15zdnd00an1n01x5 FILLER_192_1835 ();
 b15zdnd11an1n04x5 FILLER_192_1857 ();
 b15zdnd11an1n64x5 FILLER_192_1875 ();
 b15zdnd11an1n64x5 FILLER_192_1939 ();
 b15zdnd11an1n64x5 FILLER_192_2003 ();
 b15zdnd11an1n64x5 FILLER_192_2067 ();
 b15zdnd11an1n16x5 FILLER_192_2131 ();
 b15zdnd11an1n04x5 FILLER_192_2147 ();
 b15zdnd00an1n02x5 FILLER_192_2151 ();
 b15zdnd00an1n01x5 FILLER_192_2153 ();
 b15zdnd11an1n16x5 FILLER_192_2162 ();
 b15zdnd00an1n02x5 FILLER_192_2178 ();
 b15zdnd00an1n01x5 FILLER_192_2180 ();
 b15zdnd11an1n32x5 FILLER_192_2223 ();
 b15zdnd11an1n08x5 FILLER_192_2255 ();
 b15zdnd00an1n02x5 FILLER_192_2274 ();
 b15zdnd00an1n02x5 FILLER_193_0 ();
 b15zdnd11an1n16x5 FILLER_193_22 ();
 b15zdnd11an1n08x5 FILLER_193_38 ();
 b15zdnd00an1n01x5 FILLER_193_46 ();
 b15zdnd11an1n32x5 FILLER_193_50 ();
 b15zdnd00an1n01x5 FILLER_193_82 ();
 b15zdnd11an1n64x5 FILLER_193_103 ();
 b15zdnd11an1n64x5 FILLER_193_167 ();
 b15zdnd11an1n32x5 FILLER_193_231 ();
 b15zdnd11an1n04x5 FILLER_193_263 ();
 b15zdnd00an1n02x5 FILLER_193_267 ();
 b15zdnd00an1n01x5 FILLER_193_269 ();
 b15zdnd11an1n04x5 FILLER_193_273 ();
 b15zdnd11an1n08x5 FILLER_193_280 ();
 b15zdnd11an1n04x5 FILLER_193_288 ();
 b15zdnd00an1n02x5 FILLER_193_292 ();
 b15zdnd00an1n01x5 FILLER_193_294 ();
 b15zdnd11an1n64x5 FILLER_193_298 ();
 b15zdnd11an1n64x5 FILLER_193_362 ();
 b15zdnd11an1n64x5 FILLER_193_426 ();
 b15zdnd11an1n64x5 FILLER_193_490 ();
 b15zdnd11an1n32x5 FILLER_193_554 ();
 b15zdnd00an1n01x5 FILLER_193_586 ();
 b15zdnd11an1n64x5 FILLER_193_605 ();
 b15zdnd11an1n08x5 FILLER_193_669 ();
 b15zdnd11an1n64x5 FILLER_193_704 ();
 b15zdnd11an1n64x5 FILLER_193_768 ();
 b15zdnd11an1n64x5 FILLER_193_832 ();
 b15zdnd11an1n64x5 FILLER_193_896 ();
 b15zdnd11an1n32x5 FILLER_193_960 ();
 b15zdnd11an1n16x5 FILLER_193_992 ();
 b15zdnd11an1n64x5 FILLER_193_1033 ();
 b15zdnd11an1n64x5 FILLER_193_1097 ();
 b15zdnd11an1n16x5 FILLER_193_1161 ();
 b15zdnd00an1n01x5 FILLER_193_1177 ();
 b15zdnd11an1n64x5 FILLER_193_1196 ();
 b15zdnd11an1n16x5 FILLER_193_1260 ();
 b15zdnd11an1n08x5 FILLER_193_1276 ();
 b15zdnd00an1n02x5 FILLER_193_1284 ();
 b15zdnd00an1n01x5 FILLER_193_1286 ();
 b15zdnd11an1n04x5 FILLER_193_1303 ();
 b15zdnd11an1n64x5 FILLER_193_1325 ();
 b15zdnd11an1n64x5 FILLER_193_1389 ();
 b15zdnd11an1n32x5 FILLER_193_1453 ();
 b15zdnd11an1n16x5 FILLER_193_1485 ();
 b15zdnd11an1n08x5 FILLER_193_1501 ();
 b15zdnd00an1n01x5 FILLER_193_1509 ();
 b15zdnd11an1n32x5 FILLER_193_1519 ();
 b15zdnd11an1n08x5 FILLER_193_1551 ();
 b15zdnd11an1n64x5 FILLER_193_1562 ();
 b15zdnd11an1n16x5 FILLER_193_1626 ();
 b15zdnd00an1n01x5 FILLER_193_1642 ();
 b15zdnd11an1n04x5 FILLER_193_1659 ();
 b15zdnd11an1n64x5 FILLER_193_1683 ();
 b15zdnd11an1n32x5 FILLER_193_1747 ();
 b15zdnd11an1n16x5 FILLER_193_1779 ();
 b15zdnd11an1n08x5 FILLER_193_1795 ();
 b15zdnd11an1n04x5 FILLER_193_1803 ();
 b15zdnd00an1n01x5 FILLER_193_1807 ();
 b15zdnd11an1n16x5 FILLER_193_1825 ();
 b15zdnd11an1n04x5 FILLER_193_1841 ();
 b15zdnd00an1n01x5 FILLER_193_1845 ();
 b15zdnd11an1n64x5 FILLER_193_1888 ();
 b15zdnd11an1n32x5 FILLER_193_1952 ();
 b15zdnd11an1n16x5 FILLER_193_1984 ();
 b15zdnd11an1n08x5 FILLER_193_2000 ();
 b15zdnd11an1n04x5 FILLER_193_2008 ();
 b15zdnd00an1n02x5 FILLER_193_2012 ();
 b15zdnd11an1n64x5 FILLER_193_2020 ();
 b15zdnd11an1n64x5 FILLER_193_2084 ();
 b15zdnd11an1n64x5 FILLER_193_2148 ();
 b15zdnd11an1n16x5 FILLER_193_2212 ();
 b15zdnd11an1n08x5 FILLER_193_2228 ();
 b15zdnd11an1n04x5 FILLER_193_2236 ();
 b15zdnd00an1n01x5 FILLER_193_2240 ();
 b15zdnd11an1n16x5 FILLER_193_2253 ();
 b15zdnd11an1n08x5 FILLER_193_2269 ();
 b15zdnd11an1n04x5 FILLER_193_2277 ();
 b15zdnd00an1n02x5 FILLER_193_2281 ();
 b15zdnd00an1n01x5 FILLER_193_2283 ();
 b15zdnd11an1n32x5 FILLER_194_8 ();
 b15zdnd11an1n16x5 FILLER_194_40 ();
 b15zdnd11an1n08x5 FILLER_194_56 ();
 b15zdnd11an1n64x5 FILLER_194_90 ();
 b15zdnd11an1n64x5 FILLER_194_154 ();
 b15zdnd11an1n16x5 FILLER_194_218 ();
 b15zdnd11an1n08x5 FILLER_194_234 ();
 b15zdnd11an1n04x5 FILLER_194_242 ();
 b15zdnd11an1n64x5 FILLER_194_298 ();
 b15zdnd11an1n64x5 FILLER_194_362 ();
 b15zdnd11an1n64x5 FILLER_194_426 ();
 b15zdnd11an1n64x5 FILLER_194_490 ();
 b15zdnd11an1n64x5 FILLER_194_554 ();
 b15zdnd11an1n64x5 FILLER_194_618 ();
 b15zdnd00an1n01x5 FILLER_194_682 ();
 b15zdnd11an1n16x5 FILLER_194_687 ();
 b15zdnd11an1n08x5 FILLER_194_703 ();
 b15zdnd11an1n04x5 FILLER_194_711 ();
 b15zdnd00an1n02x5 FILLER_194_715 ();
 b15zdnd00an1n01x5 FILLER_194_717 ();
 b15zdnd11an1n64x5 FILLER_194_726 ();
 b15zdnd11an1n64x5 FILLER_194_790 ();
 b15zdnd11an1n64x5 FILLER_194_854 ();
 b15zdnd11an1n64x5 FILLER_194_918 ();
 b15zdnd11an1n64x5 FILLER_194_982 ();
 b15zdnd11an1n64x5 FILLER_194_1046 ();
 b15zdnd11an1n32x5 FILLER_194_1110 ();
 b15zdnd00an1n02x5 FILLER_194_1142 ();
 b15zdnd00an1n01x5 FILLER_194_1144 ();
 b15zdnd11an1n64x5 FILLER_194_1187 ();
 b15zdnd11an1n64x5 FILLER_194_1251 ();
 b15zdnd11an1n64x5 FILLER_194_1315 ();
 b15zdnd11an1n64x5 FILLER_194_1379 ();
 b15zdnd11an1n64x5 FILLER_194_1443 ();
 b15zdnd11an1n64x5 FILLER_194_1507 ();
 b15zdnd11an1n64x5 FILLER_194_1571 ();
 b15zdnd11an1n64x5 FILLER_194_1635 ();
 b15zdnd11an1n16x5 FILLER_194_1699 ();
 b15zdnd11an1n08x5 FILLER_194_1715 ();
 b15zdnd00an1n02x5 FILLER_194_1723 ();
 b15zdnd00an1n01x5 FILLER_194_1725 ();
 b15zdnd11an1n04x5 FILLER_194_1740 ();
 b15zdnd11an1n04x5 FILLER_194_1764 ();
 b15zdnd00an1n02x5 FILLER_194_1768 ();
 b15zdnd00an1n01x5 FILLER_194_1770 ();
 b15zdnd11an1n16x5 FILLER_194_1785 ();
 b15zdnd11an1n08x5 FILLER_194_1801 ();
 b15zdnd11an1n04x5 FILLER_194_1809 ();
 b15zdnd11an1n04x5 FILLER_194_1825 ();
 b15zdnd00an1n02x5 FILLER_194_1829 ();
 b15zdnd00an1n01x5 FILLER_194_1831 ();
 b15zdnd11an1n04x5 FILLER_194_1852 ();
 b15zdnd00an1n02x5 FILLER_194_1856 ();
 b15zdnd00an1n01x5 FILLER_194_1858 ();
 b15zdnd11an1n04x5 FILLER_194_1901 ();
 b15zdnd00an1n02x5 FILLER_194_1905 ();
 b15zdnd11an1n64x5 FILLER_194_1910 ();
 b15zdnd11an1n64x5 FILLER_194_1974 ();
 b15zdnd11an1n64x5 FILLER_194_2038 ();
 b15zdnd11an1n32x5 FILLER_194_2102 ();
 b15zdnd11an1n16x5 FILLER_194_2134 ();
 b15zdnd11an1n04x5 FILLER_194_2150 ();
 b15zdnd11an1n64x5 FILLER_194_2162 ();
 b15zdnd11an1n32x5 FILLER_194_2226 ();
 b15zdnd11an1n16x5 FILLER_194_2258 ();
 b15zdnd00an1n02x5 FILLER_194_2274 ();
 b15zdnd11an1n64x5 FILLER_195_0 ();
 b15zdnd11an1n64x5 FILLER_195_64 ();
 b15zdnd11an1n64x5 FILLER_195_128 ();
 b15zdnd11an1n64x5 FILLER_195_192 ();
 b15zdnd11an1n64x5 FILLER_195_256 ();
 b15zdnd11an1n64x5 FILLER_195_320 ();
 b15zdnd11an1n64x5 FILLER_195_384 ();
 b15zdnd11an1n64x5 FILLER_195_448 ();
 b15zdnd11an1n64x5 FILLER_195_512 ();
 b15zdnd00an1n01x5 FILLER_195_576 ();
 b15zdnd11an1n16x5 FILLER_195_585 ();
 b15zdnd11an1n08x5 FILLER_195_601 ();
 b15zdnd11an1n04x5 FILLER_195_609 ();
 b15zdnd00an1n02x5 FILLER_195_613 ();
 b15zdnd00an1n01x5 FILLER_195_615 ();
 b15zdnd11an1n64x5 FILLER_195_626 ();
 b15zdnd11an1n04x5 FILLER_195_690 ();
 b15zdnd00an1n02x5 FILLER_195_694 ();
 b15zdnd00an1n01x5 FILLER_195_696 ();
 b15zdnd11an1n64x5 FILLER_195_708 ();
 b15zdnd11an1n08x5 FILLER_195_772 ();
 b15zdnd11an1n04x5 FILLER_195_780 ();
 b15zdnd00an1n01x5 FILLER_195_784 ();
 b15zdnd11an1n64x5 FILLER_195_803 ();
 b15zdnd11an1n32x5 FILLER_195_867 ();
 b15zdnd00an1n01x5 FILLER_195_899 ();
 b15zdnd11an1n04x5 FILLER_195_924 ();
 b15zdnd11an1n64x5 FILLER_195_951 ();
 b15zdnd11an1n64x5 FILLER_195_1015 ();
 b15zdnd11an1n64x5 FILLER_195_1079 ();
 b15zdnd11an1n64x5 FILLER_195_1143 ();
 b15zdnd11an1n64x5 FILLER_195_1207 ();
 b15zdnd11an1n64x5 FILLER_195_1271 ();
 b15zdnd11an1n16x5 FILLER_195_1335 ();
 b15zdnd11an1n04x5 FILLER_195_1351 ();
 b15zdnd11an1n64x5 FILLER_195_1369 ();
 b15zdnd11an1n64x5 FILLER_195_1433 ();
 b15zdnd11an1n64x5 FILLER_195_1497 ();
 b15zdnd11an1n32x5 FILLER_195_1561 ();
 b15zdnd11an1n08x5 FILLER_195_1593 ();
 b15zdnd00an1n02x5 FILLER_195_1601 ();
 b15zdnd11an1n64x5 FILLER_195_1623 ();
 b15zdnd11an1n32x5 FILLER_195_1687 ();
 b15zdnd11an1n16x5 FILLER_195_1719 ();
 b15zdnd00an1n02x5 FILLER_195_1735 ();
 b15zdnd11an1n64x5 FILLER_195_1745 ();
 b15zdnd11an1n32x5 FILLER_195_1809 ();
 b15zdnd11an1n08x5 FILLER_195_1841 ();
 b15zdnd00an1n02x5 FILLER_195_1849 ();
 b15zdnd00an1n01x5 FILLER_195_1851 ();
 b15zdnd11an1n04x5 FILLER_195_1867 ();
 b15zdnd11an1n08x5 FILLER_195_1877 ();
 b15zdnd00an1n01x5 FILLER_195_1885 ();
 b15zdnd11an1n08x5 FILLER_195_1900 ();
 b15zdnd11an1n32x5 FILLER_195_1911 ();
 b15zdnd11an1n08x5 FILLER_195_1943 ();
 b15zdnd11an1n04x5 FILLER_195_1951 ();
 b15zdnd11an1n32x5 FILLER_195_1963 ();
 b15zdnd11an1n08x5 FILLER_195_1995 ();
 b15zdnd11an1n04x5 FILLER_195_2003 ();
 b15zdnd00an1n02x5 FILLER_195_2007 ();
 b15zdnd11an1n04x5 FILLER_195_2017 ();
 b15zdnd11an1n04x5 FILLER_195_2028 ();
 b15zdnd11an1n16x5 FILLER_195_2038 ();
 b15zdnd11an1n08x5 FILLER_195_2054 ();
 b15zdnd11an1n04x5 FILLER_195_2062 ();
 b15zdnd00an1n01x5 FILLER_195_2066 ();
 b15zdnd11an1n64x5 FILLER_195_2072 ();
 b15zdnd11an1n64x5 FILLER_195_2136 ();
 b15zdnd11an1n64x5 FILLER_195_2200 ();
 b15zdnd11an1n16x5 FILLER_195_2264 ();
 b15zdnd11an1n04x5 FILLER_195_2280 ();
 b15zdnd11an1n04x5 FILLER_196_8 ();
 b15zdnd11an1n64x5 FILLER_196_23 ();
 b15zdnd11an1n64x5 FILLER_196_87 ();
 b15zdnd11an1n64x5 FILLER_196_151 ();
 b15zdnd11an1n64x5 FILLER_196_215 ();
 b15zdnd11an1n64x5 FILLER_196_279 ();
 b15zdnd11an1n64x5 FILLER_196_343 ();
 b15zdnd11an1n32x5 FILLER_196_407 ();
 b15zdnd11an1n04x5 FILLER_196_439 ();
 b15zdnd00an1n02x5 FILLER_196_443 ();
 b15zdnd00an1n01x5 FILLER_196_445 ();
 b15zdnd11an1n64x5 FILLER_196_466 ();
 b15zdnd11an1n32x5 FILLER_196_530 ();
 b15zdnd11an1n16x5 FILLER_196_562 ();
 b15zdnd11an1n08x5 FILLER_196_578 ();
 b15zdnd00an1n02x5 FILLER_196_586 ();
 b15zdnd11an1n04x5 FILLER_196_611 ();
 b15zdnd11an1n64x5 FILLER_196_640 ();
 b15zdnd11an1n08x5 FILLER_196_704 ();
 b15zdnd11an1n04x5 FILLER_196_712 ();
 b15zdnd00an1n02x5 FILLER_196_716 ();
 b15zdnd11an1n64x5 FILLER_196_726 ();
 b15zdnd11an1n64x5 FILLER_196_790 ();
 b15zdnd11an1n64x5 FILLER_196_854 ();
 b15zdnd11an1n64x5 FILLER_196_918 ();
 b15zdnd11an1n32x5 FILLER_196_982 ();
 b15zdnd11an1n04x5 FILLER_196_1014 ();
 b15zdnd00an1n01x5 FILLER_196_1018 ();
 b15zdnd11an1n64x5 FILLER_196_1050 ();
 b15zdnd11an1n64x5 FILLER_196_1114 ();
 b15zdnd11an1n64x5 FILLER_196_1178 ();
 b15zdnd11an1n64x5 FILLER_196_1242 ();
 b15zdnd11an1n64x5 FILLER_196_1306 ();
 b15zdnd11an1n32x5 FILLER_196_1370 ();
 b15zdnd00an1n01x5 FILLER_196_1402 ();
 b15zdnd11an1n64x5 FILLER_196_1412 ();
 b15zdnd11an1n64x5 FILLER_196_1476 ();
 b15zdnd11an1n64x5 FILLER_196_1540 ();
 b15zdnd11an1n64x5 FILLER_196_1604 ();
 b15zdnd11an1n64x5 FILLER_196_1668 ();
 b15zdnd11an1n64x5 FILLER_196_1732 ();
 b15zdnd11an1n64x5 FILLER_196_1796 ();
 b15zdnd11an1n04x5 FILLER_196_1860 ();
 b15zdnd00an1n02x5 FILLER_196_1864 ();
 b15zdnd00an1n01x5 FILLER_196_1866 ();
 b15zdnd11an1n64x5 FILLER_196_1880 ();
 b15zdnd11an1n64x5 FILLER_196_1944 ();
 b15zdnd11an1n64x5 FILLER_196_2008 ();
 b15zdnd11an1n64x5 FILLER_196_2072 ();
 b15zdnd11an1n04x5 FILLER_196_2136 ();
 b15zdnd11an1n04x5 FILLER_196_2147 ();
 b15zdnd00an1n02x5 FILLER_196_2151 ();
 b15zdnd00an1n01x5 FILLER_196_2153 ();
 b15zdnd11an1n04x5 FILLER_196_2162 ();
 b15zdnd00an1n01x5 FILLER_196_2166 ();
 b15zdnd11an1n04x5 FILLER_196_2170 ();
 b15zdnd11an1n64x5 FILLER_196_2177 ();
 b15zdnd11an1n32x5 FILLER_196_2241 ();
 b15zdnd00an1n02x5 FILLER_196_2273 ();
 b15zdnd00an1n01x5 FILLER_196_2275 ();
 b15zdnd11an1n16x5 FILLER_197_0 ();
 b15zdnd11an1n08x5 FILLER_197_16 ();
 b15zdnd11an1n04x5 FILLER_197_24 ();
 b15zdnd00an1n01x5 FILLER_197_28 ();
 b15zdnd11an1n64x5 FILLER_197_36 ();
 b15zdnd11an1n64x5 FILLER_197_100 ();
 b15zdnd11an1n64x5 FILLER_197_164 ();
 b15zdnd11an1n08x5 FILLER_197_228 ();
 b15zdnd11an1n04x5 FILLER_197_236 ();
 b15zdnd00an1n02x5 FILLER_197_240 ();
 b15zdnd00an1n01x5 FILLER_197_242 ();
 b15zdnd11an1n64x5 FILLER_197_285 ();
 b15zdnd11an1n32x5 FILLER_197_349 ();
 b15zdnd11an1n16x5 FILLER_197_381 ();
 b15zdnd11an1n08x5 FILLER_197_397 ();
 b15zdnd11an1n04x5 FILLER_197_405 ();
 b15zdnd11an1n16x5 FILLER_197_421 ();
 b15zdnd11an1n04x5 FILLER_197_437 ();
 b15zdnd11an1n04x5 FILLER_197_461 ();
 b15zdnd11an1n64x5 FILLER_197_510 ();
 b15zdnd11an1n32x5 FILLER_197_574 ();
 b15zdnd11an1n04x5 FILLER_197_606 ();
 b15zdnd00an1n02x5 FILLER_197_610 ();
 b15zdnd11an1n64x5 FILLER_197_623 ();
 b15zdnd11an1n64x5 FILLER_197_687 ();
 b15zdnd11an1n64x5 FILLER_197_751 ();
 b15zdnd11an1n64x5 FILLER_197_815 ();
 b15zdnd11an1n64x5 FILLER_197_879 ();
 b15zdnd11an1n64x5 FILLER_197_943 ();
 b15zdnd00an1n02x5 FILLER_197_1007 ();
 b15zdnd00an1n01x5 FILLER_197_1009 ();
 b15zdnd11an1n32x5 FILLER_197_1028 ();
 b15zdnd11an1n16x5 FILLER_197_1060 ();
 b15zdnd11an1n08x5 FILLER_197_1076 ();
 b15zdnd11an1n04x5 FILLER_197_1084 ();
 b15zdnd11an1n04x5 FILLER_197_1113 ();
 b15zdnd11an1n32x5 FILLER_197_1127 ();
 b15zdnd11an1n16x5 FILLER_197_1159 ();
 b15zdnd11an1n08x5 FILLER_197_1175 ();
 b15zdnd00an1n02x5 FILLER_197_1183 ();
 b15zdnd00an1n01x5 FILLER_197_1185 ();
 b15zdnd11an1n64x5 FILLER_197_1210 ();
 b15zdnd11an1n64x5 FILLER_197_1274 ();
 b15zdnd11an1n64x5 FILLER_197_1338 ();
 b15zdnd11an1n64x5 FILLER_197_1402 ();
 b15zdnd11an1n64x5 FILLER_197_1466 ();
 b15zdnd11an1n64x5 FILLER_197_1530 ();
 b15zdnd11an1n64x5 FILLER_197_1594 ();
 b15zdnd11an1n32x5 FILLER_197_1658 ();
 b15zdnd11an1n04x5 FILLER_197_1690 ();
 b15zdnd00an1n01x5 FILLER_197_1694 ();
 b15zdnd11an1n08x5 FILLER_197_1709 ();
 b15zdnd11an1n04x5 FILLER_197_1717 ();
 b15zdnd00an1n02x5 FILLER_197_1721 ();
 b15zdnd00an1n01x5 FILLER_197_1723 ();
 b15zdnd11an1n32x5 FILLER_197_1728 ();
 b15zdnd11an1n04x5 FILLER_197_1760 ();
 b15zdnd00an1n01x5 FILLER_197_1764 ();
 b15zdnd11an1n64x5 FILLER_197_1769 ();
 b15zdnd11an1n64x5 FILLER_197_1833 ();
 b15zdnd11an1n32x5 FILLER_197_1897 ();
 b15zdnd11an1n16x5 FILLER_197_1929 ();
 b15zdnd11an1n08x5 FILLER_197_1945 ();
 b15zdnd00an1n02x5 FILLER_197_1953 ();
 b15zdnd11an1n64x5 FILLER_197_1960 ();
 b15zdnd11an1n64x5 FILLER_197_2024 ();
 b15zdnd11an1n32x5 FILLER_197_2088 ();
 b15zdnd11an1n16x5 FILLER_197_2120 ();
 b15zdnd11an1n08x5 FILLER_197_2136 ();
 b15zdnd11an1n04x5 FILLER_197_2144 ();
 b15zdnd00an1n01x5 FILLER_197_2148 ();
 b15zdnd11an1n64x5 FILLER_197_2201 ();
 b15zdnd11an1n16x5 FILLER_197_2265 ();
 b15zdnd00an1n02x5 FILLER_197_2281 ();
 b15zdnd00an1n01x5 FILLER_197_2283 ();
 b15zdnd11an1n64x5 FILLER_198_8 ();
 b15zdnd11an1n04x5 FILLER_198_72 ();
 b15zdnd11an1n64x5 FILLER_198_121 ();
 b15zdnd11an1n32x5 FILLER_198_185 ();
 b15zdnd11an1n16x5 FILLER_198_217 ();
 b15zdnd11an1n04x5 FILLER_198_233 ();
 b15zdnd11an1n64x5 FILLER_198_240 ();
 b15zdnd11an1n64x5 FILLER_198_304 ();
 b15zdnd11an1n32x5 FILLER_198_368 ();
 b15zdnd11an1n16x5 FILLER_198_400 ();
 b15zdnd11an1n04x5 FILLER_198_416 ();
 b15zdnd00an1n02x5 FILLER_198_420 ();
 b15zdnd00an1n01x5 FILLER_198_422 ();
 b15zdnd11an1n64x5 FILLER_198_443 ();
 b15zdnd11an1n64x5 FILLER_198_507 ();
 b15zdnd11an1n32x5 FILLER_198_571 ();
 b15zdnd11an1n16x5 FILLER_198_603 ();
 b15zdnd11an1n08x5 FILLER_198_619 ();
 b15zdnd11an1n04x5 FILLER_198_627 ();
 b15zdnd00an1n02x5 FILLER_198_631 ();
 b15zdnd00an1n01x5 FILLER_198_633 ();
 b15zdnd11an1n32x5 FILLER_198_640 ();
 b15zdnd11an1n16x5 FILLER_198_672 ();
 b15zdnd00an1n02x5 FILLER_198_688 ();
 b15zdnd00an1n02x5 FILLER_198_716 ();
 b15zdnd11an1n64x5 FILLER_198_726 ();
 b15zdnd11an1n64x5 FILLER_198_790 ();
 b15zdnd11an1n64x5 FILLER_198_854 ();
 b15zdnd11an1n64x5 FILLER_198_918 ();
 b15zdnd11an1n64x5 FILLER_198_982 ();
 b15zdnd11an1n64x5 FILLER_198_1046 ();
 b15zdnd11an1n64x5 FILLER_198_1110 ();
 b15zdnd11an1n64x5 FILLER_198_1174 ();
 b15zdnd11an1n64x5 FILLER_198_1238 ();
 b15zdnd11an1n64x5 FILLER_198_1302 ();
 b15zdnd11an1n64x5 FILLER_198_1366 ();
 b15zdnd11an1n64x5 FILLER_198_1430 ();
 b15zdnd11an1n64x5 FILLER_198_1494 ();
 b15zdnd11an1n64x5 FILLER_198_1558 ();
 b15zdnd11an1n64x5 FILLER_198_1622 ();
 b15zdnd11an1n64x5 FILLER_198_1686 ();
 b15zdnd11an1n16x5 FILLER_198_1750 ();
 b15zdnd11an1n04x5 FILLER_198_1766 ();
 b15zdnd00an1n02x5 FILLER_198_1770 ();
 b15zdnd00an1n01x5 FILLER_198_1772 ();
 b15zdnd11an1n64x5 FILLER_198_1777 ();
 b15zdnd11an1n64x5 FILLER_198_1841 ();
 b15zdnd11an1n32x5 FILLER_198_1905 ();
 b15zdnd11an1n04x5 FILLER_198_1937 ();
 b15zdnd11an1n64x5 FILLER_198_1948 ();
 b15zdnd11an1n32x5 FILLER_198_2012 ();
 b15zdnd11an1n16x5 FILLER_198_2044 ();
 b15zdnd00an1n01x5 FILLER_198_2060 ();
 b15zdnd11an1n64x5 FILLER_198_2064 ();
 b15zdnd11an1n16x5 FILLER_198_2128 ();
 b15zdnd11an1n08x5 FILLER_198_2144 ();
 b15zdnd00an1n02x5 FILLER_198_2152 ();
 b15zdnd11an1n08x5 FILLER_198_2162 ();
 b15zdnd11an1n04x5 FILLER_198_2170 ();
 b15zdnd11an1n64x5 FILLER_198_2177 ();
 b15zdnd11an1n08x5 FILLER_198_2241 ();
 b15zdnd11an1n04x5 FILLER_198_2269 ();
 b15zdnd00an1n02x5 FILLER_198_2273 ();
 b15zdnd00an1n01x5 FILLER_198_2275 ();
 b15zdnd11an1n16x5 FILLER_199_0 ();
 b15zdnd11an1n08x5 FILLER_199_16 ();
 b15zdnd00an1n02x5 FILLER_199_24 ();
 b15zdnd11an1n64x5 FILLER_199_34 ();
 b15zdnd11an1n64x5 FILLER_199_98 ();
 b15zdnd11an1n32x5 FILLER_199_162 ();
 b15zdnd11an1n16x5 FILLER_199_194 ();
 b15zdnd11an1n64x5 FILLER_199_262 ();
 b15zdnd00an1n01x5 FILLER_199_326 ();
 b15zdnd11an1n64x5 FILLER_199_349 ();
 b15zdnd11an1n64x5 FILLER_199_413 ();
 b15zdnd11an1n64x5 FILLER_199_477 ();
 b15zdnd11an1n64x5 FILLER_199_541 ();
 b15zdnd11an1n16x5 FILLER_199_605 ();
 b15zdnd11an1n08x5 FILLER_199_621 ();
 b15zdnd00an1n01x5 FILLER_199_629 ();
 b15zdnd11an1n32x5 FILLER_199_645 ();
 b15zdnd11an1n08x5 FILLER_199_677 ();
 b15zdnd11an1n04x5 FILLER_199_685 ();
 b15zdnd00an1n01x5 FILLER_199_689 ();
 b15zdnd11an1n64x5 FILLER_199_705 ();
 b15zdnd11an1n16x5 FILLER_199_769 ();
 b15zdnd11an1n08x5 FILLER_199_785 ();
 b15zdnd11an1n04x5 FILLER_199_793 ();
 b15zdnd00an1n02x5 FILLER_199_797 ();
 b15zdnd00an1n01x5 FILLER_199_799 ();
 b15zdnd11an1n32x5 FILLER_199_812 ();
 b15zdnd11an1n04x5 FILLER_199_844 ();
 b15zdnd00an1n02x5 FILLER_199_848 ();
 b15zdnd11an1n64x5 FILLER_199_866 ();
 b15zdnd11an1n64x5 FILLER_199_930 ();
 b15zdnd11an1n64x5 FILLER_199_994 ();
 b15zdnd11an1n64x5 FILLER_199_1058 ();
 b15zdnd11an1n64x5 FILLER_199_1122 ();
 b15zdnd00an1n02x5 FILLER_199_1186 ();
 b15zdnd00an1n01x5 FILLER_199_1188 ();
 b15zdnd11an1n64x5 FILLER_199_1220 ();
 b15zdnd11an1n64x5 FILLER_199_1284 ();
 b15zdnd11an1n64x5 FILLER_199_1348 ();
 b15zdnd11an1n64x5 FILLER_199_1412 ();
 b15zdnd11an1n64x5 FILLER_199_1476 ();
 b15zdnd11an1n08x5 FILLER_199_1540 ();
 b15zdnd11an1n08x5 FILLER_199_1568 ();
 b15zdnd11an1n04x5 FILLER_199_1576 ();
 b15zdnd00an1n02x5 FILLER_199_1580 ();
 b15zdnd00an1n01x5 FILLER_199_1582 ();
 b15zdnd11an1n64x5 FILLER_199_1593 ();
 b15zdnd11an1n16x5 FILLER_199_1657 ();
 b15zdnd11an1n08x5 FILLER_199_1673 ();
 b15zdnd11an1n64x5 FILLER_199_1689 ();
 b15zdnd11an1n16x5 FILLER_199_1753 ();
 b15zdnd11an1n04x5 FILLER_199_1769 ();
 b15zdnd11an1n64x5 FILLER_199_1777 ();
 b15zdnd11an1n64x5 FILLER_199_1841 ();
 b15zdnd11an1n64x5 FILLER_199_1905 ();
 b15zdnd11an1n64x5 FILLER_199_1969 ();
 b15zdnd11an1n16x5 FILLER_199_2033 ();
 b15zdnd11an1n08x5 FILLER_199_2049 ();
 b15zdnd11an1n04x5 FILLER_199_2057 ();
 b15zdnd11an1n32x5 FILLER_199_2064 ();
 b15zdnd11an1n64x5 FILLER_199_2101 ();
 b15zdnd11an1n64x5 FILLER_199_2165 ();
 b15zdnd11an1n32x5 FILLER_199_2229 ();
 b15zdnd11an1n16x5 FILLER_199_2261 ();
 b15zdnd11an1n04x5 FILLER_199_2277 ();
 b15zdnd00an1n02x5 FILLER_199_2281 ();
 b15zdnd00an1n01x5 FILLER_199_2283 ();
 b15zdnd11an1n16x5 FILLER_200_8 ();
 b15zdnd11an1n04x5 FILLER_200_24 ();
 b15zdnd11an1n64x5 FILLER_200_42 ();
 b15zdnd11an1n64x5 FILLER_200_106 ();
 b15zdnd11an1n16x5 FILLER_200_170 ();
 b15zdnd00an1n02x5 FILLER_200_186 ();
 b15zdnd00an1n01x5 FILLER_200_188 ();
 b15zdnd11an1n16x5 FILLER_200_197 ();
 b15zdnd11an1n08x5 FILLER_200_213 ();
 b15zdnd11an1n04x5 FILLER_200_221 ();
 b15zdnd00an1n02x5 FILLER_200_225 ();
 b15zdnd00an1n01x5 FILLER_200_227 ();
 b15zdnd11an1n04x5 FILLER_200_231 ();
 b15zdnd11an1n64x5 FILLER_200_238 ();
 b15zdnd11an1n32x5 FILLER_200_302 ();
 b15zdnd11an1n16x5 FILLER_200_334 ();
 b15zdnd11an1n08x5 FILLER_200_350 ();
 b15zdnd00an1n01x5 FILLER_200_358 ();
 b15zdnd11an1n64x5 FILLER_200_372 ();
 b15zdnd11an1n64x5 FILLER_200_436 ();
 b15zdnd11an1n32x5 FILLER_200_500 ();
 b15zdnd00an1n02x5 FILLER_200_532 ();
 b15zdnd11an1n32x5 FILLER_200_576 ();
 b15zdnd11an1n04x5 FILLER_200_608 ();
 b15zdnd00an1n02x5 FILLER_200_612 ();
 b15zdnd11an1n64x5 FILLER_200_629 ();
 b15zdnd11an1n16x5 FILLER_200_693 ();
 b15zdnd11an1n08x5 FILLER_200_709 ();
 b15zdnd00an1n01x5 FILLER_200_717 ();
 b15zdnd11an1n64x5 FILLER_200_726 ();
 b15zdnd11an1n08x5 FILLER_200_790 ();
 b15zdnd11an1n04x5 FILLER_200_798 ();
 b15zdnd11an1n64x5 FILLER_200_817 ();
 b15zdnd11an1n64x5 FILLER_200_881 ();
 b15zdnd11an1n32x5 FILLER_200_945 ();
 b15zdnd11an1n08x5 FILLER_200_977 ();
 b15zdnd11an1n04x5 FILLER_200_985 ();
 b15zdnd00an1n01x5 FILLER_200_989 ();
 b15zdnd11an1n64x5 FILLER_200_1008 ();
 b15zdnd11an1n16x5 FILLER_200_1072 ();
 b15zdnd11an1n04x5 FILLER_200_1088 ();
 b15zdnd00an1n02x5 FILLER_200_1092 ();
 b15zdnd00an1n01x5 FILLER_200_1094 ();
 b15zdnd11an1n04x5 FILLER_200_1110 ();
 b15zdnd11an1n64x5 FILLER_200_1129 ();
 b15zdnd11an1n64x5 FILLER_200_1193 ();
 b15zdnd11an1n64x5 FILLER_200_1257 ();
 b15zdnd11an1n64x5 FILLER_200_1321 ();
 b15zdnd11an1n32x5 FILLER_200_1385 ();
 b15zdnd00an1n02x5 FILLER_200_1417 ();
 b15zdnd00an1n01x5 FILLER_200_1419 ();
 b15zdnd11an1n64x5 FILLER_200_1423 ();
 b15zdnd11an1n32x5 FILLER_200_1487 ();
 b15zdnd11an1n04x5 FILLER_200_1519 ();
 b15zdnd00an1n02x5 FILLER_200_1523 ();
 b15zdnd00an1n01x5 FILLER_200_1525 ();
 b15zdnd11an1n64x5 FILLER_200_1529 ();
 b15zdnd11an1n64x5 FILLER_200_1593 ();
 b15zdnd11an1n64x5 FILLER_200_1657 ();
 b15zdnd11an1n64x5 FILLER_200_1721 ();
 b15zdnd11an1n64x5 FILLER_200_1785 ();
 b15zdnd11an1n64x5 FILLER_200_1849 ();
 b15zdnd11an1n64x5 FILLER_200_1913 ();
 b15zdnd11an1n32x5 FILLER_200_1977 ();
 b15zdnd11an1n16x5 FILLER_200_2009 ();
 b15zdnd11an1n08x5 FILLER_200_2025 ();
 b15zdnd00an1n02x5 FILLER_200_2033 ();
 b15zdnd00an1n01x5 FILLER_200_2035 ();
 b15zdnd11an1n32x5 FILLER_200_2088 ();
 b15zdnd11an1n08x5 FILLER_200_2127 ();
 b15zdnd11an1n04x5 FILLER_200_2135 ();
 b15zdnd00an1n01x5 FILLER_200_2139 ();
 b15zdnd00an1n02x5 FILLER_200_2152 ();
 b15zdnd11an1n64x5 FILLER_200_2162 ();
 b15zdnd11an1n32x5 FILLER_200_2226 ();
 b15zdnd11an1n16x5 FILLER_200_2258 ();
 b15zdnd00an1n02x5 FILLER_200_2274 ();
 b15zdnd11an1n64x5 FILLER_201_0 ();
 b15zdnd11an1n64x5 FILLER_201_64 ();
 b15zdnd11an1n32x5 FILLER_201_128 ();
 b15zdnd11an1n08x5 FILLER_201_160 ();
 b15zdnd00an1n02x5 FILLER_201_168 ();
 b15zdnd11an1n64x5 FILLER_201_197 ();
 b15zdnd11an1n64x5 FILLER_201_261 ();
 b15zdnd11an1n64x5 FILLER_201_325 ();
 b15zdnd11an1n64x5 FILLER_201_389 ();
 b15zdnd11an1n64x5 FILLER_201_453 ();
 b15zdnd11an1n16x5 FILLER_201_517 ();
 b15zdnd11an1n32x5 FILLER_201_575 ();
 b15zdnd11an1n08x5 FILLER_201_607 ();
 b15zdnd11an1n04x5 FILLER_201_615 ();
 b15zdnd00an1n01x5 FILLER_201_619 ();
 b15zdnd11an1n64x5 FILLER_201_638 ();
 b15zdnd11an1n64x5 FILLER_201_702 ();
 b15zdnd11an1n16x5 FILLER_201_766 ();
 b15zdnd11an1n08x5 FILLER_201_782 ();
 b15zdnd11an1n04x5 FILLER_201_790 ();
 b15zdnd00an1n01x5 FILLER_201_794 ();
 b15zdnd11an1n64x5 FILLER_201_821 ();
 b15zdnd11an1n64x5 FILLER_201_885 ();
 b15zdnd11an1n64x5 FILLER_201_949 ();
 b15zdnd11an1n64x5 FILLER_201_1013 ();
 b15zdnd11an1n64x5 FILLER_201_1077 ();
 b15zdnd11an1n04x5 FILLER_201_1151 ();
 b15zdnd00an1n01x5 FILLER_201_1155 ();
 b15zdnd11an1n64x5 FILLER_201_1173 ();
 b15zdnd11an1n64x5 FILLER_201_1237 ();
 b15zdnd11an1n64x5 FILLER_201_1301 ();
 b15zdnd11an1n16x5 FILLER_201_1365 ();
 b15zdnd11an1n04x5 FILLER_201_1381 ();
 b15zdnd00an1n02x5 FILLER_201_1385 ();
 b15zdnd00an1n01x5 FILLER_201_1387 ();
 b15zdnd11an1n04x5 FILLER_201_1415 ();
 b15zdnd11an1n64x5 FILLER_201_1422 ();
 b15zdnd11an1n08x5 FILLER_201_1486 ();
 b15zdnd11an1n04x5 FILLER_201_1494 ();
 b15zdnd11an1n64x5 FILLER_201_1550 ();
 b15zdnd11an1n32x5 FILLER_201_1614 ();
 b15zdnd11an1n08x5 FILLER_201_1646 ();
 b15zdnd11an1n64x5 FILLER_201_1658 ();
 b15zdnd11an1n64x5 FILLER_201_1722 ();
 b15zdnd11an1n64x5 FILLER_201_1786 ();
 b15zdnd11an1n64x5 FILLER_201_1850 ();
 b15zdnd11an1n64x5 FILLER_201_1914 ();
 b15zdnd11an1n64x5 FILLER_201_1978 ();
 b15zdnd11an1n16x5 FILLER_201_2042 ();
 b15zdnd00an1n02x5 FILLER_201_2058 ();
 b15zdnd00an1n01x5 FILLER_201_2060 ();
 b15zdnd11an1n64x5 FILLER_201_2064 ();
 b15zdnd11an1n64x5 FILLER_201_2128 ();
 b15zdnd11an1n64x5 FILLER_201_2192 ();
 b15zdnd11an1n16x5 FILLER_201_2256 ();
 b15zdnd11an1n08x5 FILLER_201_2272 ();
 b15zdnd11an1n04x5 FILLER_201_2280 ();
 b15zdnd00an1n02x5 FILLER_202_8 ();
 b15zdnd11an1n64x5 FILLER_202_21 ();
 b15zdnd11an1n64x5 FILLER_202_85 ();
 b15zdnd11an1n16x5 FILLER_202_149 ();
 b15zdnd11an1n08x5 FILLER_202_165 ();
 b15zdnd11an1n04x5 FILLER_202_173 ();
 b15zdnd11an1n64x5 FILLER_202_181 ();
 b15zdnd11an1n64x5 FILLER_202_245 ();
 b15zdnd11an1n64x5 FILLER_202_309 ();
 b15zdnd00an1n02x5 FILLER_202_373 ();
 b15zdnd11an1n04x5 FILLER_202_379 ();
 b15zdnd11an1n64x5 FILLER_202_393 ();
 b15zdnd11an1n64x5 FILLER_202_457 ();
 b15zdnd11an1n16x5 FILLER_202_521 ();
 b15zdnd00an1n02x5 FILLER_202_537 ();
 b15zdnd11an1n32x5 FILLER_202_557 ();
 b15zdnd11an1n16x5 FILLER_202_589 ();
 b15zdnd11an1n08x5 FILLER_202_605 ();
 b15zdnd11an1n04x5 FILLER_202_613 ();
 b15zdnd11an1n64x5 FILLER_202_632 ();
 b15zdnd11an1n16x5 FILLER_202_696 ();
 b15zdnd11an1n04x5 FILLER_202_712 ();
 b15zdnd00an1n02x5 FILLER_202_716 ();
 b15zdnd11an1n32x5 FILLER_202_726 ();
 b15zdnd11an1n16x5 FILLER_202_758 ();
 b15zdnd00an1n02x5 FILLER_202_774 ();
 b15zdnd11an1n16x5 FILLER_202_807 ();
 b15zdnd11an1n04x5 FILLER_202_823 ();
 b15zdnd00an1n02x5 FILLER_202_827 ();
 b15zdnd00an1n01x5 FILLER_202_829 ();
 b15zdnd11an1n64x5 FILLER_202_839 ();
 b15zdnd11an1n64x5 FILLER_202_903 ();
 b15zdnd11an1n64x5 FILLER_202_967 ();
 b15zdnd11an1n64x5 FILLER_202_1031 ();
 b15zdnd11an1n64x5 FILLER_202_1095 ();
 b15zdnd11an1n04x5 FILLER_202_1159 ();
 b15zdnd00an1n02x5 FILLER_202_1163 ();
 b15zdnd00an1n01x5 FILLER_202_1165 ();
 b15zdnd11an1n64x5 FILLER_202_1197 ();
 b15zdnd11an1n16x5 FILLER_202_1261 ();
 b15zdnd11an1n08x5 FILLER_202_1277 ();
 b15zdnd11an1n04x5 FILLER_202_1285 ();
 b15zdnd11an1n64x5 FILLER_202_1300 ();
 b15zdnd11an1n16x5 FILLER_202_1364 ();
 b15zdnd11an1n08x5 FILLER_202_1380 ();
 b15zdnd11an1n04x5 FILLER_202_1391 ();
 b15zdnd11an1n32x5 FILLER_202_1447 ();
 b15zdnd00an1n02x5 FILLER_202_1479 ();
 b15zdnd00an1n01x5 FILLER_202_1481 ();
 b15zdnd11an1n04x5 FILLER_202_1534 ();
 b15zdnd11an1n64x5 FILLER_202_1541 ();
 b15zdnd11an1n32x5 FILLER_202_1605 ();
 b15zdnd11an1n16x5 FILLER_202_1637 ();
 b15zdnd00an1n02x5 FILLER_202_1653 ();
 b15zdnd00an1n01x5 FILLER_202_1655 ();
 b15zdnd11an1n64x5 FILLER_202_1660 ();
 b15zdnd11an1n64x5 FILLER_202_1724 ();
 b15zdnd11an1n64x5 FILLER_202_1788 ();
 b15zdnd11an1n32x5 FILLER_202_1852 ();
 b15zdnd11an1n08x5 FILLER_202_1884 ();
 b15zdnd00an1n02x5 FILLER_202_1892 ();
 b15zdnd00an1n01x5 FILLER_202_1894 ();
 b15zdnd11an1n64x5 FILLER_202_1937 ();
 b15zdnd11an1n64x5 FILLER_202_2001 ();
 b15zdnd11an1n64x5 FILLER_202_2065 ();
 b15zdnd11an1n16x5 FILLER_202_2129 ();
 b15zdnd11an1n08x5 FILLER_202_2145 ();
 b15zdnd00an1n01x5 FILLER_202_2153 ();
 b15zdnd11an1n08x5 FILLER_202_2162 ();
 b15zdnd00an1n02x5 FILLER_202_2170 ();
 b15zdnd11an1n32x5 FILLER_202_2214 ();
 b15zdnd11an1n16x5 FILLER_202_2246 ();
 b15zdnd11an1n08x5 FILLER_202_2262 ();
 b15zdnd11an1n04x5 FILLER_202_2270 ();
 b15zdnd00an1n02x5 FILLER_202_2274 ();
 b15zdnd11an1n64x5 FILLER_203_0 ();
 b15zdnd11an1n64x5 FILLER_203_64 ();
 b15zdnd11an1n64x5 FILLER_203_128 ();
 b15zdnd11an1n64x5 FILLER_203_192 ();
 b15zdnd11an1n64x5 FILLER_203_256 ();
 b15zdnd11an1n64x5 FILLER_203_320 ();
 b15zdnd11an1n64x5 FILLER_203_384 ();
 b15zdnd11an1n64x5 FILLER_203_448 ();
 b15zdnd11an1n64x5 FILLER_203_512 ();
 b15zdnd11an1n32x5 FILLER_203_576 ();
 b15zdnd11an1n16x5 FILLER_203_608 ();
 b15zdnd11an1n04x5 FILLER_203_624 ();
 b15zdnd00an1n02x5 FILLER_203_628 ();
 b15zdnd11an1n64x5 FILLER_203_654 ();
 b15zdnd11an1n64x5 FILLER_203_718 ();
 b15zdnd11an1n16x5 FILLER_203_782 ();
 b15zdnd11an1n08x5 FILLER_203_798 ();
 b15zdnd11an1n04x5 FILLER_203_806 ();
 b15zdnd11an1n64x5 FILLER_203_822 ();
 b15zdnd11an1n16x5 FILLER_203_886 ();
 b15zdnd11an1n08x5 FILLER_203_902 ();
 b15zdnd11an1n04x5 FILLER_203_910 ();
 b15zdnd00an1n02x5 FILLER_203_914 ();
 b15zdnd11an1n32x5 FILLER_203_940 ();
 b15zdnd11an1n64x5 FILLER_203_992 ();
 b15zdnd11an1n64x5 FILLER_203_1056 ();
 b15zdnd11an1n64x5 FILLER_203_1120 ();
 b15zdnd11an1n64x5 FILLER_203_1184 ();
 b15zdnd11an1n64x5 FILLER_203_1248 ();
 b15zdnd11an1n64x5 FILLER_203_1312 ();
 b15zdnd11an1n32x5 FILLER_203_1376 ();
 b15zdnd11an1n08x5 FILLER_203_1408 ();
 b15zdnd11an1n04x5 FILLER_203_1416 ();
 b15zdnd11an1n64x5 FILLER_203_1423 ();
 b15zdnd11an1n08x5 FILLER_203_1487 ();
 b15zdnd11an1n04x5 FILLER_203_1495 ();
 b15zdnd00an1n01x5 FILLER_203_1499 ();
 b15zdnd11an1n04x5 FILLER_203_1503 ();
 b15zdnd11an1n08x5 FILLER_203_1510 ();
 b15zdnd00an1n02x5 FILLER_203_1518 ();
 b15zdnd00an1n01x5 FILLER_203_1520 ();
 b15zdnd11an1n64x5 FILLER_203_1524 ();
 b15zdnd11an1n64x5 FILLER_203_1588 ();
 b15zdnd11an1n16x5 FILLER_203_1652 ();
 b15zdnd00an1n01x5 FILLER_203_1668 ();
 b15zdnd11an1n16x5 FILLER_203_1683 ();
 b15zdnd11an1n08x5 FILLER_203_1699 ();
 b15zdnd00an1n01x5 FILLER_203_1707 ();
 b15zdnd11an1n64x5 FILLER_203_1750 ();
 b15zdnd11an1n64x5 FILLER_203_1814 ();
 b15zdnd11an1n64x5 FILLER_203_1878 ();
 b15zdnd11an1n64x5 FILLER_203_1942 ();
 b15zdnd11an1n64x5 FILLER_203_2006 ();
 b15zdnd11an1n64x5 FILLER_203_2070 ();
 b15zdnd11an1n16x5 FILLER_203_2134 ();
 b15zdnd00an1n01x5 FILLER_203_2150 ();
 b15zdnd11an1n64x5 FILLER_203_2193 ();
 b15zdnd11an1n16x5 FILLER_203_2257 ();
 b15zdnd11an1n04x5 FILLER_203_2273 ();
 b15zdnd00an1n02x5 FILLER_203_2281 ();
 b15zdnd00an1n01x5 FILLER_203_2283 ();
 b15zdnd11an1n64x5 FILLER_204_8 ();
 b15zdnd11an1n64x5 FILLER_204_72 ();
 b15zdnd11an1n64x5 FILLER_204_136 ();
 b15zdnd11an1n64x5 FILLER_204_200 ();
 b15zdnd11an1n64x5 FILLER_204_264 ();
 b15zdnd11an1n64x5 FILLER_204_328 ();
 b15zdnd11an1n64x5 FILLER_204_392 ();
 b15zdnd11an1n64x5 FILLER_204_456 ();
 b15zdnd11an1n64x5 FILLER_204_520 ();
 b15zdnd11an1n64x5 FILLER_204_584 ();
 b15zdnd11an1n64x5 FILLER_204_648 ();
 b15zdnd11an1n04x5 FILLER_204_712 ();
 b15zdnd00an1n02x5 FILLER_204_716 ();
 b15zdnd11an1n64x5 FILLER_204_726 ();
 b15zdnd11an1n32x5 FILLER_204_790 ();
 b15zdnd11an1n04x5 FILLER_204_822 ();
 b15zdnd00an1n02x5 FILLER_204_826 ();
 b15zdnd00an1n01x5 FILLER_204_828 ();
 b15zdnd11an1n04x5 FILLER_204_843 ();
 b15zdnd11an1n64x5 FILLER_204_857 ();
 b15zdnd11an1n16x5 FILLER_204_921 ();
 b15zdnd00an1n02x5 FILLER_204_937 ();
 b15zdnd00an1n01x5 FILLER_204_939 ();
 b15zdnd11an1n16x5 FILLER_204_950 ();
 b15zdnd11an1n08x5 FILLER_204_966 ();
 b15zdnd11an1n04x5 FILLER_204_974 ();
 b15zdnd00an1n02x5 FILLER_204_978 ();
 b15zdnd11an1n04x5 FILLER_204_998 ();
 b15zdnd11an1n16x5 FILLER_204_1017 ();
 b15zdnd11an1n08x5 FILLER_204_1033 ();
 b15zdnd00an1n01x5 FILLER_204_1041 ();
 b15zdnd11an1n64x5 FILLER_204_1052 ();
 b15zdnd11an1n64x5 FILLER_204_1116 ();
 b15zdnd11an1n64x5 FILLER_204_1180 ();
 b15zdnd11an1n08x5 FILLER_204_1244 ();
 b15zdnd11an1n04x5 FILLER_204_1252 ();
 b15zdnd00an1n02x5 FILLER_204_1256 ();
 b15zdnd11an1n04x5 FILLER_204_1261 ();
 b15zdnd11an1n64x5 FILLER_204_1268 ();
 b15zdnd11an1n64x5 FILLER_204_1332 ();
 b15zdnd11an1n64x5 FILLER_204_1396 ();
 b15zdnd11an1n32x5 FILLER_204_1460 ();
 b15zdnd11an1n08x5 FILLER_204_1492 ();
 b15zdnd00an1n02x5 FILLER_204_1500 ();
 b15zdnd11an1n64x5 FILLER_204_1505 ();
 b15zdnd11an1n64x5 FILLER_204_1569 ();
 b15zdnd11an1n64x5 FILLER_204_1633 ();
 b15zdnd11an1n16x5 FILLER_204_1697 ();
 b15zdnd11an1n08x5 FILLER_204_1713 ();
 b15zdnd11an1n04x5 FILLER_204_1721 ();
 b15zdnd11an1n04x5 FILLER_204_1767 ();
 b15zdnd11an1n64x5 FILLER_204_1775 ();
 b15zdnd11an1n64x5 FILLER_204_1839 ();
 b15zdnd11an1n64x5 FILLER_204_1903 ();
 b15zdnd11an1n64x5 FILLER_204_1967 ();
 b15zdnd11an1n64x5 FILLER_204_2031 ();
 b15zdnd11an1n16x5 FILLER_204_2095 ();
 b15zdnd11an1n04x5 FILLER_204_2111 ();
 b15zdnd00an1n02x5 FILLER_204_2115 ();
 b15zdnd11an1n08x5 FILLER_204_2144 ();
 b15zdnd00an1n02x5 FILLER_204_2152 ();
 b15zdnd11an1n64x5 FILLER_204_2162 ();
 b15zdnd11an1n16x5 FILLER_204_2226 ();
 b15zdnd11an1n08x5 FILLER_204_2242 ();
 b15zdnd11an1n04x5 FILLER_204_2250 ();
 b15zdnd00an1n02x5 FILLER_204_2254 ();
 b15zdnd11an1n04x5 FILLER_204_2260 ();
 b15zdnd00an1n02x5 FILLER_204_2264 ();
 b15zdnd00an1n02x5 FILLER_204_2274 ();
 b15zdnd11an1n64x5 FILLER_205_0 ();
 b15zdnd11an1n64x5 FILLER_205_64 ();
 b15zdnd11an1n64x5 FILLER_205_128 ();
 b15zdnd11an1n64x5 FILLER_205_192 ();
 b15zdnd11an1n64x5 FILLER_205_256 ();
 b15zdnd11an1n64x5 FILLER_205_320 ();
 b15zdnd11an1n64x5 FILLER_205_384 ();
 b15zdnd11an1n64x5 FILLER_205_448 ();
 b15zdnd11an1n64x5 FILLER_205_512 ();
 b15zdnd11an1n64x5 FILLER_205_576 ();
 b15zdnd11an1n64x5 FILLER_205_640 ();
 b15zdnd11an1n64x5 FILLER_205_704 ();
 b15zdnd11an1n16x5 FILLER_205_768 ();
 b15zdnd11an1n08x5 FILLER_205_784 ();
 b15zdnd11an1n04x5 FILLER_205_792 ();
 b15zdnd00an1n01x5 FILLER_205_796 ();
 b15zdnd11an1n04x5 FILLER_205_809 ();
 b15zdnd11an1n32x5 FILLER_205_827 ();
 b15zdnd11an1n04x5 FILLER_205_859 ();
 b15zdnd00an1n02x5 FILLER_205_863 ();
 b15zdnd11an1n16x5 FILLER_205_875 ();
 b15zdnd11an1n16x5 FILLER_205_911 ();
 b15zdnd11an1n04x5 FILLER_205_927 ();
 b15zdnd00an1n01x5 FILLER_205_931 ();
 b15zdnd11an1n64x5 FILLER_205_947 ();
 b15zdnd11an1n64x5 FILLER_205_1011 ();
 b15zdnd11an1n64x5 FILLER_205_1075 ();
 b15zdnd11an1n04x5 FILLER_205_1139 ();
 b15zdnd00an1n01x5 FILLER_205_1143 ();
 b15zdnd11an1n32x5 FILLER_205_1152 ();
 b15zdnd11an1n08x5 FILLER_205_1184 ();
 b15zdnd11an1n16x5 FILLER_205_1210 ();
 b15zdnd11an1n08x5 FILLER_205_1226 ();
 b15zdnd11an1n04x5 FILLER_205_1234 ();
 b15zdnd00an1n02x5 FILLER_205_1238 ();
 b15zdnd11an1n64x5 FILLER_205_1292 ();
 b15zdnd11an1n64x5 FILLER_205_1356 ();
 b15zdnd11an1n64x5 FILLER_205_1420 ();
 b15zdnd11an1n64x5 FILLER_205_1484 ();
 b15zdnd11an1n64x5 FILLER_205_1548 ();
 b15zdnd11an1n64x5 FILLER_205_1612 ();
 b15zdnd11an1n64x5 FILLER_205_1676 ();
 b15zdnd11an1n64x5 FILLER_205_1740 ();
 b15zdnd11an1n64x5 FILLER_205_1804 ();
 b15zdnd11an1n32x5 FILLER_205_1868 ();
 b15zdnd11an1n16x5 FILLER_205_1900 ();
 b15zdnd11an1n08x5 FILLER_205_1916 ();
 b15zdnd11an1n04x5 FILLER_205_1924 ();
 b15zdnd00an1n02x5 FILLER_205_1928 ();
 b15zdnd11an1n64x5 FILLER_205_1972 ();
 b15zdnd11an1n64x5 FILLER_205_2036 ();
 b15zdnd11an1n16x5 FILLER_205_2100 ();
 b15zdnd00an1n01x5 FILLER_205_2116 ();
 b15zdnd11an1n64x5 FILLER_205_2120 ();
 b15zdnd11an1n32x5 FILLER_205_2184 ();
 b15zdnd11an1n16x5 FILLER_205_2216 ();
 b15zdnd11an1n08x5 FILLER_205_2232 ();
 b15zdnd00an1n02x5 FILLER_205_2282 ();
 b15zdnd11an1n32x5 FILLER_206_8 ();
 b15zdnd11an1n16x5 FILLER_206_40 ();
 b15zdnd11an1n04x5 FILLER_206_56 ();
 b15zdnd00an1n02x5 FILLER_206_60 ();
 b15zdnd11an1n64x5 FILLER_206_93 ();
 b15zdnd11an1n64x5 FILLER_206_157 ();
 b15zdnd11an1n64x5 FILLER_206_221 ();
 b15zdnd11an1n64x5 FILLER_206_285 ();
 b15zdnd11an1n64x5 FILLER_206_349 ();
 b15zdnd11an1n64x5 FILLER_206_413 ();
 b15zdnd11an1n64x5 FILLER_206_477 ();
 b15zdnd11an1n64x5 FILLER_206_541 ();
 b15zdnd11an1n64x5 FILLER_206_605 ();
 b15zdnd11an1n32x5 FILLER_206_669 ();
 b15zdnd00an1n01x5 FILLER_206_701 ();
 b15zdnd11an1n08x5 FILLER_206_710 ();
 b15zdnd11an1n64x5 FILLER_206_726 ();
 b15zdnd11an1n08x5 FILLER_206_790 ();
 b15zdnd11an1n04x5 FILLER_206_798 ();
 b15zdnd00an1n02x5 FILLER_206_802 ();
 b15zdnd11an1n32x5 FILLER_206_815 ();
 b15zdnd11an1n08x5 FILLER_206_847 ();
 b15zdnd11an1n64x5 FILLER_206_865 ();
 b15zdnd11an1n32x5 FILLER_206_929 ();
 b15zdnd11an1n04x5 FILLER_206_961 ();
 b15zdnd00an1n02x5 FILLER_206_965 ();
 b15zdnd00an1n01x5 FILLER_206_967 ();
 b15zdnd11an1n64x5 FILLER_206_982 ();
 b15zdnd11an1n64x5 FILLER_206_1046 ();
 b15zdnd11an1n16x5 FILLER_206_1110 ();
 b15zdnd11an1n08x5 FILLER_206_1126 ();
 b15zdnd11an1n04x5 FILLER_206_1134 ();
 b15zdnd00an1n01x5 FILLER_206_1138 ();
 b15zdnd11an1n04x5 FILLER_206_1144 ();
 b15zdnd11an1n16x5 FILLER_206_1152 ();
 b15zdnd11an1n08x5 FILLER_206_1168 ();
 b15zdnd00an1n01x5 FILLER_206_1176 ();
 b15zdnd11an1n64x5 FILLER_206_1194 ();
 b15zdnd11an1n08x5 FILLER_206_1258 ();
 b15zdnd11an1n32x5 FILLER_206_1269 ();
 b15zdnd11an1n08x5 FILLER_206_1301 ();
 b15zdnd11an1n04x5 FILLER_206_1309 ();
 b15zdnd00an1n02x5 FILLER_206_1313 ();
 b15zdnd11an1n04x5 FILLER_206_1319 ();
 b15zdnd11an1n64x5 FILLER_206_1337 ();
 b15zdnd11an1n64x5 FILLER_206_1401 ();
 b15zdnd11an1n64x5 FILLER_206_1465 ();
 b15zdnd11an1n64x5 FILLER_206_1529 ();
 b15zdnd11an1n64x5 FILLER_206_1593 ();
 b15zdnd11an1n64x5 FILLER_206_1657 ();
 b15zdnd11an1n64x5 FILLER_206_1721 ();
 b15zdnd11an1n64x5 FILLER_206_1785 ();
 b15zdnd11an1n64x5 FILLER_206_1849 ();
 b15zdnd11an1n16x5 FILLER_206_1913 ();
 b15zdnd11an1n04x5 FILLER_206_1929 ();
 b15zdnd11an1n04x5 FILLER_206_1936 ();
 b15zdnd11an1n64x5 FILLER_206_1943 ();
 b15zdnd11an1n64x5 FILLER_206_2007 ();
 b15zdnd11an1n64x5 FILLER_206_2071 ();
 b15zdnd11an1n16x5 FILLER_206_2135 ();
 b15zdnd00an1n02x5 FILLER_206_2151 ();
 b15zdnd00an1n01x5 FILLER_206_2153 ();
 b15zdnd11an1n64x5 FILLER_206_2162 ();
 b15zdnd11an1n32x5 FILLER_206_2226 ();
 b15zdnd00an1n02x5 FILLER_206_2258 ();
 b15zdnd00an1n01x5 FILLER_206_2260 ();
 b15zdnd11an1n08x5 FILLER_206_2265 ();
 b15zdnd00an1n02x5 FILLER_206_2273 ();
 b15zdnd00an1n01x5 FILLER_206_2275 ();
 b15zdnd00an1n02x5 FILLER_207_0 ();
 b15zdnd11an1n08x5 FILLER_207_16 ();
 b15zdnd11an1n04x5 FILLER_207_24 ();
 b15zdnd00an1n01x5 FILLER_207_28 ();
 b15zdnd11an1n64x5 FILLER_207_34 ();
 b15zdnd11an1n64x5 FILLER_207_98 ();
 b15zdnd11an1n64x5 FILLER_207_162 ();
 b15zdnd11an1n64x5 FILLER_207_226 ();
 b15zdnd11an1n64x5 FILLER_207_290 ();
 b15zdnd11an1n32x5 FILLER_207_354 ();
 b15zdnd11an1n04x5 FILLER_207_386 ();
 b15zdnd00an1n01x5 FILLER_207_390 ();
 b15zdnd11an1n08x5 FILLER_207_394 ();
 b15zdnd00an1n02x5 FILLER_207_402 ();
 b15zdnd00an1n01x5 FILLER_207_404 ();
 b15zdnd11an1n64x5 FILLER_207_417 ();
 b15zdnd11an1n64x5 FILLER_207_481 ();
 b15zdnd11an1n32x5 FILLER_207_545 ();
 b15zdnd11an1n08x5 FILLER_207_577 ();
 b15zdnd11an1n04x5 FILLER_207_585 ();
 b15zdnd00an1n01x5 FILLER_207_589 ();
 b15zdnd11an1n64x5 FILLER_207_598 ();
 b15zdnd11an1n32x5 FILLER_207_662 ();
 b15zdnd11an1n16x5 FILLER_207_694 ();
 b15zdnd11an1n04x5 FILLER_207_710 ();
 b15zdnd11an1n04x5 FILLER_207_725 ();
 b15zdnd11an1n64x5 FILLER_207_736 ();
 b15zdnd11an1n08x5 FILLER_207_800 ();
 b15zdnd11an1n04x5 FILLER_207_853 ();
 b15zdnd11an1n64x5 FILLER_207_860 ();
 b15zdnd11an1n64x5 FILLER_207_924 ();
 b15zdnd11an1n04x5 FILLER_207_988 ();
 b15zdnd00an1n02x5 FILLER_207_992 ();
 b15zdnd11an1n32x5 FILLER_207_1019 ();
 b15zdnd00an1n01x5 FILLER_207_1051 ();
 b15zdnd11an1n64x5 FILLER_207_1066 ();
 b15zdnd11an1n64x5 FILLER_207_1130 ();
 b15zdnd11an1n64x5 FILLER_207_1194 ();
 b15zdnd11an1n64x5 FILLER_207_1258 ();
 b15zdnd11an1n64x5 FILLER_207_1322 ();
 b15zdnd11an1n64x5 FILLER_207_1386 ();
 b15zdnd11an1n32x5 FILLER_207_1450 ();
 b15zdnd11an1n04x5 FILLER_207_1482 ();
 b15zdnd00an1n02x5 FILLER_207_1486 ();
 b15zdnd11an1n64x5 FILLER_207_1497 ();
 b15zdnd11an1n64x5 FILLER_207_1561 ();
 b15zdnd11an1n64x5 FILLER_207_1625 ();
 b15zdnd11an1n32x5 FILLER_207_1689 ();
 b15zdnd11an1n16x5 FILLER_207_1721 ();
 b15zdnd00an1n01x5 FILLER_207_1737 ();
 b15zdnd11an1n64x5 FILLER_207_1747 ();
 b15zdnd11an1n64x5 FILLER_207_1811 ();
 b15zdnd11an1n32x5 FILLER_207_1875 ();
 b15zdnd11an1n08x5 FILLER_207_1907 ();
 b15zdnd11an1n64x5 FILLER_207_1967 ();
 b15zdnd11an1n64x5 FILLER_207_2031 ();
 b15zdnd11an1n64x5 FILLER_207_2095 ();
 b15zdnd11an1n64x5 FILLER_207_2159 ();
 b15zdnd11an1n32x5 FILLER_207_2223 ();
 b15zdnd11an1n16x5 FILLER_207_2255 ();
 b15zdnd11an1n08x5 FILLER_207_2271 ();
 b15zdnd11an1n04x5 FILLER_207_2279 ();
 b15zdnd00an1n01x5 FILLER_207_2283 ();
 b15zdnd11an1n04x5 FILLER_208_8 ();
 b15zdnd00an1n01x5 FILLER_208_12 ();
 b15zdnd11an1n64x5 FILLER_208_18 ();
 b15zdnd11an1n64x5 FILLER_208_82 ();
 b15zdnd11an1n64x5 FILLER_208_146 ();
 b15zdnd11an1n64x5 FILLER_208_210 ();
 b15zdnd11an1n64x5 FILLER_208_274 ();
 b15zdnd11an1n16x5 FILLER_208_338 ();
 b15zdnd11an1n08x5 FILLER_208_354 ();
 b15zdnd00an1n02x5 FILLER_208_362 ();
 b15zdnd11an1n64x5 FILLER_208_416 ();
 b15zdnd11an1n64x5 FILLER_208_480 ();
 b15zdnd11an1n64x5 FILLER_208_544 ();
 b15zdnd11an1n32x5 FILLER_208_608 ();
 b15zdnd11an1n16x5 FILLER_208_640 ();
 b15zdnd11an1n08x5 FILLER_208_656 ();
 b15zdnd00an1n02x5 FILLER_208_664 ();
 b15zdnd00an1n01x5 FILLER_208_666 ();
 b15zdnd11an1n32x5 FILLER_208_681 ();
 b15zdnd11an1n04x5 FILLER_208_713 ();
 b15zdnd00an1n01x5 FILLER_208_717 ();
 b15zdnd11an1n64x5 FILLER_208_726 ();
 b15zdnd11an1n64x5 FILLER_208_790 ();
 b15zdnd11an1n04x5 FILLER_208_854 ();
 b15zdnd11an1n32x5 FILLER_208_885 ();
 b15zdnd11an1n16x5 FILLER_208_917 ();
 b15zdnd11an1n08x5 FILLER_208_933 ();
 b15zdnd11an1n04x5 FILLER_208_941 ();
 b15zdnd00an1n02x5 FILLER_208_945 ();
 b15zdnd11an1n32x5 FILLER_208_961 ();
 b15zdnd11an1n04x5 FILLER_208_993 ();
 b15zdnd11an1n64x5 FILLER_208_1022 ();
 b15zdnd11an1n08x5 FILLER_208_1086 ();
 b15zdnd00an1n02x5 FILLER_208_1094 ();
 b15zdnd00an1n01x5 FILLER_208_1096 ();
 b15zdnd11an1n32x5 FILLER_208_1111 ();
 b15zdnd11an1n16x5 FILLER_208_1143 ();
 b15zdnd11an1n08x5 FILLER_208_1159 ();
 b15zdnd11an1n04x5 FILLER_208_1167 ();
 b15zdnd00an1n02x5 FILLER_208_1171 ();
 b15zdnd00an1n01x5 FILLER_208_1173 ();
 b15zdnd11an1n64x5 FILLER_208_1195 ();
 b15zdnd11an1n32x5 FILLER_208_1259 ();
 b15zdnd11an1n16x5 FILLER_208_1291 ();
 b15zdnd11an1n08x5 FILLER_208_1307 ();
 b15zdnd11an1n04x5 FILLER_208_1315 ();
 b15zdnd00an1n02x5 FILLER_208_1319 ();
 b15zdnd00an1n01x5 FILLER_208_1321 ();
 b15zdnd11an1n64x5 FILLER_208_1336 ();
 b15zdnd11an1n64x5 FILLER_208_1400 ();
 b15zdnd11an1n64x5 FILLER_208_1464 ();
 b15zdnd11an1n64x5 FILLER_208_1528 ();
 b15zdnd11an1n64x5 FILLER_208_1592 ();
 b15zdnd11an1n64x5 FILLER_208_1656 ();
 b15zdnd11an1n64x5 FILLER_208_1720 ();
 b15zdnd11an1n64x5 FILLER_208_1784 ();
 b15zdnd11an1n08x5 FILLER_208_1848 ();
 b15zdnd11an1n04x5 FILLER_208_1856 ();
 b15zdnd11an1n64x5 FILLER_208_1876 ();
 b15zdnd00an1n01x5 FILLER_208_1940 ();
 b15zdnd11an1n64x5 FILLER_208_1944 ();
 b15zdnd11an1n64x5 FILLER_208_2008 ();
 b15zdnd11an1n64x5 FILLER_208_2072 ();
 b15zdnd11an1n16x5 FILLER_208_2136 ();
 b15zdnd00an1n02x5 FILLER_208_2152 ();
 b15zdnd11an1n64x5 FILLER_208_2162 ();
 b15zdnd11an1n32x5 FILLER_208_2226 ();
 b15zdnd11an1n16x5 FILLER_208_2258 ();
 b15zdnd00an1n02x5 FILLER_208_2274 ();
 b15zdnd11an1n16x5 FILLER_209_0 ();
 b15zdnd11an1n08x5 FILLER_209_16 ();
 b15zdnd00an1n02x5 FILLER_209_24 ();
 b15zdnd00an1n01x5 FILLER_209_26 ();
 b15zdnd11an1n04x5 FILLER_209_31 ();
 b15zdnd00an1n02x5 FILLER_209_35 ();
 b15zdnd11an1n64x5 FILLER_209_41 ();
 b15zdnd11an1n64x5 FILLER_209_105 ();
 b15zdnd11an1n32x5 FILLER_209_183 ();
 b15zdnd00an1n01x5 FILLER_209_215 ();
 b15zdnd11an1n64x5 FILLER_209_221 ();
 b15zdnd11an1n64x5 FILLER_209_285 ();
 b15zdnd11an1n32x5 FILLER_209_349 ();
 b15zdnd11an1n04x5 FILLER_209_381 ();
 b15zdnd00an1n02x5 FILLER_209_385 ();
 b15zdnd00an1n01x5 FILLER_209_387 ();
 b15zdnd11an1n04x5 FILLER_209_391 ();
 b15zdnd11an1n04x5 FILLER_209_398 ();
 b15zdnd11an1n04x5 FILLER_209_407 ();
 b15zdnd11an1n64x5 FILLER_209_453 ();
 b15zdnd00an1n01x5 FILLER_209_517 ();
 b15zdnd11an1n04x5 FILLER_209_523 ();
 b15zdnd11an1n64x5 FILLER_209_536 ();
 b15zdnd11an1n64x5 FILLER_209_600 ();
 b15zdnd11an1n64x5 FILLER_209_664 ();
 b15zdnd11an1n32x5 FILLER_209_728 ();
 b15zdnd11an1n04x5 FILLER_209_760 ();
 b15zdnd00an1n02x5 FILLER_209_764 ();
 b15zdnd00an1n01x5 FILLER_209_766 ();
 b15zdnd11an1n64x5 FILLER_209_779 ();
 b15zdnd11an1n08x5 FILLER_209_843 ();
 b15zdnd11an1n04x5 FILLER_209_851 ();
 b15zdnd00an1n01x5 FILLER_209_855 ();
 b15zdnd11an1n04x5 FILLER_209_881 ();
 b15zdnd00an1n02x5 FILLER_209_885 ();
 b15zdnd11an1n16x5 FILLER_209_912 ();
 b15zdnd11an1n04x5 FILLER_209_928 ();
 b15zdnd11an1n64x5 FILLER_209_942 ();
 b15zdnd11an1n64x5 FILLER_209_1006 ();
 b15zdnd11an1n64x5 FILLER_209_1070 ();
 b15zdnd11an1n04x5 FILLER_209_1134 ();
 b15zdnd00an1n01x5 FILLER_209_1138 ();
 b15zdnd11an1n08x5 FILLER_209_1176 ();
 b15zdnd11an1n04x5 FILLER_209_1184 ();
 b15zdnd00an1n01x5 FILLER_209_1188 ();
 b15zdnd11an1n04x5 FILLER_209_1203 ();
 b15zdnd11an1n64x5 FILLER_209_1218 ();
 b15zdnd00an1n02x5 FILLER_209_1282 ();
 b15zdnd11an1n64x5 FILLER_209_1296 ();
 b15zdnd11an1n64x5 FILLER_209_1360 ();
 b15zdnd11an1n64x5 FILLER_209_1424 ();
 b15zdnd11an1n64x5 FILLER_209_1488 ();
 b15zdnd11an1n64x5 FILLER_209_1552 ();
 b15zdnd11an1n64x5 FILLER_209_1616 ();
 b15zdnd11an1n64x5 FILLER_209_1680 ();
 b15zdnd11an1n64x5 FILLER_209_1744 ();
 b15zdnd11an1n32x5 FILLER_209_1808 ();
 b15zdnd11an1n16x5 FILLER_209_1840 ();
 b15zdnd00an1n02x5 FILLER_209_1856 ();
 b15zdnd11an1n64x5 FILLER_209_1865 ();
 b15zdnd11an1n64x5 FILLER_209_1929 ();
 b15zdnd11an1n64x5 FILLER_209_1993 ();
 b15zdnd11an1n64x5 FILLER_209_2057 ();
 b15zdnd11an1n32x5 FILLER_209_2121 ();
 b15zdnd11an1n08x5 FILLER_209_2153 ();
 b15zdnd11an1n04x5 FILLER_209_2161 ();
 b15zdnd00an1n02x5 FILLER_209_2165 ();
 b15zdnd00an1n01x5 FILLER_209_2167 ();
 b15zdnd11an1n64x5 FILLER_209_2175 ();
 b15zdnd11an1n32x5 FILLER_209_2239 ();
 b15zdnd11an1n08x5 FILLER_209_2271 ();
 b15zdnd11an1n04x5 FILLER_209_2279 ();
 b15zdnd00an1n01x5 FILLER_209_2283 ();
 b15zdnd11an1n64x5 FILLER_210_8 ();
 b15zdnd11an1n64x5 FILLER_210_72 ();
 b15zdnd11an1n64x5 FILLER_210_136 ();
 b15zdnd00an1n01x5 FILLER_210_200 ();
 b15zdnd11an1n04x5 FILLER_210_204 ();
 b15zdnd11an1n64x5 FILLER_210_222 ();
 b15zdnd11an1n64x5 FILLER_210_286 ();
 b15zdnd11an1n32x5 FILLER_210_350 ();
 b15zdnd11an1n04x5 FILLER_210_382 ();
 b15zdnd11an1n64x5 FILLER_210_393 ();
 b15zdnd11an1n64x5 FILLER_210_457 ();
 b15zdnd11an1n04x5 FILLER_210_524 ();
 b15zdnd11an1n64x5 FILLER_210_532 ();
 b15zdnd11an1n64x5 FILLER_210_596 ();
 b15zdnd11an1n32x5 FILLER_210_660 ();
 b15zdnd11an1n16x5 FILLER_210_692 ();
 b15zdnd11an1n08x5 FILLER_210_708 ();
 b15zdnd00an1n02x5 FILLER_210_716 ();
 b15zdnd11an1n32x5 FILLER_210_726 ();
 b15zdnd11an1n64x5 FILLER_210_782 ();
 b15zdnd11an1n64x5 FILLER_210_846 ();
 b15zdnd11an1n64x5 FILLER_210_910 ();
 b15zdnd11an1n64x5 FILLER_210_974 ();
 b15zdnd11an1n64x5 FILLER_210_1038 ();
 b15zdnd11an1n64x5 FILLER_210_1102 ();
 b15zdnd11an1n64x5 FILLER_210_1166 ();
 b15zdnd11an1n04x5 FILLER_210_1230 ();
 b15zdnd11an1n04x5 FILLER_210_1248 ();
 b15zdnd00an1n02x5 FILLER_210_1252 ();
 b15zdnd00an1n01x5 FILLER_210_1254 ();
 b15zdnd11an1n64x5 FILLER_210_1287 ();
 b15zdnd11an1n64x5 FILLER_210_1351 ();
 b15zdnd11an1n64x5 FILLER_210_1415 ();
 b15zdnd11an1n64x5 FILLER_210_1479 ();
 b15zdnd11an1n64x5 FILLER_210_1543 ();
 b15zdnd11an1n64x5 FILLER_210_1607 ();
 b15zdnd11an1n64x5 FILLER_210_1671 ();
 b15zdnd11an1n64x5 FILLER_210_1735 ();
 b15zdnd11an1n32x5 FILLER_210_1799 ();
 b15zdnd11an1n04x5 FILLER_210_1831 ();
 b15zdnd11an1n64x5 FILLER_210_1849 ();
 b15zdnd11an1n64x5 FILLER_210_1913 ();
 b15zdnd11an1n64x5 FILLER_210_1977 ();
 b15zdnd11an1n64x5 FILLER_210_2041 ();
 b15zdnd11an1n32x5 FILLER_210_2105 ();
 b15zdnd11an1n16x5 FILLER_210_2137 ();
 b15zdnd00an1n01x5 FILLER_210_2153 ();
 b15zdnd11an1n64x5 FILLER_210_2162 ();
 b15zdnd11an1n32x5 FILLER_210_2226 ();
 b15zdnd11an1n16x5 FILLER_210_2258 ();
 b15zdnd00an1n02x5 FILLER_210_2274 ();
 b15zdnd11an1n64x5 FILLER_211_0 ();
 b15zdnd11an1n64x5 FILLER_211_64 ();
 b15zdnd11an1n64x5 FILLER_211_128 ();
 b15zdnd00an1n02x5 FILLER_211_192 ();
 b15zdnd11an1n08x5 FILLER_211_209 ();
 b15zdnd00an1n01x5 FILLER_211_217 ();
 b15zdnd11an1n16x5 FILLER_211_224 ();
 b15zdnd11an1n04x5 FILLER_211_240 ();
 b15zdnd11an1n64x5 FILLER_211_247 ();
 b15zdnd11an1n64x5 FILLER_211_311 ();
 b15zdnd11an1n08x5 FILLER_211_375 ();
 b15zdnd00an1n02x5 FILLER_211_383 ();
 b15zdnd00an1n01x5 FILLER_211_385 ();
 b15zdnd11an1n04x5 FILLER_211_389 ();
 b15zdnd11an1n64x5 FILLER_211_398 ();
 b15zdnd11an1n32x5 FILLER_211_462 ();
 b15zdnd11an1n16x5 FILLER_211_494 ();
 b15zdnd11an1n04x5 FILLER_211_510 ();
 b15zdnd00an1n01x5 FILLER_211_514 ();
 b15zdnd11an1n04x5 FILLER_211_518 ();
 b15zdnd11an1n08x5 FILLER_211_529 ();
 b15zdnd00an1n02x5 FILLER_211_537 ();
 b15zdnd00an1n01x5 FILLER_211_539 ();
 b15zdnd11an1n64x5 FILLER_211_555 ();
 b15zdnd11an1n64x5 FILLER_211_619 ();
 b15zdnd11an1n32x5 FILLER_211_683 ();
 b15zdnd11an1n08x5 FILLER_211_715 ();
 b15zdnd11an1n04x5 FILLER_211_723 ();
 b15zdnd00an1n02x5 FILLER_211_727 ();
 b15zdnd00an1n01x5 FILLER_211_729 ();
 b15zdnd11an1n08x5 FILLER_211_750 ();
 b15zdnd11an1n04x5 FILLER_211_758 ();
 b15zdnd00an1n02x5 FILLER_211_762 ();
 b15zdnd00an1n01x5 FILLER_211_764 ();
 b15zdnd11an1n64x5 FILLER_211_779 ();
 b15zdnd11an1n64x5 FILLER_211_843 ();
 b15zdnd11an1n64x5 FILLER_211_907 ();
 b15zdnd11an1n64x5 FILLER_211_971 ();
 b15zdnd11an1n64x5 FILLER_211_1035 ();
 b15zdnd11an1n64x5 FILLER_211_1099 ();
 b15zdnd11an1n64x5 FILLER_211_1163 ();
 b15zdnd11an1n64x5 FILLER_211_1227 ();
 b15zdnd11an1n64x5 FILLER_211_1291 ();
 b15zdnd11an1n64x5 FILLER_211_1355 ();
 b15zdnd11an1n08x5 FILLER_211_1419 ();
 b15zdnd11an1n04x5 FILLER_211_1427 ();
 b15zdnd00an1n01x5 FILLER_211_1431 ();
 b15zdnd11an1n16x5 FILLER_211_1441 ();
 b15zdnd11an1n08x5 FILLER_211_1457 ();
 b15zdnd11an1n04x5 FILLER_211_1465 ();
 b15zdnd00an1n02x5 FILLER_211_1469 ();
 b15zdnd00an1n01x5 FILLER_211_1471 ();
 b15zdnd11an1n64x5 FILLER_211_1481 ();
 b15zdnd11an1n64x5 FILLER_211_1545 ();
 b15zdnd11an1n16x5 FILLER_211_1609 ();
 b15zdnd11an1n04x5 FILLER_211_1625 ();
 b15zdnd00an1n02x5 FILLER_211_1629 ();
 b15zdnd00an1n01x5 FILLER_211_1631 ();
 b15zdnd11an1n64x5 FILLER_211_1684 ();
 b15zdnd11an1n16x5 FILLER_211_1748 ();
 b15zdnd11an1n04x5 FILLER_211_1764 ();
 b15zdnd00an1n02x5 FILLER_211_1768 ();
 b15zdnd00an1n01x5 FILLER_211_1770 ();
 b15zdnd11an1n64x5 FILLER_211_1774 ();
 b15zdnd11an1n04x5 FILLER_211_1838 ();
 b15zdnd11an1n64x5 FILLER_211_1849 ();
 b15zdnd11an1n16x5 FILLER_211_1913 ();
 b15zdnd11an1n08x5 FILLER_211_1929 ();
 b15zdnd11an1n16x5 FILLER_211_1979 ();
 b15zdnd11an1n08x5 FILLER_211_1995 ();
 b15zdnd11an1n04x5 FILLER_211_2003 ();
 b15zdnd00an1n01x5 FILLER_211_2007 ();
 b15zdnd11an1n64x5 FILLER_211_2023 ();
 b15zdnd11an1n64x5 FILLER_211_2087 ();
 b15zdnd11an1n64x5 FILLER_211_2151 ();
 b15zdnd11an1n64x5 FILLER_211_2215 ();
 b15zdnd11an1n04x5 FILLER_211_2279 ();
 b15zdnd00an1n01x5 FILLER_211_2283 ();
 b15zdnd11an1n64x5 FILLER_212_8 ();
 b15zdnd11an1n64x5 FILLER_212_72 ();
 b15zdnd11an1n32x5 FILLER_212_136 ();
 b15zdnd11an1n16x5 FILLER_212_168 ();
 b15zdnd00an1n02x5 FILLER_212_184 ();
 b15zdnd11an1n08x5 FILLER_212_204 ();
 b15zdnd11an1n04x5 FILLER_212_212 ();
 b15zdnd11an1n64x5 FILLER_212_248 ();
 b15zdnd11an1n64x5 FILLER_212_312 ();
 b15zdnd11an1n64x5 FILLER_212_376 ();
 b15zdnd11an1n64x5 FILLER_212_440 ();
 b15zdnd00an1n01x5 FILLER_212_504 ();
 b15zdnd11an1n04x5 FILLER_212_547 ();
 b15zdnd11an1n64x5 FILLER_212_557 ();
 b15zdnd11an1n64x5 FILLER_212_621 ();
 b15zdnd11an1n32x5 FILLER_212_685 ();
 b15zdnd00an1n01x5 FILLER_212_717 ();
 b15zdnd11an1n64x5 FILLER_212_726 ();
 b15zdnd11an1n64x5 FILLER_212_790 ();
 b15zdnd11an1n64x5 FILLER_212_854 ();
 b15zdnd11an1n64x5 FILLER_212_918 ();
 b15zdnd11an1n64x5 FILLER_212_982 ();
 b15zdnd11an1n64x5 FILLER_212_1046 ();
 b15zdnd11an1n64x5 FILLER_212_1110 ();
 b15zdnd11an1n64x5 FILLER_212_1174 ();
 b15zdnd11an1n64x5 FILLER_212_1238 ();
 b15zdnd11an1n64x5 FILLER_212_1302 ();
 b15zdnd11an1n64x5 FILLER_212_1366 ();
 b15zdnd11an1n64x5 FILLER_212_1430 ();
 b15zdnd11an1n64x5 FILLER_212_1494 ();
 b15zdnd11an1n64x5 FILLER_212_1558 ();
 b15zdnd11an1n32x5 FILLER_212_1622 ();
 b15zdnd00an1n01x5 FILLER_212_1654 ();
 b15zdnd11an1n04x5 FILLER_212_1658 ();
 b15zdnd11an1n64x5 FILLER_212_1665 ();
 b15zdnd11an1n32x5 FILLER_212_1729 ();
 b15zdnd11an1n08x5 FILLER_212_1761 ();
 b15zdnd00an1n02x5 FILLER_212_1769 ();
 b15zdnd11an1n64x5 FILLER_212_1774 ();
 b15zdnd11an1n64x5 FILLER_212_1838 ();
 b15zdnd11an1n04x5 FILLER_212_1902 ();
 b15zdnd00an1n02x5 FILLER_212_1906 ();
 b15zdnd11an1n64x5 FILLER_212_1917 ();
 b15zdnd11an1n32x5 FILLER_212_1981 ();
 b15zdnd00an1n02x5 FILLER_212_2013 ();
 b15zdnd00an1n01x5 FILLER_212_2015 ();
 b15zdnd11an1n64x5 FILLER_212_2022 ();
 b15zdnd11an1n64x5 FILLER_212_2086 ();
 b15zdnd11an1n04x5 FILLER_212_2150 ();
 b15zdnd11an1n64x5 FILLER_212_2162 ();
 b15zdnd11an1n32x5 FILLER_212_2226 ();
 b15zdnd11an1n16x5 FILLER_212_2258 ();
 b15zdnd00an1n02x5 FILLER_212_2274 ();
 b15zdnd11an1n64x5 FILLER_213_0 ();
 b15zdnd11an1n64x5 FILLER_213_64 ();
 b15zdnd11an1n64x5 FILLER_213_128 ();
 b15zdnd11an1n32x5 FILLER_213_192 ();
 b15zdnd11an1n16x5 FILLER_213_224 ();
 b15zdnd11an1n04x5 FILLER_213_240 ();
 b15zdnd11an1n64x5 FILLER_213_247 ();
 b15zdnd11an1n64x5 FILLER_213_311 ();
 b15zdnd11an1n64x5 FILLER_213_375 ();
 b15zdnd11an1n32x5 FILLER_213_439 ();
 b15zdnd11an1n16x5 FILLER_213_471 ();
 b15zdnd11an1n04x5 FILLER_213_487 ();
 b15zdnd00an1n02x5 FILLER_213_491 ();
 b15zdnd00an1n01x5 FILLER_213_493 ();
 b15zdnd11an1n64x5 FILLER_213_546 ();
 b15zdnd11an1n64x5 FILLER_213_610 ();
 b15zdnd11an1n64x5 FILLER_213_674 ();
 b15zdnd11an1n64x5 FILLER_213_738 ();
 b15zdnd11an1n64x5 FILLER_213_802 ();
 b15zdnd11an1n64x5 FILLER_213_866 ();
 b15zdnd11an1n64x5 FILLER_213_930 ();
 b15zdnd11an1n64x5 FILLER_213_994 ();
 b15zdnd11an1n64x5 FILLER_213_1058 ();
 b15zdnd11an1n64x5 FILLER_213_1122 ();
 b15zdnd11an1n64x5 FILLER_213_1186 ();
 b15zdnd11an1n64x5 FILLER_213_1250 ();
 b15zdnd11an1n64x5 FILLER_213_1314 ();
 b15zdnd11an1n64x5 FILLER_213_1378 ();
 b15zdnd11an1n64x5 FILLER_213_1442 ();
 b15zdnd11an1n64x5 FILLER_213_1506 ();
 b15zdnd11an1n64x5 FILLER_213_1570 ();
 b15zdnd11an1n16x5 FILLER_213_1634 ();
 b15zdnd11an1n04x5 FILLER_213_1650 ();
 b15zdnd00an1n02x5 FILLER_213_1654 ();
 b15zdnd00an1n01x5 FILLER_213_1656 ();
 b15zdnd11an1n64x5 FILLER_213_1660 ();
 b15zdnd11an1n16x5 FILLER_213_1724 ();
 b15zdnd11an1n04x5 FILLER_213_1740 ();
 b15zdnd00an1n02x5 FILLER_213_1744 ();
 b15zdnd11an1n16x5 FILLER_213_1798 ();
 b15zdnd11an1n04x5 FILLER_213_1814 ();
 b15zdnd00an1n02x5 FILLER_213_1818 ();
 b15zdnd00an1n01x5 FILLER_213_1820 ();
 b15zdnd11an1n32x5 FILLER_213_1863 ();
 b15zdnd00an1n02x5 FILLER_213_1895 ();
 b15zdnd11an1n08x5 FILLER_213_1903 ();
 b15zdnd11an1n64x5 FILLER_213_1919 ();
 b15zdnd11an1n32x5 FILLER_213_1983 ();
 b15zdnd11an1n04x5 FILLER_213_2015 ();
 b15zdnd00an1n02x5 FILLER_213_2019 ();
 b15zdnd11an1n64x5 FILLER_213_2063 ();
 b15zdnd11an1n32x5 FILLER_213_2127 ();
 b15zdnd11an1n04x5 FILLER_213_2159 ();
 b15zdnd11an1n08x5 FILLER_213_2174 ();
 b15zdnd11an1n64x5 FILLER_213_2190 ();
 b15zdnd11an1n16x5 FILLER_213_2254 ();
 b15zdnd11an1n08x5 FILLER_213_2270 ();
 b15zdnd11an1n04x5 FILLER_213_2278 ();
 b15zdnd00an1n02x5 FILLER_213_2282 ();
 b15zdnd11an1n64x5 FILLER_214_8 ();
 b15zdnd11an1n64x5 FILLER_214_72 ();
 b15zdnd11an1n32x5 FILLER_214_136 ();
 b15zdnd11an1n16x5 FILLER_214_168 ();
 b15zdnd11an1n08x5 FILLER_214_184 ();
 b15zdnd00an1n01x5 FILLER_214_192 ();
 b15zdnd11an1n64x5 FILLER_214_199 ();
 b15zdnd11an1n64x5 FILLER_214_263 ();
 b15zdnd11an1n64x5 FILLER_214_327 ();
 b15zdnd11an1n64x5 FILLER_214_391 ();
 b15zdnd11an1n32x5 FILLER_214_455 ();
 b15zdnd11an1n16x5 FILLER_214_487 ();
 b15zdnd11an1n08x5 FILLER_214_503 ();
 b15zdnd00an1n02x5 FILLER_214_511 ();
 b15zdnd00an1n01x5 FILLER_214_513 ();
 b15zdnd11an1n08x5 FILLER_214_517 ();
 b15zdnd00an1n02x5 FILLER_214_525 ();
 b15zdnd00an1n01x5 FILLER_214_527 ();
 b15zdnd11an1n64x5 FILLER_214_532 ();
 b15zdnd11an1n64x5 FILLER_214_596 ();
 b15zdnd11an1n32x5 FILLER_214_660 ();
 b15zdnd11an1n16x5 FILLER_214_692 ();
 b15zdnd11an1n08x5 FILLER_214_708 ();
 b15zdnd00an1n02x5 FILLER_214_716 ();
 b15zdnd11an1n64x5 FILLER_214_726 ();
 b15zdnd11an1n64x5 FILLER_214_790 ();
 b15zdnd11an1n64x5 FILLER_214_854 ();
 b15zdnd11an1n32x5 FILLER_214_918 ();
 b15zdnd11an1n08x5 FILLER_214_950 ();
 b15zdnd11an1n04x5 FILLER_214_958 ();
 b15zdnd00an1n01x5 FILLER_214_962 ();
 b15zdnd11an1n64x5 FILLER_214_988 ();
 b15zdnd11an1n08x5 FILLER_214_1052 ();
 b15zdnd11an1n04x5 FILLER_214_1060 ();
 b15zdnd00an1n02x5 FILLER_214_1064 ();
 b15zdnd00an1n01x5 FILLER_214_1066 ();
 b15zdnd11an1n32x5 FILLER_214_1091 ();
 b15zdnd11an1n04x5 FILLER_214_1123 ();
 b15zdnd11an1n64x5 FILLER_214_1136 ();
 b15zdnd11an1n64x5 FILLER_214_1200 ();
 b15zdnd11an1n64x5 FILLER_214_1264 ();
 b15zdnd11an1n64x5 FILLER_214_1328 ();
 b15zdnd11an1n64x5 FILLER_214_1392 ();
 b15zdnd11an1n16x5 FILLER_214_1456 ();
 b15zdnd11an1n64x5 FILLER_214_1483 ();
 b15zdnd11an1n64x5 FILLER_214_1547 ();
 b15zdnd11an1n16x5 FILLER_214_1611 ();
 b15zdnd00an1n02x5 FILLER_214_1627 ();
 b15zdnd00an1n01x5 FILLER_214_1629 ();
 b15zdnd11an1n64x5 FILLER_214_1657 ();
 b15zdnd11an1n32x5 FILLER_214_1721 ();
 b15zdnd11an1n08x5 FILLER_214_1753 ();
 b15zdnd11an1n04x5 FILLER_214_1761 ();
 b15zdnd11an1n04x5 FILLER_214_1768 ();
 b15zdnd11an1n64x5 FILLER_214_1775 ();
 b15zdnd11an1n16x5 FILLER_214_1839 ();
 b15zdnd11an1n04x5 FILLER_214_1855 ();
 b15zdnd00an1n02x5 FILLER_214_1859 ();
 b15zdnd11an1n04x5 FILLER_214_1866 ();
 b15zdnd11an1n16x5 FILLER_214_1876 ();
 b15zdnd11an1n04x5 FILLER_214_1892 ();
 b15zdnd00an1n02x5 FILLER_214_1896 ();
 b15zdnd11an1n04x5 FILLER_214_1904 ();
 b15zdnd11an1n32x5 FILLER_214_1914 ();
 b15zdnd11an1n16x5 FILLER_214_1946 ();
 b15zdnd11an1n08x5 FILLER_214_1962 ();
 b15zdnd00an1n01x5 FILLER_214_1970 ();
 b15zdnd11an1n04x5 FILLER_214_2015 ();
 b15zdnd11an1n64x5 FILLER_214_2059 ();
 b15zdnd11an1n16x5 FILLER_214_2123 ();
 b15zdnd11an1n08x5 FILLER_214_2139 ();
 b15zdnd11an1n04x5 FILLER_214_2147 ();
 b15zdnd00an1n02x5 FILLER_214_2151 ();
 b15zdnd00an1n01x5 FILLER_214_2153 ();
 b15zdnd11an1n64x5 FILLER_214_2162 ();
 b15zdnd11an1n32x5 FILLER_214_2226 ();
 b15zdnd11an1n16x5 FILLER_214_2258 ();
 b15zdnd00an1n02x5 FILLER_214_2274 ();
 b15zdnd11an1n64x5 FILLER_215_0 ();
 b15zdnd11an1n64x5 FILLER_215_64 ();
 b15zdnd11an1n64x5 FILLER_215_128 ();
 b15zdnd11an1n64x5 FILLER_215_192 ();
 b15zdnd11an1n04x5 FILLER_215_256 ();
 b15zdnd00an1n02x5 FILLER_215_260 ();
 b15zdnd00an1n01x5 FILLER_215_262 ();
 b15zdnd11an1n04x5 FILLER_215_305 ();
 b15zdnd00an1n02x5 FILLER_215_309 ();
 b15zdnd11an1n64x5 FILLER_215_314 ();
 b15zdnd11an1n64x5 FILLER_215_378 ();
 b15zdnd11an1n32x5 FILLER_215_442 ();
 b15zdnd11an1n16x5 FILLER_215_474 ();
 b15zdnd11an1n08x5 FILLER_215_490 ();
 b15zdnd11an1n04x5 FILLER_215_498 ();
 b15zdnd00an1n02x5 FILLER_215_502 ();
 b15zdnd00an1n01x5 FILLER_215_504 ();
 b15zdnd11an1n08x5 FILLER_215_516 ();
 b15zdnd00an1n01x5 FILLER_215_524 ();
 b15zdnd11an1n04x5 FILLER_215_529 ();
 b15zdnd11an1n04x5 FILLER_215_539 ();
 b15zdnd11an1n64x5 FILLER_215_585 ();
 b15zdnd11an1n32x5 FILLER_215_649 ();
 b15zdnd11an1n04x5 FILLER_215_681 ();
 b15zdnd11an1n08x5 FILLER_215_692 ();
 b15zdnd11an1n04x5 FILLER_215_700 ();
 b15zdnd11an1n64x5 FILLER_215_735 ();
 b15zdnd11an1n08x5 FILLER_215_799 ();
 b15zdnd11an1n04x5 FILLER_215_807 ();
 b15zdnd00an1n01x5 FILLER_215_811 ();
 b15zdnd11an1n64x5 FILLER_215_824 ();
 b15zdnd11an1n64x5 FILLER_215_888 ();
 b15zdnd11an1n32x5 FILLER_215_952 ();
 b15zdnd11an1n08x5 FILLER_215_984 ();
 b15zdnd11an1n04x5 FILLER_215_992 ();
 b15zdnd00an1n02x5 FILLER_215_996 ();
 b15zdnd11an1n32x5 FILLER_215_1029 ();
 b15zdnd11an1n08x5 FILLER_215_1061 ();
 b15zdnd11an1n04x5 FILLER_215_1069 ();
 b15zdnd11an1n08x5 FILLER_215_1104 ();
 b15zdnd11an1n04x5 FILLER_215_1112 ();
 b15zdnd00an1n01x5 FILLER_215_1116 ();
 b15zdnd11an1n32x5 FILLER_215_1136 ();
 b15zdnd11an1n04x5 FILLER_215_1168 ();
 b15zdnd00an1n01x5 FILLER_215_1172 ();
 b15zdnd11an1n64x5 FILLER_215_1184 ();
 b15zdnd11an1n16x5 FILLER_215_1248 ();
 b15zdnd11an1n04x5 FILLER_215_1264 ();
 b15zdnd00an1n02x5 FILLER_215_1268 ();
 b15zdnd11an1n08x5 FILLER_215_1281 ();
 b15zdnd11an1n04x5 FILLER_215_1298 ();
 b15zdnd11an1n64x5 FILLER_215_1316 ();
 b15zdnd11an1n64x5 FILLER_215_1380 ();
 b15zdnd11an1n64x5 FILLER_215_1444 ();
 b15zdnd11an1n64x5 FILLER_215_1508 ();
 b15zdnd11an1n32x5 FILLER_215_1572 ();
 b15zdnd11an1n16x5 FILLER_215_1604 ();
 b15zdnd11an1n04x5 FILLER_215_1620 ();
 b15zdnd00an1n02x5 FILLER_215_1624 ();
 b15zdnd00an1n01x5 FILLER_215_1626 ();
 b15zdnd11an1n64x5 FILLER_215_1630 ();
 b15zdnd11an1n32x5 FILLER_215_1694 ();
 b15zdnd11an1n16x5 FILLER_215_1726 ();
 b15zdnd11an1n04x5 FILLER_215_1742 ();
 b15zdnd11an1n64x5 FILLER_215_1798 ();
 b15zdnd11an1n32x5 FILLER_215_1862 ();
 b15zdnd00an1n02x5 FILLER_215_1894 ();
 b15zdnd00an1n01x5 FILLER_215_1896 ();
 b15zdnd11an1n04x5 FILLER_215_1903 ();
 b15zdnd11an1n04x5 FILLER_215_1949 ();
 b15zdnd11an1n04x5 FILLER_215_1995 ();
 b15zdnd11an1n04x5 FILLER_215_2002 ();
 b15zdnd11an1n32x5 FILLER_215_2009 ();
 b15zdnd11an1n08x5 FILLER_215_2041 ();
 b15zdnd11an1n04x5 FILLER_215_2049 ();
 b15zdnd11an1n04x5 FILLER_215_2056 ();
 b15zdnd11an1n64x5 FILLER_215_2063 ();
 b15zdnd11an1n64x5 FILLER_215_2127 ();
 b15zdnd11an1n64x5 FILLER_215_2191 ();
 b15zdnd11an1n16x5 FILLER_215_2255 ();
 b15zdnd11an1n08x5 FILLER_215_2271 ();
 b15zdnd11an1n04x5 FILLER_215_2279 ();
 b15zdnd00an1n01x5 FILLER_215_2283 ();
 b15zdnd11an1n64x5 FILLER_216_8 ();
 b15zdnd11an1n64x5 FILLER_216_72 ();
 b15zdnd11an1n64x5 FILLER_216_136 ();
 b15zdnd11an1n64x5 FILLER_216_200 ();
 b15zdnd11an1n16x5 FILLER_216_264 ();
 b15zdnd00an1n02x5 FILLER_216_280 ();
 b15zdnd00an1n01x5 FILLER_216_282 ();
 b15zdnd11an1n64x5 FILLER_216_315 ();
 b15zdnd11an1n64x5 FILLER_216_379 ();
 b15zdnd11an1n64x5 FILLER_216_443 ();
 b15zdnd11an1n16x5 FILLER_216_507 ();
 b15zdnd11an1n04x5 FILLER_216_523 ();
 b15zdnd00an1n02x5 FILLER_216_527 ();
 b15zdnd11an1n64x5 FILLER_216_540 ();
 b15zdnd11an1n64x5 FILLER_216_604 ();
 b15zdnd11an1n32x5 FILLER_216_668 ();
 b15zdnd11an1n16x5 FILLER_216_700 ();
 b15zdnd00an1n02x5 FILLER_216_716 ();
 b15zdnd00an1n02x5 FILLER_216_726 ();
 b15zdnd11an1n08x5 FILLER_216_748 ();
 b15zdnd11an1n64x5 FILLER_216_776 ();
 b15zdnd11an1n64x5 FILLER_216_848 ();
 b15zdnd11an1n32x5 FILLER_216_912 ();
 b15zdnd11an1n16x5 FILLER_216_944 ();
 b15zdnd11an1n08x5 FILLER_216_960 ();
 b15zdnd00an1n02x5 FILLER_216_968 ();
 b15zdnd00an1n01x5 FILLER_216_970 ();
 b15zdnd11an1n64x5 FILLER_216_988 ();
 b15zdnd11an1n64x5 FILLER_216_1052 ();
 b15zdnd11an1n64x5 FILLER_216_1116 ();
 b15zdnd11an1n64x5 FILLER_216_1180 ();
 b15zdnd11an1n16x5 FILLER_216_1244 ();
 b15zdnd11an1n08x5 FILLER_216_1260 ();
 b15zdnd00an1n02x5 FILLER_216_1268 ();
 b15zdnd11an1n64x5 FILLER_216_1282 ();
 b15zdnd11an1n32x5 FILLER_216_1346 ();
 b15zdnd11an1n16x5 FILLER_216_1378 ();
 b15zdnd11an1n04x5 FILLER_216_1394 ();
 b15zdnd00an1n01x5 FILLER_216_1398 ();
 b15zdnd11an1n04x5 FILLER_216_1402 ();
 b15zdnd11an1n64x5 FILLER_216_1409 ();
 b15zdnd11an1n64x5 FILLER_216_1482 ();
 b15zdnd11an1n64x5 FILLER_216_1546 ();
 b15zdnd11an1n64x5 FILLER_216_1610 ();
 b15zdnd11an1n08x5 FILLER_216_1674 ();
 b15zdnd11an1n32x5 FILLER_216_1691 ();
 b15zdnd11an1n08x5 FILLER_216_1723 ();
 b15zdnd11an1n04x5 FILLER_216_1731 ();
 b15zdnd00an1n02x5 FILLER_216_1735 ();
 b15zdnd00an1n01x5 FILLER_216_1737 ();
 b15zdnd11an1n16x5 FILLER_216_1747 ();
 b15zdnd00an1n01x5 FILLER_216_1763 ();
 b15zdnd11an1n04x5 FILLER_216_1767 ();
 b15zdnd11an1n16x5 FILLER_216_1774 ();
 b15zdnd11an1n08x5 FILLER_216_1790 ();
 b15zdnd11an1n04x5 FILLER_216_1798 ();
 b15zdnd11an1n64x5 FILLER_216_1809 ();
 b15zdnd11an1n64x5 FILLER_216_1873 ();
 b15zdnd11an1n32x5 FILLER_216_1937 ();
 b15zdnd11an1n16x5 FILLER_216_1969 ();
 b15zdnd11an1n08x5 FILLER_216_1985 ();
 b15zdnd11an1n04x5 FILLER_216_1993 ();
 b15zdnd00an1n02x5 FILLER_216_1997 ();
 b15zdnd11an1n64x5 FILLER_216_2002 ();
 b15zdnd11an1n64x5 FILLER_216_2066 ();
 b15zdnd11an1n16x5 FILLER_216_2130 ();
 b15zdnd11an1n08x5 FILLER_216_2146 ();
 b15zdnd11an1n64x5 FILLER_216_2162 ();
 b15zdnd11an1n32x5 FILLER_216_2226 ();
 b15zdnd11an1n16x5 FILLER_216_2258 ();
 b15zdnd00an1n02x5 FILLER_216_2274 ();
 b15zdnd11an1n64x5 FILLER_217_0 ();
 b15zdnd11an1n08x5 FILLER_217_64 ();
 b15zdnd11an1n04x5 FILLER_217_72 ();
 b15zdnd11an1n64x5 FILLER_217_96 ();
 b15zdnd11an1n16x5 FILLER_217_160 ();
 b15zdnd11an1n08x5 FILLER_217_176 ();
 b15zdnd11an1n04x5 FILLER_217_184 ();
 b15zdnd00an1n02x5 FILLER_217_188 ();
 b15zdnd00an1n01x5 FILLER_217_190 ();
 b15zdnd11an1n64x5 FILLER_217_201 ();
 b15zdnd11an1n32x5 FILLER_217_265 ();
 b15zdnd11an1n08x5 FILLER_217_297 ();
 b15zdnd11an1n04x5 FILLER_217_305 ();
 b15zdnd00an1n01x5 FILLER_217_309 ();
 b15zdnd11an1n64x5 FILLER_217_313 ();
 b15zdnd11an1n08x5 FILLER_217_377 ();
 b15zdnd00an1n01x5 FILLER_217_385 ();
 b15zdnd11an1n64x5 FILLER_217_391 ();
 b15zdnd11an1n64x5 FILLER_217_455 ();
 b15zdnd11an1n64x5 FILLER_217_519 ();
 b15zdnd11an1n32x5 FILLER_217_583 ();
 b15zdnd11an1n16x5 FILLER_217_615 ();
 b15zdnd11an1n04x5 FILLER_217_631 ();
 b15zdnd00an1n01x5 FILLER_217_635 ();
 b15zdnd11an1n08x5 FILLER_217_639 ();
 b15zdnd11an1n04x5 FILLER_217_647 ();
 b15zdnd00an1n02x5 FILLER_217_651 ();
 b15zdnd00an1n01x5 FILLER_217_653 ();
 b15zdnd11an1n64x5 FILLER_217_696 ();
 b15zdnd11an1n64x5 FILLER_217_760 ();
 b15zdnd11an1n64x5 FILLER_217_824 ();
 b15zdnd11an1n64x5 FILLER_217_888 ();
 b15zdnd11an1n64x5 FILLER_217_952 ();
 b15zdnd11an1n64x5 FILLER_217_1016 ();
 b15zdnd11an1n64x5 FILLER_217_1080 ();
 b15zdnd11an1n64x5 FILLER_217_1144 ();
 b15zdnd11an1n32x5 FILLER_217_1208 ();
 b15zdnd11an1n04x5 FILLER_217_1240 ();
 b15zdnd00an1n02x5 FILLER_217_1244 ();
 b15zdnd11an1n08x5 FILLER_217_1258 ();
 b15zdnd11an1n04x5 FILLER_217_1266 ();
 b15zdnd00an1n01x5 FILLER_217_1270 ();
 b15zdnd11an1n04x5 FILLER_217_1275 ();
 b15zdnd11an1n64x5 FILLER_217_1283 ();
 b15zdnd11an1n32x5 FILLER_217_1347 ();
 b15zdnd00an1n02x5 FILLER_217_1379 ();
 b15zdnd11an1n64x5 FILLER_217_1433 ();
 b15zdnd11an1n64x5 FILLER_217_1497 ();
 b15zdnd11an1n64x5 FILLER_217_1561 ();
 b15zdnd11an1n64x5 FILLER_217_1625 ();
 b15zdnd11an1n64x5 FILLER_217_1689 ();
 b15zdnd11an1n64x5 FILLER_217_1753 ();
 b15zdnd11an1n16x5 FILLER_217_1817 ();
 b15zdnd11an1n08x5 FILLER_217_1833 ();
 b15zdnd00an1n02x5 FILLER_217_1841 ();
 b15zdnd11an1n64x5 FILLER_217_1857 ();
 b15zdnd11an1n64x5 FILLER_217_1921 ();
 b15zdnd11an1n64x5 FILLER_217_1985 ();
 b15zdnd11an1n64x5 FILLER_217_2049 ();
 b15zdnd11an1n64x5 FILLER_217_2113 ();
 b15zdnd11an1n64x5 FILLER_217_2177 ();
 b15zdnd11an1n32x5 FILLER_217_2241 ();
 b15zdnd11an1n08x5 FILLER_217_2273 ();
 b15zdnd00an1n02x5 FILLER_217_2281 ();
 b15zdnd00an1n01x5 FILLER_217_2283 ();
 b15zdnd00an1n02x5 FILLER_218_8 ();
 b15zdnd11an1n04x5 FILLER_218_30 ();
 b15zdnd11an1n64x5 FILLER_218_38 ();
 b15zdnd11an1n64x5 FILLER_218_102 ();
 b15zdnd11an1n64x5 FILLER_218_166 ();
 b15zdnd11an1n64x5 FILLER_218_230 ();
 b15zdnd11an1n64x5 FILLER_218_294 ();
 b15zdnd11an1n16x5 FILLER_218_358 ();
 b15zdnd11an1n08x5 FILLER_218_374 ();
 b15zdnd11an1n04x5 FILLER_218_382 ();
 b15zdnd00an1n02x5 FILLER_218_386 ();
 b15zdnd00an1n01x5 FILLER_218_388 ();
 b15zdnd11an1n64x5 FILLER_218_405 ();
 b15zdnd11an1n64x5 FILLER_218_469 ();
 b15zdnd11an1n64x5 FILLER_218_533 ();
 b15zdnd11an1n08x5 FILLER_218_597 ();
 b15zdnd11an1n04x5 FILLER_218_605 ();
 b15zdnd11an1n32x5 FILLER_218_661 ();
 b15zdnd11an1n16x5 FILLER_218_693 ();
 b15zdnd11an1n08x5 FILLER_218_709 ();
 b15zdnd00an1n01x5 FILLER_218_717 ();
 b15zdnd11an1n64x5 FILLER_218_726 ();
 b15zdnd11an1n64x5 FILLER_218_790 ();
 b15zdnd11an1n64x5 FILLER_218_854 ();
 b15zdnd11an1n64x5 FILLER_218_918 ();
 b15zdnd11an1n64x5 FILLER_218_982 ();
 b15zdnd11an1n08x5 FILLER_218_1046 ();
 b15zdnd00an1n01x5 FILLER_218_1054 ();
 b15zdnd11an1n64x5 FILLER_218_1069 ();
 b15zdnd11an1n64x5 FILLER_218_1133 ();
 b15zdnd11an1n64x5 FILLER_218_1197 ();
 b15zdnd11an1n16x5 FILLER_218_1261 ();
 b15zdnd11an1n08x5 FILLER_218_1277 ();
 b15zdnd00an1n01x5 FILLER_218_1285 ();
 b15zdnd11an1n32x5 FILLER_218_1295 ();
 b15zdnd11an1n08x5 FILLER_218_1327 ();
 b15zdnd11an1n04x5 FILLER_218_1335 ();
 b15zdnd00an1n02x5 FILLER_218_1339 ();
 b15zdnd11an1n04x5 FILLER_218_1357 ();
 b15zdnd11an1n16x5 FILLER_218_1370 ();
 b15zdnd11an1n08x5 FILLER_218_1386 ();
 b15zdnd11an1n04x5 FILLER_218_1394 ();
 b15zdnd00an1n02x5 FILLER_218_1398 ();
 b15zdnd11an1n04x5 FILLER_218_1403 ();
 b15zdnd11an1n04x5 FILLER_218_1410 ();
 b15zdnd11an1n08x5 FILLER_218_1417 ();
 b15zdnd11an1n64x5 FILLER_218_1428 ();
 b15zdnd11an1n16x5 FILLER_218_1492 ();
 b15zdnd00an1n02x5 FILLER_218_1508 ();
 b15zdnd11an1n64x5 FILLER_218_1513 ();
 b15zdnd11an1n04x5 FILLER_218_1577 ();
 b15zdnd00an1n01x5 FILLER_218_1581 ();
 b15zdnd11an1n64x5 FILLER_218_1593 ();
 b15zdnd11an1n64x5 FILLER_218_1657 ();
 b15zdnd11an1n64x5 FILLER_218_1721 ();
 b15zdnd11an1n08x5 FILLER_218_1785 ();
 b15zdnd00an1n01x5 FILLER_218_1793 ();
 b15zdnd11an1n64x5 FILLER_218_1836 ();
 b15zdnd11an1n64x5 FILLER_218_1900 ();
 b15zdnd11an1n64x5 FILLER_218_1964 ();
 b15zdnd11an1n64x5 FILLER_218_2028 ();
 b15zdnd11an1n16x5 FILLER_218_2092 ();
 b15zdnd11an1n08x5 FILLER_218_2108 ();
 b15zdnd11an1n04x5 FILLER_218_2116 ();
 b15zdnd00an1n02x5 FILLER_218_2120 ();
 b15zdnd00an1n01x5 FILLER_218_2122 ();
 b15zdnd11an1n16x5 FILLER_218_2135 ();
 b15zdnd00an1n02x5 FILLER_218_2151 ();
 b15zdnd00an1n01x5 FILLER_218_2153 ();
 b15zdnd11an1n64x5 FILLER_218_2162 ();
 b15zdnd11an1n32x5 FILLER_218_2226 ();
 b15zdnd11an1n16x5 FILLER_218_2258 ();
 b15zdnd00an1n02x5 FILLER_218_2274 ();
 b15zdnd11an1n08x5 FILLER_219_0 ();
 b15zdnd11an1n04x5 FILLER_219_8 ();
 b15zdnd00an1n01x5 FILLER_219_12 ();
 b15zdnd11an1n64x5 FILLER_219_55 ();
 b15zdnd11an1n64x5 FILLER_219_119 ();
 b15zdnd00an1n02x5 FILLER_219_183 ();
 b15zdnd00an1n01x5 FILLER_219_185 ();
 b15zdnd11an1n64x5 FILLER_219_206 ();
 b15zdnd11an1n64x5 FILLER_219_270 ();
 b15zdnd11an1n08x5 FILLER_219_334 ();
 b15zdnd11an1n04x5 FILLER_219_342 ();
 b15zdnd00an1n02x5 FILLER_219_346 ();
 b15zdnd11an1n08x5 FILLER_219_390 ();
 b15zdnd00an1n01x5 FILLER_219_398 ();
 b15zdnd11an1n64x5 FILLER_219_415 ();
 b15zdnd11an1n16x5 FILLER_219_479 ();
 b15zdnd11an1n08x5 FILLER_219_495 ();
 b15zdnd00an1n01x5 FILLER_219_503 ();
 b15zdnd11an1n64x5 FILLER_219_546 ();
 b15zdnd11an1n16x5 FILLER_219_610 ();
 b15zdnd00an1n01x5 FILLER_219_626 ();
 b15zdnd11an1n04x5 FILLER_219_630 ();
 b15zdnd11an1n64x5 FILLER_219_637 ();
 b15zdnd11an1n64x5 FILLER_219_701 ();
 b15zdnd11an1n16x5 FILLER_219_765 ();
 b15zdnd11an1n08x5 FILLER_219_781 ();
 b15zdnd11an1n04x5 FILLER_219_789 ();
 b15zdnd00an1n02x5 FILLER_219_793 ();
 b15zdnd00an1n01x5 FILLER_219_795 ();
 b15zdnd11an1n64x5 FILLER_219_804 ();
 b15zdnd11an1n64x5 FILLER_219_868 ();
 b15zdnd11an1n16x5 FILLER_219_932 ();
 b15zdnd11an1n08x5 FILLER_219_948 ();
 b15zdnd11an1n04x5 FILLER_219_956 ();
 b15zdnd00an1n01x5 FILLER_219_960 ();
 b15zdnd11an1n08x5 FILLER_219_978 ();
 b15zdnd00an1n02x5 FILLER_219_986 ();
 b15zdnd11an1n16x5 FILLER_219_1002 ();
 b15zdnd11an1n04x5 FILLER_219_1018 ();
 b15zdnd00an1n02x5 FILLER_219_1022 ();
 b15zdnd00an1n01x5 FILLER_219_1024 ();
 b15zdnd11an1n64x5 FILLER_219_1030 ();
 b15zdnd11an1n64x5 FILLER_219_1094 ();
 b15zdnd11an1n64x5 FILLER_219_1158 ();
 b15zdnd11an1n64x5 FILLER_219_1222 ();
 b15zdnd11an1n64x5 FILLER_219_1286 ();
 b15zdnd11an1n32x5 FILLER_219_1350 ();
 b15zdnd11an1n32x5 FILLER_219_1434 ();
 b15zdnd11an1n16x5 FILLER_219_1466 ();
 b15zdnd00an1n02x5 FILLER_219_1482 ();
 b15zdnd11an1n64x5 FILLER_219_1536 ();
 b15zdnd11an1n64x5 FILLER_219_1600 ();
 b15zdnd11an1n32x5 FILLER_219_1664 ();
 b15zdnd11an1n16x5 FILLER_219_1696 ();
 b15zdnd00an1n02x5 FILLER_219_1712 ();
 b15zdnd00an1n01x5 FILLER_219_1714 ();
 b15zdnd11an1n64x5 FILLER_219_1724 ();
 b15zdnd11an1n64x5 FILLER_219_1788 ();
 b15zdnd11an1n04x5 FILLER_219_1852 ();
 b15zdnd11an1n64x5 FILLER_219_1870 ();
 b15zdnd11an1n64x5 FILLER_219_1934 ();
 b15zdnd11an1n64x5 FILLER_219_1998 ();
 b15zdnd11an1n64x5 FILLER_219_2062 ();
 b15zdnd11an1n32x5 FILLER_219_2126 ();
 b15zdnd11an1n16x5 FILLER_219_2158 ();
 b15zdnd11an1n08x5 FILLER_219_2174 ();
 b15zdnd00an1n02x5 FILLER_219_2182 ();
 b15zdnd00an1n01x5 FILLER_219_2184 ();
 b15zdnd11an1n04x5 FILLER_219_2188 ();
 b15zdnd11an1n64x5 FILLER_219_2195 ();
 b15zdnd11an1n16x5 FILLER_219_2259 ();
 b15zdnd11an1n08x5 FILLER_219_2275 ();
 b15zdnd00an1n01x5 FILLER_219_2283 ();
 b15zdnd11an1n16x5 FILLER_220_8 ();
 b15zdnd00an1n02x5 FILLER_220_24 ();
 b15zdnd11an1n04x5 FILLER_220_40 ();
 b15zdnd11an1n64x5 FILLER_220_55 ();
 b15zdnd11an1n64x5 FILLER_220_119 ();
 b15zdnd11an1n08x5 FILLER_220_183 ();
 b15zdnd11an1n04x5 FILLER_220_191 ();
 b15zdnd00an1n02x5 FILLER_220_195 ();
 b15zdnd11an1n64x5 FILLER_220_203 ();
 b15zdnd11an1n32x5 FILLER_220_267 ();
 b15zdnd11an1n16x5 FILLER_220_299 ();
 b15zdnd11an1n04x5 FILLER_220_315 ();
 b15zdnd00an1n02x5 FILLER_220_319 ();
 b15zdnd11an1n16x5 FILLER_220_363 ();
 b15zdnd11an1n04x5 FILLER_220_379 ();
 b15zdnd00an1n01x5 FILLER_220_383 ();
 b15zdnd11an1n64x5 FILLER_220_395 ();
 b15zdnd11an1n08x5 FILLER_220_459 ();
 b15zdnd11an1n64x5 FILLER_220_509 ();
 b15zdnd11an1n64x5 FILLER_220_573 ();
 b15zdnd11an1n64x5 FILLER_220_637 ();
 b15zdnd11an1n16x5 FILLER_220_701 ();
 b15zdnd00an1n01x5 FILLER_220_717 ();
 b15zdnd11an1n64x5 FILLER_220_726 ();
 b15zdnd11an1n64x5 FILLER_220_790 ();
 b15zdnd11an1n64x5 FILLER_220_854 ();
 b15zdnd11an1n64x5 FILLER_220_918 ();
 b15zdnd11an1n64x5 FILLER_220_982 ();
 b15zdnd11an1n64x5 FILLER_220_1046 ();
 b15zdnd11an1n64x5 FILLER_220_1110 ();
 b15zdnd11an1n64x5 FILLER_220_1174 ();
 b15zdnd11an1n32x5 FILLER_220_1238 ();
 b15zdnd11an1n64x5 FILLER_220_1274 ();
 b15zdnd11an1n32x5 FILLER_220_1338 ();
 b15zdnd11an1n16x5 FILLER_220_1370 ();
 b15zdnd11an1n08x5 FILLER_220_1386 ();
 b15zdnd11an1n04x5 FILLER_220_1394 ();
 b15zdnd11an1n08x5 FILLER_220_1450 ();
 b15zdnd11an1n04x5 FILLER_220_1458 ();
 b15zdnd00an1n01x5 FILLER_220_1462 ();
 b15zdnd11an1n08x5 FILLER_220_1474 ();
 b15zdnd00an1n01x5 FILLER_220_1482 ();
 b15zdnd11an1n64x5 FILLER_220_1535 ();
 b15zdnd11an1n64x5 FILLER_220_1599 ();
 b15zdnd11an1n64x5 FILLER_220_1663 ();
 b15zdnd11an1n64x5 FILLER_220_1727 ();
 b15zdnd11an1n64x5 FILLER_220_1791 ();
 b15zdnd11an1n64x5 FILLER_220_1855 ();
 b15zdnd11an1n64x5 FILLER_220_1919 ();
 b15zdnd11an1n64x5 FILLER_220_1983 ();
 b15zdnd11an1n32x5 FILLER_220_2047 ();
 b15zdnd11an1n04x5 FILLER_220_2079 ();
 b15zdnd00an1n02x5 FILLER_220_2083 ();
 b15zdnd11an1n32x5 FILLER_220_2093 ();
 b15zdnd11an1n16x5 FILLER_220_2125 ();
 b15zdnd11an1n08x5 FILLER_220_2141 ();
 b15zdnd11an1n04x5 FILLER_220_2149 ();
 b15zdnd00an1n01x5 FILLER_220_2153 ();
 b15zdnd11an1n04x5 FILLER_220_2162 ();
 b15zdnd00an1n01x5 FILLER_220_2166 ();
 b15zdnd11an1n32x5 FILLER_220_2219 ();
 b15zdnd11an1n16x5 FILLER_220_2251 ();
 b15zdnd11an1n08x5 FILLER_220_2267 ();
 b15zdnd00an1n01x5 FILLER_220_2275 ();
 b15zdnd11an1n08x5 FILLER_221_0 ();
 b15zdnd00an1n02x5 FILLER_221_8 ();
 b15zdnd11an1n64x5 FILLER_221_52 ();
 b15zdnd11an1n64x5 FILLER_221_116 ();
 b15zdnd11an1n64x5 FILLER_221_180 ();
 b15zdnd11an1n64x5 FILLER_221_244 ();
 b15zdnd11an1n64x5 FILLER_221_308 ();
 b15zdnd11an1n08x5 FILLER_221_372 ();
 b15zdnd11an1n04x5 FILLER_221_380 ();
 b15zdnd00an1n02x5 FILLER_221_384 ();
 b15zdnd11an1n64x5 FILLER_221_397 ();
 b15zdnd11an1n64x5 FILLER_221_461 ();
 b15zdnd11an1n32x5 FILLER_221_525 ();
 b15zdnd11an1n16x5 FILLER_221_557 ();
 b15zdnd00an1n02x5 FILLER_221_573 ();
 b15zdnd00an1n01x5 FILLER_221_575 ();
 b15zdnd11an1n64x5 FILLER_221_584 ();
 b15zdnd11an1n64x5 FILLER_221_648 ();
 b15zdnd11an1n64x5 FILLER_221_712 ();
 b15zdnd11an1n64x5 FILLER_221_776 ();
 b15zdnd11an1n64x5 FILLER_221_840 ();
 b15zdnd11an1n64x5 FILLER_221_904 ();
 b15zdnd11an1n64x5 FILLER_221_968 ();
 b15zdnd11an1n64x5 FILLER_221_1032 ();
 b15zdnd11an1n64x5 FILLER_221_1096 ();
 b15zdnd11an1n64x5 FILLER_221_1160 ();
 b15zdnd11an1n32x5 FILLER_221_1224 ();
 b15zdnd11an1n08x5 FILLER_221_1256 ();
 b15zdnd11an1n04x5 FILLER_221_1264 ();
 b15zdnd00an1n02x5 FILLER_221_1268 ();
 b15zdnd11an1n64x5 FILLER_221_1274 ();
 b15zdnd11an1n08x5 FILLER_221_1338 ();
 b15zdnd11an1n04x5 FILLER_221_1346 ();
 b15zdnd11an1n32x5 FILLER_221_1362 ();
 b15zdnd11an1n08x5 FILLER_221_1394 ();
 b15zdnd11an1n04x5 FILLER_221_1402 ();
 b15zdnd00an1n01x5 FILLER_221_1406 ();
 b15zdnd11an1n04x5 FILLER_221_1410 ();
 b15zdnd00an1n02x5 FILLER_221_1414 ();
 b15zdnd11an1n04x5 FILLER_221_1419 ();
 b15zdnd11an1n64x5 FILLER_221_1426 ();
 b15zdnd11an1n08x5 FILLER_221_1490 ();
 b15zdnd00an1n02x5 FILLER_221_1498 ();
 b15zdnd00an1n01x5 FILLER_221_1500 ();
 b15zdnd11an1n04x5 FILLER_221_1504 ();
 b15zdnd11an1n04x5 FILLER_221_1511 ();
 b15zdnd11an1n64x5 FILLER_221_1518 ();
 b15zdnd11an1n64x5 FILLER_221_1582 ();
 b15zdnd11an1n64x5 FILLER_221_1646 ();
 b15zdnd11an1n64x5 FILLER_221_1710 ();
 b15zdnd11an1n64x5 FILLER_221_1774 ();
 b15zdnd11an1n64x5 FILLER_221_1838 ();
 b15zdnd11an1n64x5 FILLER_221_1902 ();
 b15zdnd11an1n64x5 FILLER_221_1966 ();
 b15zdnd11an1n64x5 FILLER_221_2030 ();
 b15zdnd11an1n64x5 FILLER_221_2094 ();
 b15zdnd11an1n32x5 FILLER_221_2158 ();
 b15zdnd00an1n02x5 FILLER_221_2190 ();
 b15zdnd00an1n01x5 FILLER_221_2192 ();
 b15zdnd11an1n64x5 FILLER_221_2196 ();
 b15zdnd11an1n16x5 FILLER_221_2260 ();
 b15zdnd11an1n08x5 FILLER_221_2276 ();
 b15zdnd11an1n16x5 FILLER_222_8 ();
 b15zdnd00an1n02x5 FILLER_222_24 ();
 b15zdnd00an1n01x5 FILLER_222_26 ();
 b15zdnd11an1n04x5 FILLER_222_32 ();
 b15zdnd11an1n64x5 FILLER_222_40 ();
 b15zdnd11an1n64x5 FILLER_222_104 ();
 b15zdnd11an1n08x5 FILLER_222_168 ();
 b15zdnd11an1n04x5 FILLER_222_176 ();
 b15zdnd00an1n02x5 FILLER_222_180 ();
 b15zdnd11an1n64x5 FILLER_222_190 ();
 b15zdnd11an1n64x5 FILLER_222_254 ();
 b15zdnd11an1n64x5 FILLER_222_318 ();
 b15zdnd11an1n16x5 FILLER_222_382 ();
 b15zdnd00an1n02x5 FILLER_222_398 ();
 b15zdnd00an1n01x5 FILLER_222_400 ();
 b15zdnd11an1n64x5 FILLER_222_406 ();
 b15zdnd11an1n64x5 FILLER_222_470 ();
 b15zdnd11an1n64x5 FILLER_222_534 ();
 b15zdnd11an1n64x5 FILLER_222_598 ();
 b15zdnd11an1n32x5 FILLER_222_662 ();
 b15zdnd11an1n16x5 FILLER_222_694 ();
 b15zdnd11an1n08x5 FILLER_222_710 ();
 b15zdnd11an1n64x5 FILLER_222_726 ();
 b15zdnd11an1n16x5 FILLER_222_790 ();
 b15zdnd11an1n08x5 FILLER_222_806 ();
 b15zdnd11an1n04x5 FILLER_222_814 ();
 b15zdnd11an1n32x5 FILLER_222_838 ();
 b15zdnd11an1n16x5 FILLER_222_870 ();
 b15zdnd11an1n04x5 FILLER_222_886 ();
 b15zdnd00an1n01x5 FILLER_222_890 ();
 b15zdnd11an1n64x5 FILLER_222_911 ();
 b15zdnd11an1n32x5 FILLER_222_975 ();
 b15zdnd11an1n08x5 FILLER_222_1007 ();
 b15zdnd11an1n64x5 FILLER_222_1024 ();
 b15zdnd11an1n64x5 FILLER_222_1088 ();
 b15zdnd11an1n64x5 FILLER_222_1152 ();
 b15zdnd11an1n64x5 FILLER_222_1216 ();
 b15zdnd11an1n64x5 FILLER_222_1280 ();
 b15zdnd11an1n64x5 FILLER_222_1344 ();
 b15zdnd11an1n64x5 FILLER_222_1408 ();
 b15zdnd11an1n32x5 FILLER_222_1472 ();
 b15zdnd11an1n04x5 FILLER_222_1507 ();
 b15zdnd11an1n64x5 FILLER_222_1514 ();
 b15zdnd11an1n64x5 FILLER_222_1578 ();
 b15zdnd00an1n01x5 FILLER_222_1642 ();
 b15zdnd11an1n64x5 FILLER_222_1646 ();
 b15zdnd11an1n32x5 FILLER_222_1710 ();
 b15zdnd11an1n16x5 FILLER_222_1742 ();
 b15zdnd11an1n08x5 FILLER_222_1758 ();
 b15zdnd00an1n01x5 FILLER_222_1766 ();
 b15zdnd11an1n64x5 FILLER_222_1770 ();
 b15zdnd11an1n32x5 FILLER_222_1834 ();
 b15zdnd11an1n16x5 FILLER_222_1866 ();
 b15zdnd11an1n04x5 FILLER_222_1882 ();
 b15zdnd00an1n02x5 FILLER_222_1886 ();
 b15zdnd00an1n01x5 FILLER_222_1888 ();
 b15zdnd11an1n64x5 FILLER_222_1893 ();
 b15zdnd11an1n64x5 FILLER_222_1957 ();
 b15zdnd11an1n64x5 FILLER_222_2021 ();
 b15zdnd11an1n64x5 FILLER_222_2085 ();
 b15zdnd11an1n04x5 FILLER_222_2149 ();
 b15zdnd00an1n01x5 FILLER_222_2153 ();
 b15zdnd11an1n64x5 FILLER_222_2162 ();
 b15zdnd11an1n32x5 FILLER_222_2226 ();
 b15zdnd11an1n16x5 FILLER_222_2258 ();
 b15zdnd00an1n02x5 FILLER_222_2274 ();
 b15zdnd11an1n16x5 FILLER_223_0 ();
 b15zdnd11an1n08x5 FILLER_223_16 ();
 b15zdnd11an1n64x5 FILLER_223_28 ();
 b15zdnd11an1n64x5 FILLER_223_92 ();
 b15zdnd11an1n64x5 FILLER_223_156 ();
 b15zdnd11an1n64x5 FILLER_223_220 ();
 b15zdnd11an1n64x5 FILLER_223_284 ();
 b15zdnd11an1n04x5 FILLER_223_348 ();
 b15zdnd00an1n01x5 FILLER_223_352 ();
 b15zdnd11an1n04x5 FILLER_223_395 ();
 b15zdnd11an1n64x5 FILLER_223_403 ();
 b15zdnd11an1n64x5 FILLER_223_467 ();
 b15zdnd11an1n64x5 FILLER_223_531 ();
 b15zdnd11an1n64x5 FILLER_223_595 ();
 b15zdnd11an1n64x5 FILLER_223_659 ();
 b15zdnd11an1n64x5 FILLER_223_723 ();
 b15zdnd11an1n64x5 FILLER_223_787 ();
 b15zdnd11an1n64x5 FILLER_223_851 ();
 b15zdnd11an1n64x5 FILLER_223_915 ();
 b15zdnd11an1n64x5 FILLER_223_979 ();
 b15zdnd11an1n64x5 FILLER_223_1043 ();
 b15zdnd11an1n64x5 FILLER_223_1107 ();
 b15zdnd00an1n01x5 FILLER_223_1171 ();
 b15zdnd11an1n64x5 FILLER_223_1183 ();
 b15zdnd11an1n64x5 FILLER_223_1247 ();
 b15zdnd11an1n32x5 FILLER_223_1311 ();
 b15zdnd11an1n08x5 FILLER_223_1343 ();
 b15zdnd11an1n04x5 FILLER_223_1351 ();
 b15zdnd00an1n02x5 FILLER_223_1355 ();
 b15zdnd00an1n01x5 FILLER_223_1357 ();
 b15zdnd11an1n64x5 FILLER_223_1400 ();
 b15zdnd11an1n64x5 FILLER_223_1464 ();
 b15zdnd11an1n64x5 FILLER_223_1528 ();
 b15zdnd11an1n32x5 FILLER_223_1592 ();
 b15zdnd11an1n16x5 FILLER_223_1624 ();
 b15zdnd00an1n01x5 FILLER_223_1640 ();
 b15zdnd11an1n04x5 FILLER_223_1644 ();
 b15zdnd11an1n04x5 FILLER_223_1651 ();
 b15zdnd11an1n64x5 FILLER_223_1658 ();
 b15zdnd11an1n32x5 FILLER_223_1722 ();
 b15zdnd11an1n08x5 FILLER_223_1754 ();
 b15zdnd00an1n02x5 FILLER_223_1762 ();
 b15zdnd00an1n01x5 FILLER_223_1764 ();
 b15zdnd11an1n04x5 FILLER_223_1768 ();
 b15zdnd11an1n04x5 FILLER_223_1775 ();
 b15zdnd11an1n64x5 FILLER_223_1782 ();
 b15zdnd11an1n64x5 FILLER_223_1846 ();
 b15zdnd11an1n64x5 FILLER_223_1910 ();
 b15zdnd11an1n64x5 FILLER_223_1974 ();
 b15zdnd11an1n64x5 FILLER_223_2038 ();
 b15zdnd11an1n64x5 FILLER_223_2102 ();
 b15zdnd11an1n64x5 FILLER_223_2166 ();
 b15zdnd11an1n32x5 FILLER_223_2230 ();
 b15zdnd11an1n16x5 FILLER_223_2262 ();
 b15zdnd11an1n04x5 FILLER_223_2278 ();
 b15zdnd00an1n02x5 FILLER_223_2282 ();
 b15zdnd11an1n16x5 FILLER_224_8 ();
 b15zdnd11an1n64x5 FILLER_224_28 ();
 b15zdnd11an1n64x5 FILLER_224_92 ();
 b15zdnd11an1n16x5 FILLER_224_156 ();
 b15zdnd11an1n08x5 FILLER_224_172 ();
 b15zdnd11an1n64x5 FILLER_224_222 ();
 b15zdnd11an1n64x5 FILLER_224_286 ();
 b15zdnd11an1n16x5 FILLER_224_350 ();
 b15zdnd11an1n04x5 FILLER_224_366 ();
 b15zdnd00an1n02x5 FILLER_224_370 ();
 b15zdnd11an1n64x5 FILLER_224_414 ();
 b15zdnd11an1n64x5 FILLER_224_478 ();
 b15zdnd11an1n64x5 FILLER_224_542 ();
 b15zdnd11an1n32x5 FILLER_224_606 ();
 b15zdnd11an1n08x5 FILLER_224_638 ();
 b15zdnd11an1n04x5 FILLER_224_646 ();
 b15zdnd00an1n01x5 FILLER_224_650 ();
 b15zdnd11an1n32x5 FILLER_224_672 ();
 b15zdnd11an1n08x5 FILLER_224_704 ();
 b15zdnd11an1n04x5 FILLER_224_712 ();
 b15zdnd00an1n02x5 FILLER_224_716 ();
 b15zdnd11an1n64x5 FILLER_224_726 ();
 b15zdnd11an1n32x5 FILLER_224_790 ();
 b15zdnd11an1n04x5 FILLER_224_822 ();
 b15zdnd11an1n64x5 FILLER_224_840 ();
 b15zdnd11an1n64x5 FILLER_224_904 ();
 b15zdnd11an1n08x5 FILLER_224_968 ();
 b15zdnd11an1n04x5 FILLER_224_976 ();
 b15zdnd00an1n01x5 FILLER_224_980 ();
 b15zdnd11an1n04x5 FILLER_224_1017 ();
 b15zdnd11an1n64x5 FILLER_224_1032 ();
 b15zdnd11an1n64x5 FILLER_224_1096 ();
 b15zdnd11an1n04x5 FILLER_224_1160 ();
 b15zdnd11an1n64x5 FILLER_224_1168 ();
 b15zdnd11an1n64x5 FILLER_224_1232 ();
 b15zdnd11an1n64x5 FILLER_224_1296 ();
 b15zdnd00an1n02x5 FILLER_224_1360 ();
 b15zdnd11an1n64x5 FILLER_224_1371 ();
 b15zdnd11an1n64x5 FILLER_224_1435 ();
 b15zdnd11an1n64x5 FILLER_224_1499 ();
 b15zdnd11an1n32x5 FILLER_224_1563 ();
 b15zdnd11an1n16x5 FILLER_224_1595 ();
 b15zdnd11an1n08x5 FILLER_224_1611 ();
 b15zdnd11an1n04x5 FILLER_224_1619 ();
 b15zdnd11an1n64x5 FILLER_224_1675 ();
 b15zdnd11an1n08x5 FILLER_224_1739 ();
 b15zdnd11an1n64x5 FILLER_224_1799 ();
 b15zdnd11an1n64x5 FILLER_224_1863 ();
 b15zdnd11an1n64x5 FILLER_224_1927 ();
 b15zdnd11an1n64x5 FILLER_224_1991 ();
 b15zdnd11an1n64x5 FILLER_224_2055 ();
 b15zdnd11an1n32x5 FILLER_224_2119 ();
 b15zdnd00an1n02x5 FILLER_224_2151 ();
 b15zdnd00an1n01x5 FILLER_224_2153 ();
 b15zdnd11an1n64x5 FILLER_224_2162 ();
 b15zdnd11an1n32x5 FILLER_224_2226 ();
 b15zdnd11an1n16x5 FILLER_224_2258 ();
 b15zdnd00an1n02x5 FILLER_224_2274 ();
 b15zdnd11an1n64x5 FILLER_225_0 ();
 b15zdnd11an1n64x5 FILLER_225_64 ();
 b15zdnd11an1n64x5 FILLER_225_128 ();
 b15zdnd11an1n16x5 FILLER_225_192 ();
 b15zdnd11an1n64x5 FILLER_225_211 ();
 b15zdnd11an1n64x5 FILLER_225_275 ();
 b15zdnd11an1n64x5 FILLER_225_339 ();
 b15zdnd11an1n64x5 FILLER_225_403 ();
 b15zdnd11an1n64x5 FILLER_225_467 ();
 b15zdnd11an1n08x5 FILLER_225_531 ();
 b15zdnd11an1n04x5 FILLER_225_539 ();
 b15zdnd00an1n02x5 FILLER_225_543 ();
 b15zdnd00an1n01x5 FILLER_225_545 ();
 b15zdnd11an1n04x5 FILLER_225_551 ();
 b15zdnd00an1n02x5 FILLER_225_555 ();
 b15zdnd11an1n32x5 FILLER_225_599 ();
 b15zdnd11an1n16x5 FILLER_225_631 ();
 b15zdnd11an1n08x5 FILLER_225_647 ();
 b15zdnd11an1n04x5 FILLER_225_655 ();
 b15zdnd11an1n32x5 FILLER_225_673 ();
 b15zdnd11an1n16x5 FILLER_225_705 ();
 b15zdnd11an1n08x5 FILLER_225_728 ();
 b15zdnd00an1n01x5 FILLER_225_736 ();
 b15zdnd11an1n64x5 FILLER_225_743 ();
 b15zdnd11an1n64x5 FILLER_225_807 ();
 b15zdnd11an1n64x5 FILLER_225_871 ();
 b15zdnd11an1n64x5 FILLER_225_935 ();
 b15zdnd11an1n64x5 FILLER_225_999 ();
 b15zdnd11an1n08x5 FILLER_225_1063 ();
 b15zdnd00an1n02x5 FILLER_225_1071 ();
 b15zdnd11an1n64x5 FILLER_225_1084 ();
 b15zdnd11an1n64x5 FILLER_225_1148 ();
 b15zdnd11an1n64x5 FILLER_225_1212 ();
 b15zdnd11an1n64x5 FILLER_225_1276 ();
 b15zdnd11an1n64x5 FILLER_225_1340 ();
 b15zdnd11an1n64x5 FILLER_225_1404 ();
 b15zdnd11an1n64x5 FILLER_225_1468 ();
 b15zdnd11an1n64x5 FILLER_225_1532 ();
 b15zdnd11an1n16x5 FILLER_225_1596 ();
 b15zdnd11an1n04x5 FILLER_225_1612 ();
 b15zdnd00an1n02x5 FILLER_225_1616 ();
 b15zdnd00an1n01x5 FILLER_225_1618 ();
 b15zdnd11an1n64x5 FILLER_225_1671 ();
 b15zdnd00an1n02x5 FILLER_225_1735 ();
 b15zdnd00an1n01x5 FILLER_225_1737 ();
 b15zdnd11an1n64x5 FILLER_225_1790 ();
 b15zdnd11an1n64x5 FILLER_225_1854 ();
 b15zdnd11an1n64x5 FILLER_225_1918 ();
 b15zdnd11an1n64x5 FILLER_225_1982 ();
 b15zdnd11an1n64x5 FILLER_225_2046 ();
 b15zdnd11an1n64x5 FILLER_225_2110 ();
 b15zdnd11an1n64x5 FILLER_225_2174 ();
 b15zdnd11an1n32x5 FILLER_225_2238 ();
 b15zdnd11an1n08x5 FILLER_225_2270 ();
 b15zdnd11an1n04x5 FILLER_225_2278 ();
 b15zdnd00an1n02x5 FILLER_225_2282 ();
 b15zdnd11an1n32x5 FILLER_226_8 ();
 b15zdnd11an1n16x5 FILLER_226_40 ();
 b15zdnd11an1n08x5 FILLER_226_56 ();
 b15zdnd11an1n04x5 FILLER_226_64 ();
 b15zdnd11an1n64x5 FILLER_226_83 ();
 b15zdnd11an1n16x5 FILLER_226_147 ();
 b15zdnd11an1n08x5 FILLER_226_163 ();
 b15zdnd00an1n01x5 FILLER_226_171 ();
 b15zdnd11an1n04x5 FILLER_226_212 ();
 b15zdnd11an1n64x5 FILLER_226_219 ();
 b15zdnd11an1n64x5 FILLER_226_283 ();
 b15zdnd11an1n64x5 FILLER_226_347 ();
 b15zdnd11an1n64x5 FILLER_226_411 ();
 b15zdnd11an1n64x5 FILLER_226_475 ();
 b15zdnd11an1n04x5 FILLER_226_539 ();
 b15zdnd00an1n02x5 FILLER_226_543 ();
 b15zdnd11an1n16x5 FILLER_226_548 ();
 b15zdnd11an1n08x5 FILLER_226_564 ();
 b15zdnd11an1n16x5 FILLER_226_614 ();
 b15zdnd11an1n04x5 FILLER_226_630 ();
 b15zdnd00an1n02x5 FILLER_226_634 ();
 b15zdnd00an1n01x5 FILLER_226_636 ();
 b15zdnd11an1n16x5 FILLER_226_663 ();
 b15zdnd00an1n01x5 FILLER_226_679 ();
 b15zdnd11an1n16x5 FILLER_226_698 ();
 b15zdnd11an1n04x5 FILLER_226_714 ();
 b15zdnd11an1n32x5 FILLER_226_726 ();
 b15zdnd11an1n08x5 FILLER_226_758 ();
 b15zdnd11an1n64x5 FILLER_226_778 ();
 b15zdnd11an1n16x5 FILLER_226_842 ();
 b15zdnd11an1n08x5 FILLER_226_878 ();
 b15zdnd11an1n64x5 FILLER_226_893 ();
 b15zdnd11an1n64x5 FILLER_226_957 ();
 b15zdnd11an1n32x5 FILLER_226_1021 ();
 b15zdnd11an1n16x5 FILLER_226_1053 ();
 b15zdnd00an1n02x5 FILLER_226_1069 ();
 b15zdnd11an1n64x5 FILLER_226_1078 ();
 b15zdnd11an1n64x5 FILLER_226_1142 ();
 b15zdnd11an1n32x5 FILLER_226_1206 ();
 b15zdnd11an1n08x5 FILLER_226_1238 ();
 b15zdnd00an1n01x5 FILLER_226_1246 ();
 b15zdnd11an1n64x5 FILLER_226_1261 ();
 b15zdnd11an1n16x5 FILLER_226_1325 ();
 b15zdnd11an1n08x5 FILLER_226_1341 ();
 b15zdnd00an1n02x5 FILLER_226_1349 ();
 b15zdnd00an1n01x5 FILLER_226_1351 ();
 b15zdnd11an1n64x5 FILLER_226_1394 ();
 b15zdnd11an1n64x5 FILLER_226_1458 ();
 b15zdnd11an1n64x5 FILLER_226_1522 ();
 b15zdnd11an1n32x5 FILLER_226_1586 ();
 b15zdnd00an1n02x5 FILLER_226_1618 ();
 b15zdnd00an1n01x5 FILLER_226_1620 ();
 b15zdnd11an1n04x5 FILLER_226_1673 ();
 b15zdnd11an1n64x5 FILLER_226_1680 ();
 b15zdnd11an1n08x5 FILLER_226_1744 ();
 b15zdnd11an1n04x5 FILLER_226_1752 ();
 b15zdnd11an1n04x5 FILLER_226_1759 ();
 b15zdnd11an1n64x5 FILLER_226_1766 ();
 b15zdnd11an1n64x5 FILLER_226_1830 ();
 b15zdnd11an1n64x5 FILLER_226_1894 ();
 b15zdnd11an1n64x5 FILLER_226_1958 ();
 b15zdnd11an1n64x5 FILLER_226_2022 ();
 b15zdnd11an1n64x5 FILLER_226_2086 ();
 b15zdnd11an1n04x5 FILLER_226_2150 ();
 b15zdnd11an1n64x5 FILLER_226_2162 ();
 b15zdnd11an1n16x5 FILLER_226_2226 ();
 b15zdnd11an1n08x5 FILLER_226_2242 ();
 b15zdnd11an1n04x5 FILLER_226_2250 ();
 b15zdnd00an1n02x5 FILLER_226_2254 ();
 b15zdnd11an1n16x5 FILLER_226_2260 ();
 b15zdnd11an1n16x5 FILLER_227_0 ();
 b15zdnd11an1n04x5 FILLER_227_16 ();
 b15zdnd00an1n02x5 FILLER_227_20 ();
 b15zdnd11an1n64x5 FILLER_227_37 ();
 b15zdnd11an1n64x5 FILLER_227_101 ();
 b15zdnd11an1n32x5 FILLER_227_165 ();
 b15zdnd11an1n16x5 FILLER_227_197 ();
 b15zdnd11an1n04x5 FILLER_227_213 ();
 b15zdnd00an1n01x5 FILLER_227_217 ();
 b15zdnd11an1n64x5 FILLER_227_221 ();
 b15zdnd11an1n64x5 FILLER_227_285 ();
 b15zdnd11an1n64x5 FILLER_227_349 ();
 b15zdnd11an1n64x5 FILLER_227_413 ();
 b15zdnd11an1n64x5 FILLER_227_477 ();
 b15zdnd11an1n32x5 FILLER_227_541 ();
 b15zdnd11an1n16x5 FILLER_227_573 ();
 b15zdnd00an1n01x5 FILLER_227_589 ();
 b15zdnd11an1n64x5 FILLER_227_632 ();
 b15zdnd11an1n16x5 FILLER_227_696 ();
 b15zdnd00an1n02x5 FILLER_227_712 ();
 b15zdnd11an1n64x5 FILLER_227_766 ();
 b15zdnd11an1n16x5 FILLER_227_830 ();
 b15zdnd11an1n08x5 FILLER_227_846 ();
 b15zdnd11an1n16x5 FILLER_227_863 ();
 b15zdnd00an1n02x5 FILLER_227_879 ();
 b15zdnd00an1n01x5 FILLER_227_881 ();
 b15zdnd11an1n64x5 FILLER_227_902 ();
 b15zdnd11an1n08x5 FILLER_227_966 ();
 b15zdnd11an1n04x5 FILLER_227_974 ();
 b15zdnd00an1n02x5 FILLER_227_978 ();
 b15zdnd11an1n64x5 FILLER_227_990 ();
 b15zdnd11an1n08x5 FILLER_227_1054 ();
 b15zdnd11an1n04x5 FILLER_227_1062 ();
 b15zdnd00an1n02x5 FILLER_227_1066 ();
 b15zdnd00an1n01x5 FILLER_227_1068 ();
 b15zdnd11an1n64x5 FILLER_227_1082 ();
 b15zdnd11an1n64x5 FILLER_227_1146 ();
 b15zdnd11an1n64x5 FILLER_227_1210 ();
 b15zdnd11an1n64x5 FILLER_227_1274 ();
 b15zdnd11an1n64x5 FILLER_227_1338 ();
 b15zdnd11an1n64x5 FILLER_227_1402 ();
 b15zdnd11an1n64x5 FILLER_227_1466 ();
 b15zdnd11an1n64x5 FILLER_227_1530 ();
 b15zdnd11an1n32x5 FILLER_227_1594 ();
 b15zdnd11an1n08x5 FILLER_227_1626 ();
 b15zdnd00an1n02x5 FILLER_227_1634 ();
 b15zdnd00an1n01x5 FILLER_227_1636 ();
 b15zdnd11an1n04x5 FILLER_227_1640 ();
 b15zdnd11an1n04x5 FILLER_227_1647 ();
 b15zdnd11an1n64x5 FILLER_227_1654 ();
 b15zdnd11an1n64x5 FILLER_227_1718 ();
 b15zdnd11an1n64x5 FILLER_227_1782 ();
 b15zdnd11an1n64x5 FILLER_227_1846 ();
 b15zdnd11an1n64x5 FILLER_227_1910 ();
 b15zdnd11an1n64x5 FILLER_227_1974 ();
 b15zdnd11an1n64x5 FILLER_227_2038 ();
 b15zdnd11an1n64x5 FILLER_227_2102 ();
 b15zdnd11an1n32x5 FILLER_227_2166 ();
 b15zdnd11an1n16x5 FILLER_227_2215 ();
 b15zdnd11an1n08x5 FILLER_227_2231 ();
 b15zdnd11an1n04x5 FILLER_227_2239 ();
 b15zdnd00an1n01x5 FILLER_227_2243 ();
 b15zdnd11an1n16x5 FILLER_227_2248 ();
 b15zdnd11an1n04x5 FILLER_227_2264 ();
 b15zdnd00an1n01x5 FILLER_227_2268 ();
 b15zdnd11an1n08x5 FILLER_227_2273 ();
 b15zdnd00an1n02x5 FILLER_227_2281 ();
 b15zdnd00an1n01x5 FILLER_227_2283 ();
 b15zdnd11an1n64x5 FILLER_228_8 ();
 b15zdnd11an1n32x5 FILLER_228_72 ();
 b15zdnd00an1n02x5 FILLER_228_104 ();
 b15zdnd00an1n01x5 FILLER_228_106 ();
 b15zdnd11an1n32x5 FILLER_228_122 ();
 b15zdnd11an1n16x5 FILLER_228_154 ();
 b15zdnd11an1n08x5 FILLER_228_170 ();
 b15zdnd11an1n04x5 FILLER_228_178 ();
 b15zdnd00an1n02x5 FILLER_228_182 ();
 b15zdnd11an1n64x5 FILLER_228_224 ();
 b15zdnd11an1n64x5 FILLER_228_288 ();
 b15zdnd11an1n16x5 FILLER_228_352 ();
 b15zdnd11an1n32x5 FILLER_228_371 ();
 b15zdnd11an1n16x5 FILLER_228_403 ();
 b15zdnd11an1n08x5 FILLER_228_419 ();
 b15zdnd00an1n02x5 FILLER_228_427 ();
 b15zdnd00an1n01x5 FILLER_228_429 ();
 b15zdnd11an1n64x5 FILLER_228_433 ();
 b15zdnd11an1n32x5 FILLER_228_497 ();
 b15zdnd11an1n16x5 FILLER_228_529 ();
 b15zdnd11an1n64x5 FILLER_228_597 ();
 b15zdnd11an1n08x5 FILLER_228_661 ();
 b15zdnd11an1n04x5 FILLER_228_669 ();
 b15zdnd00an1n01x5 FILLER_228_673 ();
 b15zdnd00an1n02x5 FILLER_228_716 ();
 b15zdnd11an1n08x5 FILLER_228_726 ();
 b15zdnd11an1n04x5 FILLER_228_737 ();
 b15zdnd11an1n64x5 FILLER_228_744 ();
 b15zdnd11an1n08x5 FILLER_228_808 ();
 b15zdnd11an1n04x5 FILLER_228_816 ();
 b15zdnd00an1n02x5 FILLER_228_820 ();
 b15zdnd11an1n32x5 FILLER_228_825 ();
 b15zdnd11an1n08x5 FILLER_228_857 ();
 b15zdnd11an1n04x5 FILLER_228_865 ();
 b15zdnd00an1n01x5 FILLER_228_869 ();
 b15zdnd11an1n64x5 FILLER_228_876 ();
 b15zdnd11an1n64x5 FILLER_228_940 ();
 b15zdnd11an1n64x5 FILLER_228_1004 ();
 b15zdnd11an1n32x5 FILLER_228_1068 ();
 b15zdnd11an1n08x5 FILLER_228_1100 ();
 b15zdnd00an1n02x5 FILLER_228_1108 ();
 b15zdnd00an1n01x5 FILLER_228_1110 ();
 b15zdnd11an1n32x5 FILLER_228_1122 ();
 b15zdnd00an1n02x5 FILLER_228_1154 ();
 b15zdnd11an1n64x5 FILLER_228_1160 ();
 b15zdnd11an1n64x5 FILLER_228_1224 ();
 b15zdnd11an1n64x5 FILLER_228_1288 ();
 b15zdnd11an1n32x5 FILLER_228_1352 ();
 b15zdnd11an1n16x5 FILLER_228_1384 ();
 b15zdnd11an1n08x5 FILLER_228_1400 ();
 b15zdnd11an1n64x5 FILLER_228_1450 ();
 b15zdnd11an1n08x5 FILLER_228_1514 ();
 b15zdnd11an1n04x5 FILLER_228_1522 ();
 b15zdnd00an1n02x5 FILLER_228_1526 ();
 b15zdnd00an1n01x5 FILLER_228_1528 ();
 b15zdnd11an1n64x5 FILLER_228_1571 ();
 b15zdnd11an1n08x5 FILLER_228_1635 ();
 b15zdnd00an1n02x5 FILLER_228_1643 ();
 b15zdnd11an1n64x5 FILLER_228_1648 ();
 b15zdnd11an1n64x5 FILLER_228_1712 ();
 b15zdnd11an1n64x5 FILLER_228_1776 ();
 b15zdnd11an1n64x5 FILLER_228_1840 ();
 b15zdnd11an1n64x5 FILLER_228_1904 ();
 b15zdnd11an1n64x5 FILLER_228_1968 ();
 b15zdnd11an1n64x5 FILLER_228_2032 ();
 b15zdnd11an1n32x5 FILLER_228_2096 ();
 b15zdnd11an1n16x5 FILLER_228_2128 ();
 b15zdnd11an1n08x5 FILLER_228_2144 ();
 b15zdnd00an1n02x5 FILLER_228_2152 ();
 b15zdnd11an1n32x5 FILLER_228_2162 ();
 b15zdnd11an1n04x5 FILLER_228_2194 ();
 b15zdnd00an1n02x5 FILLER_228_2198 ();
 b15zdnd00an1n01x5 FILLER_228_2200 ();
 b15zdnd11an1n04x5 FILLER_228_2225 ();
 b15zdnd00an1n02x5 FILLER_228_2229 ();
 b15zdnd00an1n01x5 FILLER_228_2231 ();
 b15zdnd00an1n02x5 FILLER_228_2274 ();
 b15zdnd11an1n64x5 FILLER_229_0 ();
 b15zdnd11an1n16x5 FILLER_229_64 ();
 b15zdnd00an1n02x5 FILLER_229_80 ();
 b15zdnd00an1n01x5 FILLER_229_82 ();
 b15zdnd11an1n64x5 FILLER_229_101 ();
 b15zdnd11an1n32x5 FILLER_229_165 ();
 b15zdnd11an1n16x5 FILLER_229_197 ();
 b15zdnd11an1n04x5 FILLER_229_213 ();
 b15zdnd00an1n02x5 FILLER_229_217 ();
 b15zdnd00an1n01x5 FILLER_229_219 ();
 b15zdnd11an1n64x5 FILLER_229_223 ();
 b15zdnd11an1n32x5 FILLER_229_287 ();
 b15zdnd11an1n16x5 FILLER_229_319 ();
 b15zdnd11an1n08x5 FILLER_229_335 ();
 b15zdnd00an1n02x5 FILLER_229_343 ();
 b15zdnd00an1n01x5 FILLER_229_345 ();
 b15zdnd11an1n64x5 FILLER_229_398 ();
 b15zdnd11an1n64x5 FILLER_229_462 ();
 b15zdnd11an1n32x5 FILLER_229_526 ();
 b15zdnd00an1n02x5 FILLER_229_558 ();
 b15zdnd00an1n01x5 FILLER_229_560 ();
 b15zdnd11an1n04x5 FILLER_229_564 ();
 b15zdnd11an1n04x5 FILLER_229_571 ();
 b15zdnd11an1n04x5 FILLER_229_578 ();
 b15zdnd11an1n64x5 FILLER_229_613 ();
 b15zdnd11an1n32x5 FILLER_229_677 ();
 b15zdnd11an1n08x5 FILLER_229_709 ();
 b15zdnd00an1n02x5 FILLER_229_717 ();
 b15zdnd00an1n01x5 FILLER_229_719 ();
 b15zdnd11an1n04x5 FILLER_229_730 ();
 b15zdnd00an1n01x5 FILLER_229_734 ();
 b15zdnd11an1n32x5 FILLER_229_738 ();
 b15zdnd11an1n16x5 FILLER_229_770 ();
 b15zdnd11an1n08x5 FILLER_229_786 ();
 b15zdnd00an1n01x5 FILLER_229_794 ();
 b15zdnd11an1n64x5 FILLER_229_847 ();
 b15zdnd11an1n64x5 FILLER_229_911 ();
 b15zdnd11an1n16x5 FILLER_229_975 ();
 b15zdnd11an1n08x5 FILLER_229_991 ();
 b15zdnd11an1n04x5 FILLER_229_999 ();
 b15zdnd11an1n64x5 FILLER_229_1023 ();
 b15zdnd11an1n64x5 FILLER_229_1087 ();
 b15zdnd11an1n64x5 FILLER_229_1151 ();
 b15zdnd11an1n64x5 FILLER_229_1215 ();
 b15zdnd11an1n64x5 FILLER_229_1279 ();
 b15zdnd11an1n64x5 FILLER_229_1343 ();
 b15zdnd11an1n64x5 FILLER_229_1407 ();
 b15zdnd11an1n64x5 FILLER_229_1471 ();
 b15zdnd11an1n64x5 FILLER_229_1535 ();
 b15zdnd11an1n64x5 FILLER_229_1599 ();
 b15zdnd11an1n64x5 FILLER_229_1663 ();
 b15zdnd11an1n64x5 FILLER_229_1727 ();
 b15zdnd11an1n64x5 FILLER_229_1791 ();
 b15zdnd11an1n64x5 FILLER_229_1855 ();
 b15zdnd11an1n64x5 FILLER_229_1919 ();
 b15zdnd11an1n64x5 FILLER_229_1983 ();
 b15zdnd11an1n64x5 FILLER_229_2047 ();
 b15zdnd11an1n64x5 FILLER_229_2111 ();
 b15zdnd11an1n32x5 FILLER_229_2175 ();
 b15zdnd11an1n16x5 FILLER_229_2207 ();
 b15zdnd11an1n08x5 FILLER_229_2223 ();
 b15zdnd00an1n01x5 FILLER_229_2231 ();
 b15zdnd11an1n04x5 FILLER_229_2236 ();
 b15zdnd00an1n02x5 FILLER_229_2282 ();
 b15zdnd11an1n64x5 FILLER_230_8 ();
 b15zdnd11an1n64x5 FILLER_230_72 ();
 b15zdnd11an1n64x5 FILLER_230_136 ();
 b15zdnd11an1n64x5 FILLER_230_200 ();
 b15zdnd11an1n64x5 FILLER_230_264 ();
 b15zdnd11an1n32x5 FILLER_230_328 ();
 b15zdnd00an1n02x5 FILLER_230_360 ();
 b15zdnd00an1n01x5 FILLER_230_362 ();
 b15zdnd11an1n04x5 FILLER_230_366 ();
 b15zdnd11an1n16x5 FILLER_230_373 ();
 b15zdnd11an1n04x5 FILLER_230_389 ();
 b15zdnd00an1n02x5 FILLER_230_393 ();
 b15zdnd11an1n04x5 FILLER_230_427 ();
 b15zdnd11an1n64x5 FILLER_230_434 ();
 b15zdnd11an1n64x5 FILLER_230_498 ();
 b15zdnd11an1n64x5 FILLER_230_562 ();
 b15zdnd11an1n32x5 FILLER_230_626 ();
 b15zdnd11an1n04x5 FILLER_230_658 ();
 b15zdnd00an1n01x5 FILLER_230_662 ();
 b15zdnd11an1n08x5 FILLER_230_677 ();
 b15zdnd11an1n04x5 FILLER_230_685 ();
 b15zdnd00an1n01x5 FILLER_230_689 ();
 b15zdnd00an1n02x5 FILLER_230_716 ();
 b15zdnd00an1n02x5 FILLER_230_726 ();
 b15zdnd11an1n64x5 FILLER_230_741 ();
 b15zdnd11an1n08x5 FILLER_230_805 ();
 b15zdnd11an1n04x5 FILLER_230_816 ();
 b15zdnd11an1n16x5 FILLER_230_823 ();
 b15zdnd11an1n04x5 FILLER_230_839 ();
 b15zdnd11an1n04x5 FILLER_230_850 ();
 b15zdnd11an1n64x5 FILLER_230_861 ();
 b15zdnd11an1n16x5 FILLER_230_925 ();
 b15zdnd11an1n08x5 FILLER_230_941 ();
 b15zdnd11an1n04x5 FILLER_230_949 ();
 b15zdnd00an1n02x5 FILLER_230_953 ();
 b15zdnd00an1n01x5 FILLER_230_955 ();
 b15zdnd11an1n32x5 FILLER_230_970 ();
 b15zdnd11an1n04x5 FILLER_230_1002 ();
 b15zdnd11an1n32x5 FILLER_230_1014 ();
 b15zdnd11an1n08x5 FILLER_230_1046 ();
 b15zdnd11an1n04x5 FILLER_230_1054 ();
 b15zdnd11an1n16x5 FILLER_230_1061 ();
 b15zdnd00an1n01x5 FILLER_230_1077 ();
 b15zdnd11an1n64x5 FILLER_230_1097 ();
 b15zdnd11an1n16x5 FILLER_230_1161 ();
 b15zdnd11an1n08x5 FILLER_230_1177 ();
 b15zdnd00an1n02x5 FILLER_230_1185 ();
 b15zdnd00an1n01x5 FILLER_230_1187 ();
 b15zdnd11an1n64x5 FILLER_230_1191 ();
 b15zdnd11an1n16x5 FILLER_230_1255 ();
 b15zdnd00an1n01x5 FILLER_230_1271 ();
 b15zdnd11an1n64x5 FILLER_230_1275 ();
 b15zdnd11an1n64x5 FILLER_230_1339 ();
 b15zdnd11an1n64x5 FILLER_230_1403 ();
 b15zdnd11an1n16x5 FILLER_230_1467 ();
 b15zdnd11an1n08x5 FILLER_230_1483 ();
 b15zdnd11an1n04x5 FILLER_230_1491 ();
 b15zdnd00an1n01x5 FILLER_230_1495 ();
 b15zdnd11an1n64x5 FILLER_230_1505 ();
 b15zdnd11an1n64x5 FILLER_230_1569 ();
 b15zdnd11an1n64x5 FILLER_230_1633 ();
 b15zdnd11an1n64x5 FILLER_230_1697 ();
 b15zdnd11an1n32x5 FILLER_230_1761 ();
 b15zdnd11an1n08x5 FILLER_230_1793 ();
 b15zdnd00an1n02x5 FILLER_230_1801 ();
 b15zdnd00an1n01x5 FILLER_230_1803 ();
 b15zdnd11an1n64x5 FILLER_230_1846 ();
 b15zdnd11an1n64x5 FILLER_230_1910 ();
 b15zdnd11an1n64x5 FILLER_230_1974 ();
 b15zdnd11an1n64x5 FILLER_230_2038 ();
 b15zdnd11an1n32x5 FILLER_230_2102 ();
 b15zdnd11an1n16x5 FILLER_230_2134 ();
 b15zdnd11an1n04x5 FILLER_230_2150 ();
 b15zdnd11an1n64x5 FILLER_230_2162 ();
 b15zdnd11an1n04x5 FILLER_230_2226 ();
 b15zdnd00an1n02x5 FILLER_230_2230 ();
 b15zdnd00an1n02x5 FILLER_230_2274 ();
 b15zdnd11an1n64x5 FILLER_231_0 ();
 b15zdnd11an1n64x5 FILLER_231_64 ();
 b15zdnd11an1n64x5 FILLER_231_128 ();
 b15zdnd11an1n64x5 FILLER_231_192 ();
 b15zdnd11an1n64x5 FILLER_231_256 ();
 b15zdnd11an1n64x5 FILLER_231_320 ();
 b15zdnd11an1n64x5 FILLER_231_384 ();
 b15zdnd11an1n64x5 FILLER_231_448 ();
 b15zdnd11an1n64x5 FILLER_231_512 ();
 b15zdnd11an1n64x5 FILLER_231_576 ();
 b15zdnd11an1n16x5 FILLER_231_640 ();
 b15zdnd11an1n04x5 FILLER_231_682 ();
 b15zdnd11an1n08x5 FILLER_231_700 ();
 b15zdnd11an1n04x5 FILLER_231_708 ();
 b15zdnd11an1n64x5 FILLER_231_734 ();
 b15zdnd11an1n32x5 FILLER_231_798 ();
 b15zdnd11an1n16x5 FILLER_231_830 ();
 b15zdnd11an1n04x5 FILLER_231_846 ();
 b15zdnd11an1n32x5 FILLER_231_862 ();
 b15zdnd11an1n64x5 FILLER_231_912 ();
 b15zdnd11an1n32x5 FILLER_231_976 ();
 b15zdnd11an1n16x5 FILLER_231_1008 ();
 b15zdnd11an1n04x5 FILLER_231_1024 ();
 b15zdnd00an1n02x5 FILLER_231_1028 ();
 b15zdnd00an1n01x5 FILLER_231_1030 ();
 b15zdnd11an1n64x5 FILLER_231_1083 ();
 b15zdnd11an1n32x5 FILLER_231_1147 ();
 b15zdnd00an1n02x5 FILLER_231_1179 ();
 b15zdnd00an1n01x5 FILLER_231_1181 ();
 b15zdnd11an1n04x5 FILLER_231_1185 ();
 b15zdnd11an1n64x5 FILLER_231_1192 ();
 b15zdnd11an1n08x5 FILLER_231_1256 ();
 b15zdnd11an1n04x5 FILLER_231_1264 ();
 b15zdnd00an1n02x5 FILLER_231_1268 ();
 b15zdnd11an1n04x5 FILLER_231_1273 ();
 b15zdnd11an1n64x5 FILLER_231_1280 ();
 b15zdnd11an1n64x5 FILLER_231_1344 ();
 b15zdnd11an1n64x5 FILLER_231_1408 ();
 b15zdnd11an1n64x5 FILLER_231_1472 ();
 b15zdnd11an1n64x5 FILLER_231_1536 ();
 b15zdnd11an1n64x5 FILLER_231_1600 ();
 b15zdnd11an1n64x5 FILLER_231_1664 ();
 b15zdnd11an1n64x5 FILLER_231_1728 ();
 b15zdnd11an1n64x5 FILLER_231_1792 ();
 b15zdnd11an1n64x5 FILLER_231_1856 ();
 b15zdnd11an1n64x5 FILLER_231_1920 ();
 b15zdnd11an1n64x5 FILLER_231_1984 ();
 b15zdnd11an1n64x5 FILLER_231_2048 ();
 b15zdnd11an1n64x5 FILLER_231_2112 ();
 b15zdnd11an1n64x5 FILLER_231_2176 ();
 b15zdnd00an1n02x5 FILLER_231_2282 ();
 b15zdnd00an1n02x5 FILLER_232_8 ();
 b15zdnd11an1n64x5 FILLER_232_30 ();
 b15zdnd11an1n64x5 FILLER_232_94 ();
 b15zdnd11an1n64x5 FILLER_232_158 ();
 b15zdnd11an1n64x5 FILLER_232_222 ();
 b15zdnd11an1n64x5 FILLER_232_286 ();
 b15zdnd11an1n64x5 FILLER_232_350 ();
 b15zdnd11an1n32x5 FILLER_232_414 ();
 b15zdnd11an1n08x5 FILLER_232_446 ();
 b15zdnd11an1n16x5 FILLER_232_463 ();
 b15zdnd11an1n64x5 FILLER_232_482 ();
 b15zdnd11an1n32x5 FILLER_232_546 ();
 b15zdnd11an1n04x5 FILLER_232_578 ();
 b15zdnd00an1n02x5 FILLER_232_582 ();
 b15zdnd11an1n64x5 FILLER_232_626 ();
 b15zdnd11an1n16x5 FILLER_232_690 ();
 b15zdnd11an1n08x5 FILLER_232_706 ();
 b15zdnd11an1n04x5 FILLER_232_714 ();
 b15zdnd11an1n32x5 FILLER_232_726 ();
 b15zdnd11an1n08x5 FILLER_232_758 ();
 b15zdnd11an1n04x5 FILLER_232_766 ();
 b15zdnd00an1n01x5 FILLER_232_770 ();
 b15zdnd11an1n16x5 FILLER_232_783 ();
 b15zdnd11an1n04x5 FILLER_232_799 ();
 b15zdnd00an1n02x5 FILLER_232_803 ();
 b15zdnd11an1n64x5 FILLER_232_821 ();
 b15zdnd11an1n16x5 FILLER_232_885 ();
 b15zdnd00an1n02x5 FILLER_232_901 ();
 b15zdnd00an1n01x5 FILLER_232_903 ();
 b15zdnd11an1n64x5 FILLER_232_918 ();
 b15zdnd11an1n32x5 FILLER_232_982 ();
 b15zdnd11an1n04x5 FILLER_232_1014 ();
 b15zdnd00an1n01x5 FILLER_232_1018 ();
 b15zdnd11an1n16x5 FILLER_232_1033 ();
 b15zdnd11an1n04x5 FILLER_232_1052 ();
 b15zdnd11an1n64x5 FILLER_232_1059 ();
 b15zdnd11an1n32x5 FILLER_232_1123 ();
 b15zdnd11an1n08x5 FILLER_232_1155 ();
 b15zdnd00an1n01x5 FILLER_232_1163 ();
 b15zdnd11an1n32x5 FILLER_232_1216 ();
 b15zdnd11an1n04x5 FILLER_232_1248 ();
 b15zdnd11an1n64x5 FILLER_232_1304 ();
 b15zdnd11an1n64x5 FILLER_232_1368 ();
 b15zdnd11an1n64x5 FILLER_232_1432 ();
 b15zdnd11an1n16x5 FILLER_232_1496 ();
 b15zdnd00an1n02x5 FILLER_232_1512 ();
 b15zdnd00an1n01x5 FILLER_232_1514 ();
 b15zdnd11an1n64x5 FILLER_232_1524 ();
 b15zdnd11an1n64x5 FILLER_232_1588 ();
 b15zdnd11an1n64x5 FILLER_232_1652 ();
 b15zdnd11an1n64x5 FILLER_232_1716 ();
 b15zdnd11an1n64x5 FILLER_232_1780 ();
 b15zdnd11an1n64x5 FILLER_232_1844 ();
 b15zdnd11an1n64x5 FILLER_232_1908 ();
 b15zdnd11an1n64x5 FILLER_232_1972 ();
 b15zdnd11an1n64x5 FILLER_232_2036 ();
 b15zdnd11an1n32x5 FILLER_232_2100 ();
 b15zdnd11an1n16x5 FILLER_232_2132 ();
 b15zdnd11an1n04x5 FILLER_232_2148 ();
 b15zdnd00an1n02x5 FILLER_232_2152 ();
 b15zdnd11an1n32x5 FILLER_232_2162 ();
 b15zdnd11an1n08x5 FILLER_232_2194 ();
 b15zdnd11an1n04x5 FILLER_232_2202 ();
 b15zdnd11an1n16x5 FILLER_232_2248 ();
 b15zdnd11an1n08x5 FILLER_232_2264 ();
 b15zdnd11an1n04x5 FILLER_232_2272 ();
 b15zdnd11an1n64x5 FILLER_233_0 ();
 b15zdnd11an1n64x5 FILLER_233_64 ();
 b15zdnd11an1n64x5 FILLER_233_128 ();
 b15zdnd11an1n64x5 FILLER_233_192 ();
 b15zdnd11an1n64x5 FILLER_233_256 ();
 b15zdnd00an1n02x5 FILLER_233_320 ();
 b15zdnd11an1n64x5 FILLER_233_333 ();
 b15zdnd11an1n32x5 FILLER_233_397 ();
 b15zdnd11an1n16x5 FILLER_233_429 ();
 b15zdnd11an1n04x5 FILLER_233_445 ();
 b15zdnd00an1n02x5 FILLER_233_449 ();
 b15zdnd00an1n01x5 FILLER_233_451 ();
 b15zdnd11an1n64x5 FILLER_233_504 ();
 b15zdnd11an1n64x5 FILLER_233_568 ();
 b15zdnd11an1n64x5 FILLER_233_632 ();
 b15zdnd11an1n32x5 FILLER_233_696 ();
 b15zdnd11an1n08x5 FILLER_233_728 ();
 b15zdnd11an1n04x5 FILLER_233_736 ();
 b15zdnd00an1n02x5 FILLER_233_740 ();
 b15zdnd00an1n01x5 FILLER_233_742 ();
 b15zdnd11an1n08x5 FILLER_233_767 ();
 b15zdnd00an1n01x5 FILLER_233_775 ();
 b15zdnd11an1n64x5 FILLER_233_818 ();
 b15zdnd11an1n16x5 FILLER_233_882 ();
 b15zdnd00an1n02x5 FILLER_233_898 ();
 b15zdnd11an1n64x5 FILLER_233_926 ();
 b15zdnd11an1n64x5 FILLER_233_990 ();
 b15zdnd11an1n64x5 FILLER_233_1054 ();
 b15zdnd11an1n32x5 FILLER_233_1118 ();
 b15zdnd11an1n16x5 FILLER_233_1150 ();
 b15zdnd11an1n08x5 FILLER_233_1166 ();
 b15zdnd11an1n04x5 FILLER_233_1174 ();
 b15zdnd00an1n01x5 FILLER_233_1178 ();
 b15zdnd11an1n32x5 FILLER_233_1206 ();
 b15zdnd11an1n08x5 FILLER_233_1238 ();
 b15zdnd11an1n04x5 FILLER_233_1246 ();
 b15zdnd00an1n02x5 FILLER_233_1250 ();
 b15zdnd11an1n64x5 FILLER_233_1304 ();
 b15zdnd11an1n64x5 FILLER_233_1368 ();
 b15zdnd11an1n64x5 FILLER_233_1432 ();
 b15zdnd11an1n64x5 FILLER_233_1496 ();
 b15zdnd11an1n08x5 FILLER_233_1560 ();
 b15zdnd00an1n01x5 FILLER_233_1568 ();
 b15zdnd11an1n64x5 FILLER_233_1580 ();
 b15zdnd11an1n64x5 FILLER_233_1644 ();
 b15zdnd11an1n64x5 FILLER_233_1708 ();
 b15zdnd00an1n02x5 FILLER_233_1772 ();
 b15zdnd00an1n01x5 FILLER_233_1774 ();
 b15zdnd11an1n16x5 FILLER_233_1779 ();
 b15zdnd00an1n01x5 FILLER_233_1795 ();
 b15zdnd11an1n64x5 FILLER_233_1816 ();
 b15zdnd11an1n64x5 FILLER_233_1880 ();
 b15zdnd11an1n64x5 FILLER_233_1944 ();
 b15zdnd11an1n64x5 FILLER_233_2008 ();
 b15zdnd11an1n64x5 FILLER_233_2072 ();
 b15zdnd11an1n32x5 FILLER_233_2136 ();
 b15zdnd11an1n16x5 FILLER_233_2168 ();
 b15zdnd11an1n04x5 FILLER_233_2184 ();
 b15zdnd11an1n08x5 FILLER_233_2230 ();
 b15zdnd00an1n02x5 FILLER_233_2238 ();
 b15zdnd00an1n02x5 FILLER_233_2282 ();
 b15zdnd11an1n32x5 FILLER_234_8 ();
 b15zdnd11an1n08x5 FILLER_234_40 ();
 b15zdnd11an1n04x5 FILLER_234_48 ();
 b15zdnd00an1n02x5 FILLER_234_52 ();
 b15zdnd11an1n16x5 FILLER_234_72 ();
 b15zdnd11an1n08x5 FILLER_234_88 ();
 b15zdnd00an1n02x5 FILLER_234_96 ();
 b15zdnd11an1n64x5 FILLER_234_113 ();
 b15zdnd11an1n64x5 FILLER_234_177 ();
 b15zdnd11an1n64x5 FILLER_234_241 ();
 b15zdnd11an1n64x5 FILLER_234_305 ();
 b15zdnd11an1n64x5 FILLER_234_369 ();
 b15zdnd11an1n16x5 FILLER_234_433 ();
 b15zdnd11an1n04x5 FILLER_234_449 ();
 b15zdnd00an1n02x5 FILLER_234_453 ();
 b15zdnd11an1n04x5 FILLER_234_466 ();
 b15zdnd11an1n04x5 FILLER_234_473 ();
 b15zdnd11an1n64x5 FILLER_234_480 ();
 b15zdnd11an1n64x5 FILLER_234_544 ();
 b15zdnd11an1n64x5 FILLER_234_608 ();
 b15zdnd11an1n16x5 FILLER_234_672 ();
 b15zdnd11an1n08x5 FILLER_234_688 ();
 b15zdnd00an1n01x5 FILLER_234_696 ();
 b15zdnd11an1n04x5 FILLER_234_711 ();
 b15zdnd00an1n02x5 FILLER_234_715 ();
 b15zdnd00an1n01x5 FILLER_234_717 ();
 b15zdnd11an1n04x5 FILLER_234_726 ();
 b15zdnd00an1n01x5 FILLER_234_730 ();
 b15zdnd11an1n04x5 FILLER_234_751 ();
 b15zdnd11an1n04x5 FILLER_234_769 ();
 b15zdnd11an1n32x5 FILLER_234_784 ();
 b15zdnd11an1n16x5 FILLER_234_816 ();
 b15zdnd00an1n01x5 FILLER_234_832 ();
 b15zdnd11an1n32x5 FILLER_234_844 ();
 b15zdnd11an1n16x5 FILLER_234_876 ();
 b15zdnd11an1n08x5 FILLER_234_892 ();
 b15zdnd11an1n04x5 FILLER_234_900 ();
 b15zdnd11an1n64x5 FILLER_234_908 ();
 b15zdnd11an1n64x5 FILLER_234_972 ();
 b15zdnd11an1n32x5 FILLER_234_1036 ();
 b15zdnd11an1n08x5 FILLER_234_1068 ();
 b15zdnd11an1n04x5 FILLER_234_1076 ();
 b15zdnd00an1n01x5 FILLER_234_1080 ();
 b15zdnd11an1n32x5 FILLER_234_1123 ();
 b15zdnd11an1n16x5 FILLER_234_1155 ();
 b15zdnd11an1n08x5 FILLER_234_1171 ();
 b15zdnd00an1n01x5 FILLER_234_1179 ();
 b15zdnd11an1n64x5 FILLER_234_1183 ();
 b15zdnd11an1n16x5 FILLER_234_1247 ();
 b15zdnd11an1n04x5 FILLER_234_1263 ();
 b15zdnd00an1n02x5 FILLER_234_1267 ();
 b15zdnd00an1n01x5 FILLER_234_1269 ();
 b15zdnd11an1n04x5 FILLER_234_1273 ();
 b15zdnd11an1n64x5 FILLER_234_1280 ();
 b15zdnd11an1n32x5 FILLER_234_1344 ();
 b15zdnd11an1n08x5 FILLER_234_1376 ();
 b15zdnd11an1n04x5 FILLER_234_1384 ();
 b15zdnd00an1n02x5 FILLER_234_1388 ();
 b15zdnd00an1n01x5 FILLER_234_1390 ();
 b15zdnd11an1n64x5 FILLER_234_1400 ();
 b15zdnd11an1n64x5 FILLER_234_1464 ();
 b15zdnd11an1n32x5 FILLER_234_1528 ();
 b15zdnd11an1n08x5 FILLER_234_1560 ();
 b15zdnd11an1n04x5 FILLER_234_1568 ();
 b15zdnd00an1n02x5 FILLER_234_1572 ();
 b15zdnd11an1n04x5 FILLER_234_1591 ();
 b15zdnd11an1n64x5 FILLER_234_1601 ();
 b15zdnd11an1n64x5 FILLER_234_1665 ();
 b15zdnd11an1n64x5 FILLER_234_1729 ();
 b15zdnd11an1n64x5 FILLER_234_1793 ();
 b15zdnd11an1n64x5 FILLER_234_1857 ();
 b15zdnd11an1n64x5 FILLER_234_1921 ();
 b15zdnd11an1n64x5 FILLER_234_1985 ();
 b15zdnd11an1n64x5 FILLER_234_2049 ();
 b15zdnd11an1n32x5 FILLER_234_2113 ();
 b15zdnd11an1n08x5 FILLER_234_2145 ();
 b15zdnd00an1n01x5 FILLER_234_2153 ();
 b15zdnd11an1n04x5 FILLER_234_2162 ();
 b15zdnd11an1n08x5 FILLER_234_2218 ();
 b15zdnd11an1n04x5 FILLER_234_2226 ();
 b15zdnd11an1n04x5 FILLER_234_2272 ();
 b15zdnd11an1n64x5 FILLER_235_0 ();
 b15zdnd11an1n32x5 FILLER_235_64 ();
 b15zdnd11an1n64x5 FILLER_235_127 ();
 b15zdnd11an1n64x5 FILLER_235_191 ();
 b15zdnd11an1n64x5 FILLER_235_255 ();
 b15zdnd11an1n64x5 FILLER_235_319 ();
 b15zdnd11an1n64x5 FILLER_235_383 ();
 b15zdnd11an1n64x5 FILLER_235_447 ();
 b15zdnd11an1n64x5 FILLER_235_511 ();
 b15zdnd11an1n64x5 FILLER_235_575 ();
 b15zdnd11an1n64x5 FILLER_235_639 ();
 b15zdnd11an1n16x5 FILLER_235_703 ();
 b15zdnd11an1n08x5 FILLER_235_719 ();
 b15zdnd11an1n04x5 FILLER_235_727 ();
 b15zdnd00an1n02x5 FILLER_235_731 ();
 b15zdnd00an1n01x5 FILLER_235_733 ();
 b15zdnd11an1n64x5 FILLER_235_776 ();
 b15zdnd11an1n64x5 FILLER_235_840 ();
 b15zdnd11an1n64x5 FILLER_235_904 ();
 b15zdnd11an1n08x5 FILLER_235_968 ();
 b15zdnd11an1n04x5 FILLER_235_976 ();
 b15zdnd00an1n01x5 FILLER_235_980 ();
 b15zdnd11an1n04x5 FILLER_235_1004 ();
 b15zdnd11an1n04x5 FILLER_235_1034 ();
 b15zdnd11an1n64x5 FILLER_235_1052 ();
 b15zdnd11an1n08x5 FILLER_235_1116 ();
 b15zdnd00an1n02x5 FILLER_235_1124 ();
 b15zdnd00an1n01x5 FILLER_235_1126 ();
 b15zdnd11an1n32x5 FILLER_235_1136 ();
 b15zdnd11an1n08x5 FILLER_235_1168 ();
 b15zdnd11an1n04x5 FILLER_235_1176 ();
 b15zdnd00an1n02x5 FILLER_235_1180 ();
 b15zdnd11an1n32x5 FILLER_235_1191 ();
 b15zdnd11an1n08x5 FILLER_235_1223 ();
 b15zdnd11an1n04x5 FILLER_235_1231 ();
 b15zdnd00an1n02x5 FILLER_235_1235 ();
 b15zdnd00an1n01x5 FILLER_235_1237 ();
 b15zdnd11an1n16x5 FILLER_235_1247 ();
 b15zdnd11an1n08x5 FILLER_235_1263 ();
 b15zdnd11an1n04x5 FILLER_235_1271 ();
 b15zdnd00an1n02x5 FILLER_235_1275 ();
 b15zdnd11an1n64x5 FILLER_235_1280 ();
 b15zdnd11an1n64x5 FILLER_235_1344 ();
 b15zdnd11an1n64x5 FILLER_235_1408 ();
 b15zdnd11an1n64x5 FILLER_235_1472 ();
 b15zdnd11an1n64x5 FILLER_235_1536 ();
 b15zdnd11an1n32x5 FILLER_235_1600 ();
 b15zdnd11an1n08x5 FILLER_235_1632 ();
 b15zdnd00an1n02x5 FILLER_235_1640 ();
 b15zdnd11an1n64x5 FILLER_235_1650 ();
 b15zdnd11an1n64x5 FILLER_235_1714 ();
 b15zdnd11an1n32x5 FILLER_235_1778 ();
 b15zdnd11an1n16x5 FILLER_235_1810 ();
 b15zdnd11an1n08x5 FILLER_235_1826 ();
 b15zdnd11an1n04x5 FILLER_235_1834 ();
 b15zdnd00an1n01x5 FILLER_235_1838 ();
 b15zdnd11an1n64x5 FILLER_235_1845 ();
 b15zdnd11an1n64x5 FILLER_235_1909 ();
 b15zdnd11an1n64x5 FILLER_235_1973 ();
 b15zdnd11an1n64x5 FILLER_235_2037 ();
 b15zdnd11an1n64x5 FILLER_235_2101 ();
 b15zdnd11an1n16x5 FILLER_235_2165 ();
 b15zdnd00an1n02x5 FILLER_235_2181 ();
 b15zdnd00an1n01x5 FILLER_235_2183 ();
 b15zdnd11an1n04x5 FILLER_235_2187 ();
 b15zdnd11an1n32x5 FILLER_235_2194 ();
 b15zdnd11an1n16x5 FILLER_235_2226 ();
 b15zdnd11an1n08x5 FILLER_235_2242 ();
 b15zdnd11an1n04x5 FILLER_235_2250 ();
 b15zdnd00an1n02x5 FILLER_235_2254 ();
 b15zdnd11an1n16x5 FILLER_235_2260 ();
 b15zdnd11an1n08x5 FILLER_235_2276 ();
 b15zdnd11an1n64x5 FILLER_236_8 ();
 b15zdnd11an1n64x5 FILLER_236_72 ();
 b15zdnd11an1n64x5 FILLER_236_136 ();
 b15zdnd11an1n64x5 FILLER_236_200 ();
 b15zdnd11an1n08x5 FILLER_236_264 ();
 b15zdnd00an1n02x5 FILLER_236_272 ();
 b15zdnd11an1n64x5 FILLER_236_280 ();
 b15zdnd11an1n32x5 FILLER_236_344 ();
 b15zdnd00an1n01x5 FILLER_236_376 ();
 b15zdnd11an1n64x5 FILLER_236_387 ();
 b15zdnd11an1n64x5 FILLER_236_451 ();
 b15zdnd11an1n64x5 FILLER_236_515 ();
 b15zdnd11an1n64x5 FILLER_236_579 ();
 b15zdnd11an1n64x5 FILLER_236_643 ();
 b15zdnd11an1n08x5 FILLER_236_707 ();
 b15zdnd00an1n02x5 FILLER_236_715 ();
 b15zdnd00an1n01x5 FILLER_236_717 ();
 b15zdnd11an1n64x5 FILLER_236_726 ();
 b15zdnd11an1n64x5 FILLER_236_790 ();
 b15zdnd11an1n64x5 FILLER_236_854 ();
 b15zdnd11an1n32x5 FILLER_236_918 ();
 b15zdnd00an1n01x5 FILLER_236_950 ();
 b15zdnd11an1n64x5 FILLER_236_971 ();
 b15zdnd11an1n32x5 FILLER_236_1035 ();
 b15zdnd11an1n16x5 FILLER_236_1067 ();
 b15zdnd11an1n08x5 FILLER_236_1083 ();
 b15zdnd00an1n01x5 FILLER_236_1091 ();
 b15zdnd11an1n16x5 FILLER_236_1106 ();
 b15zdnd00an1n02x5 FILLER_236_1122 ();
 b15zdnd11an1n64x5 FILLER_236_1138 ();
 b15zdnd11an1n64x5 FILLER_236_1202 ();
 b15zdnd11an1n64x5 FILLER_236_1266 ();
 b15zdnd11an1n64x5 FILLER_236_1330 ();
 b15zdnd11an1n64x5 FILLER_236_1394 ();
 b15zdnd11an1n64x5 FILLER_236_1458 ();
 b15zdnd11an1n64x5 FILLER_236_1522 ();
 b15zdnd11an1n64x5 FILLER_236_1586 ();
 b15zdnd11an1n64x5 FILLER_236_1650 ();
 b15zdnd11an1n32x5 FILLER_236_1714 ();
 b15zdnd11an1n16x5 FILLER_236_1746 ();
 b15zdnd11an1n08x5 FILLER_236_1762 ();
 b15zdnd00an1n02x5 FILLER_236_1770 ();
 b15zdnd00an1n01x5 FILLER_236_1772 ();
 b15zdnd11an1n64x5 FILLER_236_1777 ();
 b15zdnd11an1n64x5 FILLER_236_1841 ();
 b15zdnd11an1n16x5 FILLER_236_1905 ();
 b15zdnd11an1n04x5 FILLER_236_1921 ();
 b15zdnd00an1n02x5 FILLER_236_1925 ();
 b15zdnd11an1n64x5 FILLER_236_1930 ();
 b15zdnd11an1n64x5 FILLER_236_1994 ();
 b15zdnd11an1n64x5 FILLER_236_2058 ();
 b15zdnd11an1n32x5 FILLER_236_2122 ();
 b15zdnd11an1n16x5 FILLER_236_2162 ();
 b15zdnd11an1n08x5 FILLER_236_2178 ();
 b15zdnd11an1n04x5 FILLER_236_2186 ();
 b15zdnd11an1n64x5 FILLER_236_2193 ();
 b15zdnd11an1n16x5 FILLER_236_2257 ();
 b15zdnd00an1n02x5 FILLER_236_2273 ();
 b15zdnd00an1n01x5 FILLER_236_2275 ();
 b15zdnd11an1n08x5 FILLER_237_0 ();
 b15zdnd11an1n64x5 FILLER_237_13 ();
 b15zdnd11an1n64x5 FILLER_237_77 ();
 b15zdnd11an1n64x5 FILLER_237_141 ();
 b15zdnd11an1n64x5 FILLER_237_205 ();
 b15zdnd11an1n64x5 FILLER_237_269 ();
 b15zdnd11an1n64x5 FILLER_237_333 ();
 b15zdnd11an1n64x5 FILLER_237_397 ();
 b15zdnd11an1n64x5 FILLER_237_461 ();
 b15zdnd11an1n64x5 FILLER_237_525 ();
 b15zdnd11an1n64x5 FILLER_237_589 ();
 b15zdnd11an1n64x5 FILLER_237_653 ();
 b15zdnd11an1n64x5 FILLER_237_717 ();
 b15zdnd11an1n64x5 FILLER_237_781 ();
 b15zdnd11an1n64x5 FILLER_237_845 ();
 b15zdnd11an1n64x5 FILLER_237_909 ();
 b15zdnd11an1n32x5 FILLER_237_973 ();
 b15zdnd11an1n08x5 FILLER_237_1005 ();
 b15zdnd00an1n02x5 FILLER_237_1013 ();
 b15zdnd00an1n01x5 FILLER_237_1015 ();
 b15zdnd11an1n08x5 FILLER_237_1030 ();
 b15zdnd11an1n04x5 FILLER_237_1038 ();
 b15zdnd00an1n02x5 FILLER_237_1042 ();
 b15zdnd00an1n01x5 FILLER_237_1044 ();
 b15zdnd11an1n16x5 FILLER_237_1059 ();
 b15zdnd00an1n01x5 FILLER_237_1075 ();
 b15zdnd11an1n64x5 FILLER_237_1082 ();
 b15zdnd11an1n64x5 FILLER_237_1146 ();
 b15zdnd11an1n64x5 FILLER_237_1210 ();
 b15zdnd11an1n64x5 FILLER_237_1274 ();
 b15zdnd11an1n64x5 FILLER_237_1338 ();
 b15zdnd11an1n64x5 FILLER_237_1402 ();
 b15zdnd11an1n32x5 FILLER_237_1466 ();
 b15zdnd11an1n16x5 FILLER_237_1498 ();
 b15zdnd00an1n02x5 FILLER_237_1514 ();
 b15zdnd11an1n04x5 FILLER_237_1525 ();
 b15zdnd11an1n64x5 FILLER_237_1538 ();
 b15zdnd11an1n64x5 FILLER_237_1602 ();
 b15zdnd11an1n64x5 FILLER_237_1666 ();
 b15zdnd11an1n64x5 FILLER_237_1730 ();
 b15zdnd11an1n64x5 FILLER_237_1794 ();
 b15zdnd11an1n64x5 FILLER_237_1858 ();
 b15zdnd11an1n04x5 FILLER_237_1922 ();
 b15zdnd00an1n02x5 FILLER_237_1926 ();
 b15zdnd11an1n16x5 FILLER_237_1931 ();
 b15zdnd11an1n08x5 FILLER_237_1947 ();
 b15zdnd11an1n04x5 FILLER_237_1955 ();
 b15zdnd00an1n02x5 FILLER_237_1959 ();
 b15zdnd00an1n01x5 FILLER_237_1961 ();
 b15zdnd11an1n64x5 FILLER_237_1965 ();
 b15zdnd11an1n64x5 FILLER_237_2029 ();
 b15zdnd11an1n64x5 FILLER_237_2093 ();
 b15zdnd11an1n64x5 FILLER_237_2157 ();
 b15zdnd11an1n32x5 FILLER_237_2221 ();
 b15zdnd11an1n16x5 FILLER_237_2253 ();
 b15zdnd11an1n08x5 FILLER_237_2269 ();
 b15zdnd11an1n04x5 FILLER_237_2277 ();
 b15zdnd00an1n02x5 FILLER_237_2281 ();
 b15zdnd00an1n01x5 FILLER_237_2283 ();
 b15zdnd11an1n64x5 FILLER_238_8 ();
 b15zdnd11an1n64x5 FILLER_238_72 ();
 b15zdnd11an1n64x5 FILLER_238_136 ();
 b15zdnd11an1n64x5 FILLER_238_200 ();
 b15zdnd11an1n64x5 FILLER_238_264 ();
 b15zdnd11an1n64x5 FILLER_238_328 ();
 b15zdnd11an1n64x5 FILLER_238_392 ();
 b15zdnd11an1n64x5 FILLER_238_456 ();
 b15zdnd11an1n64x5 FILLER_238_520 ();
 b15zdnd11an1n32x5 FILLER_238_584 ();
 b15zdnd11an1n16x5 FILLER_238_616 ();
 b15zdnd11an1n08x5 FILLER_238_632 ();
 b15zdnd00an1n02x5 FILLER_238_640 ();
 b15zdnd11an1n32x5 FILLER_238_665 ();
 b15zdnd11an1n16x5 FILLER_238_697 ();
 b15zdnd11an1n04x5 FILLER_238_713 ();
 b15zdnd00an1n01x5 FILLER_238_717 ();
 b15zdnd11an1n64x5 FILLER_238_726 ();
 b15zdnd11an1n64x5 FILLER_238_790 ();
 b15zdnd11an1n64x5 FILLER_238_854 ();
 b15zdnd11an1n64x5 FILLER_238_918 ();
 b15zdnd11an1n16x5 FILLER_238_982 ();
 b15zdnd00an1n02x5 FILLER_238_998 ();
 b15zdnd00an1n01x5 FILLER_238_1000 ();
 b15zdnd11an1n64x5 FILLER_238_1027 ();
 b15zdnd11an1n64x5 FILLER_238_1091 ();
 b15zdnd11an1n64x5 FILLER_238_1155 ();
 b15zdnd11an1n64x5 FILLER_238_1219 ();
 b15zdnd11an1n64x5 FILLER_238_1283 ();
 b15zdnd11an1n64x5 FILLER_238_1347 ();
 b15zdnd11an1n16x5 FILLER_238_1411 ();
 b15zdnd11an1n04x5 FILLER_238_1427 ();
 b15zdnd00an1n01x5 FILLER_238_1431 ();
 b15zdnd11an1n64x5 FILLER_238_1441 ();
 b15zdnd11an1n64x5 FILLER_238_1505 ();
 b15zdnd11an1n64x5 FILLER_238_1569 ();
 b15zdnd11an1n64x5 FILLER_238_1633 ();
 b15zdnd11an1n64x5 FILLER_238_1697 ();
 b15zdnd11an1n32x5 FILLER_238_1761 ();
 b15zdnd11an1n16x5 FILLER_238_1793 ();
 b15zdnd11an1n04x5 FILLER_238_1809 ();
 b15zdnd00an1n01x5 FILLER_238_1813 ();
 b15zdnd11an1n64x5 FILLER_238_1818 ();
 b15zdnd11an1n16x5 FILLER_238_1882 ();
 b15zdnd11an1n04x5 FILLER_238_1898 ();
 b15zdnd00an1n02x5 FILLER_238_1902 ();
 b15zdnd00an1n01x5 FILLER_238_1904 ();
 b15zdnd11an1n04x5 FILLER_238_1957 ();
 b15zdnd11an1n04x5 FILLER_238_1964 ();
 b15zdnd00an1n01x5 FILLER_238_1968 ();
 b15zdnd11an1n64x5 FILLER_238_1972 ();
 b15zdnd11an1n16x5 FILLER_238_2036 ();
 b15zdnd00an1n02x5 FILLER_238_2052 ();
 b15zdnd00an1n01x5 FILLER_238_2054 ();
 b15zdnd11an1n64x5 FILLER_238_2060 ();
 b15zdnd11an1n16x5 FILLER_238_2124 ();
 b15zdnd11an1n08x5 FILLER_238_2140 ();
 b15zdnd11an1n04x5 FILLER_238_2148 ();
 b15zdnd00an1n02x5 FILLER_238_2152 ();
 b15zdnd11an1n64x5 FILLER_238_2162 ();
 b15zdnd11an1n32x5 FILLER_238_2226 ();
 b15zdnd11an1n16x5 FILLER_238_2258 ();
 b15zdnd00an1n02x5 FILLER_238_2274 ();
 b15zdnd11an1n08x5 FILLER_239_0 ();
 b15zdnd00an1n02x5 FILLER_239_8 ();
 b15zdnd11an1n04x5 FILLER_239_14 ();
 b15zdnd11an1n16x5 FILLER_239_22 ();
 b15zdnd11an1n08x5 FILLER_239_38 ();
 b15zdnd00an1n02x5 FILLER_239_46 ();
 b15zdnd11an1n16x5 FILLER_239_79 ();
 b15zdnd11an1n08x5 FILLER_239_95 ();
 b15zdnd11an1n04x5 FILLER_239_103 ();
 b15zdnd00an1n02x5 FILLER_239_107 ();
 b15zdnd00an1n01x5 FILLER_239_109 ();
 b15zdnd11an1n64x5 FILLER_239_125 ();
 b15zdnd11an1n64x5 FILLER_239_189 ();
 b15zdnd11an1n16x5 FILLER_239_253 ();
 b15zdnd11an1n04x5 FILLER_239_269 ();
 b15zdnd00an1n02x5 FILLER_239_273 ();
 b15zdnd11an1n08x5 FILLER_239_281 ();
 b15zdnd00an1n01x5 FILLER_239_289 ();
 b15zdnd11an1n32x5 FILLER_239_313 ();
 b15zdnd11an1n08x5 FILLER_239_345 ();
 b15zdnd11an1n04x5 FILLER_239_353 ();
 b15zdnd00an1n02x5 FILLER_239_357 ();
 b15zdnd00an1n01x5 FILLER_239_359 ();
 b15zdnd11an1n64x5 FILLER_239_380 ();
 b15zdnd11an1n16x5 FILLER_239_444 ();
 b15zdnd11an1n08x5 FILLER_239_460 ();
 b15zdnd11an1n64x5 FILLER_239_491 ();
 b15zdnd11an1n64x5 FILLER_239_555 ();
 b15zdnd11an1n16x5 FILLER_239_619 ();
 b15zdnd11an1n08x5 FILLER_239_635 ();
 b15zdnd11an1n04x5 FILLER_239_643 ();
 b15zdnd00an1n02x5 FILLER_239_647 ();
 b15zdnd11an1n64x5 FILLER_239_653 ();
 b15zdnd11an1n64x5 FILLER_239_717 ();
 b15zdnd11an1n04x5 FILLER_239_781 ();
 b15zdnd00an1n02x5 FILLER_239_785 ();
 b15zdnd11an1n32x5 FILLER_239_794 ();
 b15zdnd00an1n01x5 FILLER_239_826 ();
 b15zdnd11an1n64x5 FILLER_239_847 ();
 b15zdnd11an1n64x5 FILLER_239_911 ();
 b15zdnd11an1n32x5 FILLER_239_975 ();
 b15zdnd11an1n16x5 FILLER_239_1007 ();
 b15zdnd11an1n64x5 FILLER_239_1043 ();
 b15zdnd11an1n64x5 FILLER_239_1107 ();
 b15zdnd11an1n64x5 FILLER_239_1171 ();
 b15zdnd11an1n64x5 FILLER_239_1235 ();
 b15zdnd11an1n64x5 FILLER_239_1299 ();
 b15zdnd11an1n64x5 FILLER_239_1363 ();
 b15zdnd11an1n64x5 FILLER_239_1427 ();
 b15zdnd00an1n02x5 FILLER_239_1491 ();
 b15zdnd11an1n04x5 FILLER_239_1502 ();
 b15zdnd11an1n16x5 FILLER_239_1520 ();
 b15zdnd11an1n08x5 FILLER_239_1536 ();
 b15zdnd11an1n04x5 FILLER_239_1544 ();
 b15zdnd00an1n01x5 FILLER_239_1548 ();
 b15zdnd11an1n64x5 FILLER_239_1556 ();
 b15zdnd00an1n01x5 FILLER_239_1620 ();
 b15zdnd11an1n04x5 FILLER_239_1628 ();
 b15zdnd00an1n01x5 FILLER_239_1632 ();
 b15zdnd11an1n04x5 FILLER_239_1637 ();
 b15zdnd11an1n04x5 FILLER_239_1645 ();
 b15zdnd11an1n64x5 FILLER_239_1653 ();
 b15zdnd11an1n64x5 FILLER_239_1717 ();
 b15zdnd11an1n32x5 FILLER_239_1781 ();
 b15zdnd11an1n04x5 FILLER_239_1813 ();
 b15zdnd00an1n01x5 FILLER_239_1817 ();
 b15zdnd11an1n32x5 FILLER_239_1822 ();
 b15zdnd11an1n64x5 FILLER_239_1858 ();
 b15zdnd00an1n01x5 FILLER_239_1922 ();
 b15zdnd11an1n04x5 FILLER_239_1975 ();
 b15zdnd11an1n64x5 FILLER_239_1982 ();
 b15zdnd11an1n32x5 FILLER_239_2046 ();
 b15zdnd11an1n08x5 FILLER_239_2078 ();
 b15zdnd11an1n04x5 FILLER_239_2086 ();
 b15zdnd00an1n02x5 FILLER_239_2090 ();
 b15zdnd11an1n32x5 FILLER_239_2097 ();
 b15zdnd11an1n08x5 FILLER_239_2129 ();
 b15zdnd11an1n64x5 FILLER_239_2148 ();
 b15zdnd11an1n64x5 FILLER_239_2212 ();
 b15zdnd11an1n08x5 FILLER_239_2276 ();
 b15zdnd00an1n02x5 FILLER_240_8 ();
 b15zdnd11an1n04x5 FILLER_240_30 ();
 b15zdnd11an1n64x5 FILLER_240_59 ();
 b15zdnd11an1n64x5 FILLER_240_123 ();
 b15zdnd11an1n64x5 FILLER_240_187 ();
 b15zdnd11an1n64x5 FILLER_240_251 ();
 b15zdnd11an1n64x5 FILLER_240_315 ();
 b15zdnd11an1n08x5 FILLER_240_379 ();
 b15zdnd00an1n02x5 FILLER_240_387 ();
 b15zdnd00an1n01x5 FILLER_240_389 ();
 b15zdnd11an1n64x5 FILLER_240_401 ();
 b15zdnd11an1n32x5 FILLER_240_465 ();
 b15zdnd11an1n64x5 FILLER_240_509 ();
 b15zdnd11an1n64x5 FILLER_240_573 ();
 b15zdnd11an1n16x5 FILLER_240_637 ();
 b15zdnd11an1n08x5 FILLER_240_653 ();
 b15zdnd11an1n32x5 FILLER_240_681 ();
 b15zdnd11an1n04x5 FILLER_240_713 ();
 b15zdnd00an1n01x5 FILLER_240_717 ();
 b15zdnd11an1n64x5 FILLER_240_726 ();
 b15zdnd11an1n32x5 FILLER_240_790 ();
 b15zdnd11an1n32x5 FILLER_240_839 ();
 b15zdnd11an1n04x5 FILLER_240_871 ();
 b15zdnd00an1n02x5 FILLER_240_875 ();
 b15zdnd11an1n64x5 FILLER_240_885 ();
 b15zdnd11an1n08x5 FILLER_240_949 ();
 b15zdnd11an1n04x5 FILLER_240_957 ();
 b15zdnd00an1n02x5 FILLER_240_961 ();
 b15zdnd00an1n01x5 FILLER_240_963 ();
 b15zdnd11an1n08x5 FILLER_240_1006 ();
 b15zdnd11an1n04x5 FILLER_240_1014 ();
 b15zdnd11an1n64x5 FILLER_240_1032 ();
 b15zdnd11an1n64x5 FILLER_240_1096 ();
 b15zdnd11an1n64x5 FILLER_240_1160 ();
 b15zdnd11an1n64x5 FILLER_240_1224 ();
 b15zdnd11an1n64x5 FILLER_240_1288 ();
 b15zdnd11an1n64x5 FILLER_240_1352 ();
 b15zdnd11an1n64x5 FILLER_240_1416 ();
 b15zdnd11an1n32x5 FILLER_240_1480 ();
 b15zdnd11an1n16x5 FILLER_240_1512 ();
 b15zdnd11an1n04x5 FILLER_240_1528 ();
 b15zdnd00an1n01x5 FILLER_240_1532 ();
 b15zdnd11an1n64x5 FILLER_240_1547 ();
 b15zdnd11an1n64x5 FILLER_240_1611 ();
 b15zdnd11an1n64x5 FILLER_240_1675 ();
 b15zdnd11an1n64x5 FILLER_240_1739 ();
 b15zdnd11an1n16x5 FILLER_240_1803 ();
 b15zdnd11an1n08x5 FILLER_240_1819 ();
 b15zdnd11an1n04x5 FILLER_240_1827 ();
 b15zdnd11an1n32x5 FILLER_240_1835 ();
 b15zdnd11an1n08x5 FILLER_240_1867 ();
 b15zdnd00an1n01x5 FILLER_240_1875 ();
 b15zdnd11an1n32x5 FILLER_240_1880 ();
 b15zdnd11an1n08x5 FILLER_240_1912 ();
 b15zdnd11an1n04x5 FILLER_240_1920 ();
 b15zdnd11an1n04x5 FILLER_240_1976 ();
 b15zdnd11an1n04x5 FILLER_240_1983 ();
 b15zdnd11an1n64x5 FILLER_240_1990 ();
 b15zdnd11an1n64x5 FILLER_240_2054 ();
 b15zdnd11an1n32x5 FILLER_240_2118 ();
 b15zdnd11an1n04x5 FILLER_240_2150 ();
 b15zdnd11an1n32x5 FILLER_240_2162 ();
 b15zdnd11an1n16x5 FILLER_240_2194 ();
 b15zdnd00an1n02x5 FILLER_240_2210 ();
 b15zdnd00an1n01x5 FILLER_240_2212 ();
 b15zdnd11an1n32x5 FILLER_240_2222 ();
 b15zdnd11an1n16x5 FILLER_240_2254 ();
 b15zdnd11an1n04x5 FILLER_240_2270 ();
 b15zdnd00an1n02x5 FILLER_240_2274 ();
 b15zdnd11an1n64x5 FILLER_241_0 ();
 b15zdnd11an1n64x5 FILLER_241_64 ();
 b15zdnd11an1n64x5 FILLER_241_128 ();
 b15zdnd11an1n64x5 FILLER_241_192 ();
 b15zdnd11an1n64x5 FILLER_241_256 ();
 b15zdnd11an1n64x5 FILLER_241_320 ();
 b15zdnd11an1n64x5 FILLER_241_384 ();
 b15zdnd11an1n32x5 FILLER_241_448 ();
 b15zdnd11an1n16x5 FILLER_241_480 ();
 b15zdnd11an1n04x5 FILLER_241_496 ();
 b15zdnd00an1n02x5 FILLER_241_500 ();
 b15zdnd11an1n32x5 FILLER_241_522 ();
 b15zdnd11an1n04x5 FILLER_241_554 ();
 b15zdnd00an1n01x5 FILLER_241_558 ();
 b15zdnd11an1n64x5 FILLER_241_580 ();
 b15zdnd11an1n08x5 FILLER_241_644 ();
 b15zdnd00an1n02x5 FILLER_241_652 ();
 b15zdnd11an1n08x5 FILLER_241_670 ();
 b15zdnd11an1n64x5 FILLER_241_694 ();
 b15zdnd11an1n16x5 FILLER_241_758 ();
 b15zdnd11an1n04x5 FILLER_241_774 ();
 b15zdnd00an1n02x5 FILLER_241_778 ();
 b15zdnd11an1n64x5 FILLER_241_788 ();
 b15zdnd11an1n64x5 FILLER_241_852 ();
 b15zdnd11an1n64x5 FILLER_241_916 ();
 b15zdnd11an1n64x5 FILLER_241_980 ();
 b15zdnd11an1n64x5 FILLER_241_1044 ();
 b15zdnd11an1n64x5 FILLER_241_1108 ();
 b15zdnd11an1n64x5 FILLER_241_1172 ();
 b15zdnd11an1n64x5 FILLER_241_1236 ();
 b15zdnd11an1n64x5 FILLER_241_1300 ();
 b15zdnd11an1n32x5 FILLER_241_1364 ();
 b15zdnd11an1n08x5 FILLER_241_1396 ();
 b15zdnd11an1n04x5 FILLER_241_1404 ();
 b15zdnd00an1n02x5 FILLER_241_1408 ();
 b15zdnd00an1n01x5 FILLER_241_1410 ();
 b15zdnd11an1n64x5 FILLER_241_1431 ();
 b15zdnd11an1n64x5 FILLER_241_1495 ();
 b15zdnd11an1n64x5 FILLER_241_1559 ();
 b15zdnd11an1n64x5 FILLER_241_1623 ();
 b15zdnd11an1n64x5 FILLER_241_1687 ();
 b15zdnd00an1n02x5 FILLER_241_1751 ();
 b15zdnd00an1n01x5 FILLER_241_1753 ();
 b15zdnd11an1n64x5 FILLER_241_1757 ();
 b15zdnd11an1n64x5 FILLER_241_1821 ();
 b15zdnd11an1n16x5 FILLER_241_1885 ();
 b15zdnd11an1n04x5 FILLER_241_1901 ();
 b15zdnd00an1n01x5 FILLER_241_1905 ();
 b15zdnd11an1n04x5 FILLER_241_1933 ();
 b15zdnd11an1n64x5 FILLER_241_1989 ();
 b15zdnd11an1n16x5 FILLER_241_2053 ();
 b15zdnd11an1n08x5 FILLER_241_2069 ();
 b15zdnd00an1n02x5 FILLER_241_2077 ();
 b15zdnd11an1n64x5 FILLER_241_2103 ();
 b15zdnd11an1n64x5 FILLER_241_2167 ();
 b15zdnd11an1n32x5 FILLER_241_2231 ();
 b15zdnd11an1n16x5 FILLER_241_2263 ();
 b15zdnd11an1n04x5 FILLER_241_2279 ();
 b15zdnd00an1n01x5 FILLER_241_2283 ();
 b15zdnd11an1n64x5 FILLER_242_8 ();
 b15zdnd11an1n64x5 FILLER_242_72 ();
 b15zdnd11an1n64x5 FILLER_242_136 ();
 b15zdnd11an1n64x5 FILLER_242_200 ();
 b15zdnd11an1n64x5 FILLER_242_264 ();
 b15zdnd11an1n64x5 FILLER_242_328 ();
 b15zdnd11an1n64x5 FILLER_242_392 ();
 b15zdnd11an1n32x5 FILLER_242_456 ();
 b15zdnd11an1n04x5 FILLER_242_488 ();
 b15zdnd00an1n02x5 FILLER_242_492 ();
 b15zdnd11an1n32x5 FILLER_242_512 ();
 b15zdnd11an1n16x5 FILLER_242_544 ();
 b15zdnd00an1n01x5 FILLER_242_560 ();
 b15zdnd11an1n64x5 FILLER_242_565 ();
 b15zdnd11an1n16x5 FILLER_242_629 ();
 b15zdnd11an1n08x5 FILLER_242_645 ();
 b15zdnd00an1n02x5 FILLER_242_653 ();
 b15zdnd00an1n01x5 FILLER_242_655 ();
 b15zdnd11an1n04x5 FILLER_242_661 ();
 b15zdnd11an1n08x5 FILLER_242_688 ();
 b15zdnd11an1n08x5 FILLER_242_710 ();
 b15zdnd11an1n64x5 FILLER_242_726 ();
 b15zdnd11an1n64x5 FILLER_242_790 ();
 b15zdnd11an1n64x5 FILLER_242_854 ();
 b15zdnd11an1n64x5 FILLER_242_918 ();
 b15zdnd11an1n64x5 FILLER_242_982 ();
 b15zdnd11an1n64x5 FILLER_242_1046 ();
 b15zdnd11an1n64x5 FILLER_242_1110 ();
 b15zdnd11an1n64x5 FILLER_242_1174 ();
 b15zdnd11an1n64x5 FILLER_242_1247 ();
 b15zdnd11an1n64x5 FILLER_242_1311 ();
 b15zdnd11an1n64x5 FILLER_242_1375 ();
 b15zdnd11an1n64x5 FILLER_242_1439 ();
 b15zdnd11an1n64x5 FILLER_242_1503 ();
 b15zdnd11an1n64x5 FILLER_242_1567 ();
 b15zdnd11an1n64x5 FILLER_242_1631 ();
 b15zdnd11an1n32x5 FILLER_242_1695 ();
 b15zdnd00an1n02x5 FILLER_242_1727 ();
 b15zdnd11an1n16x5 FILLER_242_1781 ();
 b15zdnd11an1n08x5 FILLER_242_1797 ();
 b15zdnd00an1n02x5 FILLER_242_1805 ();
 b15zdnd00an1n01x5 FILLER_242_1807 ();
 b15zdnd11an1n32x5 FILLER_242_1850 ();
 b15zdnd11an1n16x5 FILLER_242_1882 ();
 b15zdnd11an1n08x5 FILLER_242_1898 ();
 b15zdnd00an1n01x5 FILLER_242_1906 ();
 b15zdnd11an1n32x5 FILLER_242_1910 ();
 b15zdnd11an1n04x5 FILLER_242_1942 ();
 b15zdnd00an1n01x5 FILLER_242_1946 ();
 b15zdnd11an1n04x5 FILLER_242_1950 ();
 b15zdnd11an1n04x5 FILLER_242_1957 ();
 b15zdnd11an1n64x5 FILLER_242_1964 ();
 b15zdnd11an1n64x5 FILLER_242_2028 ();
 b15zdnd11an1n32x5 FILLER_242_2092 ();
 b15zdnd11an1n16x5 FILLER_242_2124 ();
 b15zdnd11an1n08x5 FILLER_242_2140 ();
 b15zdnd11an1n04x5 FILLER_242_2148 ();
 b15zdnd00an1n02x5 FILLER_242_2152 ();
 b15zdnd11an1n64x5 FILLER_242_2162 ();
 b15zdnd11an1n32x5 FILLER_242_2226 ();
 b15zdnd11an1n16x5 FILLER_242_2258 ();
 b15zdnd00an1n02x5 FILLER_242_2274 ();
 b15zdnd11an1n08x5 FILLER_243_0 ();
 b15zdnd11an1n32x5 FILLER_243_13 ();
 b15zdnd11an1n16x5 FILLER_243_45 ();
 b15zdnd11an1n04x5 FILLER_243_61 ();
 b15zdnd00an1n01x5 FILLER_243_65 ();
 b15zdnd11an1n04x5 FILLER_243_73 ();
 b15zdnd11an1n04x5 FILLER_243_116 ();
 b15zdnd00an1n02x5 FILLER_243_120 ();
 b15zdnd11an1n64x5 FILLER_243_146 ();
 b15zdnd11an1n64x5 FILLER_243_210 ();
 b15zdnd11an1n64x5 FILLER_243_274 ();
 b15zdnd11an1n32x5 FILLER_243_338 ();
 b15zdnd11an1n16x5 FILLER_243_370 ();
 b15zdnd11an1n08x5 FILLER_243_386 ();
 b15zdnd00an1n02x5 FILLER_243_394 ();
 b15zdnd11an1n16x5 FILLER_243_412 ();
 b15zdnd11an1n04x5 FILLER_243_428 ();
 b15zdnd00an1n02x5 FILLER_243_432 ();
 b15zdnd11an1n64x5 FILLER_243_458 ();
 b15zdnd11an1n32x5 FILLER_243_522 ();
 b15zdnd11an1n16x5 FILLER_243_554 ();
 b15zdnd00an1n02x5 FILLER_243_570 ();
 b15zdnd11an1n32x5 FILLER_243_578 ();
 b15zdnd00an1n02x5 FILLER_243_610 ();
 b15zdnd11an1n64x5 FILLER_243_624 ();
 b15zdnd11an1n64x5 FILLER_243_688 ();
 b15zdnd11an1n64x5 FILLER_243_752 ();
 b15zdnd11an1n64x5 FILLER_243_816 ();
 b15zdnd11an1n64x5 FILLER_243_880 ();
 b15zdnd11an1n64x5 FILLER_243_944 ();
 b15zdnd11an1n64x5 FILLER_243_1008 ();
 b15zdnd11an1n64x5 FILLER_243_1072 ();
 b15zdnd11an1n64x5 FILLER_243_1136 ();
 b15zdnd11an1n64x5 FILLER_243_1200 ();
 b15zdnd11an1n64x5 FILLER_243_1264 ();
 b15zdnd11an1n64x5 FILLER_243_1328 ();
 b15zdnd11an1n64x5 FILLER_243_1392 ();
 b15zdnd11an1n64x5 FILLER_243_1456 ();
 b15zdnd11an1n64x5 FILLER_243_1520 ();
 b15zdnd11an1n64x5 FILLER_243_1584 ();
 b15zdnd11an1n64x5 FILLER_243_1648 ();
 b15zdnd11an1n16x5 FILLER_243_1712 ();
 b15zdnd11an1n04x5 FILLER_243_1728 ();
 b15zdnd00an1n02x5 FILLER_243_1732 ();
 b15zdnd11an1n04x5 FILLER_243_1776 ();
 b15zdnd00an1n02x5 FILLER_243_1780 ();
 b15zdnd00an1n01x5 FILLER_243_1782 ();
 b15zdnd11an1n08x5 FILLER_243_1825 ();
 b15zdnd00an1n02x5 FILLER_243_1833 ();
 b15zdnd00an1n01x5 FILLER_243_1835 ();
 b15zdnd11an1n16x5 FILLER_243_1844 ();
 b15zdnd11an1n08x5 FILLER_243_1860 ();
 b15zdnd11an1n04x5 FILLER_243_1868 ();
 b15zdnd00an1n02x5 FILLER_243_1872 ();
 b15zdnd00an1n01x5 FILLER_243_1874 ();
 b15zdnd11an1n32x5 FILLER_243_1917 ();
 b15zdnd00an1n02x5 FILLER_243_1949 ();
 b15zdnd11an1n04x5 FILLER_243_1954 ();
 b15zdnd11an1n04x5 FILLER_243_2003 ();
 b15zdnd11an1n64x5 FILLER_243_2014 ();
 b15zdnd11an1n64x5 FILLER_243_2078 ();
 b15zdnd11an1n64x5 FILLER_243_2142 ();
 b15zdnd11an1n64x5 FILLER_243_2206 ();
 b15zdnd11an1n08x5 FILLER_243_2270 ();
 b15zdnd11an1n04x5 FILLER_243_2278 ();
 b15zdnd00an1n02x5 FILLER_243_2282 ();
 b15zdnd11an1n08x5 FILLER_244_8 ();
 b15zdnd00an1n02x5 FILLER_244_16 ();
 b15zdnd00an1n01x5 FILLER_244_18 ();
 b15zdnd11an1n04x5 FILLER_244_25 ();
 b15zdnd11an1n32x5 FILLER_244_34 ();
 b15zdnd11an1n08x5 FILLER_244_66 ();
 b15zdnd11an1n04x5 FILLER_244_74 ();
 b15zdnd00an1n02x5 FILLER_244_78 ();
 b15zdnd00an1n01x5 FILLER_244_80 ();
 b15zdnd11an1n64x5 FILLER_244_107 ();
 b15zdnd11an1n64x5 FILLER_244_171 ();
 b15zdnd11an1n64x5 FILLER_244_235 ();
 b15zdnd11an1n64x5 FILLER_244_299 ();
 b15zdnd11an1n64x5 FILLER_244_363 ();
 b15zdnd11an1n64x5 FILLER_244_427 ();
 b15zdnd11an1n64x5 FILLER_244_491 ();
 b15zdnd11an1n08x5 FILLER_244_555 ();
 b15zdnd11an1n04x5 FILLER_244_563 ();
 b15zdnd00an1n01x5 FILLER_244_567 ();
 b15zdnd11an1n08x5 FILLER_244_578 ();
 b15zdnd11an1n04x5 FILLER_244_586 ();
 b15zdnd00an1n02x5 FILLER_244_590 ();
 b15zdnd00an1n01x5 FILLER_244_592 ();
 b15zdnd11an1n64x5 FILLER_244_600 ();
 b15zdnd11an1n32x5 FILLER_244_664 ();
 b15zdnd11an1n16x5 FILLER_244_696 ();
 b15zdnd11an1n04x5 FILLER_244_712 ();
 b15zdnd00an1n02x5 FILLER_244_716 ();
 b15zdnd11an1n64x5 FILLER_244_726 ();
 b15zdnd11an1n16x5 FILLER_244_790 ();
 b15zdnd11an1n08x5 FILLER_244_806 ();
 b15zdnd11an1n04x5 FILLER_244_814 ();
 b15zdnd11an1n64x5 FILLER_244_824 ();
 b15zdnd11an1n64x5 FILLER_244_888 ();
 b15zdnd11an1n64x5 FILLER_244_952 ();
 b15zdnd11an1n64x5 FILLER_244_1016 ();
 b15zdnd11an1n32x5 FILLER_244_1080 ();
 b15zdnd11an1n08x5 FILLER_244_1112 ();
 b15zdnd11an1n04x5 FILLER_244_1120 ();
 b15zdnd00an1n01x5 FILLER_244_1124 ();
 b15zdnd11an1n64x5 FILLER_244_1167 ();
 b15zdnd11an1n04x5 FILLER_244_1231 ();
 b15zdnd00an1n02x5 FILLER_244_1235 ();
 b15zdnd00an1n01x5 FILLER_244_1237 ();
 b15zdnd11an1n64x5 FILLER_244_1247 ();
 b15zdnd11an1n64x5 FILLER_244_1311 ();
 b15zdnd11an1n64x5 FILLER_244_1375 ();
 b15zdnd11an1n32x5 FILLER_244_1439 ();
 b15zdnd11an1n16x5 FILLER_244_1471 ();
 b15zdnd11an1n64x5 FILLER_244_1493 ();
 b15zdnd11an1n64x5 FILLER_244_1557 ();
 b15zdnd11an1n16x5 FILLER_244_1621 ();
 b15zdnd11an1n16x5 FILLER_244_1641 ();
 b15zdnd00an1n02x5 FILLER_244_1657 ();
 b15zdnd11an1n64x5 FILLER_244_1667 ();
 b15zdnd11an1n04x5 FILLER_244_1731 ();
 b15zdnd00an1n01x5 FILLER_244_1735 ();
 b15zdnd11an1n04x5 FILLER_244_1743 ();
 b15zdnd00an1n01x5 FILLER_244_1747 ();
 b15zdnd11an1n04x5 FILLER_244_1751 ();
 b15zdnd11an1n08x5 FILLER_244_1758 ();
 b15zdnd00an1n02x5 FILLER_244_1766 ();
 b15zdnd11an1n64x5 FILLER_244_1794 ();
 b15zdnd11an1n64x5 FILLER_244_1858 ();
 b15zdnd11an1n64x5 FILLER_244_1922 ();
 b15zdnd11an1n64x5 FILLER_244_1986 ();
 b15zdnd11an1n64x5 FILLER_244_2050 ();
 b15zdnd11an1n04x5 FILLER_244_2114 ();
 b15zdnd11an1n16x5 FILLER_244_2129 ();
 b15zdnd11an1n08x5 FILLER_244_2145 ();
 b15zdnd00an1n01x5 FILLER_244_2153 ();
 b15zdnd11an1n64x5 FILLER_244_2162 ();
 b15zdnd11an1n16x5 FILLER_244_2226 ();
 b15zdnd11an1n08x5 FILLER_244_2242 ();
 b15zdnd11an1n16x5 FILLER_244_2256 ();
 b15zdnd11an1n04x5 FILLER_244_2272 ();
 b15zdnd11an1n16x5 FILLER_245_0 ();
 b15zdnd11an1n04x5 FILLER_245_16 ();
 b15zdnd00an1n01x5 FILLER_245_20 ();
 b15zdnd11an1n32x5 FILLER_245_26 ();
 b15zdnd11an1n16x5 FILLER_245_58 ();
 b15zdnd11an1n64x5 FILLER_245_105 ();
 b15zdnd11an1n64x5 FILLER_245_169 ();
 b15zdnd11an1n64x5 FILLER_245_233 ();
 b15zdnd11an1n64x5 FILLER_245_297 ();
 b15zdnd11an1n64x5 FILLER_245_361 ();
 b15zdnd11an1n64x5 FILLER_245_425 ();
 b15zdnd11an1n16x5 FILLER_245_489 ();
 b15zdnd11an1n08x5 FILLER_245_505 ();
 b15zdnd00an1n02x5 FILLER_245_513 ();
 b15zdnd00an1n01x5 FILLER_245_515 ();
 b15zdnd11an1n32x5 FILLER_245_532 ();
 b15zdnd11an1n08x5 FILLER_245_564 ();
 b15zdnd11an1n04x5 FILLER_245_572 ();
 b15zdnd00an1n02x5 FILLER_245_576 ();
 b15zdnd00an1n01x5 FILLER_245_578 ();
 b15zdnd11an1n16x5 FILLER_245_602 ();
 b15zdnd11an1n08x5 FILLER_245_618 ();
 b15zdnd11an1n04x5 FILLER_245_626 ();
 b15zdnd00an1n02x5 FILLER_245_630 ();
 b15zdnd11an1n16x5 FILLER_245_644 ();
 b15zdnd11an1n08x5 FILLER_245_660 ();
 b15zdnd11an1n64x5 FILLER_245_684 ();
 b15zdnd11an1n32x5 FILLER_245_748 ();
 b15zdnd11an1n16x5 FILLER_245_780 ();
 b15zdnd11an1n16x5 FILLER_245_803 ();
 b15zdnd00an1n01x5 FILLER_245_819 ();
 b15zdnd11an1n08x5 FILLER_245_827 ();
 b15zdnd00an1n02x5 FILLER_245_835 ();
 b15zdnd11an1n64x5 FILLER_245_857 ();
 b15zdnd11an1n64x5 FILLER_245_921 ();
 b15zdnd11an1n08x5 FILLER_245_985 ();
 b15zdnd11an1n04x5 FILLER_245_993 ();
 b15zdnd00an1n02x5 FILLER_245_997 ();
 b15zdnd00an1n01x5 FILLER_245_999 ();
 b15zdnd11an1n32x5 FILLER_245_1006 ();
 b15zdnd11an1n04x5 FILLER_245_1038 ();
 b15zdnd00an1n02x5 FILLER_245_1042 ();
 b15zdnd11an1n64x5 FILLER_245_1064 ();
 b15zdnd11an1n64x5 FILLER_245_1128 ();
 b15zdnd11an1n32x5 FILLER_245_1192 ();
 b15zdnd11an1n04x5 FILLER_245_1224 ();
 b15zdnd00an1n01x5 FILLER_245_1228 ();
 b15zdnd11an1n64x5 FILLER_245_1271 ();
 b15zdnd11an1n32x5 FILLER_245_1335 ();
 b15zdnd11an1n16x5 FILLER_245_1367 ();
 b15zdnd11an1n08x5 FILLER_245_1383 ();
 b15zdnd11an1n04x5 FILLER_245_1391 ();
 b15zdnd00an1n02x5 FILLER_245_1395 ();
 b15zdnd00an1n01x5 FILLER_245_1397 ();
 b15zdnd11an1n64x5 FILLER_245_1418 ();
 b15zdnd11an1n64x5 FILLER_245_1482 ();
 b15zdnd11an1n64x5 FILLER_245_1546 ();
 b15zdnd11an1n16x5 FILLER_245_1610 ();
 b15zdnd11an1n08x5 FILLER_245_1626 ();
 b15zdnd00an1n01x5 FILLER_245_1634 ();
 b15zdnd11an1n32x5 FILLER_245_1645 ();
 b15zdnd00an1n02x5 FILLER_245_1677 ();
 b15zdnd11an1n16x5 FILLER_245_1691 ();
 b15zdnd11an1n08x5 FILLER_245_1707 ();
 b15zdnd00an1n01x5 FILLER_245_1715 ();
 b15zdnd11an1n16x5 FILLER_245_1725 ();
 b15zdnd11an1n08x5 FILLER_245_1741 ();
 b15zdnd00an1n01x5 FILLER_245_1749 ();
 b15zdnd11an1n64x5 FILLER_245_1762 ();
 b15zdnd11an1n64x5 FILLER_245_1826 ();
 b15zdnd11an1n32x5 FILLER_245_1890 ();
 b15zdnd11an1n08x5 FILLER_245_1922 ();
 b15zdnd00an1n02x5 FILLER_245_1930 ();
 b15zdnd11an1n64x5 FILLER_245_1941 ();
 b15zdnd11an1n32x5 FILLER_245_2005 ();
 b15zdnd11an1n08x5 FILLER_245_2037 ();
 b15zdnd00an1n02x5 FILLER_245_2045 ();
 b15zdnd00an1n01x5 FILLER_245_2047 ();
 b15zdnd11an1n64x5 FILLER_245_2090 ();
 b15zdnd11an1n64x5 FILLER_245_2154 ();
 b15zdnd11an1n64x5 FILLER_245_2218 ();
 b15zdnd00an1n02x5 FILLER_245_2282 ();
 b15zdnd11an1n16x5 FILLER_246_8 ();
 b15zdnd11an1n64x5 FILLER_246_30 ();
 b15zdnd11an1n64x5 FILLER_246_94 ();
 b15zdnd11an1n64x5 FILLER_246_158 ();
 b15zdnd11an1n64x5 FILLER_246_222 ();
 b15zdnd11an1n64x5 FILLER_246_286 ();
 b15zdnd11an1n64x5 FILLER_246_350 ();
 b15zdnd11an1n32x5 FILLER_246_414 ();
 b15zdnd11an1n08x5 FILLER_246_446 ();
 b15zdnd11an1n32x5 FILLER_246_477 ();
 b15zdnd11an1n04x5 FILLER_246_525 ();
 b15zdnd11an1n16x5 FILLER_246_549 ();
 b15zdnd11an1n08x5 FILLER_246_565 ();
 b15zdnd00an1n02x5 FILLER_246_573 ();
 b15zdnd00an1n01x5 FILLER_246_575 ();
 b15zdnd11an1n04x5 FILLER_246_592 ();
 b15zdnd00an1n01x5 FILLER_246_596 ();
 b15zdnd11an1n64x5 FILLER_246_620 ();
 b15zdnd11an1n32x5 FILLER_246_684 ();
 b15zdnd00an1n02x5 FILLER_246_716 ();
 b15zdnd11an1n64x5 FILLER_246_726 ();
 b15zdnd11an1n16x5 FILLER_246_790 ();
 b15zdnd11an1n04x5 FILLER_246_806 ();
 b15zdnd00an1n01x5 FILLER_246_810 ();
 b15zdnd11an1n04x5 FILLER_246_817 ();
 b15zdnd11an1n64x5 FILLER_246_847 ();
 b15zdnd11an1n64x5 FILLER_246_911 ();
 b15zdnd11an1n32x5 FILLER_246_975 ();
 b15zdnd11an1n08x5 FILLER_246_1007 ();
 b15zdnd00an1n02x5 FILLER_246_1015 ();
 b15zdnd00an1n01x5 FILLER_246_1017 ();
 b15zdnd11an1n64x5 FILLER_246_1038 ();
 b15zdnd11an1n64x5 FILLER_246_1102 ();
 b15zdnd11an1n64x5 FILLER_246_1166 ();
 b15zdnd11an1n64x5 FILLER_246_1230 ();
 b15zdnd11an1n64x5 FILLER_246_1294 ();
 b15zdnd11an1n32x5 FILLER_246_1358 ();
 b15zdnd11an1n16x5 FILLER_246_1390 ();
 b15zdnd11an1n08x5 FILLER_246_1406 ();
 b15zdnd00an1n02x5 FILLER_246_1414 ();
 b15zdnd11an1n64x5 FILLER_246_1432 ();
 b15zdnd11an1n64x5 FILLER_246_1496 ();
 b15zdnd11an1n64x5 FILLER_246_1560 ();
 b15zdnd11an1n08x5 FILLER_246_1624 ();
 b15zdnd11an1n04x5 FILLER_246_1632 ();
 b15zdnd00an1n02x5 FILLER_246_1636 ();
 b15zdnd11an1n32x5 FILLER_246_1642 ();
 b15zdnd11an1n04x5 FILLER_246_1674 ();
 b15zdnd11an1n64x5 FILLER_246_1698 ();
 b15zdnd11an1n64x5 FILLER_246_1762 ();
 b15zdnd11an1n64x5 FILLER_246_1826 ();
 b15zdnd11an1n64x5 FILLER_246_1890 ();
 b15zdnd11an1n64x5 FILLER_246_1954 ();
 b15zdnd11an1n64x5 FILLER_246_2018 ();
 b15zdnd11an1n64x5 FILLER_246_2082 ();
 b15zdnd11an1n08x5 FILLER_246_2146 ();
 b15zdnd11an1n64x5 FILLER_246_2162 ();
 b15zdnd11an1n16x5 FILLER_246_2226 ();
 b15zdnd11an1n08x5 FILLER_246_2242 ();
 b15zdnd11an1n04x5 FILLER_246_2250 ();
 b15zdnd11an1n08x5 FILLER_246_2258 ();
 b15zdnd11an1n04x5 FILLER_246_2266 ();
 b15zdnd00an1n02x5 FILLER_246_2274 ();
 b15zdnd11an1n08x5 FILLER_247_0 ();
 b15zdnd11an1n04x5 FILLER_247_8 ();
 b15zdnd00an1n02x5 FILLER_247_12 ();
 b15zdnd11an1n32x5 FILLER_247_18 ();
 b15zdnd11an1n16x5 FILLER_247_50 ();
 b15zdnd00an1n02x5 FILLER_247_66 ();
 b15zdnd00an1n01x5 FILLER_247_68 ();
 b15zdnd11an1n16x5 FILLER_247_77 ();
 b15zdnd11an1n08x5 FILLER_247_93 ();
 b15zdnd11an1n04x5 FILLER_247_101 ();
 b15zdnd11an1n64x5 FILLER_247_129 ();
 b15zdnd11an1n08x5 FILLER_247_193 ();
 b15zdnd11an1n04x5 FILLER_247_201 ();
 b15zdnd11an1n64x5 FILLER_247_225 ();
 b15zdnd11an1n08x5 FILLER_247_289 ();
 b15zdnd00an1n01x5 FILLER_247_297 ();
 b15zdnd11an1n64x5 FILLER_247_308 ();
 b15zdnd11an1n16x5 FILLER_247_372 ();
 b15zdnd11an1n08x5 FILLER_247_388 ();
 b15zdnd11an1n04x5 FILLER_247_396 ();
 b15zdnd00an1n01x5 FILLER_247_400 ();
 b15zdnd11an1n16x5 FILLER_247_416 ();
 b15zdnd11an1n04x5 FILLER_247_432 ();
 b15zdnd00an1n02x5 FILLER_247_436 ();
 b15zdnd00an1n01x5 FILLER_247_438 ();
 b15zdnd11an1n16x5 FILLER_247_459 ();
 b15zdnd11an1n08x5 FILLER_247_475 ();
 b15zdnd00an1n02x5 FILLER_247_483 ();
 b15zdnd11an1n64x5 FILLER_247_495 ();
 b15zdnd11an1n16x5 FILLER_247_559 ();
 b15zdnd11an1n08x5 FILLER_247_575 ();
 b15zdnd00an1n02x5 FILLER_247_583 ();
 b15zdnd00an1n01x5 FILLER_247_585 ();
 b15zdnd11an1n08x5 FILLER_247_598 ();
 b15zdnd11an1n04x5 FILLER_247_606 ();
 b15zdnd00an1n01x5 FILLER_247_610 ();
 b15zdnd11an1n64x5 FILLER_247_621 ();
 b15zdnd11an1n64x5 FILLER_247_685 ();
 b15zdnd11an1n64x5 FILLER_247_749 ();
 b15zdnd11an1n04x5 FILLER_247_813 ();
 b15zdnd00an1n02x5 FILLER_247_817 ();
 b15zdnd00an1n01x5 FILLER_247_819 ();
 b15zdnd11an1n64x5 FILLER_247_827 ();
 b15zdnd11an1n32x5 FILLER_247_891 ();
 b15zdnd00an1n02x5 FILLER_247_923 ();
 b15zdnd11an1n04x5 FILLER_247_931 ();
 b15zdnd11an1n04x5 FILLER_247_938 ();
 b15zdnd11an1n64x5 FILLER_247_945 ();
 b15zdnd11an1n08x5 FILLER_247_1009 ();
 b15zdnd00an1n01x5 FILLER_247_1017 ();
 b15zdnd11an1n04x5 FILLER_247_1044 ();
 b15zdnd11an1n04x5 FILLER_247_1060 ();
 b15zdnd00an1n01x5 FILLER_247_1064 ();
 b15zdnd11an1n08x5 FILLER_247_1081 ();
 b15zdnd11an1n04x5 FILLER_247_1089 ();
 b15zdnd00an1n01x5 FILLER_247_1093 ();
 b15zdnd11an1n64x5 FILLER_247_1114 ();
 b15zdnd00an1n01x5 FILLER_247_1178 ();
 b15zdnd11an1n04x5 FILLER_247_1182 ();
 b15zdnd11an1n64x5 FILLER_247_1189 ();
 b15zdnd11an1n64x5 FILLER_247_1253 ();
 b15zdnd11an1n64x5 FILLER_247_1317 ();
 b15zdnd11an1n32x5 FILLER_247_1381 ();
 b15zdnd00an1n02x5 FILLER_247_1413 ();
 b15zdnd00an1n01x5 FILLER_247_1415 ();
 b15zdnd11an1n16x5 FILLER_247_1419 ();
 b15zdnd00an1n02x5 FILLER_247_1435 ();
 b15zdnd00an1n01x5 FILLER_247_1437 ();
 b15zdnd11an1n16x5 FILLER_247_1448 ();
 b15zdnd11an1n04x5 FILLER_247_1464 ();
 b15zdnd00an1n02x5 FILLER_247_1468 ();
 b15zdnd00an1n01x5 FILLER_247_1470 ();
 b15zdnd11an1n32x5 FILLER_247_1491 ();
 b15zdnd11an1n08x5 FILLER_247_1523 ();
 b15zdnd11an1n64x5 FILLER_247_1547 ();
 b15zdnd11an1n16x5 FILLER_247_1611 ();
 b15zdnd11an1n08x5 FILLER_247_1627 ();
 b15zdnd11an1n04x5 FILLER_247_1635 ();
 b15zdnd00an1n01x5 FILLER_247_1639 ();
 b15zdnd11an1n32x5 FILLER_247_1646 ();
 b15zdnd11an1n04x5 FILLER_247_1678 ();
 b15zdnd00an1n02x5 FILLER_247_1682 ();
 b15zdnd00an1n01x5 FILLER_247_1684 ();
 b15zdnd11an1n64x5 FILLER_247_1696 ();
 b15zdnd11an1n64x5 FILLER_247_1760 ();
 b15zdnd11an1n64x5 FILLER_247_1824 ();
 b15zdnd11an1n64x5 FILLER_247_1888 ();
 b15zdnd11an1n64x5 FILLER_247_1952 ();
 b15zdnd11an1n64x5 FILLER_247_2016 ();
 b15zdnd11an1n64x5 FILLER_247_2080 ();
 b15zdnd11an1n64x5 FILLER_247_2144 ();
 b15zdnd11an1n32x5 FILLER_247_2208 ();
 b15zdnd11an1n08x5 FILLER_247_2240 ();
 b15zdnd11an1n04x5 FILLER_247_2248 ();
 b15zdnd11an1n16x5 FILLER_247_2256 ();
 b15zdnd11an1n08x5 FILLER_247_2272 ();
 b15zdnd11an1n04x5 FILLER_247_2280 ();
 b15zdnd11an1n04x5 FILLER_248_8 ();
 b15zdnd00an1n01x5 FILLER_248_12 ();
 b15zdnd11an1n08x5 FILLER_248_19 ();
 b15zdnd11an1n04x5 FILLER_248_27 ();
 b15zdnd00an1n01x5 FILLER_248_31 ();
 b15zdnd11an1n08x5 FILLER_248_36 ();
 b15zdnd11an1n04x5 FILLER_248_44 ();
 b15zdnd00an1n02x5 FILLER_248_48 ();
 b15zdnd11an1n04x5 FILLER_248_70 ();
 b15zdnd11an1n64x5 FILLER_248_78 ();
 b15zdnd11an1n64x5 FILLER_248_142 ();
 b15zdnd11an1n64x5 FILLER_248_216 ();
 b15zdnd11an1n64x5 FILLER_248_280 ();
 b15zdnd11an1n64x5 FILLER_248_344 ();
 b15zdnd11an1n64x5 FILLER_248_408 ();
 b15zdnd11an1n64x5 FILLER_248_472 ();
 b15zdnd11an1n64x5 FILLER_248_536 ();
 b15zdnd11an1n64x5 FILLER_248_600 ();
 b15zdnd11an1n32x5 FILLER_248_664 ();
 b15zdnd11an1n16x5 FILLER_248_696 ();
 b15zdnd11an1n04x5 FILLER_248_712 ();
 b15zdnd00an1n02x5 FILLER_248_716 ();
 b15zdnd11an1n64x5 FILLER_248_726 ();
 b15zdnd11an1n32x5 FILLER_248_790 ();
 b15zdnd00an1n02x5 FILLER_248_822 ();
 b15zdnd11an1n32x5 FILLER_248_866 ();
 b15zdnd11an1n08x5 FILLER_248_898 ();
 b15zdnd11an1n32x5 FILLER_248_946 ();
 b15zdnd11an1n16x5 FILLER_248_978 ();
 b15zdnd11an1n04x5 FILLER_248_1015 ();
 b15zdnd11an1n08x5 FILLER_248_1039 ();
 b15zdnd11an1n64x5 FILLER_248_1057 ();
 b15zdnd11an1n32x5 FILLER_248_1121 ();
 b15zdnd11an1n08x5 FILLER_248_1153 ();
 b15zdnd11an1n64x5 FILLER_248_1213 ();
 b15zdnd11an1n64x5 FILLER_248_1277 ();
 b15zdnd11an1n64x5 FILLER_248_1341 ();
 b15zdnd00an1n02x5 FILLER_248_1405 ();
 b15zdnd11an1n16x5 FILLER_248_1420 ();
 b15zdnd00an1n01x5 FILLER_248_1436 ();
 b15zdnd11an1n32x5 FILLER_248_1440 ();
 b15zdnd00an1n02x5 FILLER_248_1472 ();
 b15zdnd00an1n01x5 FILLER_248_1474 ();
 b15zdnd11an1n08x5 FILLER_248_1517 ();
 b15zdnd00an1n01x5 FILLER_248_1525 ();
 b15zdnd11an1n64x5 FILLER_248_1533 ();
 b15zdnd11an1n64x5 FILLER_248_1597 ();
 b15zdnd11an1n64x5 FILLER_248_1661 ();
 b15zdnd11an1n64x5 FILLER_248_1725 ();
 b15zdnd11an1n04x5 FILLER_248_1795 ();
 b15zdnd00an1n01x5 FILLER_248_1799 ();
 b15zdnd11an1n32x5 FILLER_248_1806 ();
 b15zdnd00an1n02x5 FILLER_248_1838 ();
 b15zdnd11an1n64x5 FILLER_248_1860 ();
 b15zdnd11an1n64x5 FILLER_248_1924 ();
 b15zdnd11an1n64x5 FILLER_248_1988 ();
 b15zdnd11an1n64x5 FILLER_248_2052 ();
 b15zdnd11an1n32x5 FILLER_248_2116 ();
 b15zdnd11an1n04x5 FILLER_248_2148 ();
 b15zdnd00an1n02x5 FILLER_248_2152 ();
 b15zdnd11an1n32x5 FILLER_248_2162 ();
 b15zdnd11an1n08x5 FILLER_248_2194 ();
 b15zdnd00an1n02x5 FILLER_248_2202 ();
 b15zdnd11an1n64x5 FILLER_248_2208 ();
 b15zdnd11an1n04x5 FILLER_248_2272 ();
 b15zdnd11an1n04x5 FILLER_249_0 ();
 b15zdnd00an1n02x5 FILLER_249_4 ();
 b15zdnd11an1n04x5 FILLER_249_20 ();
 b15zdnd11an1n64x5 FILLER_249_76 ();
 b15zdnd11an1n64x5 FILLER_249_140 ();
 b15zdnd11an1n64x5 FILLER_249_204 ();
 b15zdnd11an1n32x5 FILLER_249_268 ();
 b15zdnd11an1n04x5 FILLER_249_300 ();
 b15zdnd00an1n02x5 FILLER_249_304 ();
 b15zdnd11an1n04x5 FILLER_249_318 ();
 b15zdnd11an1n08x5 FILLER_249_340 ();
 b15zdnd11an1n04x5 FILLER_249_348 ();
 b15zdnd00an1n01x5 FILLER_249_352 ();
 b15zdnd11an1n64x5 FILLER_249_371 ();
 b15zdnd11an1n32x5 FILLER_249_435 ();
 b15zdnd11an1n16x5 FILLER_249_467 ();
 b15zdnd00an1n01x5 FILLER_249_483 ();
 b15zdnd11an1n64x5 FILLER_249_506 ();
 b15zdnd11an1n64x5 FILLER_249_570 ();
 b15zdnd11an1n64x5 FILLER_249_634 ();
 b15zdnd11an1n64x5 FILLER_249_698 ();
 b15zdnd11an1n64x5 FILLER_249_762 ();
 b15zdnd11an1n08x5 FILLER_249_826 ();
 b15zdnd00an1n02x5 FILLER_249_834 ();
 b15zdnd00an1n01x5 FILLER_249_836 ();
 b15zdnd11an1n64x5 FILLER_249_879 ();
 b15zdnd00an1n01x5 FILLER_249_943 ();
 b15zdnd11an1n32x5 FILLER_249_948 ();
 b15zdnd11an1n16x5 FILLER_249_980 ();
 b15zdnd00an1n01x5 FILLER_249_996 ();
 b15zdnd11an1n16x5 FILLER_249_1029 ();
 b15zdnd11an1n64x5 FILLER_249_1077 ();
 b15zdnd11an1n32x5 FILLER_249_1141 ();
 b15zdnd11an1n08x5 FILLER_249_1173 ();
 b15zdnd11an1n04x5 FILLER_249_1181 ();
 b15zdnd00an1n02x5 FILLER_249_1185 ();
 b15zdnd11an1n04x5 FILLER_249_1190 ();
 b15zdnd00an1n02x5 FILLER_249_1194 ();
 b15zdnd00an1n01x5 FILLER_249_1196 ();
 b15zdnd11an1n04x5 FILLER_249_1200 ();
 b15zdnd11an1n64x5 FILLER_249_1207 ();
 b15zdnd11an1n16x5 FILLER_249_1271 ();
 b15zdnd11an1n04x5 FILLER_249_1290 ();
 b15zdnd11an1n64x5 FILLER_249_1297 ();
 b15zdnd11an1n64x5 FILLER_249_1361 ();
 b15zdnd11an1n32x5 FILLER_249_1425 ();
 b15zdnd11an1n08x5 FILLER_249_1457 ();
 b15zdnd11an1n04x5 FILLER_249_1465 ();
 b15zdnd00an1n02x5 FILLER_249_1469 ();
 b15zdnd11an1n16x5 FILLER_249_1483 ();
 b15zdnd00an1n02x5 FILLER_249_1499 ();
 b15zdnd00an1n01x5 FILLER_249_1501 ();
 b15zdnd11an1n64x5 FILLER_249_1513 ();
 b15zdnd11an1n64x5 FILLER_249_1577 ();
 b15zdnd11an1n64x5 FILLER_249_1641 ();
 b15zdnd11an1n64x5 FILLER_249_1705 ();
 b15zdnd11an1n64x5 FILLER_249_1769 ();
 b15zdnd11an1n64x5 FILLER_249_1833 ();
 b15zdnd11an1n64x5 FILLER_249_1897 ();
 b15zdnd11an1n64x5 FILLER_249_1961 ();
 b15zdnd11an1n64x5 FILLER_249_2025 ();
 b15zdnd11an1n64x5 FILLER_249_2089 ();
 b15zdnd11an1n64x5 FILLER_249_2153 ();
 b15zdnd11an1n64x5 FILLER_249_2217 ();
 b15zdnd00an1n02x5 FILLER_249_2281 ();
 b15zdnd00an1n01x5 FILLER_249_2283 ();
 b15zdnd11an1n16x5 FILLER_250_8 ();
 b15zdnd11an1n04x5 FILLER_250_24 ();
 b15zdnd00an1n01x5 FILLER_250_28 ();
 b15zdnd11an1n04x5 FILLER_250_36 ();
 b15zdnd11an1n04x5 FILLER_250_43 ();
 b15zdnd11an1n04x5 FILLER_250_50 ();
 b15zdnd11an1n64x5 FILLER_250_57 ();
 b15zdnd11an1n64x5 FILLER_250_121 ();
 b15zdnd00an1n02x5 FILLER_250_185 ();
 b15zdnd00an1n01x5 FILLER_250_187 ();
 b15zdnd11an1n64x5 FILLER_250_203 ();
 b15zdnd11an1n32x5 FILLER_250_267 ();
 b15zdnd11an1n16x5 FILLER_250_299 ();
 b15zdnd00an1n02x5 FILLER_250_315 ();
 b15zdnd11an1n64x5 FILLER_250_336 ();
 b15zdnd11an1n32x5 FILLER_250_400 ();
 b15zdnd11an1n16x5 FILLER_250_432 ();
 b15zdnd11an1n08x5 FILLER_250_448 ();
 b15zdnd11an1n04x5 FILLER_250_456 ();
 b15zdnd00an1n02x5 FILLER_250_460 ();
 b15zdnd00an1n01x5 FILLER_250_462 ();
 b15zdnd11an1n64x5 FILLER_250_485 ();
 b15zdnd11an1n64x5 FILLER_250_549 ();
 b15zdnd11an1n64x5 FILLER_250_613 ();
 b15zdnd11an1n32x5 FILLER_250_677 ();
 b15zdnd11an1n08x5 FILLER_250_709 ();
 b15zdnd00an1n01x5 FILLER_250_717 ();
 b15zdnd11an1n64x5 FILLER_250_726 ();
 b15zdnd11an1n16x5 FILLER_250_790 ();
 b15zdnd11an1n04x5 FILLER_250_806 ();
 b15zdnd11an1n64x5 FILLER_250_852 ();
 b15zdnd11an1n04x5 FILLER_250_916 ();
 b15zdnd00an1n01x5 FILLER_250_920 ();
 b15zdnd11an1n32x5 FILLER_250_963 ();
 b15zdnd11an1n08x5 FILLER_250_995 ();
 b15zdnd11an1n04x5 FILLER_250_1029 ();
 b15zdnd11an1n64x5 FILLER_250_1059 ();
 b15zdnd11an1n32x5 FILLER_250_1123 ();
 b15zdnd11an1n16x5 FILLER_250_1155 ();
 b15zdnd00an1n01x5 FILLER_250_1171 ();
 b15zdnd11an1n32x5 FILLER_250_1224 ();
 b15zdnd11an1n08x5 FILLER_250_1256 ();
 b15zdnd11an1n04x5 FILLER_250_1264 ();
 b15zdnd00an1n01x5 FILLER_250_1268 ();
 b15zdnd11an1n64x5 FILLER_250_1321 ();
 b15zdnd11an1n32x5 FILLER_250_1385 ();
 b15zdnd11an1n04x5 FILLER_250_1417 ();
 b15zdnd11an1n04x5 FILLER_250_1424 ();
 b15zdnd11an1n04x5 FILLER_250_1431 ();
 b15zdnd11an1n16x5 FILLER_250_1455 ();
 b15zdnd11an1n08x5 FILLER_250_1471 ();
 b15zdnd00an1n01x5 FILLER_250_1479 ();
 b15zdnd11an1n64x5 FILLER_250_1501 ();
 b15zdnd11an1n64x5 FILLER_250_1565 ();
 b15zdnd11an1n64x5 FILLER_250_1629 ();
 b15zdnd11an1n64x5 FILLER_250_1693 ();
 b15zdnd11an1n64x5 FILLER_250_1757 ();
 b15zdnd11an1n64x5 FILLER_250_1821 ();
 b15zdnd11an1n64x5 FILLER_250_1885 ();
 b15zdnd11an1n64x5 FILLER_250_1949 ();
 b15zdnd11an1n64x5 FILLER_250_2013 ();
 b15zdnd11an1n64x5 FILLER_250_2077 ();
 b15zdnd11an1n08x5 FILLER_250_2141 ();
 b15zdnd11an1n04x5 FILLER_250_2149 ();
 b15zdnd00an1n01x5 FILLER_250_2153 ();
 b15zdnd11an1n64x5 FILLER_250_2162 ();
 b15zdnd11an1n32x5 FILLER_250_2226 ();
 b15zdnd11an1n16x5 FILLER_250_2258 ();
 b15zdnd00an1n02x5 FILLER_250_2274 ();
 b15zdnd11an1n08x5 FILLER_251_0 ();
 b15zdnd00an1n02x5 FILLER_251_8 ();
 b15zdnd11an1n08x5 FILLER_251_17 ();
 b15zdnd00an1n02x5 FILLER_251_25 ();
 b15zdnd11an1n32x5 FILLER_251_41 ();
 b15zdnd11an1n16x5 FILLER_251_73 ();
 b15zdnd11an1n08x5 FILLER_251_89 ();
 b15zdnd11an1n32x5 FILLER_251_128 ();
 b15zdnd11an1n16x5 FILLER_251_160 ();
 b15zdnd11an1n04x5 FILLER_251_176 ();
 b15zdnd00an1n02x5 FILLER_251_180 ();
 b15zdnd00an1n01x5 FILLER_251_182 ();
 b15zdnd11an1n64x5 FILLER_251_208 ();
 b15zdnd11an1n64x5 FILLER_251_272 ();
 b15zdnd11an1n32x5 FILLER_251_336 ();
 b15zdnd00an1n02x5 FILLER_251_368 ();
 b15zdnd11an1n32x5 FILLER_251_375 ();
 b15zdnd00an1n02x5 FILLER_251_407 ();
 b15zdnd00an1n01x5 FILLER_251_409 ();
 b15zdnd11an1n64x5 FILLER_251_452 ();
 b15zdnd11an1n64x5 FILLER_251_516 ();
 b15zdnd11an1n64x5 FILLER_251_580 ();
 b15zdnd11an1n64x5 FILLER_251_644 ();
 b15zdnd11an1n64x5 FILLER_251_708 ();
 b15zdnd11an1n32x5 FILLER_251_772 ();
 b15zdnd11an1n08x5 FILLER_251_804 ();
 b15zdnd11an1n04x5 FILLER_251_812 ();
 b15zdnd00an1n02x5 FILLER_251_816 ();
 b15zdnd00an1n01x5 FILLER_251_818 ();
 b15zdnd11an1n04x5 FILLER_251_822 ();
 b15zdnd00an1n02x5 FILLER_251_826 ();
 b15zdnd11an1n64x5 FILLER_251_831 ();
 b15zdnd11an1n16x5 FILLER_251_895 ();
 b15zdnd11an1n08x5 FILLER_251_911 ();
 b15zdnd11an1n04x5 FILLER_251_919 ();
 b15zdnd00an1n02x5 FILLER_251_923 ();
 b15zdnd00an1n01x5 FILLER_251_925 ();
 b15zdnd11an1n64x5 FILLER_251_937 ();
 b15zdnd11an1n04x5 FILLER_251_1001 ();
 b15zdnd00an1n02x5 FILLER_251_1005 ();
 b15zdnd11an1n16x5 FILLER_251_1027 ();
 b15zdnd00an1n02x5 FILLER_251_1043 ();
 b15zdnd11an1n04x5 FILLER_251_1048 ();
 b15zdnd00an1n02x5 FILLER_251_1052 ();
 b15zdnd11an1n04x5 FILLER_251_1057 ();
 b15zdnd11an1n64x5 FILLER_251_1071 ();
 b15zdnd11an1n32x5 FILLER_251_1135 ();
 b15zdnd11an1n16x5 FILLER_251_1167 ();
 b15zdnd11an1n08x5 FILLER_251_1183 ();
 b15zdnd11an1n04x5 FILLER_251_1191 ();
 b15zdnd00an1n02x5 FILLER_251_1195 ();
 b15zdnd11an1n32x5 FILLER_251_1200 ();
 b15zdnd11an1n16x5 FILLER_251_1232 ();
 b15zdnd11an1n08x5 FILLER_251_1248 ();
 b15zdnd11an1n04x5 FILLER_251_1256 ();
 b15zdnd00an1n01x5 FILLER_251_1260 ();
 b15zdnd11an1n04x5 FILLER_251_1313 ();
 b15zdnd11an1n64x5 FILLER_251_1320 ();
 b15zdnd11an1n08x5 FILLER_251_1384 ();
 b15zdnd11an1n04x5 FILLER_251_1392 ();
 b15zdnd00an1n02x5 FILLER_251_1396 ();
 b15zdnd00an1n01x5 FILLER_251_1398 ();
 b15zdnd11an1n64x5 FILLER_251_1443 ();
 b15zdnd11an1n04x5 FILLER_251_1507 ();
 b15zdnd11an1n04x5 FILLER_251_1525 ();
 b15zdnd11an1n04x5 FILLER_251_1534 ();
 b15zdnd11an1n64x5 FILLER_251_1547 ();
 b15zdnd11an1n64x5 FILLER_251_1611 ();
 b15zdnd11an1n64x5 FILLER_251_1675 ();
 b15zdnd11an1n08x5 FILLER_251_1739 ();
 b15zdnd11an1n04x5 FILLER_251_1747 ();
 b15zdnd11an1n64x5 FILLER_251_1761 ();
 b15zdnd11an1n64x5 FILLER_251_1825 ();
 b15zdnd11an1n64x5 FILLER_251_1889 ();
 b15zdnd00an1n02x5 FILLER_251_1953 ();
 b15zdnd00an1n01x5 FILLER_251_1955 ();
 b15zdnd11an1n64x5 FILLER_251_1965 ();
 b15zdnd11an1n64x5 FILLER_251_2029 ();
 b15zdnd11an1n64x5 FILLER_251_2093 ();
 b15zdnd11an1n64x5 FILLER_251_2157 ();
 b15zdnd11an1n32x5 FILLER_251_2221 ();
 b15zdnd11an1n16x5 FILLER_251_2253 ();
 b15zdnd11an1n08x5 FILLER_251_2269 ();
 b15zdnd11an1n04x5 FILLER_251_2277 ();
 b15zdnd00an1n02x5 FILLER_251_2281 ();
 b15zdnd00an1n01x5 FILLER_251_2283 ();
 b15zdnd11an1n64x5 FILLER_252_8 ();
 b15zdnd11an1n64x5 FILLER_252_72 ();
 b15zdnd11an1n64x5 FILLER_252_136 ();
 b15zdnd11an1n64x5 FILLER_252_200 ();
 b15zdnd11an1n64x5 FILLER_252_264 ();
 b15zdnd11an1n64x5 FILLER_252_328 ();
 b15zdnd11an1n16x5 FILLER_252_392 ();
 b15zdnd11an1n08x5 FILLER_252_408 ();
 b15zdnd11an1n64x5 FILLER_252_458 ();
 b15zdnd11an1n64x5 FILLER_252_522 ();
 b15zdnd11an1n64x5 FILLER_252_586 ();
 b15zdnd11an1n64x5 FILLER_252_650 ();
 b15zdnd11an1n04x5 FILLER_252_714 ();
 b15zdnd11an1n32x5 FILLER_252_726 ();
 b15zdnd11an1n16x5 FILLER_252_758 ();
 b15zdnd11an1n08x5 FILLER_252_774 ();
 b15zdnd11an1n04x5 FILLER_252_782 ();
 b15zdnd00an1n01x5 FILLER_252_786 ();
 b15zdnd11an1n08x5 FILLER_252_790 ();
 b15zdnd00an1n02x5 FILLER_252_798 ();
 b15zdnd00an1n01x5 FILLER_252_800 ();
 b15zdnd11an1n64x5 FILLER_252_853 ();
 b15zdnd11an1n08x5 FILLER_252_917 ();
 b15zdnd11an1n04x5 FILLER_252_925 ();
 b15zdnd11an1n04x5 FILLER_252_936 ();
 b15zdnd11an1n64x5 FILLER_252_979 ();
 b15zdnd00an1n01x5 FILLER_252_1043 ();
 b15zdnd11an1n64x5 FILLER_252_1058 ();
 b15zdnd11an1n64x5 FILLER_252_1122 ();
 b15zdnd11an1n64x5 FILLER_252_1186 ();
 b15zdnd11an1n08x5 FILLER_252_1250 ();
 b15zdnd11an1n04x5 FILLER_252_1258 ();
 b15zdnd11an1n64x5 FILLER_252_1314 ();
 b15zdnd11an1n32x5 FILLER_252_1378 ();
 b15zdnd11an1n08x5 FILLER_252_1410 ();
 b15zdnd11an1n04x5 FILLER_252_1418 ();
 b15zdnd11an1n64x5 FILLER_252_1425 ();
 b15zdnd11an1n64x5 FILLER_252_1489 ();
 b15zdnd11an1n16x5 FILLER_252_1553 ();
 b15zdnd11an1n08x5 FILLER_252_1569 ();
 b15zdnd11an1n04x5 FILLER_252_1577 ();
 b15zdnd00an1n02x5 FILLER_252_1581 ();
 b15zdnd11an1n64x5 FILLER_252_1589 ();
 b15zdnd11an1n64x5 FILLER_252_1653 ();
 b15zdnd11an1n64x5 FILLER_252_1717 ();
 b15zdnd11an1n64x5 FILLER_252_1781 ();
 b15zdnd11an1n64x5 FILLER_252_1845 ();
 b15zdnd11an1n64x5 FILLER_252_1909 ();
 b15zdnd11an1n64x5 FILLER_252_1973 ();
 b15zdnd11an1n64x5 FILLER_252_2037 ();
 b15zdnd11an1n32x5 FILLER_252_2101 ();
 b15zdnd11an1n16x5 FILLER_252_2133 ();
 b15zdnd11an1n04x5 FILLER_252_2149 ();
 b15zdnd00an1n01x5 FILLER_252_2153 ();
 b15zdnd11an1n64x5 FILLER_252_2162 ();
 b15zdnd11an1n32x5 FILLER_252_2226 ();
 b15zdnd11an1n16x5 FILLER_252_2258 ();
 b15zdnd00an1n02x5 FILLER_252_2274 ();
 b15zdnd11an1n64x5 FILLER_253_0 ();
 b15zdnd11an1n32x5 FILLER_253_64 ();
 b15zdnd11an1n16x5 FILLER_253_96 ();
 b15zdnd11an1n08x5 FILLER_253_112 ();
 b15zdnd00an1n02x5 FILLER_253_120 ();
 b15zdnd00an1n01x5 FILLER_253_122 ();
 b15zdnd11an1n16x5 FILLER_253_141 ();
 b15zdnd11an1n08x5 FILLER_253_157 ();
 b15zdnd00an1n02x5 FILLER_253_165 ();
 b15zdnd11an1n32x5 FILLER_253_178 ();
 b15zdnd11an1n08x5 FILLER_253_210 ();
 b15zdnd00an1n02x5 FILLER_253_218 ();
 b15zdnd11an1n64x5 FILLER_253_229 ();
 b15zdnd11an1n64x5 FILLER_253_293 ();
 b15zdnd11an1n32x5 FILLER_253_357 ();
 b15zdnd11an1n16x5 FILLER_253_389 ();
 b15zdnd11an1n08x5 FILLER_253_405 ();
 b15zdnd11an1n04x5 FILLER_253_413 ();
 b15zdnd00an1n02x5 FILLER_253_417 ();
 b15zdnd00an1n01x5 FILLER_253_419 ();
 b15zdnd11an1n64x5 FILLER_253_428 ();
 b15zdnd11an1n64x5 FILLER_253_492 ();
 b15zdnd11an1n08x5 FILLER_253_556 ();
 b15zdnd11an1n64x5 FILLER_253_606 ();
 b15zdnd11an1n64x5 FILLER_253_670 ();
 b15zdnd11an1n16x5 FILLER_253_734 ();
 b15zdnd11an1n08x5 FILLER_253_750 ();
 b15zdnd00an1n02x5 FILLER_253_758 ();
 b15zdnd11an1n08x5 FILLER_253_812 ();
 b15zdnd00an1n01x5 FILLER_253_820 ();
 b15zdnd11an1n04x5 FILLER_253_837 ();
 b15zdnd11an1n64x5 FILLER_253_844 ();
 b15zdnd00an1n02x5 FILLER_253_908 ();
 b15zdnd11an1n64x5 FILLER_253_916 ();
 b15zdnd11an1n64x5 FILLER_253_980 ();
 b15zdnd11an1n64x5 FILLER_253_1044 ();
 b15zdnd11an1n16x5 FILLER_253_1108 ();
 b15zdnd11an1n08x5 FILLER_253_1124 ();
 b15zdnd11an1n04x5 FILLER_253_1136 ();
 b15zdnd00an1n02x5 FILLER_253_1140 ();
 b15zdnd11an1n64x5 FILLER_253_1148 ();
 b15zdnd11an1n64x5 FILLER_253_1212 ();
 b15zdnd00an1n02x5 FILLER_253_1276 ();
 b15zdnd00an1n01x5 FILLER_253_1278 ();
 b15zdnd11an1n04x5 FILLER_253_1282 ();
 b15zdnd11an1n04x5 FILLER_253_1289 ();
 b15zdnd11an1n64x5 FILLER_253_1296 ();
 b15zdnd11an1n64x5 FILLER_253_1360 ();
 b15zdnd11an1n64x5 FILLER_253_1424 ();
 b15zdnd11an1n64x5 FILLER_253_1488 ();
 b15zdnd11an1n32x5 FILLER_253_1552 ();
 b15zdnd00an1n02x5 FILLER_253_1584 ();
 b15zdnd00an1n01x5 FILLER_253_1586 ();
 b15zdnd11an1n64x5 FILLER_253_1603 ();
 b15zdnd11an1n64x5 FILLER_253_1667 ();
 b15zdnd11an1n64x5 FILLER_253_1731 ();
 b15zdnd11an1n64x5 FILLER_253_1795 ();
 b15zdnd11an1n32x5 FILLER_253_1859 ();
 b15zdnd11an1n16x5 FILLER_253_1891 ();
 b15zdnd11an1n08x5 FILLER_253_1907 ();
 b15zdnd11an1n04x5 FILLER_253_1915 ();
 b15zdnd11an1n64x5 FILLER_253_1933 ();
 b15zdnd11an1n64x5 FILLER_253_1997 ();
 b15zdnd11an1n32x5 FILLER_253_2061 ();
 b15zdnd11an1n04x5 FILLER_253_2093 ();
 b15zdnd11an1n64x5 FILLER_253_2100 ();
 b15zdnd11an1n64x5 FILLER_253_2164 ();
 b15zdnd11an1n32x5 FILLER_253_2228 ();
 b15zdnd11an1n16x5 FILLER_253_2260 ();
 b15zdnd11an1n08x5 FILLER_253_2276 ();
 b15zdnd11an1n64x5 FILLER_254_8 ();
 b15zdnd11an1n64x5 FILLER_254_72 ();
 b15zdnd11an1n64x5 FILLER_254_136 ();
 b15zdnd11an1n16x5 FILLER_254_200 ();
 b15zdnd11an1n04x5 FILLER_254_216 ();
 b15zdnd00an1n02x5 FILLER_254_220 ();
 b15zdnd00an1n01x5 FILLER_254_222 ();
 b15zdnd11an1n64x5 FILLER_254_238 ();
 b15zdnd11an1n16x5 FILLER_254_302 ();
 b15zdnd11an1n08x5 FILLER_254_318 ();
 b15zdnd11an1n04x5 FILLER_254_326 ();
 b15zdnd00an1n02x5 FILLER_254_330 ();
 b15zdnd11an1n64x5 FILLER_254_356 ();
 b15zdnd11an1n64x5 FILLER_254_420 ();
 b15zdnd11an1n64x5 FILLER_254_484 ();
 b15zdnd11an1n64x5 FILLER_254_548 ();
 b15zdnd11an1n64x5 FILLER_254_612 ();
 b15zdnd11an1n32x5 FILLER_254_676 ();
 b15zdnd11an1n08x5 FILLER_254_708 ();
 b15zdnd00an1n02x5 FILLER_254_716 ();
 b15zdnd11an1n32x5 FILLER_254_726 ();
 b15zdnd11an1n16x5 FILLER_254_758 ();
 b15zdnd11an1n04x5 FILLER_254_777 ();
 b15zdnd11an1n04x5 FILLER_254_784 ();
 b15zdnd11an1n04x5 FILLER_254_795 ();
 b15zdnd11an1n04x5 FILLER_254_806 ();
 b15zdnd11an1n04x5 FILLER_254_852 ();
 b15zdnd11an1n64x5 FILLER_254_863 ();
 b15zdnd11an1n64x5 FILLER_254_927 ();
 b15zdnd11an1n64x5 FILLER_254_991 ();
 b15zdnd11an1n64x5 FILLER_254_1055 ();
 b15zdnd11an1n32x5 FILLER_254_1119 ();
 b15zdnd11an1n04x5 FILLER_254_1151 ();
 b15zdnd00an1n01x5 FILLER_254_1155 ();
 b15zdnd11an1n64x5 FILLER_254_1160 ();
 b15zdnd11an1n32x5 FILLER_254_1224 ();
 b15zdnd11an1n16x5 FILLER_254_1256 ();
 b15zdnd11an1n08x5 FILLER_254_1272 ();
 b15zdnd11an1n04x5 FILLER_254_1283 ();
 b15zdnd11an1n04x5 FILLER_254_1290 ();
 b15zdnd11an1n64x5 FILLER_254_1297 ();
 b15zdnd11an1n32x5 FILLER_254_1361 ();
 b15zdnd11an1n16x5 FILLER_254_1393 ();
 b15zdnd11an1n64x5 FILLER_254_1429 ();
 b15zdnd11an1n64x5 FILLER_254_1493 ();
 b15zdnd11an1n64x5 FILLER_254_1557 ();
 b15zdnd11an1n64x5 FILLER_254_1621 ();
 b15zdnd11an1n64x5 FILLER_254_1685 ();
 b15zdnd11an1n64x5 FILLER_254_1749 ();
 b15zdnd11an1n64x5 FILLER_254_1813 ();
 b15zdnd11an1n32x5 FILLER_254_1877 ();
 b15zdnd11an1n16x5 FILLER_254_1909 ();
 b15zdnd11an1n04x5 FILLER_254_1925 ();
 b15zdnd00an1n02x5 FILLER_254_1929 ();
 b15zdnd00an1n01x5 FILLER_254_1931 ();
 b15zdnd11an1n64x5 FILLER_254_1941 ();
 b15zdnd11an1n64x5 FILLER_254_2005 ();
 b15zdnd11an1n16x5 FILLER_254_2069 ();
 b15zdnd11an1n08x5 FILLER_254_2085 ();
 b15zdnd11an1n04x5 FILLER_254_2093 ();
 b15zdnd11an1n32x5 FILLER_254_2100 ();
 b15zdnd11an1n16x5 FILLER_254_2132 ();
 b15zdnd11an1n04x5 FILLER_254_2148 ();
 b15zdnd00an1n02x5 FILLER_254_2152 ();
 b15zdnd11an1n64x5 FILLER_254_2162 ();
 b15zdnd11an1n32x5 FILLER_254_2226 ();
 b15zdnd11an1n16x5 FILLER_254_2258 ();
 b15zdnd00an1n02x5 FILLER_254_2274 ();
 b15zdnd11an1n64x5 FILLER_255_0 ();
 b15zdnd11an1n64x5 FILLER_255_64 ();
 b15zdnd11an1n64x5 FILLER_255_128 ();
 b15zdnd11an1n64x5 FILLER_255_192 ();
 b15zdnd11an1n64x5 FILLER_255_256 ();
 b15zdnd11an1n32x5 FILLER_255_320 ();
 b15zdnd11an1n08x5 FILLER_255_352 ();
 b15zdnd00an1n02x5 FILLER_255_360 ();
 b15zdnd11an1n64x5 FILLER_255_372 ();
 b15zdnd11an1n64x5 FILLER_255_436 ();
 b15zdnd11an1n64x5 FILLER_255_500 ();
 b15zdnd11an1n64x5 FILLER_255_564 ();
 b15zdnd11an1n64x5 FILLER_255_628 ();
 b15zdnd11an1n64x5 FILLER_255_692 ();
 b15zdnd11an1n32x5 FILLER_255_756 ();
 b15zdnd11an1n08x5 FILLER_255_788 ();
 b15zdnd11an1n04x5 FILLER_255_796 ();
 b15zdnd00an1n02x5 FILLER_255_800 ();
 b15zdnd11an1n64x5 FILLER_255_844 ();
 b15zdnd11an1n64x5 FILLER_255_908 ();
 b15zdnd11an1n64x5 FILLER_255_972 ();
 b15zdnd11an1n64x5 FILLER_255_1036 ();
 b15zdnd11an1n32x5 FILLER_255_1100 ();
 b15zdnd11an1n16x5 FILLER_255_1132 ();
 b15zdnd11an1n16x5 FILLER_255_1152 ();
 b15zdnd11an1n04x5 FILLER_255_1168 ();
 b15zdnd00an1n02x5 FILLER_255_1172 ();
 b15zdnd00an1n01x5 FILLER_255_1174 ();
 b15zdnd11an1n64x5 FILLER_255_1179 ();
 b15zdnd11an1n64x5 FILLER_255_1243 ();
 b15zdnd11an1n64x5 FILLER_255_1307 ();
 b15zdnd11an1n64x5 FILLER_255_1371 ();
 b15zdnd11an1n64x5 FILLER_255_1435 ();
 b15zdnd11an1n64x5 FILLER_255_1499 ();
 b15zdnd11an1n64x5 FILLER_255_1563 ();
 b15zdnd11an1n64x5 FILLER_255_1627 ();
 b15zdnd11an1n08x5 FILLER_255_1691 ();
 b15zdnd00an1n02x5 FILLER_255_1699 ();
 b15zdnd00an1n01x5 FILLER_255_1701 ();
 b15zdnd11an1n64x5 FILLER_255_1718 ();
 b15zdnd11an1n32x5 FILLER_255_1782 ();
 b15zdnd11an1n16x5 FILLER_255_1814 ();
 b15zdnd11an1n04x5 FILLER_255_1830 ();
 b15zdnd00an1n02x5 FILLER_255_1834 ();
 b15zdnd11an1n64x5 FILLER_255_1846 ();
 b15zdnd11an1n64x5 FILLER_255_1910 ();
 b15zdnd11an1n64x5 FILLER_255_1974 ();
 b15zdnd11an1n32x5 FILLER_255_2038 ();
 b15zdnd00an1n02x5 FILLER_255_2070 ();
 b15zdnd11an1n64x5 FILLER_255_2124 ();
 b15zdnd11an1n64x5 FILLER_255_2188 ();
 b15zdnd11an1n32x5 FILLER_255_2252 ();
 b15zdnd11an1n16x5 FILLER_256_8 ();
 b15zdnd11an1n04x5 FILLER_256_24 ();
 b15zdnd00an1n02x5 FILLER_256_28 ();
 b15zdnd11an1n32x5 FILLER_256_37 ();
 b15zdnd11an1n16x5 FILLER_256_69 ();
 b15zdnd11an1n08x5 FILLER_256_85 ();
 b15zdnd11an1n64x5 FILLER_256_133 ();
 b15zdnd11an1n64x5 FILLER_256_197 ();
 b15zdnd11an1n64x5 FILLER_256_261 ();
 b15zdnd11an1n32x5 FILLER_256_325 ();
 b15zdnd11an1n08x5 FILLER_256_357 ();
 b15zdnd11an1n04x5 FILLER_256_365 ();
 b15zdnd11an1n64x5 FILLER_256_375 ();
 b15zdnd11an1n64x5 FILLER_256_439 ();
 b15zdnd11an1n64x5 FILLER_256_503 ();
 b15zdnd11an1n64x5 FILLER_256_567 ();
 b15zdnd11an1n64x5 FILLER_256_631 ();
 b15zdnd11an1n16x5 FILLER_256_695 ();
 b15zdnd11an1n04x5 FILLER_256_711 ();
 b15zdnd00an1n02x5 FILLER_256_715 ();
 b15zdnd00an1n01x5 FILLER_256_717 ();
 b15zdnd11an1n64x5 FILLER_256_726 ();
 b15zdnd11an1n08x5 FILLER_256_790 ();
 b15zdnd11an1n64x5 FILLER_256_840 ();
 b15zdnd11an1n32x5 FILLER_256_904 ();
 b15zdnd11an1n08x5 FILLER_256_936 ();
 b15zdnd11an1n04x5 FILLER_256_944 ();
 b15zdnd00an1n02x5 FILLER_256_948 ();
 b15zdnd00an1n01x5 FILLER_256_950 ();
 b15zdnd11an1n16x5 FILLER_256_957 ();
 b15zdnd11an1n08x5 FILLER_256_973 ();
 b15zdnd11an1n04x5 FILLER_256_981 ();
 b15zdnd00an1n02x5 FILLER_256_985 ();
 b15zdnd00an1n01x5 FILLER_256_987 ();
 b15zdnd11an1n64x5 FILLER_256_1030 ();
 b15zdnd11an1n32x5 FILLER_256_1094 ();
 b15zdnd11an1n16x5 FILLER_256_1126 ();
 b15zdnd11an1n08x5 FILLER_256_1142 ();
 b15zdnd11an1n04x5 FILLER_256_1150 ();
 b15zdnd00an1n02x5 FILLER_256_1154 ();
 b15zdnd11an1n04x5 FILLER_256_1162 ();
 b15zdnd00an1n01x5 FILLER_256_1166 ();
 b15zdnd11an1n04x5 FILLER_256_1175 ();
 b15zdnd11an1n64x5 FILLER_256_1183 ();
 b15zdnd11an1n64x5 FILLER_256_1247 ();
 b15zdnd11an1n64x5 FILLER_256_1311 ();
 b15zdnd11an1n64x5 FILLER_256_1375 ();
 b15zdnd00an1n02x5 FILLER_256_1439 ();
 b15zdnd00an1n01x5 FILLER_256_1441 ();
 b15zdnd11an1n64x5 FILLER_256_1458 ();
 b15zdnd11an1n64x5 FILLER_256_1522 ();
 b15zdnd11an1n64x5 FILLER_256_1586 ();
 b15zdnd11an1n64x5 FILLER_256_1650 ();
 b15zdnd11an1n64x5 FILLER_256_1714 ();
 b15zdnd11an1n64x5 FILLER_256_1778 ();
 b15zdnd11an1n64x5 FILLER_256_1842 ();
 b15zdnd11an1n64x5 FILLER_256_1906 ();
 b15zdnd11an1n64x5 FILLER_256_1970 ();
 b15zdnd11an1n32x5 FILLER_256_2034 ();
 b15zdnd11an1n16x5 FILLER_256_2066 ();
 b15zdnd11an1n08x5 FILLER_256_2082 ();
 b15zdnd11an1n04x5 FILLER_256_2090 ();
 b15zdnd00an1n02x5 FILLER_256_2094 ();
 b15zdnd00an1n01x5 FILLER_256_2096 ();
 b15zdnd11an1n32x5 FILLER_256_2100 ();
 b15zdnd11an1n16x5 FILLER_256_2132 ();
 b15zdnd11an1n04x5 FILLER_256_2148 ();
 b15zdnd00an1n02x5 FILLER_256_2152 ();
 b15zdnd11an1n64x5 FILLER_256_2162 ();
 b15zdnd11an1n32x5 FILLER_256_2226 ();
 b15zdnd11an1n16x5 FILLER_256_2258 ();
 b15zdnd00an1n02x5 FILLER_256_2274 ();
 b15zdnd11an1n16x5 FILLER_257_0 ();
 b15zdnd11an1n08x5 FILLER_257_16 ();
 b15zdnd11an1n04x5 FILLER_257_24 ();
 b15zdnd00an1n02x5 FILLER_257_28 ();
 b15zdnd11an1n08x5 FILLER_257_34 ();
 b15zdnd11an1n04x5 FILLER_257_42 ();
 b15zdnd00an1n01x5 FILLER_257_46 ();
 b15zdnd11an1n64x5 FILLER_257_51 ();
 b15zdnd11an1n64x5 FILLER_257_115 ();
 b15zdnd11an1n64x5 FILLER_257_179 ();
 b15zdnd11an1n64x5 FILLER_257_243 ();
 b15zdnd11an1n64x5 FILLER_257_307 ();
 b15zdnd11an1n64x5 FILLER_257_371 ();
 b15zdnd11an1n64x5 FILLER_257_435 ();
 b15zdnd11an1n64x5 FILLER_257_499 ();
 b15zdnd11an1n64x5 FILLER_257_563 ();
 b15zdnd11an1n16x5 FILLER_257_627 ();
 b15zdnd11an1n08x5 FILLER_257_643 ();
 b15zdnd00an1n01x5 FILLER_257_651 ();
 b15zdnd11an1n08x5 FILLER_257_684 ();
 b15zdnd00an1n02x5 FILLER_257_692 ();
 b15zdnd11an1n64x5 FILLER_257_717 ();
 b15zdnd11an1n64x5 FILLER_257_781 ();
 b15zdnd11an1n04x5 FILLER_257_845 ();
 b15zdnd00an1n01x5 FILLER_257_849 ();
 b15zdnd11an1n08x5 FILLER_257_853 ();
 b15zdnd11an1n04x5 FILLER_257_861 ();
 b15zdnd11an1n64x5 FILLER_257_868 ();
 b15zdnd11an1n16x5 FILLER_257_932 ();
 b15zdnd11an1n04x5 FILLER_257_948 ();
 b15zdnd00an1n02x5 FILLER_257_952 ();
 b15zdnd11an1n64x5 FILLER_257_958 ();
 b15zdnd11an1n64x5 FILLER_257_1022 ();
 b15zdnd11an1n08x5 FILLER_257_1086 ();
 b15zdnd11an1n04x5 FILLER_257_1094 ();
 b15zdnd00an1n02x5 FILLER_257_1098 ();
 b15zdnd00an1n01x5 FILLER_257_1100 ();
 b15zdnd11an1n64x5 FILLER_257_1108 ();
 b15zdnd11an1n64x5 FILLER_257_1172 ();
 b15zdnd11an1n64x5 FILLER_257_1236 ();
 b15zdnd11an1n64x5 FILLER_257_1300 ();
 b15zdnd11an1n64x5 FILLER_257_1364 ();
 b15zdnd11an1n64x5 FILLER_257_1428 ();
 b15zdnd11an1n64x5 FILLER_257_1492 ();
 b15zdnd11an1n32x5 FILLER_257_1556 ();
 b15zdnd11an1n04x5 FILLER_257_1588 ();
 b15zdnd00an1n02x5 FILLER_257_1592 ();
 b15zdnd00an1n01x5 FILLER_257_1594 ();
 b15zdnd11an1n08x5 FILLER_257_1605 ();
 b15zdnd11an1n64x5 FILLER_257_1616 ();
 b15zdnd11an1n64x5 FILLER_257_1680 ();
 b15zdnd11an1n64x5 FILLER_257_1744 ();
 b15zdnd11an1n64x5 FILLER_257_1808 ();
 b15zdnd11an1n64x5 FILLER_257_1872 ();
 b15zdnd11an1n64x5 FILLER_257_1936 ();
 b15zdnd11an1n64x5 FILLER_257_2000 ();
 b15zdnd11an1n64x5 FILLER_257_2064 ();
 b15zdnd11an1n64x5 FILLER_257_2128 ();
 b15zdnd11an1n08x5 FILLER_257_2192 ();
 b15zdnd11an1n64x5 FILLER_257_2203 ();
 b15zdnd11an1n16x5 FILLER_257_2267 ();
 b15zdnd00an1n01x5 FILLER_257_2283 ();
 b15zdnd11an1n08x5 FILLER_258_8 ();
 b15zdnd00an1n02x5 FILLER_258_16 ();
 b15zdnd11an1n64x5 FILLER_258_38 ();
 b15zdnd11an1n64x5 FILLER_258_102 ();
 b15zdnd11an1n64x5 FILLER_258_166 ();
 b15zdnd11an1n64x5 FILLER_258_230 ();
 b15zdnd11an1n64x5 FILLER_258_294 ();
 b15zdnd11an1n64x5 FILLER_258_358 ();
 b15zdnd11an1n64x5 FILLER_258_422 ();
 b15zdnd11an1n64x5 FILLER_258_486 ();
 b15zdnd11an1n64x5 FILLER_258_550 ();
 b15zdnd11an1n64x5 FILLER_258_614 ();
 b15zdnd11an1n32x5 FILLER_258_678 ();
 b15zdnd11an1n08x5 FILLER_258_710 ();
 b15zdnd11an1n64x5 FILLER_258_726 ();
 b15zdnd11an1n32x5 FILLER_258_790 ();
 b15zdnd11an1n16x5 FILLER_258_822 ();
 b15zdnd00an1n02x5 FILLER_258_838 ();
 b15zdnd11an1n32x5 FILLER_258_884 ();
 b15zdnd11an1n08x5 FILLER_258_916 ();
 b15zdnd00an1n01x5 FILLER_258_924 ();
 b15zdnd11an1n64x5 FILLER_258_931 ();
 b15zdnd11an1n64x5 FILLER_258_995 ();
 b15zdnd11an1n32x5 FILLER_258_1059 ();
 b15zdnd11an1n16x5 FILLER_258_1091 ();
 b15zdnd11an1n08x5 FILLER_258_1107 ();
 b15zdnd11an1n16x5 FILLER_258_1160 ();
 b15zdnd11an1n08x5 FILLER_258_1176 ();
 b15zdnd00an1n02x5 FILLER_258_1184 ();
 b15zdnd11an1n64x5 FILLER_258_1190 ();
 b15zdnd11an1n64x5 FILLER_258_1254 ();
 b15zdnd11an1n64x5 FILLER_258_1318 ();
 b15zdnd11an1n64x5 FILLER_258_1382 ();
 b15zdnd11an1n64x5 FILLER_258_1446 ();
 b15zdnd11an1n64x5 FILLER_258_1510 ();
 b15zdnd11an1n32x5 FILLER_258_1574 ();
 b15zdnd11an1n08x5 FILLER_258_1606 ();
 b15zdnd00an1n01x5 FILLER_258_1614 ();
 b15zdnd11an1n08x5 FILLER_258_1626 ();
 b15zdnd00an1n02x5 FILLER_258_1634 ();
 b15zdnd11an1n04x5 FILLER_258_1639 ();
 b15zdnd11an1n04x5 FILLER_258_1656 ();
 b15zdnd11an1n64x5 FILLER_258_1681 ();
 b15zdnd11an1n64x5 FILLER_258_1745 ();
 b15zdnd11an1n64x5 FILLER_258_1809 ();
 b15zdnd11an1n64x5 FILLER_258_1873 ();
 b15zdnd11an1n64x5 FILLER_258_1937 ();
 b15zdnd11an1n64x5 FILLER_258_2001 ();
 b15zdnd11an1n64x5 FILLER_258_2065 ();
 b15zdnd11an1n16x5 FILLER_258_2129 ();
 b15zdnd11an1n08x5 FILLER_258_2145 ();
 b15zdnd00an1n01x5 FILLER_258_2153 ();
 b15zdnd00an1n02x5 FILLER_258_2162 ();
 b15zdnd11an1n04x5 FILLER_258_2206 ();
 b15zdnd11an1n32x5 FILLER_258_2213 ();
 b15zdnd11an1n16x5 FILLER_258_2245 ();
 b15zdnd11an1n08x5 FILLER_258_2261 ();
 b15zdnd11an1n04x5 FILLER_258_2269 ();
 b15zdnd00an1n02x5 FILLER_258_2273 ();
 b15zdnd00an1n01x5 FILLER_258_2275 ();
 b15zdnd11an1n08x5 FILLER_259_0 ();
 b15zdnd00an1n02x5 FILLER_259_8 ();
 b15zdnd11an1n16x5 FILLER_259_16 ();
 b15zdnd11an1n04x5 FILLER_259_32 ();
 b15zdnd00an1n01x5 FILLER_259_36 ();
 b15zdnd11an1n04x5 FILLER_259_68 ();
 b15zdnd00an1n01x5 FILLER_259_72 ();
 b15zdnd11an1n64x5 FILLER_259_104 ();
 b15zdnd11an1n64x5 FILLER_259_168 ();
 b15zdnd11an1n64x5 FILLER_259_232 ();
 b15zdnd11an1n64x5 FILLER_259_296 ();
 b15zdnd11an1n64x5 FILLER_259_360 ();
 b15zdnd11an1n64x5 FILLER_259_424 ();
 b15zdnd11an1n64x5 FILLER_259_488 ();
 b15zdnd11an1n64x5 FILLER_259_552 ();
 b15zdnd11an1n64x5 FILLER_259_616 ();
 b15zdnd11an1n64x5 FILLER_259_680 ();
 b15zdnd11an1n32x5 FILLER_259_744 ();
 b15zdnd11an1n08x5 FILLER_259_776 ();
 b15zdnd11an1n04x5 FILLER_259_784 ();
 b15zdnd11an1n64x5 FILLER_259_796 ();
 b15zdnd00an1n01x5 FILLER_259_860 ();
 b15zdnd11an1n16x5 FILLER_259_864 ();
 b15zdnd11an1n04x5 FILLER_259_880 ();
 b15zdnd00an1n02x5 FILLER_259_884 ();
 b15zdnd00an1n01x5 FILLER_259_886 ();
 b15zdnd11an1n64x5 FILLER_259_898 ();
 b15zdnd11an1n32x5 FILLER_259_962 ();
 b15zdnd11an1n16x5 FILLER_259_994 ();
 b15zdnd00an1n02x5 FILLER_259_1010 ();
 b15zdnd11an1n64x5 FILLER_259_1026 ();
 b15zdnd11an1n32x5 FILLER_259_1090 ();
 b15zdnd11an1n08x5 FILLER_259_1122 ();
 b15zdnd11an1n64x5 FILLER_259_1136 ();
 b15zdnd11an1n64x5 FILLER_259_1200 ();
 b15zdnd11an1n64x5 FILLER_259_1264 ();
 b15zdnd11an1n64x5 FILLER_259_1328 ();
 b15zdnd11an1n64x5 FILLER_259_1392 ();
 b15zdnd11an1n64x5 FILLER_259_1456 ();
 b15zdnd11an1n64x5 FILLER_259_1520 ();
 b15zdnd11an1n64x5 FILLER_259_1584 ();
 b15zdnd11an1n64x5 FILLER_259_1648 ();
 b15zdnd11an1n08x5 FILLER_259_1712 ();
 b15zdnd11an1n32x5 FILLER_259_1734 ();
 b15zdnd00an1n02x5 FILLER_259_1766 ();
 b15zdnd00an1n01x5 FILLER_259_1768 ();
 b15zdnd11an1n04x5 FILLER_259_1783 ();
 b15zdnd00an1n01x5 FILLER_259_1787 ();
 b15zdnd11an1n64x5 FILLER_259_1791 ();
 b15zdnd11an1n64x5 FILLER_259_1855 ();
 b15zdnd11an1n32x5 FILLER_259_1919 ();
 b15zdnd00an1n02x5 FILLER_259_1951 ();
 b15zdnd11an1n64x5 FILLER_259_1995 ();
 b15zdnd11an1n64x5 FILLER_259_2059 ();
 b15zdnd11an1n32x5 FILLER_259_2123 ();
 b15zdnd11an1n16x5 FILLER_259_2155 ();
 b15zdnd11an1n08x5 FILLER_259_2171 ();
 b15zdnd00an1n02x5 FILLER_259_2179 ();
 b15zdnd00an1n01x5 FILLER_259_2181 ();
 b15zdnd11an1n32x5 FILLER_259_2234 ();
 b15zdnd11an1n16x5 FILLER_259_2266 ();
 b15zdnd00an1n02x5 FILLER_259_2282 ();
 b15zdnd11an1n32x5 FILLER_260_8 ();
 b15zdnd11an1n16x5 FILLER_260_40 ();
 b15zdnd11an1n04x5 FILLER_260_56 ();
 b15zdnd11an1n64x5 FILLER_260_85 ();
 b15zdnd11an1n64x5 FILLER_260_149 ();
 b15zdnd11an1n64x5 FILLER_260_213 ();
 b15zdnd11an1n64x5 FILLER_260_277 ();
 b15zdnd11an1n64x5 FILLER_260_341 ();
 b15zdnd11an1n64x5 FILLER_260_405 ();
 b15zdnd11an1n64x5 FILLER_260_469 ();
 b15zdnd11an1n64x5 FILLER_260_533 ();
 b15zdnd11an1n64x5 FILLER_260_597 ();
 b15zdnd11an1n32x5 FILLER_260_661 ();
 b15zdnd11an1n16x5 FILLER_260_693 ();
 b15zdnd11an1n08x5 FILLER_260_709 ();
 b15zdnd00an1n01x5 FILLER_260_717 ();
 b15zdnd11an1n64x5 FILLER_260_726 ();
 b15zdnd11an1n64x5 FILLER_260_790 ();
 b15zdnd11an1n64x5 FILLER_260_854 ();
 b15zdnd11an1n64x5 FILLER_260_918 ();
 b15zdnd11an1n64x5 FILLER_260_982 ();
 b15zdnd11an1n64x5 FILLER_260_1046 ();
 b15zdnd11an1n64x5 FILLER_260_1110 ();
 b15zdnd11an1n64x5 FILLER_260_1174 ();
 b15zdnd11an1n64x5 FILLER_260_1238 ();
 b15zdnd11an1n64x5 FILLER_260_1302 ();
 b15zdnd11an1n64x5 FILLER_260_1366 ();
 b15zdnd11an1n64x5 FILLER_260_1430 ();
 b15zdnd11an1n32x5 FILLER_260_1494 ();
 b15zdnd11an1n08x5 FILLER_260_1526 ();
 b15zdnd00an1n01x5 FILLER_260_1534 ();
 b15zdnd11an1n64x5 FILLER_260_1549 ();
 b15zdnd11an1n64x5 FILLER_260_1613 ();
 b15zdnd11an1n64x5 FILLER_260_1677 ();
 b15zdnd11an1n32x5 FILLER_260_1741 ();
 b15zdnd11an1n08x5 FILLER_260_1773 ();
 b15zdnd11an1n64x5 FILLER_260_1784 ();
 b15zdnd11an1n64x5 FILLER_260_1848 ();
 b15zdnd11an1n32x5 FILLER_260_1912 ();
 b15zdnd00an1n01x5 FILLER_260_1944 ();
 b15zdnd11an1n04x5 FILLER_260_1948 ();
 b15zdnd11an1n64x5 FILLER_260_1955 ();
 b15zdnd11an1n64x5 FILLER_260_2019 ();
 b15zdnd11an1n64x5 FILLER_260_2083 ();
 b15zdnd11an1n04x5 FILLER_260_2147 ();
 b15zdnd00an1n02x5 FILLER_260_2151 ();
 b15zdnd00an1n01x5 FILLER_260_2153 ();
 b15zdnd11an1n32x5 FILLER_260_2162 ();
 b15zdnd11an1n08x5 FILLER_260_2194 ();
 b15zdnd11an1n04x5 FILLER_260_2202 ();
 b15zdnd00an1n01x5 FILLER_260_2206 ();
 b15zdnd11an1n64x5 FILLER_260_2210 ();
 b15zdnd00an1n02x5 FILLER_260_2274 ();
 b15zdnd00an1n02x5 FILLER_261_0 ();
 b15zdnd11an1n64x5 FILLER_261_7 ();
 b15zdnd11an1n64x5 FILLER_261_71 ();
 b15zdnd11an1n64x5 FILLER_261_135 ();
 b15zdnd11an1n32x5 FILLER_261_199 ();
 b15zdnd00an1n02x5 FILLER_261_231 ();
 b15zdnd00an1n01x5 FILLER_261_233 ();
 b15zdnd11an1n64x5 FILLER_261_248 ();
 b15zdnd11an1n64x5 FILLER_261_312 ();
 b15zdnd11an1n64x5 FILLER_261_376 ();
 b15zdnd11an1n64x5 FILLER_261_440 ();
 b15zdnd11an1n64x5 FILLER_261_504 ();
 b15zdnd11an1n64x5 FILLER_261_568 ();
 b15zdnd11an1n64x5 FILLER_261_632 ();
 b15zdnd11an1n64x5 FILLER_261_696 ();
 b15zdnd11an1n16x5 FILLER_261_760 ();
 b15zdnd11an1n08x5 FILLER_261_776 ();
 b15zdnd11an1n04x5 FILLER_261_784 ();
 b15zdnd00an1n02x5 FILLER_261_788 ();
 b15zdnd00an1n01x5 FILLER_261_790 ();
 b15zdnd11an1n64x5 FILLER_261_799 ();
 b15zdnd11an1n64x5 FILLER_261_863 ();
 b15zdnd11an1n64x5 FILLER_261_927 ();
 b15zdnd11an1n64x5 FILLER_261_991 ();
 b15zdnd11an1n32x5 FILLER_261_1055 ();
 b15zdnd11an1n08x5 FILLER_261_1087 ();
 b15zdnd00an1n02x5 FILLER_261_1095 ();
 b15zdnd11an1n64x5 FILLER_261_1128 ();
 b15zdnd11an1n04x5 FILLER_261_1192 ();
 b15zdnd00an1n02x5 FILLER_261_1196 ();
 b15zdnd00an1n01x5 FILLER_261_1198 ();
 b15zdnd11an1n64x5 FILLER_261_1203 ();
 b15zdnd11an1n64x5 FILLER_261_1267 ();
 b15zdnd11an1n64x5 FILLER_261_1331 ();
 b15zdnd11an1n64x5 FILLER_261_1395 ();
 b15zdnd11an1n64x5 FILLER_261_1459 ();
 b15zdnd11an1n64x5 FILLER_261_1523 ();
 b15zdnd11an1n08x5 FILLER_261_1587 ();
 b15zdnd00an1n01x5 FILLER_261_1595 ();
 b15zdnd11an1n64x5 FILLER_261_1616 ();
 b15zdnd11an1n64x5 FILLER_261_1680 ();
 b15zdnd11an1n32x5 FILLER_261_1744 ();
 b15zdnd00an1n02x5 FILLER_261_1776 ();
 b15zdnd11an1n32x5 FILLER_261_1792 ();
 b15zdnd11an1n04x5 FILLER_261_1824 ();
 b15zdnd00an1n02x5 FILLER_261_1828 ();
 b15zdnd00an1n01x5 FILLER_261_1830 ();
 b15zdnd11an1n64x5 FILLER_261_1845 ();
 b15zdnd11an1n16x5 FILLER_261_1909 ();
 b15zdnd11an1n08x5 FILLER_261_1925 ();
 b15zdnd00an1n02x5 FILLER_261_1933 ();
 b15zdnd11an1n04x5 FILLER_261_1938 ();
 b15zdnd11an1n32x5 FILLER_261_1994 ();
 b15zdnd11an1n16x5 FILLER_261_2026 ();
 b15zdnd11an1n08x5 FILLER_261_2042 ();
 b15zdnd11an1n64x5 FILLER_261_2054 ();
 b15zdnd11an1n64x5 FILLER_261_2118 ();
 b15zdnd11an1n64x5 FILLER_261_2182 ();
 b15zdnd11an1n32x5 FILLER_261_2246 ();
 b15zdnd11an1n04x5 FILLER_261_2278 ();
 b15zdnd00an1n02x5 FILLER_261_2282 ();
 b15zdnd11an1n16x5 FILLER_262_8 ();
 b15zdnd00an1n02x5 FILLER_262_24 ();
 b15zdnd00an1n01x5 FILLER_262_26 ();
 b15zdnd11an1n32x5 FILLER_262_32 ();
 b15zdnd11an1n04x5 FILLER_262_64 ();
 b15zdnd00an1n02x5 FILLER_262_68 ();
 b15zdnd00an1n01x5 FILLER_262_70 ();
 b15zdnd11an1n64x5 FILLER_262_91 ();
 b15zdnd11an1n32x5 FILLER_262_155 ();
 b15zdnd11an1n08x5 FILLER_262_187 ();
 b15zdnd00an1n01x5 FILLER_262_195 ();
 b15zdnd11an1n08x5 FILLER_262_238 ();
 b15zdnd11an1n04x5 FILLER_262_246 ();
 b15zdnd00an1n02x5 FILLER_262_250 ();
 b15zdnd11an1n04x5 FILLER_262_270 ();
 b15zdnd00an1n02x5 FILLER_262_274 ();
 b15zdnd00an1n01x5 FILLER_262_276 ();
 b15zdnd11an1n04x5 FILLER_262_295 ();
 b15zdnd11an1n04x5 FILLER_262_313 ();
 b15zdnd11an1n64x5 FILLER_262_321 ();
 b15zdnd11an1n64x5 FILLER_262_385 ();
 b15zdnd11an1n64x5 FILLER_262_449 ();
 b15zdnd11an1n64x5 FILLER_262_513 ();
 b15zdnd00an1n01x5 FILLER_262_577 ();
 b15zdnd11an1n64x5 FILLER_262_581 ();
 b15zdnd11an1n64x5 FILLER_262_645 ();
 b15zdnd11an1n08x5 FILLER_262_709 ();
 b15zdnd00an1n01x5 FILLER_262_717 ();
 b15zdnd11an1n64x5 FILLER_262_726 ();
 b15zdnd11an1n64x5 FILLER_262_790 ();
 b15zdnd11an1n64x5 FILLER_262_854 ();
 b15zdnd11an1n64x5 FILLER_262_918 ();
 b15zdnd11an1n64x5 FILLER_262_982 ();
 b15zdnd11an1n64x5 FILLER_262_1046 ();
 b15zdnd11an1n64x5 FILLER_262_1110 ();
 b15zdnd11an1n64x5 FILLER_262_1174 ();
 b15zdnd11an1n64x5 FILLER_262_1238 ();
 b15zdnd11an1n64x5 FILLER_262_1302 ();
 b15zdnd11an1n64x5 FILLER_262_1366 ();
 b15zdnd11an1n16x5 FILLER_262_1430 ();
 b15zdnd11an1n64x5 FILLER_262_1450 ();
 b15zdnd11an1n64x5 FILLER_262_1514 ();
 b15zdnd11an1n64x5 FILLER_262_1578 ();
 b15zdnd11an1n04x5 FILLER_262_1642 ();
 b15zdnd11an1n16x5 FILLER_262_1653 ();
 b15zdnd11an1n08x5 FILLER_262_1669 ();
 b15zdnd11an1n64x5 FILLER_262_1697 ();
 b15zdnd00an1n02x5 FILLER_262_1761 ();
 b15zdnd00an1n01x5 FILLER_262_1763 ();
 b15zdnd11an1n04x5 FILLER_262_1778 ();
 b15zdnd11an1n64x5 FILLER_262_1799 ();
 b15zdnd11an1n04x5 FILLER_262_1863 ();
 b15zdnd11an1n32x5 FILLER_262_1873 ();
 b15zdnd11an1n16x5 FILLER_262_1905 ();
 b15zdnd11an1n04x5 FILLER_262_1973 ();
 b15zdnd11an1n64x5 FILLER_262_2019 ();
 b15zdnd11an1n64x5 FILLER_262_2083 ();
 b15zdnd11an1n04x5 FILLER_262_2147 ();
 b15zdnd00an1n02x5 FILLER_262_2151 ();
 b15zdnd00an1n01x5 FILLER_262_2153 ();
 b15zdnd11an1n64x5 FILLER_262_2162 ();
 b15zdnd11an1n08x5 FILLER_262_2226 ();
 b15zdnd00an1n02x5 FILLER_262_2234 ();
 b15zdnd11an1n08x5 FILLER_262_2267 ();
 b15zdnd00an1n01x5 FILLER_262_2275 ();
 b15zdnd11an1n16x5 FILLER_263_0 ();
 b15zdnd11an1n04x5 FILLER_263_16 ();
 b15zdnd11an1n16x5 FILLER_263_26 ();
 b15zdnd11an1n08x5 FILLER_263_42 ();
 b15zdnd00an1n02x5 FILLER_263_50 ();
 b15zdnd11an1n08x5 FILLER_263_58 ();
 b15zdnd00an1n02x5 FILLER_263_66 ();
 b15zdnd11an1n32x5 FILLER_263_89 ();
 b15zdnd11an1n16x5 FILLER_263_121 ();
 b15zdnd11an1n08x5 FILLER_263_137 ();
 b15zdnd11an1n32x5 FILLER_263_176 ();
 b15zdnd11an1n16x5 FILLER_263_208 ();
 b15zdnd11an1n08x5 FILLER_263_224 ();
 b15zdnd00an1n02x5 FILLER_263_232 ();
 b15zdnd11an1n08x5 FILLER_263_276 ();
 b15zdnd11an1n04x5 FILLER_263_284 ();
 b15zdnd00an1n02x5 FILLER_263_288 ();
 b15zdnd11an1n04x5 FILLER_263_294 ();
 b15zdnd11an1n64x5 FILLER_263_318 ();
 b15zdnd11an1n64x5 FILLER_263_382 ();
 b15zdnd11an1n64x5 FILLER_263_446 ();
 b15zdnd11an1n32x5 FILLER_263_510 ();
 b15zdnd11an1n04x5 FILLER_263_542 ();
 b15zdnd00an1n02x5 FILLER_263_546 ();
 b15zdnd11an1n04x5 FILLER_263_588 ();
 b15zdnd11an1n64x5 FILLER_263_595 ();
 b15zdnd11an1n64x5 FILLER_263_659 ();
 b15zdnd11an1n64x5 FILLER_263_723 ();
 b15zdnd11an1n64x5 FILLER_263_787 ();
 b15zdnd11an1n64x5 FILLER_263_851 ();
 b15zdnd11an1n32x5 FILLER_263_915 ();
 b15zdnd11an1n16x5 FILLER_263_947 ();
 b15zdnd11an1n08x5 FILLER_263_963 ();
 b15zdnd00an1n02x5 FILLER_263_971 ();
 b15zdnd00an1n01x5 FILLER_263_973 ();
 b15zdnd11an1n64x5 FILLER_263_978 ();
 b15zdnd11an1n32x5 FILLER_263_1042 ();
 b15zdnd11an1n04x5 FILLER_263_1074 ();
 b15zdnd00an1n02x5 FILLER_263_1078 ();
 b15zdnd00an1n01x5 FILLER_263_1080 ();
 b15zdnd11an1n04x5 FILLER_263_1088 ();
 b15zdnd11an1n64x5 FILLER_263_1101 ();
 b15zdnd11an1n32x5 FILLER_263_1165 ();
 b15zdnd00an1n02x5 FILLER_263_1197 ();
 b15zdnd00an1n01x5 FILLER_263_1199 ();
 b15zdnd11an1n64x5 FILLER_263_1214 ();
 b15zdnd11an1n64x5 FILLER_263_1278 ();
 b15zdnd11an1n64x5 FILLER_263_1342 ();
 b15zdnd11an1n16x5 FILLER_263_1406 ();
 b15zdnd11an1n08x5 FILLER_263_1422 ();
 b15zdnd00an1n02x5 FILLER_263_1430 ();
 b15zdnd11an1n64x5 FILLER_263_1438 ();
 b15zdnd11an1n64x5 FILLER_263_1502 ();
 b15zdnd11an1n64x5 FILLER_263_1566 ();
 b15zdnd11an1n32x5 FILLER_263_1630 ();
 b15zdnd11an1n16x5 FILLER_263_1662 ();
 b15zdnd11an1n08x5 FILLER_263_1678 ();
 b15zdnd11an1n32x5 FILLER_263_1697 ();
 b15zdnd11an1n08x5 FILLER_263_1729 ();
 b15zdnd11an1n04x5 FILLER_263_1737 ();
 b15zdnd11an1n16x5 FILLER_263_1747 ();
 b15zdnd11an1n08x5 FILLER_263_1763 ();
 b15zdnd11an1n04x5 FILLER_263_1771 ();
 b15zdnd00an1n02x5 FILLER_263_1775 ();
 b15zdnd00an1n01x5 FILLER_263_1777 ();
 b15zdnd11an1n64x5 FILLER_263_1784 ();
 b15zdnd11an1n16x5 FILLER_263_1848 ();
 b15zdnd11an1n08x5 FILLER_263_1864 ();
 b15zdnd00an1n02x5 FILLER_263_1872 ();
 b15zdnd11an1n32x5 FILLER_263_1882 ();
 b15zdnd11an1n04x5 FILLER_263_1914 ();
 b15zdnd00an1n01x5 FILLER_263_1918 ();
 b15zdnd11an1n04x5 FILLER_263_1971 ();
 b15zdnd00an1n02x5 FILLER_263_1975 ();
 b15zdnd11an1n04x5 FILLER_263_1980 ();
 b15zdnd11an1n04x5 FILLER_263_1987 ();
 b15zdnd11an1n64x5 FILLER_263_1994 ();
 b15zdnd00an1n02x5 FILLER_263_2058 ();
 b15zdnd00an1n01x5 FILLER_263_2060 ();
 b15zdnd11an1n04x5 FILLER_263_2064 ();
 b15zdnd11an1n64x5 FILLER_263_2071 ();
 b15zdnd11an1n64x5 FILLER_263_2135 ();
 b15zdnd11an1n64x5 FILLER_263_2199 ();
 b15zdnd11an1n16x5 FILLER_263_2263 ();
 b15zdnd11an1n04x5 FILLER_263_2279 ();
 b15zdnd00an1n01x5 FILLER_263_2283 ();
 b15zdnd11an1n16x5 FILLER_264_8 ();
 b15zdnd00an1n02x5 FILLER_264_24 ();
 b15zdnd00an1n01x5 FILLER_264_26 ();
 b15zdnd11an1n04x5 FILLER_264_31 ();
 b15zdnd11an1n08x5 FILLER_264_60 ();
 b15zdnd11an1n04x5 FILLER_264_68 ();
 b15zdnd00an1n02x5 FILLER_264_72 ();
 b15zdnd00an1n01x5 FILLER_264_74 ();
 b15zdnd11an1n64x5 FILLER_264_82 ();
 b15zdnd11an1n64x5 FILLER_264_146 ();
 b15zdnd11an1n32x5 FILLER_264_210 ();
 b15zdnd11an1n16x5 FILLER_264_242 ();
 b15zdnd11an1n08x5 FILLER_264_258 ();
 b15zdnd11an1n04x5 FILLER_264_266 ();
 b15zdnd00an1n01x5 FILLER_264_270 ();
 b15zdnd11an1n64x5 FILLER_264_286 ();
 b15zdnd11an1n64x5 FILLER_264_350 ();
 b15zdnd11an1n64x5 FILLER_264_414 ();
 b15zdnd11an1n16x5 FILLER_264_478 ();
 b15zdnd00an1n02x5 FILLER_264_494 ();
 b15zdnd00an1n01x5 FILLER_264_496 ();
 b15zdnd11an1n32x5 FILLER_264_503 ();
 b15zdnd11an1n08x5 FILLER_264_535 ();
 b15zdnd00an1n02x5 FILLER_264_543 ();
 b15zdnd11an1n64x5 FILLER_264_548 ();
 b15zdnd11an1n64x5 FILLER_264_612 ();
 b15zdnd11an1n32x5 FILLER_264_676 ();
 b15zdnd11an1n08x5 FILLER_264_708 ();
 b15zdnd00an1n02x5 FILLER_264_716 ();
 b15zdnd11an1n16x5 FILLER_264_726 ();
 b15zdnd00an1n02x5 FILLER_264_742 ();
 b15zdnd11an1n64x5 FILLER_264_747 ();
 b15zdnd11an1n64x5 FILLER_264_811 ();
 b15zdnd11an1n64x5 FILLER_264_875 ();
 b15zdnd11an1n64x5 FILLER_264_939 ();
 b15zdnd11an1n04x5 FILLER_264_1003 ();
 b15zdnd00an1n02x5 FILLER_264_1007 ();
 b15zdnd00an1n01x5 FILLER_264_1009 ();
 b15zdnd11an1n64x5 FILLER_264_1018 ();
 b15zdnd11an1n08x5 FILLER_264_1082 ();
 b15zdnd00an1n01x5 FILLER_264_1090 ();
 b15zdnd11an1n64x5 FILLER_264_1101 ();
 b15zdnd11an1n64x5 FILLER_264_1165 ();
 b15zdnd11an1n64x5 FILLER_264_1229 ();
 b15zdnd11an1n64x5 FILLER_264_1293 ();
 b15zdnd11an1n64x5 FILLER_264_1357 ();
 b15zdnd11an1n64x5 FILLER_264_1421 ();
 b15zdnd11an1n64x5 FILLER_264_1485 ();
 b15zdnd11an1n64x5 FILLER_264_1549 ();
 b15zdnd11an1n64x5 FILLER_264_1613 ();
 b15zdnd11an1n16x5 FILLER_264_1677 ();
 b15zdnd11an1n08x5 FILLER_264_1693 ();
 b15zdnd00an1n02x5 FILLER_264_1701 ();
 b15zdnd11an1n32x5 FILLER_264_1709 ();
 b15zdnd11an1n16x5 FILLER_264_1741 ();
 b15zdnd11an1n08x5 FILLER_264_1757 ();
 b15zdnd11an1n32x5 FILLER_264_1773 ();
 b15zdnd11an1n16x5 FILLER_264_1805 ();
 b15zdnd11an1n08x5 FILLER_264_1821 ();
 b15zdnd11an1n04x5 FILLER_264_1829 ();
 b15zdnd11an1n64x5 FILLER_264_1837 ();
 b15zdnd11an1n16x5 FILLER_264_1901 ();
 b15zdnd00an1n02x5 FILLER_264_1917 ();
 b15zdnd00an1n01x5 FILLER_264_1919 ();
 b15zdnd11an1n08x5 FILLER_264_1972 ();
 b15zdnd00an1n02x5 FILLER_264_1980 ();
 b15zdnd11an1n32x5 FILLER_264_1985 ();
 b15zdnd11an1n16x5 FILLER_264_2017 ();
 b15zdnd11an1n08x5 FILLER_264_2033 ();
 b15zdnd11an1n64x5 FILLER_264_2085 ();
 b15zdnd11an1n04x5 FILLER_264_2149 ();
 b15zdnd00an1n01x5 FILLER_264_2153 ();
 b15zdnd11an1n64x5 FILLER_264_2162 ();
 b15zdnd11an1n32x5 FILLER_264_2226 ();
 b15zdnd11an1n16x5 FILLER_264_2258 ();
 b15zdnd00an1n02x5 FILLER_264_2274 ();
 b15zdnd11an1n16x5 FILLER_265_0 ();
 b15zdnd00an1n02x5 FILLER_265_16 ();
 b15zdnd11an1n04x5 FILLER_265_29 ();
 b15zdnd11an1n64x5 FILLER_265_38 ();
 b15zdnd11an1n64x5 FILLER_265_102 ();
 b15zdnd11an1n32x5 FILLER_265_166 ();
 b15zdnd11an1n16x5 FILLER_265_198 ();
 b15zdnd11an1n08x5 FILLER_265_214 ();
 b15zdnd11an1n04x5 FILLER_265_222 ();
 b15zdnd00an1n02x5 FILLER_265_226 ();
 b15zdnd00an1n01x5 FILLER_265_228 ();
 b15zdnd11an1n32x5 FILLER_265_241 ();
 b15zdnd11an1n16x5 FILLER_265_273 ();
 b15zdnd11an1n64x5 FILLER_265_331 ();
 b15zdnd11an1n64x5 FILLER_265_395 ();
 b15zdnd11an1n32x5 FILLER_265_459 ();
 b15zdnd11an1n16x5 FILLER_265_491 ();
 b15zdnd00an1n02x5 FILLER_265_507 ();
 b15zdnd00an1n01x5 FILLER_265_509 ();
 b15zdnd11an1n64x5 FILLER_265_552 ();
 b15zdnd11an1n64x5 FILLER_265_616 ();
 b15zdnd11an1n16x5 FILLER_265_680 ();
 b15zdnd11an1n08x5 FILLER_265_696 ();
 b15zdnd11an1n04x5 FILLER_265_704 ();
 b15zdnd11an1n08x5 FILLER_265_748 ();
 b15zdnd11an1n04x5 FILLER_265_756 ();
 b15zdnd11an1n64x5 FILLER_265_771 ();
 b15zdnd11an1n64x5 FILLER_265_835 ();
 b15zdnd11an1n64x5 FILLER_265_899 ();
 b15zdnd11an1n64x5 FILLER_265_963 ();
 b15zdnd11an1n64x5 FILLER_265_1027 ();
 b15zdnd11an1n64x5 FILLER_265_1091 ();
 b15zdnd11an1n64x5 FILLER_265_1155 ();
 b15zdnd11an1n64x5 FILLER_265_1219 ();
 b15zdnd11an1n64x5 FILLER_265_1283 ();
 b15zdnd11an1n64x5 FILLER_265_1347 ();
 b15zdnd11an1n64x5 FILLER_265_1411 ();
 b15zdnd11an1n32x5 FILLER_265_1475 ();
 b15zdnd11an1n16x5 FILLER_265_1507 ();
 b15zdnd11an1n08x5 FILLER_265_1523 ();
 b15zdnd00an1n02x5 FILLER_265_1531 ();
 b15zdnd11an1n08x5 FILLER_265_1537 ();
 b15zdnd11an1n04x5 FILLER_265_1545 ();
 b15zdnd00an1n01x5 FILLER_265_1549 ();
 b15zdnd11an1n64x5 FILLER_265_1554 ();
 b15zdnd11an1n64x5 FILLER_265_1618 ();
 b15zdnd11an1n08x5 FILLER_265_1682 ();
 b15zdnd00an1n01x5 FILLER_265_1690 ();
 b15zdnd11an1n64x5 FILLER_265_1697 ();
 b15zdnd11an1n16x5 FILLER_265_1761 ();
 b15zdnd11an1n04x5 FILLER_265_1777 ();
 b15zdnd00an1n02x5 FILLER_265_1781 ();
 b15zdnd11an1n64x5 FILLER_265_1825 ();
 b15zdnd11an1n32x5 FILLER_265_1889 ();
 b15zdnd00an1n01x5 FILLER_265_1921 ();
 b15zdnd11an1n64x5 FILLER_265_1964 ();
 b15zdnd11an1n32x5 FILLER_265_2028 ();
 b15zdnd00an1n02x5 FILLER_265_2060 ();
 b15zdnd00an1n01x5 FILLER_265_2062 ();
 b15zdnd11an1n64x5 FILLER_265_2066 ();
 b15zdnd11an1n64x5 FILLER_265_2130 ();
 b15zdnd11an1n64x5 FILLER_265_2194 ();
 b15zdnd11an1n16x5 FILLER_265_2258 ();
 b15zdnd11an1n08x5 FILLER_265_2274 ();
 b15zdnd00an1n02x5 FILLER_265_2282 ();
 b15zdnd00an1n02x5 FILLER_266_8 ();
 b15zdnd11an1n04x5 FILLER_266_16 ();
 b15zdnd00an1n01x5 FILLER_266_20 ();
 b15zdnd11an1n32x5 FILLER_266_25 ();
 b15zdnd11an1n16x5 FILLER_266_57 ();
 b15zdnd11an1n04x5 FILLER_266_73 ();
 b15zdnd00an1n01x5 FILLER_266_77 ();
 b15zdnd11an1n16x5 FILLER_266_87 ();
 b15zdnd11an1n08x5 FILLER_266_103 ();
 b15zdnd11an1n64x5 FILLER_266_129 ();
 b15zdnd11an1n64x5 FILLER_266_193 ();
 b15zdnd11an1n64x5 FILLER_266_257 ();
 b15zdnd11an1n64x5 FILLER_266_321 ();
 b15zdnd11an1n64x5 FILLER_266_385 ();
 b15zdnd11an1n64x5 FILLER_266_449 ();
 b15zdnd11an1n04x5 FILLER_266_513 ();
 b15zdnd00an1n01x5 FILLER_266_517 ();
 b15zdnd11an1n64x5 FILLER_266_570 ();
 b15zdnd11an1n64x5 FILLER_266_634 ();
 b15zdnd11an1n16x5 FILLER_266_698 ();
 b15zdnd11an1n04x5 FILLER_266_714 ();
 b15zdnd00an1n02x5 FILLER_266_726 ();
 b15zdnd11an1n08x5 FILLER_266_738 ();
 b15zdnd11an1n64x5 FILLER_266_749 ();
 b15zdnd11an1n64x5 FILLER_266_813 ();
 b15zdnd11an1n64x5 FILLER_266_877 ();
 b15zdnd11an1n64x5 FILLER_266_941 ();
 b15zdnd11an1n64x5 FILLER_266_1005 ();
 b15zdnd11an1n16x5 FILLER_266_1069 ();
 b15zdnd11an1n32x5 FILLER_266_1089 ();
 b15zdnd11an1n04x5 FILLER_266_1121 ();
 b15zdnd11an1n08x5 FILLER_266_1132 ();
 b15zdnd11an1n04x5 FILLER_266_1140 ();
 b15zdnd11an1n64x5 FILLER_266_1158 ();
 b15zdnd11an1n64x5 FILLER_266_1222 ();
 b15zdnd11an1n64x5 FILLER_266_1286 ();
 b15zdnd11an1n08x5 FILLER_266_1350 ();
 b15zdnd11an1n32x5 FILLER_266_1361 ();
 b15zdnd11an1n16x5 FILLER_266_1393 ();
 b15zdnd11an1n08x5 FILLER_266_1409 ();
 b15zdnd00an1n02x5 FILLER_266_1417 ();
 b15zdnd11an1n04x5 FILLER_266_1423 ();
 b15zdnd11an1n64x5 FILLER_266_1431 ();
 b15zdnd11an1n64x5 FILLER_266_1495 ();
 b15zdnd11an1n32x5 FILLER_266_1559 ();
 b15zdnd00an1n02x5 FILLER_266_1591 ();
 b15zdnd00an1n01x5 FILLER_266_1593 ();
 b15zdnd11an1n64x5 FILLER_266_1608 ();
 b15zdnd11an1n16x5 FILLER_266_1672 ();
 b15zdnd11an1n08x5 FILLER_266_1688 ();
 b15zdnd00an1n02x5 FILLER_266_1696 ();
 b15zdnd11an1n32x5 FILLER_266_1706 ();
 b15zdnd11an1n04x5 FILLER_266_1738 ();
 b15zdnd00an1n01x5 FILLER_266_1742 ();
 b15zdnd11an1n08x5 FILLER_266_1751 ();
 b15zdnd00an1n02x5 FILLER_266_1759 ();
 b15zdnd11an1n04x5 FILLER_266_1781 ();
 b15zdnd11an1n64x5 FILLER_266_1803 ();
 b15zdnd11an1n64x5 FILLER_266_1867 ();
 b15zdnd11an1n04x5 FILLER_266_1931 ();
 b15zdnd00an1n02x5 FILLER_266_1935 ();
 b15zdnd11an1n04x5 FILLER_266_1940 ();
 b15zdnd11an1n04x5 FILLER_266_1947 ();
 b15zdnd11an1n04x5 FILLER_266_1954 ();
 b15zdnd11an1n64x5 FILLER_266_1961 ();
 b15zdnd11an1n64x5 FILLER_266_2025 ();
 b15zdnd11an1n64x5 FILLER_266_2089 ();
 b15zdnd00an1n01x5 FILLER_266_2153 ();
 b15zdnd11an1n64x5 FILLER_266_2162 ();
 b15zdnd11an1n32x5 FILLER_266_2226 ();
 b15zdnd11an1n16x5 FILLER_266_2258 ();
 b15zdnd00an1n02x5 FILLER_266_2274 ();
 b15zdnd11an1n32x5 FILLER_267_0 ();
 b15zdnd11an1n04x5 FILLER_267_32 ();
 b15zdnd00an1n02x5 FILLER_267_36 ();
 b15zdnd11an1n64x5 FILLER_267_44 ();
 b15zdnd11an1n64x5 FILLER_267_108 ();
 b15zdnd11an1n32x5 FILLER_267_172 ();
 b15zdnd11an1n08x5 FILLER_267_204 ();
 b15zdnd00an1n02x5 FILLER_267_212 ();
 b15zdnd00an1n01x5 FILLER_267_214 ();
 b15zdnd11an1n32x5 FILLER_267_227 ();
 b15zdnd11an1n04x5 FILLER_267_259 ();
 b15zdnd00an1n02x5 FILLER_267_263 ();
 b15zdnd00an1n01x5 FILLER_267_265 ();
 b15zdnd11an1n04x5 FILLER_267_308 ();
 b15zdnd00an1n02x5 FILLER_267_312 ();
 b15zdnd00an1n01x5 FILLER_267_314 ();
 b15zdnd11an1n64x5 FILLER_267_319 ();
 b15zdnd11an1n64x5 FILLER_267_383 ();
 b15zdnd11an1n32x5 FILLER_267_447 ();
 b15zdnd11an1n16x5 FILLER_267_479 ();
 b15zdnd11an1n08x5 FILLER_267_495 ();
 b15zdnd00an1n01x5 FILLER_267_503 ();
 b15zdnd11an1n16x5 FILLER_267_512 ();
 b15zdnd11an1n08x5 FILLER_267_528 ();
 b15zdnd00an1n01x5 FILLER_267_536 ();
 b15zdnd11an1n04x5 FILLER_267_579 ();
 b15zdnd11an1n64x5 FILLER_267_590 ();
 b15zdnd11an1n64x5 FILLER_267_654 ();
 b15zdnd11an1n64x5 FILLER_267_718 ();
 b15zdnd11an1n16x5 FILLER_267_782 ();
 b15zdnd11an1n08x5 FILLER_267_798 ();
 b15zdnd11an1n04x5 FILLER_267_806 ();
 b15zdnd11an1n16x5 FILLER_267_821 ();
 b15zdnd11an1n64x5 FILLER_267_841 ();
 b15zdnd11an1n64x5 FILLER_267_905 ();
 b15zdnd11an1n64x5 FILLER_267_969 ();
 b15zdnd11an1n32x5 FILLER_267_1033 ();
 b15zdnd11an1n08x5 FILLER_267_1065 ();
 b15zdnd11an1n04x5 FILLER_267_1073 ();
 b15zdnd00an1n02x5 FILLER_267_1077 ();
 b15zdnd00an1n01x5 FILLER_267_1079 ();
 b15zdnd11an1n16x5 FILLER_267_1106 ();
 b15zdnd11an1n08x5 FILLER_267_1122 ();
 b15zdnd00an1n02x5 FILLER_267_1130 ();
 b15zdnd11an1n64x5 FILLER_267_1174 ();
 b15zdnd11an1n64x5 FILLER_267_1238 ();
 b15zdnd11an1n32x5 FILLER_267_1302 ();
 b15zdnd11an1n08x5 FILLER_267_1334 ();
 b15zdnd11an1n04x5 FILLER_267_1342 ();
 b15zdnd00an1n02x5 FILLER_267_1346 ();
 b15zdnd11an1n04x5 FILLER_267_1351 ();
 b15zdnd00an1n02x5 FILLER_267_1355 ();
 b15zdnd11an1n32x5 FILLER_267_1373 ();
 b15zdnd11an1n16x5 FILLER_267_1405 ();
 b15zdnd11an1n08x5 FILLER_267_1421 ();
 b15zdnd11an1n04x5 FILLER_267_1429 ();
 b15zdnd00an1n02x5 FILLER_267_1433 ();
 b15zdnd11an1n64x5 FILLER_267_1439 ();
 b15zdnd11an1n16x5 FILLER_267_1503 ();
 b15zdnd11an1n08x5 FILLER_267_1519 ();
 b15zdnd00an1n01x5 FILLER_267_1527 ();
 b15zdnd11an1n32x5 FILLER_267_1532 ();
 b15zdnd00an1n01x5 FILLER_267_1564 ();
 b15zdnd11an1n32x5 FILLER_267_1571 ();
 b15zdnd11an1n16x5 FILLER_267_1603 ();
 b15zdnd11an1n08x5 FILLER_267_1619 ();
 b15zdnd00an1n02x5 FILLER_267_1627 ();
 b15zdnd11an1n32x5 FILLER_267_1636 ();
 b15zdnd11an1n16x5 FILLER_267_1668 ();
 b15zdnd11an1n04x5 FILLER_267_1684 ();
 b15zdnd11an1n64x5 FILLER_267_1694 ();
 b15zdnd11an1n64x5 FILLER_267_1758 ();
 b15zdnd11an1n64x5 FILLER_267_1822 ();
 b15zdnd11an1n32x5 FILLER_267_1886 ();
 b15zdnd11an1n16x5 FILLER_267_1918 ();
 b15zdnd11an1n08x5 FILLER_267_1934 ();
 b15zdnd00an1n02x5 FILLER_267_1942 ();
 b15zdnd00an1n01x5 FILLER_267_1944 ();
 b15zdnd11an1n64x5 FILLER_267_1948 ();
 b15zdnd11an1n64x5 FILLER_267_2012 ();
 b15zdnd11an1n64x5 FILLER_267_2076 ();
 b15zdnd11an1n64x5 FILLER_267_2140 ();
 b15zdnd11an1n64x5 FILLER_267_2204 ();
 b15zdnd11an1n16x5 FILLER_267_2268 ();
 b15zdnd11an1n64x5 FILLER_268_8 ();
 b15zdnd11an1n16x5 FILLER_268_72 ();
 b15zdnd11an1n64x5 FILLER_268_113 ();
 b15zdnd11an1n64x5 FILLER_268_177 ();
 b15zdnd11an1n64x5 FILLER_268_241 ();
 b15zdnd11an1n32x5 FILLER_268_305 ();
 b15zdnd11an1n08x5 FILLER_268_337 ();
 b15zdnd11an1n04x5 FILLER_268_345 ();
 b15zdnd00an1n02x5 FILLER_268_349 ();
 b15zdnd11an1n04x5 FILLER_268_372 ();
 b15zdnd11an1n08x5 FILLER_268_428 ();
 b15zdnd00an1n02x5 FILLER_268_436 ();
 b15zdnd11an1n64x5 FILLER_268_446 ();
 b15zdnd11an1n16x5 FILLER_268_510 ();
 b15zdnd11an1n08x5 FILLER_268_526 ();
 b15zdnd00an1n02x5 FILLER_268_534 ();
 b15zdnd11an1n04x5 FILLER_268_539 ();
 b15zdnd11an1n64x5 FILLER_268_546 ();
 b15zdnd11an1n64x5 FILLER_268_610 ();
 b15zdnd11an1n32x5 FILLER_268_674 ();
 b15zdnd11an1n08x5 FILLER_268_706 ();
 b15zdnd11an1n04x5 FILLER_268_714 ();
 b15zdnd00an1n02x5 FILLER_268_726 ();
 b15zdnd11an1n04x5 FILLER_268_754 ();
 b15zdnd11an1n64x5 FILLER_268_772 ();
 b15zdnd11an1n64x5 FILLER_268_836 ();
 b15zdnd11an1n64x5 FILLER_268_900 ();
 b15zdnd11an1n64x5 FILLER_268_964 ();
 b15zdnd11an1n64x5 FILLER_268_1028 ();
 b15zdnd11an1n64x5 FILLER_268_1092 ();
 b15zdnd11an1n64x5 FILLER_268_1156 ();
 b15zdnd11an1n64x5 FILLER_268_1220 ();
 b15zdnd11an1n32x5 FILLER_268_1284 ();
 b15zdnd11an1n04x5 FILLER_268_1316 ();
 b15zdnd00an1n02x5 FILLER_268_1320 ();
 b15zdnd11an1n04x5 FILLER_268_1342 ();
 b15zdnd11an1n04x5 FILLER_268_1359 ();
 b15zdnd11an1n64x5 FILLER_268_1373 ();
 b15zdnd11an1n64x5 FILLER_268_1437 ();
 b15zdnd11an1n32x5 FILLER_268_1501 ();
 b15zdnd11an1n08x5 FILLER_268_1533 ();
 b15zdnd00an1n01x5 FILLER_268_1541 ();
 b15zdnd11an1n08x5 FILLER_268_1546 ();
 b15zdnd00an1n02x5 FILLER_268_1554 ();
 b15zdnd11an1n64x5 FILLER_268_1560 ();
 b15zdnd11an1n64x5 FILLER_268_1624 ();
 b15zdnd11an1n64x5 FILLER_268_1688 ();
 b15zdnd11an1n64x5 FILLER_268_1752 ();
 b15zdnd11an1n16x5 FILLER_268_1816 ();
 b15zdnd00an1n02x5 FILLER_268_1832 ();
 b15zdnd00an1n01x5 FILLER_268_1834 ();
 b15zdnd11an1n64x5 FILLER_268_1877 ();
 b15zdnd11an1n64x5 FILLER_268_1941 ();
 b15zdnd11an1n64x5 FILLER_268_2005 ();
 b15zdnd11an1n64x5 FILLER_268_2069 ();
 b15zdnd11an1n16x5 FILLER_268_2133 ();
 b15zdnd11an1n04x5 FILLER_268_2149 ();
 b15zdnd00an1n01x5 FILLER_268_2153 ();
 b15zdnd11an1n64x5 FILLER_268_2162 ();
 b15zdnd11an1n32x5 FILLER_268_2226 ();
 b15zdnd11an1n16x5 FILLER_268_2258 ();
 b15zdnd00an1n02x5 FILLER_268_2274 ();
 b15zdnd11an1n16x5 FILLER_269_0 ();
 b15zdnd11an1n64x5 FILLER_269_23 ();
 b15zdnd11an1n64x5 FILLER_269_87 ();
 b15zdnd11an1n64x5 FILLER_269_151 ();
 b15zdnd11an1n64x5 FILLER_269_215 ();
 b15zdnd11an1n64x5 FILLER_269_279 ();
 b15zdnd11an1n08x5 FILLER_269_343 ();
 b15zdnd00an1n02x5 FILLER_269_351 ();
 b15zdnd00an1n01x5 FILLER_269_353 ();
 b15zdnd11an1n04x5 FILLER_269_361 ();
 b15zdnd00an1n02x5 FILLER_269_365 ();
 b15zdnd11an1n04x5 FILLER_269_409 ();
 b15zdnd11an1n04x5 FILLER_269_416 ();
 b15zdnd11an1n64x5 FILLER_269_462 ();
 b15zdnd11an1n64x5 FILLER_269_526 ();
 b15zdnd11an1n64x5 FILLER_269_590 ();
 b15zdnd11an1n64x5 FILLER_269_654 ();
 b15zdnd11an1n16x5 FILLER_269_718 ();
 b15zdnd11an1n08x5 FILLER_269_734 ();
 b15zdnd11an1n04x5 FILLER_269_742 ();
 b15zdnd00an1n01x5 FILLER_269_746 ();
 b15zdnd11an1n64x5 FILLER_269_761 ();
 b15zdnd11an1n16x5 FILLER_269_825 ();
 b15zdnd11an1n04x5 FILLER_269_841 ();
 b15zdnd00an1n02x5 FILLER_269_845 ();
 b15zdnd11an1n64x5 FILLER_269_851 ();
 b15zdnd11an1n64x5 FILLER_269_915 ();
 b15zdnd11an1n32x5 FILLER_269_979 ();
 b15zdnd11an1n04x5 FILLER_269_1011 ();
 b15zdnd00an1n01x5 FILLER_269_1015 ();
 b15zdnd11an1n64x5 FILLER_269_1036 ();
 b15zdnd11an1n64x5 FILLER_269_1100 ();
 b15zdnd11an1n32x5 FILLER_269_1164 ();
 b15zdnd00an1n02x5 FILLER_269_1196 ();
 b15zdnd00an1n01x5 FILLER_269_1198 ();
 b15zdnd11an1n64x5 FILLER_269_1202 ();
 b15zdnd11an1n64x5 FILLER_269_1266 ();
 b15zdnd11an1n32x5 FILLER_269_1330 ();
 b15zdnd11an1n08x5 FILLER_269_1362 ();
 b15zdnd00an1n01x5 FILLER_269_1370 ();
 b15zdnd11an1n64x5 FILLER_269_1397 ();
 b15zdnd11an1n64x5 FILLER_269_1461 ();
 b15zdnd11an1n64x5 FILLER_269_1525 ();
 b15zdnd11an1n64x5 FILLER_269_1589 ();
 b15zdnd11an1n64x5 FILLER_269_1653 ();
 b15zdnd11an1n64x5 FILLER_269_1717 ();
 b15zdnd00an1n01x5 FILLER_269_1781 ();
 b15zdnd11an1n64x5 FILLER_269_1786 ();
 b15zdnd11an1n64x5 FILLER_269_1850 ();
 b15zdnd11an1n64x5 FILLER_269_1914 ();
 b15zdnd11an1n64x5 FILLER_269_1978 ();
 b15zdnd11an1n64x5 FILLER_269_2042 ();
 b15zdnd11an1n64x5 FILLER_269_2106 ();
 b15zdnd11an1n64x5 FILLER_269_2170 ();
 b15zdnd11an1n32x5 FILLER_269_2234 ();
 b15zdnd11an1n16x5 FILLER_269_2266 ();
 b15zdnd00an1n02x5 FILLER_269_2282 ();
 b15zdnd11an1n04x5 FILLER_270_8 ();
 b15zdnd11an1n32x5 FILLER_270_19 ();
 b15zdnd11an1n08x5 FILLER_270_51 ();
 b15zdnd11an1n04x5 FILLER_270_59 ();
 b15zdnd00an1n02x5 FILLER_270_63 ();
 b15zdnd11an1n32x5 FILLER_270_96 ();
 b15zdnd11an1n16x5 FILLER_270_128 ();
 b15zdnd11an1n04x5 FILLER_270_144 ();
 b15zdnd00an1n02x5 FILLER_270_148 ();
 b15zdnd00an1n01x5 FILLER_270_150 ();
 b15zdnd11an1n64x5 FILLER_270_177 ();
 b15zdnd11an1n64x5 FILLER_270_241 ();
 b15zdnd11an1n32x5 FILLER_270_305 ();
 b15zdnd11an1n16x5 FILLER_270_337 ();
 b15zdnd11an1n08x5 FILLER_270_353 ();
 b15zdnd11an1n04x5 FILLER_270_361 ();
 b15zdnd11an1n04x5 FILLER_270_383 ();
 b15zdnd11an1n04x5 FILLER_270_394 ();
 b15zdnd11an1n04x5 FILLER_270_401 ();
 b15zdnd11an1n04x5 FILLER_270_408 ();
 b15zdnd00an1n01x5 FILLER_270_412 ();
 b15zdnd11an1n64x5 FILLER_270_420 ();
 b15zdnd11an1n64x5 FILLER_270_484 ();
 b15zdnd11an1n64x5 FILLER_270_548 ();
 b15zdnd11an1n64x5 FILLER_270_612 ();
 b15zdnd11an1n32x5 FILLER_270_676 ();
 b15zdnd11an1n08x5 FILLER_270_708 ();
 b15zdnd00an1n02x5 FILLER_270_716 ();
 b15zdnd11an1n64x5 FILLER_270_726 ();
 b15zdnd11an1n64x5 FILLER_270_790 ();
 b15zdnd11an1n64x5 FILLER_270_854 ();
 b15zdnd11an1n64x5 FILLER_270_918 ();
 b15zdnd11an1n64x5 FILLER_270_982 ();
 b15zdnd11an1n64x5 FILLER_270_1046 ();
 b15zdnd11an1n64x5 FILLER_270_1110 ();
 b15zdnd11an1n16x5 FILLER_270_1174 ();
 b15zdnd11an1n04x5 FILLER_270_1190 ();
 b15zdnd00an1n02x5 FILLER_270_1194 ();
 b15zdnd00an1n01x5 FILLER_270_1196 ();
 b15zdnd11an1n04x5 FILLER_270_1200 ();
 b15zdnd11an1n64x5 FILLER_270_1207 ();
 b15zdnd11an1n32x5 FILLER_270_1271 ();
 b15zdnd11an1n16x5 FILLER_270_1303 ();
 b15zdnd11an1n08x5 FILLER_270_1319 ();
 b15zdnd11an1n04x5 FILLER_270_1327 ();
 b15zdnd00an1n02x5 FILLER_270_1331 ();
 b15zdnd11an1n64x5 FILLER_270_1346 ();
 b15zdnd11an1n64x5 FILLER_270_1410 ();
 b15zdnd11an1n32x5 FILLER_270_1474 ();
 b15zdnd11an1n16x5 FILLER_270_1506 ();
 b15zdnd11an1n08x5 FILLER_270_1522 ();
 b15zdnd11an1n04x5 FILLER_270_1530 ();
 b15zdnd00an1n01x5 FILLER_270_1534 ();
 b15zdnd11an1n64x5 FILLER_270_1577 ();
 b15zdnd11an1n32x5 FILLER_270_1641 ();
 b15zdnd11an1n16x5 FILLER_270_1673 ();
 b15zdnd11an1n08x5 FILLER_270_1689 ();
 b15zdnd11an1n64x5 FILLER_270_1703 ();
 b15zdnd11an1n64x5 FILLER_270_1767 ();
 b15zdnd11an1n64x5 FILLER_270_1831 ();
 b15zdnd11an1n64x5 FILLER_270_1895 ();
 b15zdnd11an1n64x5 FILLER_270_1959 ();
 b15zdnd11an1n32x5 FILLER_270_2023 ();
 b15zdnd11an1n04x5 FILLER_270_2055 ();
 b15zdnd00an1n01x5 FILLER_270_2059 ();
 b15zdnd11an1n64x5 FILLER_270_2075 ();
 b15zdnd11an1n08x5 FILLER_270_2139 ();
 b15zdnd11an1n04x5 FILLER_270_2147 ();
 b15zdnd00an1n02x5 FILLER_270_2151 ();
 b15zdnd00an1n01x5 FILLER_270_2153 ();
 b15zdnd11an1n64x5 FILLER_270_2162 ();
 b15zdnd11an1n32x5 FILLER_270_2226 ();
 b15zdnd11an1n04x5 FILLER_270_2258 ();
 b15zdnd11an1n08x5 FILLER_270_2266 ();
 b15zdnd00an1n02x5 FILLER_270_2274 ();
 b15zdnd11an1n64x5 FILLER_271_0 ();
 b15zdnd11an1n64x5 FILLER_271_64 ();
 b15zdnd11an1n16x5 FILLER_271_128 ();
 b15zdnd11an1n08x5 FILLER_271_144 ();
 b15zdnd00an1n01x5 FILLER_271_152 ();
 b15zdnd11an1n16x5 FILLER_271_165 ();
 b15zdnd11an1n64x5 FILLER_271_206 ();
 b15zdnd11an1n16x5 FILLER_271_270 ();
 b15zdnd11an1n32x5 FILLER_271_311 ();
 b15zdnd11an1n16x5 FILLER_271_343 ();
 b15zdnd11an1n04x5 FILLER_271_359 ();
 b15zdnd00an1n02x5 FILLER_271_363 ();
 b15zdnd00an1n01x5 FILLER_271_365 ();
 b15zdnd11an1n64x5 FILLER_271_376 ();
 b15zdnd11an1n64x5 FILLER_271_440 ();
 b15zdnd11an1n64x5 FILLER_271_504 ();
 b15zdnd11an1n64x5 FILLER_271_568 ();
 b15zdnd11an1n64x5 FILLER_271_632 ();
 b15zdnd11an1n64x5 FILLER_271_696 ();
 b15zdnd11an1n64x5 FILLER_271_760 ();
 b15zdnd11an1n64x5 FILLER_271_824 ();
 b15zdnd11an1n64x5 FILLER_271_888 ();
 b15zdnd11an1n64x5 FILLER_271_952 ();
 b15zdnd11an1n16x5 FILLER_271_1016 ();
 b15zdnd11an1n08x5 FILLER_271_1032 ();
 b15zdnd00an1n01x5 FILLER_271_1040 ();
 b15zdnd11an1n64x5 FILLER_271_1045 ();
 b15zdnd11an1n64x5 FILLER_271_1109 ();
 b15zdnd11an1n04x5 FILLER_271_1173 ();
 b15zdnd00an1n02x5 FILLER_271_1177 ();
 b15zdnd11an1n64x5 FILLER_271_1231 ();
 b15zdnd11an1n32x5 FILLER_271_1295 ();
 b15zdnd11an1n08x5 FILLER_271_1327 ();
 b15zdnd11an1n04x5 FILLER_271_1335 ();
 b15zdnd00an1n02x5 FILLER_271_1339 ();
 b15zdnd11an1n64x5 FILLER_271_1357 ();
 b15zdnd11an1n64x5 FILLER_271_1421 ();
 b15zdnd11an1n64x5 FILLER_271_1485 ();
 b15zdnd11an1n64x5 FILLER_271_1549 ();
 b15zdnd11an1n64x5 FILLER_271_1613 ();
 b15zdnd11an1n64x5 FILLER_271_1677 ();
 b15zdnd11an1n32x5 FILLER_271_1741 ();
 b15zdnd11an1n04x5 FILLER_271_1773 ();
 b15zdnd11an1n64x5 FILLER_271_1783 ();
 b15zdnd11an1n64x5 FILLER_271_1847 ();
 b15zdnd11an1n64x5 FILLER_271_1911 ();
 b15zdnd11an1n64x5 FILLER_271_1975 ();
 b15zdnd11an1n64x5 FILLER_271_2039 ();
 b15zdnd11an1n64x5 FILLER_271_2103 ();
 b15zdnd11an1n64x5 FILLER_271_2167 ();
 b15zdnd11an1n32x5 FILLER_271_2231 ();
 b15zdnd11an1n16x5 FILLER_271_2263 ();
 b15zdnd11an1n04x5 FILLER_271_2279 ();
 b15zdnd00an1n01x5 FILLER_271_2283 ();
 b15zdnd11an1n16x5 FILLER_272_8 ();
 b15zdnd00an1n02x5 FILLER_272_24 ();
 b15zdnd00an1n01x5 FILLER_272_26 ();
 b15zdnd11an1n04x5 FILLER_272_33 ();
 b15zdnd11an1n64x5 FILLER_272_43 ();
 b15zdnd11an1n64x5 FILLER_272_107 ();
 b15zdnd11an1n64x5 FILLER_272_171 ();
 b15zdnd11an1n32x5 FILLER_272_235 ();
 b15zdnd11an1n16x5 FILLER_272_267 ();
 b15zdnd11an1n08x5 FILLER_272_283 ();
 b15zdnd11an1n04x5 FILLER_272_291 ();
 b15zdnd11an1n32x5 FILLER_272_320 ();
 b15zdnd11an1n08x5 FILLER_272_352 ();
 b15zdnd11an1n04x5 FILLER_272_360 ();
 b15zdnd00an1n02x5 FILLER_272_364 ();
 b15zdnd00an1n01x5 FILLER_272_366 ();
 b15zdnd11an1n64x5 FILLER_272_374 ();
 b15zdnd11an1n64x5 FILLER_272_438 ();
 b15zdnd11an1n64x5 FILLER_272_502 ();
 b15zdnd11an1n16x5 FILLER_272_566 ();
 b15zdnd11an1n04x5 FILLER_272_582 ();
 b15zdnd00an1n01x5 FILLER_272_586 ();
 b15zdnd11an1n04x5 FILLER_272_590 ();
 b15zdnd11an1n64x5 FILLER_272_597 ();
 b15zdnd11an1n32x5 FILLER_272_661 ();
 b15zdnd11an1n16x5 FILLER_272_693 ();
 b15zdnd11an1n08x5 FILLER_272_709 ();
 b15zdnd00an1n01x5 FILLER_272_717 ();
 b15zdnd11an1n64x5 FILLER_272_726 ();
 b15zdnd11an1n64x5 FILLER_272_790 ();
 b15zdnd11an1n64x5 FILLER_272_854 ();
 b15zdnd11an1n16x5 FILLER_272_918 ();
 b15zdnd11an1n08x5 FILLER_272_934 ();
 b15zdnd00an1n02x5 FILLER_272_942 ();
 b15zdnd11an1n64x5 FILLER_272_947 ();
 b15zdnd11an1n32x5 FILLER_272_1011 ();
 b15zdnd11an1n16x5 FILLER_272_1043 ();
 b15zdnd00an1n02x5 FILLER_272_1059 ();
 b15zdnd00an1n01x5 FILLER_272_1061 ();
 b15zdnd11an1n04x5 FILLER_272_1066 ();
 b15zdnd11an1n64x5 FILLER_272_1088 ();
 b15zdnd11an1n64x5 FILLER_272_1152 ();
 b15zdnd11an1n64x5 FILLER_272_1216 ();
 b15zdnd11an1n32x5 FILLER_272_1280 ();
 b15zdnd11an1n16x5 FILLER_272_1312 ();
 b15zdnd11an1n04x5 FILLER_272_1328 ();
 b15zdnd11an1n04x5 FILLER_272_1347 ();
 b15zdnd00an1n01x5 FILLER_272_1351 ();
 b15zdnd11an1n32x5 FILLER_272_1364 ();
 b15zdnd11an1n04x5 FILLER_272_1396 ();
 b15zdnd00an1n02x5 FILLER_272_1400 ();
 b15zdnd00an1n01x5 FILLER_272_1402 ();
 b15zdnd11an1n64x5 FILLER_272_1414 ();
 b15zdnd11an1n64x5 FILLER_272_1478 ();
 b15zdnd11an1n64x5 FILLER_272_1542 ();
 b15zdnd11an1n64x5 FILLER_272_1606 ();
 b15zdnd11an1n32x5 FILLER_272_1670 ();
 b15zdnd11an1n08x5 FILLER_272_1706 ();
 b15zdnd11an1n04x5 FILLER_272_1714 ();
 b15zdnd00an1n02x5 FILLER_272_1718 ();
 b15zdnd00an1n01x5 FILLER_272_1720 ();
 b15zdnd11an1n04x5 FILLER_272_1741 ();
 b15zdnd11an1n32x5 FILLER_272_1753 ();
 b15zdnd11an1n04x5 FILLER_272_1785 ();
 b15zdnd00an1n02x5 FILLER_272_1789 ();
 b15zdnd00an1n01x5 FILLER_272_1791 ();
 b15zdnd11an1n64x5 FILLER_272_1796 ();
 b15zdnd11an1n64x5 FILLER_272_1860 ();
 b15zdnd11an1n64x5 FILLER_272_1924 ();
 b15zdnd11an1n64x5 FILLER_272_1988 ();
 b15zdnd11an1n08x5 FILLER_272_2052 ();
 b15zdnd11an1n04x5 FILLER_272_2060 ();
 b15zdnd11an1n04x5 FILLER_272_2070 ();
 b15zdnd00an1n02x5 FILLER_272_2074 ();
 b15zdnd00an1n01x5 FILLER_272_2076 ();
 b15zdnd11an1n64x5 FILLER_272_2080 ();
 b15zdnd11an1n08x5 FILLER_272_2144 ();
 b15zdnd00an1n02x5 FILLER_272_2152 ();
 b15zdnd11an1n64x5 FILLER_272_2162 ();
 b15zdnd11an1n32x5 FILLER_272_2226 ();
 b15zdnd11an1n16x5 FILLER_272_2258 ();
 b15zdnd00an1n02x5 FILLER_272_2274 ();
 b15zdnd11an1n64x5 FILLER_273_0 ();
 b15zdnd11an1n64x5 FILLER_273_64 ();
 b15zdnd11an1n64x5 FILLER_273_128 ();
 b15zdnd11an1n64x5 FILLER_273_192 ();
 b15zdnd11an1n64x5 FILLER_273_256 ();
 b15zdnd11an1n64x5 FILLER_273_320 ();
 b15zdnd11an1n64x5 FILLER_273_384 ();
 b15zdnd11an1n64x5 FILLER_273_448 ();
 b15zdnd11an1n32x5 FILLER_273_512 ();
 b15zdnd11an1n16x5 FILLER_273_544 ();
 b15zdnd11an1n04x5 FILLER_273_560 ();
 b15zdnd00an1n02x5 FILLER_273_564 ();
 b15zdnd00an1n01x5 FILLER_273_566 ();
 b15zdnd11an1n04x5 FILLER_273_619 ();
 b15zdnd11an1n64x5 FILLER_273_641 ();
 b15zdnd11an1n64x5 FILLER_273_705 ();
 b15zdnd11an1n64x5 FILLER_273_769 ();
 b15zdnd11an1n32x5 FILLER_273_833 ();
 b15zdnd11an1n16x5 FILLER_273_865 ();
 b15zdnd00an1n02x5 FILLER_273_881 ();
 b15zdnd11an1n04x5 FILLER_273_935 ();
 b15zdnd00an1n02x5 FILLER_273_939 ();
 b15zdnd11an1n04x5 FILLER_273_944 ();
 b15zdnd11an1n04x5 FILLER_273_951 ();
 b15zdnd11an1n32x5 FILLER_273_958 ();
 b15zdnd11an1n08x5 FILLER_273_990 ();
 b15zdnd00an1n02x5 FILLER_273_998 ();
 b15zdnd11an1n64x5 FILLER_273_1007 ();
 b15zdnd11an1n16x5 FILLER_273_1071 ();
 b15zdnd11an1n08x5 FILLER_273_1087 ();
 b15zdnd00an1n01x5 FILLER_273_1095 ();
 b15zdnd11an1n04x5 FILLER_273_1101 ();
 b15zdnd11an1n64x5 FILLER_273_1125 ();
 b15zdnd11an1n32x5 FILLER_273_1189 ();
 b15zdnd11an1n08x5 FILLER_273_1221 ();
 b15zdnd00an1n01x5 FILLER_273_1229 ();
 b15zdnd11an1n64x5 FILLER_273_1250 ();
 b15zdnd11an1n64x5 FILLER_273_1314 ();
 b15zdnd11an1n64x5 FILLER_273_1378 ();
 b15zdnd11an1n64x5 FILLER_273_1442 ();
 b15zdnd11an1n64x5 FILLER_273_1506 ();
 b15zdnd11an1n64x5 FILLER_273_1570 ();
 b15zdnd11an1n64x5 FILLER_273_1634 ();
 b15zdnd11an1n04x5 FILLER_273_1698 ();
 b15zdnd00an1n01x5 FILLER_273_1702 ();
 b15zdnd11an1n04x5 FILLER_273_1707 ();
 b15zdnd11an1n64x5 FILLER_273_1715 ();
 b15zdnd11an1n08x5 FILLER_273_1779 ();
 b15zdnd00an1n02x5 FILLER_273_1787 ();
 b15zdnd11an1n64x5 FILLER_273_1793 ();
 b15zdnd11an1n64x5 FILLER_273_1857 ();
 b15zdnd11an1n64x5 FILLER_273_1921 ();
 b15zdnd11an1n64x5 FILLER_273_1985 ();
 b15zdnd11an1n64x5 FILLER_273_2049 ();
 b15zdnd11an1n64x5 FILLER_273_2113 ();
 b15zdnd11an1n16x5 FILLER_273_2177 ();
 b15zdnd11an1n04x5 FILLER_273_2193 ();
 b15zdnd00an1n02x5 FILLER_273_2197 ();
 b15zdnd00an1n01x5 FILLER_273_2199 ();
 b15zdnd11an1n32x5 FILLER_273_2242 ();
 b15zdnd11an1n08x5 FILLER_273_2274 ();
 b15zdnd00an1n02x5 FILLER_273_2282 ();
 b15zdnd11an1n64x5 FILLER_274_8 ();
 b15zdnd11an1n64x5 FILLER_274_72 ();
 b15zdnd11an1n64x5 FILLER_274_136 ();
 b15zdnd11an1n64x5 FILLER_274_200 ();
 b15zdnd11an1n16x5 FILLER_274_264 ();
 b15zdnd11an1n64x5 FILLER_274_286 ();
 b15zdnd11an1n64x5 FILLER_274_350 ();
 b15zdnd11an1n64x5 FILLER_274_414 ();
 b15zdnd11an1n64x5 FILLER_274_478 ();
 b15zdnd11an1n32x5 FILLER_274_542 ();
 b15zdnd11an1n16x5 FILLER_274_574 ();
 b15zdnd00an1n02x5 FILLER_274_590 ();
 b15zdnd11an1n16x5 FILLER_274_595 ();
 b15zdnd11an1n08x5 FILLER_274_611 ();
 b15zdnd00an1n02x5 FILLER_274_619 ();
 b15zdnd11an1n32x5 FILLER_274_663 ();
 b15zdnd11an1n16x5 FILLER_274_695 ();
 b15zdnd11an1n04x5 FILLER_274_711 ();
 b15zdnd00an1n02x5 FILLER_274_715 ();
 b15zdnd00an1n01x5 FILLER_274_717 ();
 b15zdnd11an1n64x5 FILLER_274_726 ();
 b15zdnd00an1n02x5 FILLER_274_790 ();
 b15zdnd11an1n64x5 FILLER_274_795 ();
 b15zdnd11an1n32x5 FILLER_274_859 ();
 b15zdnd11an1n08x5 FILLER_274_891 ();
 b15zdnd11an1n04x5 FILLER_274_899 ();
 b15zdnd00an1n02x5 FILLER_274_903 ();
 b15zdnd00an1n01x5 FILLER_274_905 ();
 b15zdnd11an1n04x5 FILLER_274_909 ();
 b15zdnd11an1n04x5 FILLER_274_916 ();
 b15zdnd00an1n01x5 FILLER_274_920 ();
 b15zdnd11an1n08x5 FILLER_274_973 ();
 b15zdnd11an1n08x5 FILLER_274_1001 ();
 b15zdnd00an1n02x5 FILLER_274_1009 ();
 b15zdnd00an1n01x5 FILLER_274_1011 ();
 b15zdnd11an1n64x5 FILLER_274_1019 ();
 b15zdnd11an1n16x5 FILLER_274_1083 ();
 b15zdnd11an1n08x5 FILLER_274_1099 ();
 b15zdnd11an1n04x5 FILLER_274_1107 ();
 b15zdnd11an1n04x5 FILLER_274_1117 ();
 b15zdnd00an1n02x5 FILLER_274_1121 ();
 b15zdnd00an1n01x5 FILLER_274_1123 ();
 b15zdnd11an1n04x5 FILLER_274_1127 ();
 b15zdnd11an1n64x5 FILLER_274_1134 ();
 b15zdnd11an1n64x5 FILLER_274_1198 ();
 b15zdnd11an1n64x5 FILLER_274_1262 ();
 b15zdnd11an1n64x5 FILLER_274_1326 ();
 b15zdnd11an1n64x5 FILLER_274_1390 ();
 b15zdnd11an1n64x5 FILLER_274_1454 ();
 b15zdnd11an1n64x5 FILLER_274_1518 ();
 b15zdnd11an1n64x5 FILLER_274_1582 ();
 b15zdnd11an1n64x5 FILLER_274_1646 ();
 b15zdnd11an1n64x5 FILLER_274_1710 ();
 b15zdnd11an1n64x5 FILLER_274_1774 ();
 b15zdnd11an1n64x5 FILLER_274_1838 ();
 b15zdnd11an1n64x5 FILLER_274_1902 ();
 b15zdnd11an1n64x5 FILLER_274_1966 ();
 b15zdnd11an1n64x5 FILLER_274_2030 ();
 b15zdnd11an1n32x5 FILLER_274_2094 ();
 b15zdnd11an1n16x5 FILLER_274_2126 ();
 b15zdnd11an1n08x5 FILLER_274_2142 ();
 b15zdnd11an1n04x5 FILLER_274_2150 ();
 b15zdnd11an1n64x5 FILLER_274_2162 ();
 b15zdnd11an1n32x5 FILLER_274_2226 ();
 b15zdnd11an1n16x5 FILLER_274_2258 ();
 b15zdnd00an1n02x5 FILLER_274_2274 ();
 b15zdnd11an1n16x5 FILLER_275_0 ();
 b15zdnd11an1n04x5 FILLER_275_16 ();
 b15zdnd00an1n02x5 FILLER_275_20 ();
 b15zdnd11an1n16x5 FILLER_275_28 ();
 b15zdnd11an1n08x5 FILLER_275_44 ();
 b15zdnd11an1n64x5 FILLER_275_97 ();
 b15zdnd11an1n64x5 FILLER_275_161 ();
 b15zdnd11an1n64x5 FILLER_275_225 ();
 b15zdnd11an1n64x5 FILLER_275_289 ();
 b15zdnd11an1n32x5 FILLER_275_353 ();
 b15zdnd11an1n04x5 FILLER_275_385 ();
 b15zdnd00an1n02x5 FILLER_275_389 ();
 b15zdnd00an1n01x5 FILLER_275_391 ();
 b15zdnd11an1n64x5 FILLER_275_406 ();
 b15zdnd11an1n64x5 FILLER_275_470 ();
 b15zdnd11an1n64x5 FILLER_275_534 ();
 b15zdnd11an1n64x5 FILLER_275_598 ();
 b15zdnd11an1n64x5 FILLER_275_662 ();
 b15zdnd11an1n32x5 FILLER_275_726 ();
 b15zdnd11an1n08x5 FILLER_275_758 ();
 b15zdnd11an1n04x5 FILLER_275_766 ();
 b15zdnd00an1n02x5 FILLER_275_770 ();
 b15zdnd00an1n01x5 FILLER_275_772 ();
 b15zdnd11an1n64x5 FILLER_275_801 ();
 b15zdnd11an1n32x5 FILLER_275_865 ();
 b15zdnd11an1n04x5 FILLER_275_897 ();
 b15zdnd00an1n01x5 FILLER_275_901 ();
 b15zdnd11an1n04x5 FILLER_275_905 ();
 b15zdnd11an1n04x5 FILLER_275_915 ();
 b15zdnd00an1n01x5 FILLER_275_919 ();
 b15zdnd11an1n04x5 FILLER_275_927 ();
 b15zdnd11an1n64x5 FILLER_275_983 ();
 b15zdnd11an1n16x5 FILLER_275_1047 ();
 b15zdnd11an1n08x5 FILLER_275_1063 ();
 b15zdnd11an1n04x5 FILLER_275_1071 ();
 b15zdnd00an1n01x5 FILLER_275_1075 ();
 b15zdnd11an1n16x5 FILLER_275_1080 ();
 b15zdnd11an1n08x5 FILLER_275_1096 ();
 b15zdnd11an1n16x5 FILLER_275_1156 ();
 b15zdnd11an1n04x5 FILLER_275_1172 ();
 b15zdnd11an1n64x5 FILLER_275_1193 ();
 b15zdnd11an1n64x5 FILLER_275_1257 ();
 b15zdnd11an1n64x5 FILLER_275_1321 ();
 b15zdnd11an1n64x5 FILLER_275_1385 ();
 b15zdnd11an1n64x5 FILLER_275_1449 ();
 b15zdnd11an1n64x5 FILLER_275_1513 ();
 b15zdnd11an1n64x5 FILLER_275_1577 ();
 b15zdnd11an1n32x5 FILLER_275_1641 ();
 b15zdnd11an1n16x5 FILLER_275_1673 ();
 b15zdnd11an1n08x5 FILLER_275_1689 ();
 b15zdnd11an1n04x5 FILLER_275_1697 ();
 b15zdnd11an1n04x5 FILLER_275_1705 ();
 b15zdnd00an1n02x5 FILLER_275_1709 ();
 b15zdnd11an1n64x5 FILLER_275_1715 ();
 b15zdnd11an1n64x5 FILLER_275_1779 ();
 b15zdnd11an1n64x5 FILLER_275_1843 ();
 b15zdnd11an1n64x5 FILLER_275_1907 ();
 b15zdnd00an1n02x5 FILLER_275_1971 ();
 b15zdnd11an1n32x5 FILLER_275_2015 ();
 b15zdnd11an1n16x5 FILLER_275_2047 ();
 b15zdnd00an1n02x5 FILLER_275_2063 ();
 b15zdnd00an1n01x5 FILLER_275_2065 ();
 b15zdnd11an1n64x5 FILLER_275_2108 ();
 b15zdnd11an1n64x5 FILLER_275_2172 ();
 b15zdnd11an1n32x5 FILLER_275_2236 ();
 b15zdnd11an1n16x5 FILLER_275_2268 ();
 b15zdnd11an1n64x5 FILLER_276_8 ();
 b15zdnd11an1n04x5 FILLER_276_72 ();
 b15zdnd00an1n01x5 FILLER_276_76 ();
 b15zdnd11an1n16x5 FILLER_276_92 ();
 b15zdnd11an1n08x5 FILLER_276_108 ();
 b15zdnd11an1n04x5 FILLER_276_116 ();
 b15zdnd00an1n02x5 FILLER_276_120 ();
 b15zdnd00an1n01x5 FILLER_276_122 ();
 b15zdnd11an1n64x5 FILLER_276_148 ();
 b15zdnd11an1n64x5 FILLER_276_212 ();
 b15zdnd11an1n64x5 FILLER_276_276 ();
 b15zdnd11an1n16x5 FILLER_276_340 ();
 b15zdnd11an1n08x5 FILLER_276_356 ();
 b15zdnd11an1n04x5 FILLER_276_364 ();
 b15zdnd00an1n01x5 FILLER_276_368 ();
 b15zdnd11an1n64x5 FILLER_276_414 ();
 b15zdnd11an1n64x5 FILLER_276_478 ();
 b15zdnd11an1n64x5 FILLER_276_542 ();
 b15zdnd11an1n64x5 FILLER_276_606 ();
 b15zdnd11an1n32x5 FILLER_276_670 ();
 b15zdnd11an1n16x5 FILLER_276_702 ();
 b15zdnd11an1n64x5 FILLER_276_726 ();
 b15zdnd11an1n08x5 FILLER_276_790 ();
 b15zdnd11an1n64x5 FILLER_276_801 ();
 b15zdnd11an1n16x5 FILLER_276_865 ();
 b15zdnd11an1n04x5 FILLER_276_881 ();
 b15zdnd00an1n02x5 FILLER_276_885 ();
 b15zdnd00an1n01x5 FILLER_276_887 ();
 b15zdnd11an1n04x5 FILLER_276_915 ();
 b15zdnd00an1n02x5 FILLER_276_919 ();
 b15zdnd00an1n01x5 FILLER_276_921 ();
 b15zdnd11an1n04x5 FILLER_276_929 ();
 b15zdnd00an1n02x5 FILLER_276_933 ();
 b15zdnd00an1n01x5 FILLER_276_935 ();
 b15zdnd11an1n64x5 FILLER_276_988 ();
 b15zdnd11an1n32x5 FILLER_276_1052 ();
 b15zdnd11an1n08x5 FILLER_276_1084 ();
 b15zdnd11an1n04x5 FILLER_276_1092 ();
 b15zdnd00an1n01x5 FILLER_276_1096 ();
 b15zdnd11an1n04x5 FILLER_276_1105 ();
 b15zdnd11an1n04x5 FILLER_276_1151 ();
 b15zdnd11an1n32x5 FILLER_276_1197 ();
 b15zdnd11an1n16x5 FILLER_276_1229 ();
 b15zdnd11an1n08x5 FILLER_276_1245 ();
 b15zdnd00an1n02x5 FILLER_276_1253 ();
 b15zdnd11an1n04x5 FILLER_276_1297 ();
 b15zdnd11an1n64x5 FILLER_276_1317 ();
 b15zdnd11an1n64x5 FILLER_276_1381 ();
 b15zdnd11an1n64x5 FILLER_276_1445 ();
 b15zdnd11an1n64x5 FILLER_276_1509 ();
 b15zdnd11an1n64x5 FILLER_276_1573 ();
 b15zdnd11an1n64x5 FILLER_276_1637 ();
 b15zdnd11an1n64x5 FILLER_276_1701 ();
 b15zdnd11an1n64x5 FILLER_276_1765 ();
 b15zdnd11an1n64x5 FILLER_276_1829 ();
 b15zdnd11an1n64x5 FILLER_276_1893 ();
 b15zdnd11an1n64x5 FILLER_276_1957 ();
 b15zdnd11an1n64x5 FILLER_276_2021 ();
 b15zdnd11an1n64x5 FILLER_276_2085 ();
 b15zdnd11an1n04x5 FILLER_276_2149 ();
 b15zdnd00an1n01x5 FILLER_276_2153 ();
 b15zdnd11an1n64x5 FILLER_276_2162 ();
 b15zdnd11an1n32x5 FILLER_276_2226 ();
 b15zdnd11an1n16x5 FILLER_276_2258 ();
 b15zdnd00an1n02x5 FILLER_276_2274 ();
 b15zdnd00an1n02x5 FILLER_277_0 ();
 b15zdnd11an1n08x5 FILLER_277_10 ();
 b15zdnd11an1n04x5 FILLER_277_18 ();
 b15zdnd00an1n02x5 FILLER_277_22 ();
 b15zdnd11an1n32x5 FILLER_277_31 ();
 b15zdnd11an1n08x5 FILLER_277_63 ();
 b15zdnd11an1n64x5 FILLER_277_96 ();
 b15zdnd11an1n64x5 FILLER_277_160 ();
 b15zdnd11an1n64x5 FILLER_277_224 ();
 b15zdnd11an1n64x5 FILLER_277_288 ();
 b15zdnd00an1n02x5 FILLER_277_352 ();
 b15zdnd00an1n01x5 FILLER_277_354 ();
 b15zdnd11an1n04x5 FILLER_277_395 ();
 b15zdnd11an1n64x5 FILLER_277_403 ();
 b15zdnd11an1n64x5 FILLER_277_467 ();
 b15zdnd11an1n64x5 FILLER_277_531 ();
 b15zdnd11an1n64x5 FILLER_277_595 ();
 b15zdnd11an1n64x5 FILLER_277_659 ();
 b15zdnd11an1n64x5 FILLER_277_723 ();
 b15zdnd11an1n64x5 FILLER_277_787 ();
 b15zdnd11an1n32x5 FILLER_277_851 ();
 b15zdnd11an1n04x5 FILLER_277_883 ();
 b15zdnd00an1n02x5 FILLER_277_887 ();
 b15zdnd11an1n32x5 FILLER_277_892 ();
 b15zdnd11an1n08x5 FILLER_277_924 ();
 b15zdnd00an1n02x5 FILLER_277_932 ();
 b15zdnd11an1n04x5 FILLER_277_942 ();
 b15zdnd00an1n01x5 FILLER_277_946 ();
 b15zdnd11an1n04x5 FILLER_277_950 ();
 b15zdnd11an1n04x5 FILLER_277_957 ();
 b15zdnd11an1n64x5 FILLER_277_964 ();
 b15zdnd11an1n64x5 FILLER_277_1028 ();
 b15zdnd11an1n04x5 FILLER_277_1092 ();
 b15zdnd00an1n02x5 FILLER_277_1096 ();
 b15zdnd00an1n01x5 FILLER_277_1098 ();
 b15zdnd11an1n04x5 FILLER_277_1106 ();
 b15zdnd11an1n04x5 FILLER_277_1152 ();
 b15zdnd11an1n64x5 FILLER_277_1163 ();
 b15zdnd11an1n64x5 FILLER_277_1227 ();
 b15zdnd11an1n64x5 FILLER_277_1291 ();
 b15zdnd11an1n64x5 FILLER_277_1355 ();
 b15zdnd11an1n64x5 FILLER_277_1419 ();
 b15zdnd11an1n64x5 FILLER_277_1483 ();
 b15zdnd11an1n32x5 FILLER_277_1547 ();
 b15zdnd11an1n08x5 FILLER_277_1579 ();
 b15zdnd00an1n01x5 FILLER_277_1587 ();
 b15zdnd11an1n64x5 FILLER_277_1596 ();
 b15zdnd11an1n64x5 FILLER_277_1660 ();
 b15zdnd11an1n64x5 FILLER_277_1724 ();
 b15zdnd11an1n64x5 FILLER_277_1788 ();
 b15zdnd11an1n64x5 FILLER_277_1852 ();
 b15zdnd11an1n64x5 FILLER_277_1916 ();
 b15zdnd11an1n64x5 FILLER_277_1980 ();
 b15zdnd11an1n32x5 FILLER_277_2044 ();
 b15zdnd11an1n16x5 FILLER_277_2076 ();
 b15zdnd00an1n01x5 FILLER_277_2092 ();
 b15zdnd11an1n64x5 FILLER_277_2096 ();
 b15zdnd11an1n64x5 FILLER_277_2160 ();
 b15zdnd11an1n32x5 FILLER_277_2224 ();
 b15zdnd11an1n16x5 FILLER_277_2256 ();
 b15zdnd11an1n08x5 FILLER_277_2272 ();
 b15zdnd11an1n04x5 FILLER_277_2280 ();
 b15zdnd11an1n64x5 FILLER_278_8 ();
 b15zdnd11an1n64x5 FILLER_278_80 ();
 b15zdnd11an1n64x5 FILLER_278_144 ();
 b15zdnd11an1n64x5 FILLER_278_208 ();
 b15zdnd11an1n64x5 FILLER_278_272 ();
 b15zdnd11an1n64x5 FILLER_278_336 ();
 b15zdnd11an1n64x5 FILLER_278_400 ();
 b15zdnd11an1n64x5 FILLER_278_464 ();
 b15zdnd11an1n64x5 FILLER_278_528 ();
 b15zdnd11an1n08x5 FILLER_278_592 ();
 b15zdnd00an1n02x5 FILLER_278_600 ();
 b15zdnd00an1n01x5 FILLER_278_602 ();
 b15zdnd11an1n64x5 FILLER_278_617 ();
 b15zdnd11an1n32x5 FILLER_278_681 ();
 b15zdnd11an1n04x5 FILLER_278_713 ();
 b15zdnd00an1n01x5 FILLER_278_717 ();
 b15zdnd11an1n08x5 FILLER_278_726 ();
 b15zdnd11an1n04x5 FILLER_278_734 ();
 b15zdnd11an1n64x5 FILLER_278_747 ();
 b15zdnd11an1n64x5 FILLER_278_811 ();
 b15zdnd11an1n32x5 FILLER_278_875 ();
 b15zdnd11an1n16x5 FILLER_278_907 ();
 b15zdnd11an1n08x5 FILLER_278_923 ();
 b15zdnd00an1n01x5 FILLER_278_931 ();
 b15zdnd11an1n16x5 FILLER_278_941 ();
 b15zdnd11an1n04x5 FILLER_278_960 ();
 b15zdnd11an1n64x5 FILLER_278_967 ();
 b15zdnd11an1n64x5 FILLER_278_1031 ();
 b15zdnd00an1n01x5 FILLER_278_1095 ();
 b15zdnd11an1n08x5 FILLER_278_1116 ();
 b15zdnd00an1n02x5 FILLER_278_1124 ();
 b15zdnd00an1n01x5 FILLER_278_1126 ();
 b15zdnd11an1n32x5 FILLER_278_1130 ();
 b15zdnd11an1n16x5 FILLER_278_1162 ();
 b15zdnd11an1n08x5 FILLER_278_1178 ();
 b15zdnd11an1n04x5 FILLER_278_1186 ();
 b15zdnd00an1n01x5 FILLER_278_1190 ();
 b15zdnd11an1n64x5 FILLER_278_1199 ();
 b15zdnd11an1n32x5 FILLER_278_1263 ();
 b15zdnd11an1n64x5 FILLER_278_1307 ();
 b15zdnd11an1n64x5 FILLER_278_1371 ();
 b15zdnd11an1n64x5 FILLER_278_1435 ();
 b15zdnd11an1n64x5 FILLER_278_1499 ();
 b15zdnd11an1n64x5 FILLER_278_1563 ();
 b15zdnd11an1n64x5 FILLER_278_1627 ();
 b15zdnd11an1n64x5 FILLER_278_1691 ();
 b15zdnd11an1n64x5 FILLER_278_1755 ();
 b15zdnd11an1n64x5 FILLER_278_1819 ();
 b15zdnd11an1n64x5 FILLER_278_1883 ();
 b15zdnd11an1n64x5 FILLER_278_1947 ();
 b15zdnd11an1n32x5 FILLER_278_2011 ();
 b15zdnd11an1n16x5 FILLER_278_2043 ();
 b15zdnd00an1n02x5 FILLER_278_2059 ();
 b15zdnd11an1n04x5 FILLER_278_2101 ();
 b15zdnd11an1n32x5 FILLER_278_2108 ();
 b15zdnd11an1n08x5 FILLER_278_2140 ();
 b15zdnd11an1n04x5 FILLER_278_2148 ();
 b15zdnd00an1n02x5 FILLER_278_2152 ();
 b15zdnd11an1n32x5 FILLER_278_2162 ();
 b15zdnd11an1n04x5 FILLER_278_2194 ();
 b15zdnd00an1n02x5 FILLER_278_2198 ();
 b15zdnd11an1n04x5 FILLER_278_2203 ();
 b15zdnd11an1n64x5 FILLER_278_2210 ();
 b15zdnd00an1n02x5 FILLER_278_2274 ();
 b15zdnd11an1n64x5 FILLER_279_0 ();
 b15zdnd11an1n64x5 FILLER_279_64 ();
 b15zdnd11an1n64x5 FILLER_279_128 ();
 b15zdnd11an1n64x5 FILLER_279_192 ();
 b15zdnd11an1n64x5 FILLER_279_256 ();
 b15zdnd11an1n64x5 FILLER_279_320 ();
 b15zdnd11an1n64x5 FILLER_279_384 ();
 b15zdnd11an1n08x5 FILLER_279_448 ();
 b15zdnd11an1n04x5 FILLER_279_456 ();
 b15zdnd00an1n02x5 FILLER_279_460 ();
 b15zdnd00an1n01x5 FILLER_279_462 ();
 b15zdnd11an1n64x5 FILLER_279_515 ();
 b15zdnd11an1n64x5 FILLER_279_579 ();
 b15zdnd11an1n64x5 FILLER_279_643 ();
 b15zdnd11an1n64x5 FILLER_279_707 ();
 b15zdnd11an1n32x5 FILLER_279_771 ();
 b15zdnd11an1n16x5 FILLER_279_803 ();
 b15zdnd11an1n08x5 FILLER_279_819 ();
 b15zdnd00an1n02x5 FILLER_279_827 ();
 b15zdnd11an1n64x5 FILLER_279_871 ();
 b15zdnd11an1n64x5 FILLER_279_935 ();
 b15zdnd11an1n64x5 FILLER_279_999 ();
 b15zdnd11an1n64x5 FILLER_279_1063 ();
 b15zdnd11an1n64x5 FILLER_279_1127 ();
 b15zdnd11an1n16x5 FILLER_279_1191 ();
 b15zdnd11an1n64x5 FILLER_279_1219 ();
 b15zdnd11an1n04x5 FILLER_279_1283 ();
 b15zdnd00an1n02x5 FILLER_279_1287 ();
 b15zdnd00an1n01x5 FILLER_279_1289 ();
 b15zdnd11an1n64x5 FILLER_279_1304 ();
 b15zdnd11an1n32x5 FILLER_279_1368 ();
 b15zdnd11an1n16x5 FILLER_279_1400 ();
 b15zdnd11an1n08x5 FILLER_279_1416 ();
 b15zdnd11an1n04x5 FILLER_279_1424 ();
 b15zdnd11an1n04x5 FILLER_279_1431 ();
 b15zdnd11an1n64x5 FILLER_279_1438 ();
 b15zdnd11an1n16x5 FILLER_279_1502 ();
 b15zdnd11an1n08x5 FILLER_279_1518 ();
 b15zdnd11an1n64x5 FILLER_279_1578 ();
 b15zdnd11an1n64x5 FILLER_279_1642 ();
 b15zdnd11an1n64x5 FILLER_279_1706 ();
 b15zdnd11an1n64x5 FILLER_279_1770 ();
 b15zdnd11an1n16x5 FILLER_279_1834 ();
 b15zdnd11an1n08x5 FILLER_279_1850 ();
 b15zdnd11an1n04x5 FILLER_279_1858 ();
 b15zdnd11an1n64x5 FILLER_279_1878 ();
 b15zdnd11an1n64x5 FILLER_279_1942 ();
 b15zdnd11an1n64x5 FILLER_279_2006 ();
 b15zdnd11an1n64x5 FILLER_279_2070 ();
 b15zdnd11an1n32x5 FILLER_279_2134 ();
 b15zdnd11an1n16x5 FILLER_279_2166 ();
 b15zdnd11an1n32x5 FILLER_279_2234 ();
 b15zdnd11an1n16x5 FILLER_279_2266 ();
 b15zdnd00an1n02x5 FILLER_279_2282 ();
 b15zdnd11an1n64x5 FILLER_280_8 ();
 b15zdnd11an1n64x5 FILLER_280_72 ();
 b15zdnd11an1n64x5 FILLER_280_136 ();
 b15zdnd11an1n64x5 FILLER_280_200 ();
 b15zdnd11an1n64x5 FILLER_280_264 ();
 b15zdnd11an1n08x5 FILLER_280_328 ();
 b15zdnd00an1n02x5 FILLER_280_336 ();
 b15zdnd00an1n01x5 FILLER_280_338 ();
 b15zdnd11an1n64x5 FILLER_280_347 ();
 b15zdnd11an1n64x5 FILLER_280_411 ();
 b15zdnd11an1n08x5 FILLER_280_475 ();
 b15zdnd11an1n04x5 FILLER_280_486 ();
 b15zdnd11an1n16x5 FILLER_280_493 ();
 b15zdnd11an1n04x5 FILLER_280_509 ();
 b15zdnd11an1n64x5 FILLER_280_555 ();
 b15zdnd11an1n16x5 FILLER_280_619 ();
 b15zdnd11an1n04x5 FILLER_280_635 ();
 b15zdnd00an1n02x5 FILLER_280_639 ();
 b15zdnd00an1n01x5 FILLER_280_641 ();
 b15zdnd11an1n64x5 FILLER_280_648 ();
 b15zdnd11an1n04x5 FILLER_280_712 ();
 b15zdnd00an1n02x5 FILLER_280_716 ();
 b15zdnd11an1n64x5 FILLER_280_726 ();
 b15zdnd11an1n08x5 FILLER_280_790 ();
 b15zdnd11an1n04x5 FILLER_280_798 ();
 b15zdnd11an1n64x5 FILLER_280_817 ();
 b15zdnd11an1n64x5 FILLER_280_881 ();
 b15zdnd11an1n64x5 FILLER_280_945 ();
 b15zdnd11an1n64x5 FILLER_280_1009 ();
 b15zdnd11an1n64x5 FILLER_280_1073 ();
 b15zdnd11an1n64x5 FILLER_280_1137 ();
 b15zdnd00an1n01x5 FILLER_280_1201 ();
 b15zdnd11an1n64x5 FILLER_280_1216 ();
 b15zdnd11an1n64x5 FILLER_280_1287 ();
 b15zdnd11an1n32x5 FILLER_280_1351 ();
 b15zdnd11an1n08x5 FILLER_280_1383 ();
 b15zdnd00an1n01x5 FILLER_280_1391 ();
 b15zdnd11an1n08x5 FILLER_280_1396 ();
 b15zdnd11an1n04x5 FILLER_280_1404 ();
 b15zdnd00an1n02x5 FILLER_280_1408 ();
 b15zdnd11an1n64x5 FILLER_280_1462 ();
 b15zdnd11an1n04x5 FILLER_280_1526 ();
 b15zdnd00an1n02x5 FILLER_280_1530 ();
 b15zdnd11an1n64x5 FILLER_280_1584 ();
 b15zdnd11an1n64x5 FILLER_280_1648 ();
 b15zdnd11an1n64x5 FILLER_280_1712 ();
 b15zdnd11an1n64x5 FILLER_280_1776 ();
 b15zdnd11an1n64x5 FILLER_280_1840 ();
 b15zdnd11an1n64x5 FILLER_280_1904 ();
 b15zdnd11an1n64x5 FILLER_280_1968 ();
 b15zdnd11an1n64x5 FILLER_280_2032 ();
 b15zdnd11an1n32x5 FILLER_280_2096 ();
 b15zdnd11an1n16x5 FILLER_280_2128 ();
 b15zdnd11an1n08x5 FILLER_280_2144 ();
 b15zdnd00an1n02x5 FILLER_280_2152 ();
 b15zdnd11an1n32x5 FILLER_280_2162 ();
 b15zdnd11an1n04x5 FILLER_280_2194 ();
 b15zdnd11an1n32x5 FILLER_280_2240 ();
 b15zdnd11an1n04x5 FILLER_280_2272 ();
 b15zdnd11an1n64x5 FILLER_281_0 ();
 b15zdnd11an1n64x5 FILLER_281_64 ();
 b15zdnd11an1n64x5 FILLER_281_128 ();
 b15zdnd11an1n64x5 FILLER_281_192 ();
 b15zdnd11an1n04x5 FILLER_281_256 ();
 b15zdnd00an1n02x5 FILLER_281_260 ();
 b15zdnd00an1n01x5 FILLER_281_262 ();
 b15zdnd11an1n64x5 FILLER_281_281 ();
 b15zdnd11an1n64x5 FILLER_281_345 ();
 b15zdnd11an1n64x5 FILLER_281_409 ();
 b15zdnd11an1n08x5 FILLER_281_473 ();
 b15zdnd00an1n02x5 FILLER_281_481 ();
 b15zdnd00an1n01x5 FILLER_281_483 ();
 b15zdnd11an1n16x5 FILLER_281_487 ();
 b15zdnd11an1n04x5 FILLER_281_503 ();
 b15zdnd00an1n02x5 FILLER_281_507 ();
 b15zdnd11an1n64x5 FILLER_281_540 ();
 b15zdnd11an1n64x5 FILLER_281_604 ();
 b15zdnd11an1n64x5 FILLER_281_668 ();
 b15zdnd11an1n64x5 FILLER_281_732 ();
 b15zdnd11an1n16x5 FILLER_281_796 ();
 b15zdnd00an1n02x5 FILLER_281_812 ();
 b15zdnd11an1n64x5 FILLER_281_822 ();
 b15zdnd11an1n64x5 FILLER_281_886 ();
 b15zdnd11an1n64x5 FILLER_281_950 ();
 b15zdnd11an1n64x5 FILLER_281_1014 ();
 b15zdnd11an1n08x5 FILLER_281_1078 ();
 b15zdnd11an1n04x5 FILLER_281_1086 ();
 b15zdnd11an1n64x5 FILLER_281_1114 ();
 b15zdnd11an1n32x5 FILLER_281_1178 ();
 b15zdnd11an1n16x5 FILLER_281_1210 ();
 b15zdnd00an1n01x5 FILLER_281_1226 ();
 b15zdnd11an1n64x5 FILLER_281_1243 ();
 b15zdnd11an1n32x5 FILLER_281_1307 ();
 b15zdnd11an1n16x5 FILLER_281_1339 ();
 b15zdnd11an1n32x5 FILLER_281_1363 ();
 b15zdnd11an1n08x5 FILLER_281_1395 ();
 b15zdnd11an1n04x5 FILLER_281_1403 ();
 b15zdnd00an1n01x5 FILLER_281_1407 ();
 b15zdnd11an1n04x5 FILLER_281_1460 ();
 b15zdnd11an1n64x5 FILLER_281_1472 ();
 b15zdnd11an1n08x5 FILLER_281_1536 ();
 b15zdnd11an1n04x5 FILLER_281_1547 ();
 b15zdnd11an1n04x5 FILLER_281_1554 ();
 b15zdnd11an1n04x5 FILLER_281_1561 ();
 b15zdnd00an1n01x5 FILLER_281_1565 ();
 b15zdnd11an1n64x5 FILLER_281_1580 ();
 b15zdnd11an1n64x5 FILLER_281_1644 ();
 b15zdnd11an1n64x5 FILLER_281_1708 ();
 b15zdnd11an1n08x5 FILLER_281_1772 ();
 b15zdnd00an1n01x5 FILLER_281_1780 ();
 b15zdnd11an1n64x5 FILLER_281_1785 ();
 b15zdnd11an1n16x5 FILLER_281_1849 ();
 b15zdnd11an1n08x5 FILLER_281_1865 ();
 b15zdnd11an1n04x5 FILLER_281_1873 ();
 b15zdnd00an1n02x5 FILLER_281_1877 ();
 b15zdnd11an1n64x5 FILLER_281_1895 ();
 b15zdnd11an1n64x5 FILLER_281_1959 ();
 b15zdnd11an1n64x5 FILLER_281_2023 ();
 b15zdnd00an1n01x5 FILLER_281_2087 ();
 b15zdnd11an1n64x5 FILLER_281_2097 ();
 b15zdnd11an1n32x5 FILLER_281_2161 ();
 b15zdnd11an1n08x5 FILLER_281_2193 ();
 b15zdnd11an1n04x5 FILLER_281_2201 ();
 b15zdnd00an1n02x5 FILLER_281_2205 ();
 b15zdnd00an1n01x5 FILLER_281_2207 ();
 b15zdnd11an1n64x5 FILLER_281_2211 ();
 b15zdnd11an1n08x5 FILLER_281_2275 ();
 b15zdnd00an1n01x5 FILLER_281_2283 ();
 b15zdnd11an1n16x5 FILLER_282_8 ();
 b15zdnd00an1n01x5 FILLER_282_24 ();
 b15zdnd11an1n64x5 FILLER_282_31 ();
 b15zdnd11an1n64x5 FILLER_282_95 ();
 b15zdnd11an1n64x5 FILLER_282_159 ();
 b15zdnd11an1n16x5 FILLER_282_223 ();
 b15zdnd11an1n08x5 FILLER_282_239 ();
 b15zdnd11an1n64x5 FILLER_282_265 ();
 b15zdnd00an1n01x5 FILLER_282_329 ();
 b15zdnd11an1n64x5 FILLER_282_340 ();
 b15zdnd11an1n64x5 FILLER_282_404 ();
 b15zdnd11an1n64x5 FILLER_282_468 ();
 b15zdnd11an1n64x5 FILLER_282_532 ();
 b15zdnd11an1n64x5 FILLER_282_596 ();
 b15zdnd11an1n32x5 FILLER_282_660 ();
 b15zdnd11an1n16x5 FILLER_282_692 ();
 b15zdnd11an1n08x5 FILLER_282_708 ();
 b15zdnd00an1n02x5 FILLER_282_716 ();
 b15zdnd11an1n64x5 FILLER_282_726 ();
 b15zdnd11an1n64x5 FILLER_282_790 ();
 b15zdnd11an1n64x5 FILLER_282_854 ();
 b15zdnd11an1n64x5 FILLER_282_918 ();
 b15zdnd11an1n64x5 FILLER_282_982 ();
 b15zdnd11an1n32x5 FILLER_282_1046 ();
 b15zdnd11an1n16x5 FILLER_282_1078 ();
 b15zdnd11an1n08x5 FILLER_282_1094 ();
 b15zdnd11an1n04x5 FILLER_282_1102 ();
 b15zdnd00an1n01x5 FILLER_282_1106 ();
 b15zdnd11an1n64x5 FILLER_282_1124 ();
 b15zdnd11an1n64x5 FILLER_282_1188 ();
 b15zdnd11an1n64x5 FILLER_282_1252 ();
 b15zdnd11an1n64x5 FILLER_282_1316 ();
 b15zdnd11an1n32x5 FILLER_282_1380 ();
 b15zdnd11an1n08x5 FILLER_282_1412 ();
 b15zdnd11an1n04x5 FILLER_282_1420 ();
 b15zdnd00an1n02x5 FILLER_282_1424 ();
 b15zdnd11an1n04x5 FILLER_282_1429 ();
 b15zdnd11an1n04x5 FILLER_282_1436 ();
 b15zdnd11an1n64x5 FILLER_282_1443 ();
 b15zdnd11an1n32x5 FILLER_282_1507 ();
 b15zdnd11an1n08x5 FILLER_282_1539 ();
 b15zdnd00an1n02x5 FILLER_282_1547 ();
 b15zdnd00an1n01x5 FILLER_282_1549 ();
 b15zdnd11an1n04x5 FILLER_282_1553 ();
 b15zdnd11an1n64x5 FILLER_282_1560 ();
 b15zdnd11an1n64x5 FILLER_282_1624 ();
 b15zdnd11an1n64x5 FILLER_282_1688 ();
 b15zdnd11an1n64x5 FILLER_282_1752 ();
 b15zdnd11an1n64x5 FILLER_282_1816 ();
 b15zdnd11an1n64x5 FILLER_282_1880 ();
 b15zdnd11an1n64x5 FILLER_282_1944 ();
 b15zdnd11an1n64x5 FILLER_282_2008 ();
 b15zdnd11an1n64x5 FILLER_282_2072 ();
 b15zdnd11an1n16x5 FILLER_282_2136 ();
 b15zdnd00an1n02x5 FILLER_282_2152 ();
 b15zdnd11an1n64x5 FILLER_282_2162 ();
 b15zdnd11an1n32x5 FILLER_282_2226 ();
 b15zdnd11an1n16x5 FILLER_282_2258 ();
 b15zdnd00an1n02x5 FILLER_282_2274 ();
 b15zdnd11an1n32x5 FILLER_283_0 ();
 b15zdnd11an1n08x5 FILLER_283_38 ();
 b15zdnd11an1n04x5 FILLER_283_46 ();
 b15zdnd00an1n01x5 FILLER_283_50 ();
 b15zdnd11an1n04x5 FILLER_283_75 ();
 b15zdnd11an1n64x5 FILLER_283_91 ();
 b15zdnd11an1n64x5 FILLER_283_155 ();
 b15zdnd11an1n64x5 FILLER_283_219 ();
 b15zdnd11an1n32x5 FILLER_283_283 ();
 b15zdnd11an1n08x5 FILLER_283_315 ();
 b15zdnd11an1n04x5 FILLER_283_323 ();
 b15zdnd00an1n01x5 FILLER_283_327 ();
 b15zdnd11an1n64x5 FILLER_283_338 ();
 b15zdnd11an1n64x5 FILLER_283_402 ();
 b15zdnd11an1n64x5 FILLER_283_466 ();
 b15zdnd11an1n64x5 FILLER_283_530 ();
 b15zdnd11an1n32x5 FILLER_283_594 ();
 b15zdnd11an1n16x5 FILLER_283_626 ();
 b15zdnd11an1n08x5 FILLER_283_642 ();
 b15zdnd11an1n64x5 FILLER_283_659 ();
 b15zdnd11an1n64x5 FILLER_283_723 ();
 b15zdnd11an1n64x5 FILLER_283_787 ();
 b15zdnd11an1n64x5 FILLER_283_851 ();
 b15zdnd11an1n64x5 FILLER_283_915 ();
 b15zdnd11an1n64x5 FILLER_283_979 ();
 b15zdnd11an1n64x5 FILLER_283_1043 ();
 b15zdnd11an1n64x5 FILLER_283_1107 ();
 b15zdnd11an1n64x5 FILLER_283_1171 ();
 b15zdnd11an1n64x5 FILLER_283_1235 ();
 b15zdnd11an1n64x5 FILLER_283_1299 ();
 b15zdnd11an1n64x5 FILLER_283_1363 ();
 b15zdnd11an1n04x5 FILLER_283_1427 ();
 b15zdnd11an1n16x5 FILLER_283_1434 ();
 b15zdnd11an1n08x5 FILLER_283_1450 ();
 b15zdnd00an1n02x5 FILLER_283_1458 ();
 b15zdnd11an1n32x5 FILLER_283_1469 ();
 b15zdnd11an1n08x5 FILLER_283_1501 ();
 b15zdnd11an1n04x5 FILLER_283_1509 ();
 b15zdnd00an1n02x5 FILLER_283_1513 ();
 b15zdnd00an1n01x5 FILLER_283_1515 ();
 b15zdnd11an1n16x5 FILLER_283_1525 ();
 b15zdnd11an1n08x5 FILLER_283_1541 ();
 b15zdnd11an1n04x5 FILLER_283_1549 ();
 b15zdnd00an1n02x5 FILLER_283_1553 ();
 b15zdnd00an1n01x5 FILLER_283_1555 ();
 b15zdnd11an1n64x5 FILLER_283_1559 ();
 b15zdnd11an1n64x5 FILLER_283_1623 ();
 b15zdnd11an1n64x5 FILLER_283_1687 ();
 b15zdnd11an1n64x5 FILLER_283_1751 ();
 b15zdnd11an1n64x5 FILLER_283_1815 ();
 b15zdnd11an1n64x5 FILLER_283_1879 ();
 b15zdnd11an1n64x5 FILLER_283_1943 ();
 b15zdnd11an1n64x5 FILLER_283_2007 ();
 b15zdnd11an1n64x5 FILLER_283_2071 ();
 b15zdnd11an1n64x5 FILLER_283_2135 ();
 b15zdnd11an1n64x5 FILLER_283_2199 ();
 b15zdnd11an1n16x5 FILLER_283_2263 ();
 b15zdnd11an1n04x5 FILLER_283_2279 ();
 b15zdnd00an1n01x5 FILLER_283_2283 ();
 b15zdnd11an1n16x5 FILLER_284_8 ();
 b15zdnd11an1n16x5 FILLER_284_31 ();
 b15zdnd11an1n08x5 FILLER_284_47 ();
 b15zdnd11an1n04x5 FILLER_284_55 ();
 b15zdnd11an1n64x5 FILLER_284_92 ();
 b15zdnd11an1n64x5 FILLER_284_156 ();
 b15zdnd11an1n64x5 FILLER_284_220 ();
 b15zdnd11an1n16x5 FILLER_284_284 ();
 b15zdnd11an1n04x5 FILLER_284_300 ();
 b15zdnd11an1n64x5 FILLER_284_314 ();
 b15zdnd11an1n64x5 FILLER_284_378 ();
 b15zdnd11an1n64x5 FILLER_284_442 ();
 b15zdnd11an1n64x5 FILLER_284_506 ();
 b15zdnd11an1n64x5 FILLER_284_570 ();
 b15zdnd11an1n16x5 FILLER_284_634 ();
 b15zdnd11an1n08x5 FILLER_284_650 ();
 b15zdnd11an1n32x5 FILLER_284_661 ();
 b15zdnd11an1n16x5 FILLER_284_693 ();
 b15zdnd11an1n08x5 FILLER_284_709 ();
 b15zdnd00an1n01x5 FILLER_284_717 ();
 b15zdnd11an1n64x5 FILLER_284_726 ();
 b15zdnd11an1n64x5 FILLER_284_790 ();
 b15zdnd11an1n64x5 FILLER_284_854 ();
 b15zdnd11an1n64x5 FILLER_284_918 ();
 b15zdnd11an1n64x5 FILLER_284_982 ();
 b15zdnd11an1n64x5 FILLER_284_1046 ();
 b15zdnd11an1n64x5 FILLER_284_1110 ();
 b15zdnd11an1n64x5 FILLER_284_1174 ();
 b15zdnd11an1n64x5 FILLER_284_1238 ();
 b15zdnd11an1n64x5 FILLER_284_1302 ();
 b15zdnd11an1n64x5 FILLER_284_1366 ();
 b15zdnd11an1n64x5 FILLER_284_1430 ();
 b15zdnd11an1n64x5 FILLER_284_1494 ();
 b15zdnd11an1n64x5 FILLER_284_1558 ();
 b15zdnd11an1n64x5 FILLER_284_1622 ();
 b15zdnd11an1n64x5 FILLER_284_1686 ();
 b15zdnd11an1n64x5 FILLER_284_1750 ();
 b15zdnd11an1n32x5 FILLER_284_1814 ();
 b15zdnd11an1n16x5 FILLER_284_1846 ();
 b15zdnd11an1n08x5 FILLER_284_1862 ();
 b15zdnd00an1n01x5 FILLER_284_1870 ();
 b15zdnd11an1n04x5 FILLER_284_1877 ();
 b15zdnd00an1n01x5 FILLER_284_1881 ();
 b15zdnd11an1n04x5 FILLER_284_1888 ();
 b15zdnd11an1n04x5 FILLER_284_1905 ();
 b15zdnd11an1n32x5 FILLER_284_1923 ();
 b15zdnd11an1n16x5 FILLER_284_1955 ();
 b15zdnd00an1n02x5 FILLER_284_1971 ();
 b15zdnd11an1n64x5 FILLER_284_1978 ();
 b15zdnd11an1n64x5 FILLER_284_2042 ();
 b15zdnd11an1n32x5 FILLER_284_2106 ();
 b15zdnd11an1n16x5 FILLER_284_2138 ();
 b15zdnd11an1n64x5 FILLER_284_2162 ();
 b15zdnd11an1n04x5 FILLER_284_2226 ();
 b15zdnd00an1n02x5 FILLER_284_2230 ();
 b15zdnd00an1n02x5 FILLER_284_2274 ();
 b15zdnd11an1n32x5 FILLER_285_0 ();
 b15zdnd00an1n02x5 FILLER_285_32 ();
 b15zdnd11an1n04x5 FILLER_285_38 ();
 b15zdnd11an1n08x5 FILLER_285_48 ();
 b15zdnd11an1n04x5 FILLER_285_56 ();
 b15zdnd00an1n02x5 FILLER_285_60 ();
 b15zdnd00an1n01x5 FILLER_285_62 ();
 b15zdnd11an1n64x5 FILLER_285_94 ();
 b15zdnd11an1n64x5 FILLER_285_158 ();
 b15zdnd11an1n32x5 FILLER_285_222 ();
 b15zdnd11an1n16x5 FILLER_285_254 ();
 b15zdnd00an1n01x5 FILLER_285_270 ();
 b15zdnd11an1n16x5 FILLER_285_275 ();
 b15zdnd00an1n01x5 FILLER_285_291 ();
 b15zdnd11an1n64x5 FILLER_285_304 ();
 b15zdnd11an1n64x5 FILLER_285_368 ();
 b15zdnd11an1n64x5 FILLER_285_432 ();
 b15zdnd00an1n01x5 FILLER_285_496 ();
 b15zdnd11an1n64x5 FILLER_285_539 ();
 b15zdnd11an1n32x5 FILLER_285_603 ();
 b15zdnd11an1n08x5 FILLER_285_635 ();
 b15zdnd11an1n04x5 FILLER_285_643 ();
 b15zdnd00an1n02x5 FILLER_285_647 ();
 b15zdnd00an1n01x5 FILLER_285_649 ();
 b15zdnd11an1n04x5 FILLER_285_657 ();
 b15zdnd11an1n64x5 FILLER_285_703 ();
 b15zdnd11an1n32x5 FILLER_285_767 ();
 b15zdnd11an1n04x5 FILLER_285_799 ();
 b15zdnd11an1n64x5 FILLER_285_806 ();
 b15zdnd11an1n64x5 FILLER_285_870 ();
 b15zdnd11an1n64x5 FILLER_285_934 ();
 b15zdnd11an1n64x5 FILLER_285_998 ();
 b15zdnd11an1n64x5 FILLER_285_1062 ();
 b15zdnd11an1n08x5 FILLER_285_1126 ();
 b15zdnd11an1n04x5 FILLER_285_1134 ();
 b15zdnd00an1n01x5 FILLER_285_1138 ();
 b15zdnd11an1n64x5 FILLER_285_1151 ();
 b15zdnd11an1n64x5 FILLER_285_1215 ();
 b15zdnd11an1n64x5 FILLER_285_1279 ();
 b15zdnd11an1n64x5 FILLER_285_1343 ();
 b15zdnd11an1n64x5 FILLER_285_1407 ();
 b15zdnd11an1n64x5 FILLER_285_1471 ();
 b15zdnd11an1n64x5 FILLER_285_1535 ();
 b15zdnd11an1n64x5 FILLER_285_1599 ();
 b15zdnd11an1n64x5 FILLER_285_1663 ();
 b15zdnd11an1n64x5 FILLER_285_1727 ();
 b15zdnd11an1n64x5 FILLER_285_1791 ();
 b15zdnd11an1n08x5 FILLER_285_1855 ();
 b15zdnd11an1n04x5 FILLER_285_1863 ();
 b15zdnd11an1n08x5 FILLER_285_1881 ();
 b15zdnd00an1n02x5 FILLER_285_1889 ();
 b15zdnd11an1n04x5 FILLER_285_1894 ();
 b15zdnd11an1n64x5 FILLER_285_1901 ();
 b15zdnd11an1n64x5 FILLER_285_1965 ();
 b15zdnd11an1n64x5 FILLER_285_2029 ();
 b15zdnd11an1n64x5 FILLER_285_2093 ();
 b15zdnd11an1n32x5 FILLER_285_2157 ();
 b15zdnd11an1n16x5 FILLER_285_2189 ();
 b15zdnd11an1n04x5 FILLER_285_2205 ();
 b15zdnd00an1n01x5 FILLER_285_2209 ();
 b15zdnd11an1n04x5 FILLER_285_2213 ();
 b15zdnd11an1n16x5 FILLER_285_2220 ();
 b15zdnd11an1n04x5 FILLER_285_2236 ();
 b15zdnd00an1n02x5 FILLER_285_2282 ();
 b15zdnd00an1n02x5 FILLER_286_8 ();
 b15zdnd11an1n04x5 FILLER_286_14 ();
 b15zdnd00an1n02x5 FILLER_286_18 ();
 b15zdnd00an1n01x5 FILLER_286_20 ();
 b15zdnd11an1n64x5 FILLER_286_25 ();
 b15zdnd11an1n64x5 FILLER_286_89 ();
 b15zdnd11an1n64x5 FILLER_286_153 ();
 b15zdnd11an1n16x5 FILLER_286_217 ();
 b15zdnd00an1n02x5 FILLER_286_233 ();
 b15zdnd11an1n64x5 FILLER_286_238 ();
 b15zdnd11an1n64x5 FILLER_286_302 ();
 b15zdnd11an1n64x5 FILLER_286_366 ();
 b15zdnd11an1n64x5 FILLER_286_430 ();
 b15zdnd11an1n64x5 FILLER_286_494 ();
 b15zdnd11an1n64x5 FILLER_286_558 ();
 b15zdnd11an1n16x5 FILLER_286_622 ();
 b15zdnd11an1n08x5 FILLER_286_638 ();
 b15zdnd11an1n04x5 FILLER_286_646 ();
 b15zdnd00an1n02x5 FILLER_286_650 ();
 b15zdnd00an1n01x5 FILLER_286_652 ();
 b15zdnd11an1n04x5 FILLER_286_658 ();
 b15zdnd00an1n02x5 FILLER_286_662 ();
 b15zdnd00an1n01x5 FILLER_286_664 ();
 b15zdnd11an1n08x5 FILLER_286_707 ();
 b15zdnd00an1n02x5 FILLER_286_715 ();
 b15zdnd00an1n01x5 FILLER_286_717 ();
 b15zdnd11an1n64x5 FILLER_286_726 ();
 b15zdnd11an1n04x5 FILLER_286_790 ();
 b15zdnd00an1n02x5 FILLER_286_794 ();
 b15zdnd00an1n01x5 FILLER_286_796 ();
 b15zdnd11an1n64x5 FILLER_286_839 ();
 b15zdnd11an1n32x5 FILLER_286_903 ();
 b15zdnd11an1n08x5 FILLER_286_935 ();
 b15zdnd00an1n02x5 FILLER_286_943 ();
 b15zdnd11an1n64x5 FILLER_286_954 ();
 b15zdnd11an1n64x5 FILLER_286_1018 ();
 b15zdnd11an1n64x5 FILLER_286_1082 ();
 b15zdnd11an1n64x5 FILLER_286_1146 ();
 b15zdnd11an1n64x5 FILLER_286_1210 ();
 b15zdnd11an1n32x5 FILLER_286_1274 ();
 b15zdnd11an1n16x5 FILLER_286_1306 ();
 b15zdnd11an1n04x5 FILLER_286_1322 ();
 b15zdnd00an1n02x5 FILLER_286_1326 ();
 b15zdnd11an1n64x5 FILLER_286_1336 ();
 b15zdnd11an1n64x5 FILLER_286_1400 ();
 b15zdnd11an1n32x5 FILLER_286_1464 ();
 b15zdnd11an1n08x5 FILLER_286_1496 ();
 b15zdnd00an1n01x5 FILLER_286_1504 ();
 b15zdnd11an1n16x5 FILLER_286_1514 ();
 b15zdnd11an1n08x5 FILLER_286_1530 ();
 b15zdnd11an1n64x5 FILLER_286_1590 ();
 b15zdnd11an1n32x5 FILLER_286_1654 ();
 b15zdnd11an1n16x5 FILLER_286_1686 ();
 b15zdnd00an1n01x5 FILLER_286_1702 ();
 b15zdnd11an1n64x5 FILLER_286_1706 ();
 b15zdnd11an1n64x5 FILLER_286_1770 ();
 b15zdnd11an1n32x5 FILLER_286_1834 ();
 b15zdnd11an1n04x5 FILLER_286_1866 ();
 b15zdnd00an1n02x5 FILLER_286_1870 ();
 b15zdnd00an1n01x5 FILLER_286_1872 ();
 b15zdnd11an1n64x5 FILLER_286_1891 ();
 b15zdnd11an1n64x5 FILLER_286_1955 ();
 b15zdnd11an1n32x5 FILLER_286_2019 ();
 b15zdnd11an1n16x5 FILLER_286_2051 ();
 b15zdnd00an1n02x5 FILLER_286_2067 ();
 b15zdnd00an1n01x5 FILLER_286_2069 ();
 b15zdnd11an1n32x5 FILLER_286_2122 ();
 b15zdnd11an1n16x5 FILLER_286_2162 ();
 b15zdnd11an1n04x5 FILLER_286_2178 ();
 b15zdnd00an1n02x5 FILLER_286_2182 ();
 b15zdnd00an1n01x5 FILLER_286_2184 ();
 b15zdnd11an1n04x5 FILLER_286_2237 ();
 b15zdnd00an1n01x5 FILLER_286_2241 ();
 b15zdnd11an1n16x5 FILLER_286_2246 ();
 b15zdnd11an1n08x5 FILLER_286_2262 ();
 b15zdnd00an1n02x5 FILLER_286_2274 ();
 b15zdnd00an1n02x5 FILLER_287_0 ();
 b15zdnd11an1n64x5 FILLER_287_44 ();
 b15zdnd11an1n64x5 FILLER_287_108 ();
 b15zdnd11an1n32x5 FILLER_287_172 ();
 b15zdnd11an1n04x5 FILLER_287_204 ();
 b15zdnd00an1n01x5 FILLER_287_208 ();
 b15zdnd11an1n04x5 FILLER_287_225 ();
 b15zdnd11an1n64x5 FILLER_287_253 ();
 b15zdnd11an1n32x5 FILLER_287_317 ();
 b15zdnd11an1n08x5 FILLER_287_349 ();
 b15zdnd00an1n01x5 FILLER_287_357 ();
 b15zdnd11an1n64x5 FILLER_287_372 ();
 b15zdnd11an1n64x5 FILLER_287_436 ();
 b15zdnd11an1n64x5 FILLER_287_500 ();
 b15zdnd11an1n64x5 FILLER_287_564 ();
 b15zdnd11an1n16x5 FILLER_287_628 ();
 b15zdnd11an1n04x5 FILLER_287_644 ();
 b15zdnd11an1n04x5 FILLER_287_652 ();
 b15zdnd11an1n08x5 FILLER_287_663 ();
 b15zdnd00an1n02x5 FILLER_287_671 ();
 b15zdnd11an1n64x5 FILLER_287_725 ();
 b15zdnd11an1n16x5 FILLER_287_789 ();
 b15zdnd11an1n08x5 FILLER_287_805 ();
 b15zdnd11an1n04x5 FILLER_287_813 ();
 b15zdnd11an1n64x5 FILLER_287_825 ();
 b15zdnd11an1n32x5 FILLER_287_889 ();
 b15zdnd11an1n08x5 FILLER_287_921 ();
 b15zdnd00an1n02x5 FILLER_287_929 ();
 b15zdnd00an1n01x5 FILLER_287_931 ();
 b15zdnd11an1n64x5 FILLER_287_941 ();
 b15zdnd11an1n64x5 FILLER_287_1005 ();
 b15zdnd11an1n64x5 FILLER_287_1069 ();
 b15zdnd11an1n64x5 FILLER_287_1133 ();
 b15zdnd11an1n64x5 FILLER_287_1197 ();
 b15zdnd11an1n64x5 FILLER_287_1261 ();
 b15zdnd11an1n64x5 FILLER_287_1325 ();
 b15zdnd11an1n64x5 FILLER_287_1389 ();
 b15zdnd11an1n64x5 FILLER_287_1453 ();
 b15zdnd11an1n32x5 FILLER_287_1517 ();
 b15zdnd11an1n04x5 FILLER_287_1549 ();
 b15zdnd00an1n02x5 FILLER_287_1553 ();
 b15zdnd00an1n01x5 FILLER_287_1555 ();
 b15zdnd11an1n04x5 FILLER_287_1559 ();
 b15zdnd11an1n64x5 FILLER_287_1566 ();
 b15zdnd11an1n32x5 FILLER_287_1630 ();
 b15zdnd11an1n16x5 FILLER_287_1662 ();
 b15zdnd11an1n04x5 FILLER_287_1678 ();
 b15zdnd00an1n02x5 FILLER_287_1682 ();
 b15zdnd11an1n32x5 FILLER_287_1736 ();
 b15zdnd11an1n08x5 FILLER_287_1768 ();
 b15zdnd11an1n04x5 FILLER_287_1776 ();
 b15zdnd11an1n64x5 FILLER_287_1783 ();
 b15zdnd11an1n32x5 FILLER_287_1847 ();
 b15zdnd11an1n04x5 FILLER_287_1879 ();
 b15zdnd00an1n01x5 FILLER_287_1883 ();
 b15zdnd11an1n32x5 FILLER_287_1904 ();
 b15zdnd11an1n16x5 FILLER_287_1936 ();
 b15zdnd00an1n01x5 FILLER_287_1952 ();
 b15zdnd11an1n16x5 FILLER_287_1965 ();
 b15zdnd11an1n04x5 FILLER_287_1981 ();
 b15zdnd00an1n01x5 FILLER_287_1985 ();
 b15zdnd11an1n64x5 FILLER_287_1991 ();
 b15zdnd11an1n32x5 FILLER_287_2055 ();
 b15zdnd00an1n01x5 FILLER_287_2087 ();
 b15zdnd11an1n04x5 FILLER_287_2091 ();
 b15zdnd11an1n16x5 FILLER_287_2098 ();
 b15zdnd00an1n02x5 FILLER_287_2114 ();
 b15zdnd11an1n04x5 FILLER_287_2158 ();
 b15zdnd11an1n04x5 FILLER_287_2204 ();
 b15zdnd11an1n16x5 FILLER_287_2250 ();
 b15zdnd00an1n02x5 FILLER_287_2266 ();
 b15zdnd11an1n08x5 FILLER_287_2272 ();
 b15zdnd11an1n04x5 FILLER_287_2280 ();
 b15zdnd11an1n04x5 FILLER_288_8 ();
 b15zdnd11an1n04x5 FILLER_288_19 ();
 b15zdnd00an1n02x5 FILLER_288_23 ();
 b15zdnd00an1n01x5 FILLER_288_25 ();
 b15zdnd11an1n64x5 FILLER_288_31 ();
 b15zdnd11an1n64x5 FILLER_288_95 ();
 b15zdnd11an1n32x5 FILLER_288_159 ();
 b15zdnd11an1n16x5 FILLER_288_191 ();
 b15zdnd11an1n08x5 FILLER_288_207 ();
 b15zdnd11an1n04x5 FILLER_288_215 ();
 b15zdnd00an1n02x5 FILLER_288_219 ();
 b15zdnd00an1n01x5 FILLER_288_221 ();
 b15zdnd11an1n16x5 FILLER_288_225 ();
 b15zdnd11an1n04x5 FILLER_288_241 ();
 b15zdnd00an1n02x5 FILLER_288_245 ();
 b15zdnd11an1n64x5 FILLER_288_257 ();
 b15zdnd11an1n64x5 FILLER_288_321 ();
 b15zdnd11an1n64x5 FILLER_288_385 ();
 b15zdnd11an1n64x5 FILLER_288_449 ();
 b15zdnd11an1n64x5 FILLER_288_513 ();
 b15zdnd11an1n64x5 FILLER_288_577 ();
 b15zdnd11an1n04x5 FILLER_288_641 ();
 b15zdnd00an1n02x5 FILLER_288_645 ();
 b15zdnd00an1n01x5 FILLER_288_647 ();
 b15zdnd11an1n08x5 FILLER_288_657 ();
 b15zdnd00an1n02x5 FILLER_288_665 ();
 b15zdnd00an1n01x5 FILLER_288_667 ();
 b15zdnd11an1n08x5 FILLER_288_710 ();
 b15zdnd00an1n02x5 FILLER_288_726 ();
 b15zdnd11an1n64x5 FILLER_288_731 ();
 b15zdnd11an1n08x5 FILLER_288_795 ();
 b15zdnd00an1n01x5 FILLER_288_803 ();
 b15zdnd11an1n64x5 FILLER_288_818 ();
 b15zdnd11an1n64x5 FILLER_288_882 ();
 b15zdnd11an1n64x5 FILLER_288_946 ();
 b15zdnd11an1n64x5 FILLER_288_1010 ();
 b15zdnd11an1n64x5 FILLER_288_1074 ();
 b15zdnd11an1n64x5 FILLER_288_1138 ();
 b15zdnd11an1n16x5 FILLER_288_1202 ();
 b15zdnd11an1n04x5 FILLER_288_1218 ();
 b15zdnd00an1n01x5 FILLER_288_1222 ();
 b15zdnd11an1n04x5 FILLER_288_1236 ();
 b15zdnd11an1n64x5 FILLER_288_1243 ();
 b15zdnd11an1n64x5 FILLER_288_1307 ();
 b15zdnd11an1n64x5 FILLER_288_1371 ();
 b15zdnd11an1n64x5 FILLER_288_1435 ();
 b15zdnd11an1n64x5 FILLER_288_1499 ();
 b15zdnd00an1n01x5 FILLER_288_1563 ();
 b15zdnd11an1n64x5 FILLER_288_1567 ();
 b15zdnd11an1n32x5 FILLER_288_1631 ();
 b15zdnd11an1n16x5 FILLER_288_1663 ();
 b15zdnd00an1n01x5 FILLER_288_1679 ();
 b15zdnd11an1n04x5 FILLER_288_1732 ();
 b15zdnd00an1n02x5 FILLER_288_1736 ();
 b15zdnd11an1n32x5 FILLER_288_1746 ();
 b15zdnd00an1n02x5 FILLER_288_1778 ();
 b15zdnd11an1n64x5 FILLER_288_1783 ();
 b15zdnd11an1n64x5 FILLER_288_1847 ();
 b15zdnd11an1n64x5 FILLER_288_1911 ();
 b15zdnd11an1n64x5 FILLER_288_1975 ();
 b15zdnd11an1n32x5 FILLER_288_2039 ();
 b15zdnd11an1n16x5 FILLER_288_2071 ();
 b15zdnd11an1n08x5 FILLER_288_2087 ();
 b15zdnd11an1n32x5 FILLER_288_2098 ();
 b15zdnd11an1n16x5 FILLER_288_2130 ();
 b15zdnd11an1n08x5 FILLER_288_2146 ();
 b15zdnd00an1n02x5 FILLER_288_2162 ();
 b15zdnd11an1n04x5 FILLER_288_2206 ();
 b15zdnd11an1n04x5 FILLER_288_2213 ();
 b15zdnd00an1n01x5 FILLER_288_2217 ();
 b15zdnd11an1n04x5 FILLER_288_2260 ();
 b15zdnd11an1n08x5 FILLER_288_2268 ();
 b15zdnd11an1n08x5 FILLER_289_0 ();
 b15zdnd00an1n01x5 FILLER_289_8 ();
 b15zdnd11an1n64x5 FILLER_289_15 ();
 b15zdnd11an1n64x5 FILLER_289_79 ();
 b15zdnd11an1n16x5 FILLER_289_143 ();
 b15zdnd11an1n08x5 FILLER_289_159 ();
 b15zdnd00an1n02x5 FILLER_289_167 ();
 b15zdnd00an1n01x5 FILLER_289_169 ();
 b15zdnd11an1n32x5 FILLER_289_185 ();
 b15zdnd11an1n08x5 FILLER_289_217 ();
 b15zdnd11an1n04x5 FILLER_289_225 ();
 b15zdnd00an1n02x5 FILLER_289_229 ();
 b15zdnd00an1n01x5 FILLER_289_231 ();
 b15zdnd11an1n64x5 FILLER_289_250 ();
 b15zdnd11an1n32x5 FILLER_289_314 ();
 b15zdnd11an1n16x5 FILLER_289_346 ();
 b15zdnd11an1n04x5 FILLER_289_362 ();
 b15zdnd00an1n01x5 FILLER_289_366 ();
 b15zdnd11an1n64x5 FILLER_289_378 ();
 b15zdnd11an1n64x5 FILLER_289_442 ();
 b15zdnd11an1n32x5 FILLER_289_506 ();
 b15zdnd11an1n16x5 FILLER_289_538 ();
 b15zdnd11an1n08x5 FILLER_289_554 ();
 b15zdnd00an1n01x5 FILLER_289_562 ();
 b15zdnd11an1n64x5 FILLER_289_570 ();
 b15zdnd11an1n16x5 FILLER_289_634 ();
 b15zdnd00an1n01x5 FILLER_289_650 ();
 b15zdnd11an1n04x5 FILLER_289_656 ();
 b15zdnd00an1n01x5 FILLER_289_660 ();
 b15zdnd11an1n08x5 FILLER_289_666 ();
 b15zdnd11an1n04x5 FILLER_289_674 ();
 b15zdnd00an1n02x5 FILLER_289_678 ();
 b15zdnd11an1n04x5 FILLER_289_683 ();
 b15zdnd11an1n04x5 FILLER_289_690 ();
 b15zdnd11an1n64x5 FILLER_289_736 ();
 b15zdnd11an1n64x5 FILLER_289_800 ();
 b15zdnd11an1n64x5 FILLER_289_864 ();
 b15zdnd11an1n64x5 FILLER_289_928 ();
 b15zdnd11an1n32x5 FILLER_289_992 ();
 b15zdnd11an1n16x5 FILLER_289_1024 ();
 b15zdnd00an1n01x5 FILLER_289_1040 ();
 b15zdnd11an1n64x5 FILLER_289_1047 ();
 b15zdnd11an1n64x5 FILLER_289_1111 ();
 b15zdnd11an1n32x5 FILLER_289_1175 ();
 b15zdnd11an1n16x5 FILLER_289_1207 ();
 b15zdnd11an1n04x5 FILLER_289_1223 ();
 b15zdnd00an1n01x5 FILLER_289_1227 ();
 b15zdnd11an1n64x5 FILLER_289_1242 ();
 b15zdnd11an1n64x5 FILLER_289_1306 ();
 b15zdnd11an1n32x5 FILLER_289_1370 ();
 b15zdnd11an1n08x5 FILLER_289_1402 ();
 b15zdnd11an1n04x5 FILLER_289_1410 ();
 b15zdnd00an1n02x5 FILLER_289_1414 ();
 b15zdnd00an1n01x5 FILLER_289_1416 ();
 b15zdnd11an1n64x5 FILLER_289_1444 ();
 b15zdnd11an1n64x5 FILLER_289_1508 ();
 b15zdnd11an1n64x5 FILLER_289_1572 ();
 b15zdnd11an1n32x5 FILLER_289_1636 ();
 b15zdnd11an1n16x5 FILLER_289_1668 ();
 b15zdnd11an1n16x5 FILLER_289_1736 ();
 b15zdnd00an1n02x5 FILLER_289_1752 ();
 b15zdnd00an1n01x5 FILLER_289_1754 ();
 b15zdnd11an1n64x5 FILLER_289_1807 ();
 b15zdnd11an1n32x5 FILLER_289_1871 ();
 b15zdnd11an1n16x5 FILLER_289_1903 ();
 b15zdnd00an1n01x5 FILLER_289_1919 ();
 b15zdnd11an1n64x5 FILLER_289_1934 ();
 b15zdnd11an1n64x5 FILLER_289_1998 ();
 b15zdnd11an1n64x5 FILLER_289_2062 ();
 b15zdnd11an1n64x5 FILLER_289_2126 ();
 b15zdnd11an1n16x5 FILLER_289_2190 ();
 b15zdnd11an1n08x5 FILLER_289_2206 ();
 b15zdnd00an1n02x5 FILLER_289_2214 ();
 b15zdnd00an1n01x5 FILLER_289_2216 ();
 b15zdnd11an1n04x5 FILLER_289_2225 ();
 b15zdnd11an1n08x5 FILLER_289_2271 ();
 b15zdnd11an1n04x5 FILLER_289_2279 ();
 b15zdnd00an1n01x5 FILLER_289_2283 ();
 b15zdnd11an1n08x5 FILLER_290_8 ();
 b15zdnd11an1n04x5 FILLER_290_16 ();
 b15zdnd00an1n02x5 FILLER_290_20 ();
 b15zdnd11an1n64x5 FILLER_290_28 ();
 b15zdnd11an1n64x5 FILLER_290_92 ();
 b15zdnd11an1n16x5 FILLER_290_156 ();
 b15zdnd11an1n04x5 FILLER_290_172 ();
 b15zdnd11an1n64x5 FILLER_290_194 ();
 b15zdnd11an1n64x5 FILLER_290_258 ();
 b15zdnd11an1n64x5 FILLER_290_322 ();
 b15zdnd11an1n64x5 FILLER_290_386 ();
 b15zdnd11an1n32x5 FILLER_290_450 ();
 b15zdnd11an1n16x5 FILLER_290_482 ();
 b15zdnd11an1n08x5 FILLER_290_498 ();
 b15zdnd00an1n02x5 FILLER_290_506 ();
 b15zdnd00an1n01x5 FILLER_290_508 ();
 b15zdnd11an1n64x5 FILLER_290_516 ();
 b15zdnd11an1n32x5 FILLER_290_580 ();
 b15zdnd11an1n16x5 FILLER_290_612 ();
 b15zdnd11an1n08x5 FILLER_290_628 ();
 b15zdnd00an1n02x5 FILLER_290_636 ();
 b15zdnd11an1n08x5 FILLER_290_643 ();
 b15zdnd11an1n04x5 FILLER_290_651 ();
 b15zdnd00an1n01x5 FILLER_290_655 ();
 b15zdnd11an1n04x5 FILLER_290_660 ();
 b15zdnd11an1n08x5 FILLER_290_706 ();
 b15zdnd11an1n04x5 FILLER_290_714 ();
 b15zdnd11an1n64x5 FILLER_290_726 ();
 b15zdnd11an1n16x5 FILLER_290_790 ();
 b15zdnd00an1n01x5 FILLER_290_806 ();
 b15zdnd11an1n64x5 FILLER_290_810 ();
 b15zdnd11an1n64x5 FILLER_290_874 ();
 b15zdnd11an1n64x5 FILLER_290_938 ();
 b15zdnd11an1n64x5 FILLER_290_1002 ();
 b15zdnd11an1n64x5 FILLER_290_1066 ();
 b15zdnd11an1n64x5 FILLER_290_1130 ();
 b15zdnd11an1n32x5 FILLER_290_1194 ();
 b15zdnd00an1n02x5 FILLER_290_1226 ();
 b15zdnd11an1n08x5 FILLER_290_1231 ();
 b15zdnd11an1n64x5 FILLER_290_1254 ();
 b15zdnd11an1n64x5 FILLER_290_1318 ();
 b15zdnd11an1n32x5 FILLER_290_1382 ();
 b15zdnd11an1n04x5 FILLER_290_1414 ();
 b15zdnd00an1n02x5 FILLER_290_1418 ();
 b15zdnd00an1n01x5 FILLER_290_1420 ();
 b15zdnd11an1n64x5 FILLER_290_1424 ();
 b15zdnd11an1n64x5 FILLER_290_1488 ();
 b15zdnd00an1n02x5 FILLER_290_1552 ();
 b15zdnd00an1n01x5 FILLER_290_1554 ();
 b15zdnd11an1n64x5 FILLER_290_1559 ();
 b15zdnd11an1n64x5 FILLER_290_1623 ();
 b15zdnd11an1n08x5 FILLER_290_1687 ();
 b15zdnd11an1n04x5 FILLER_290_1695 ();
 b15zdnd00an1n01x5 FILLER_290_1699 ();
 b15zdnd11an1n04x5 FILLER_290_1703 ();
 b15zdnd11an1n04x5 FILLER_290_1710 ();
 b15zdnd11an1n04x5 FILLER_290_1717 ();
 b15zdnd11an1n04x5 FILLER_290_1724 ();
 b15zdnd11an1n32x5 FILLER_290_1731 ();
 b15zdnd11an1n16x5 FILLER_290_1763 ();
 b15zdnd00an1n02x5 FILLER_290_1779 ();
 b15zdnd11an1n04x5 FILLER_290_1784 ();
 b15zdnd11an1n64x5 FILLER_290_1791 ();
 b15zdnd11an1n32x5 FILLER_290_1855 ();
 b15zdnd11an1n16x5 FILLER_290_1887 ();
 b15zdnd00an1n02x5 FILLER_290_1903 ();
 b15zdnd11an1n04x5 FILLER_290_1919 ();
 b15zdnd11an1n08x5 FILLER_290_1926 ();
 b15zdnd00an1n02x5 FILLER_290_1934 ();
 b15zdnd11an1n64x5 FILLER_290_1956 ();
 b15zdnd11an1n64x5 FILLER_290_2020 ();
 b15zdnd11an1n64x5 FILLER_290_2084 ();
 b15zdnd11an1n04x5 FILLER_290_2148 ();
 b15zdnd00an1n02x5 FILLER_290_2152 ();
 b15zdnd11an1n64x5 FILLER_290_2162 ();
 b15zdnd11an1n04x5 FILLER_290_2226 ();
 b15zdnd00an1n02x5 FILLER_290_2230 ();
 b15zdnd00an1n02x5 FILLER_290_2274 ();
 b15zdnd11an1n64x5 FILLER_291_0 ();
 b15zdnd11an1n32x5 FILLER_291_64 ();
 b15zdnd11an1n16x5 FILLER_291_96 ();
 b15zdnd11an1n08x5 FILLER_291_112 ();
 b15zdnd11an1n04x5 FILLER_291_120 ();
 b15zdnd00an1n01x5 FILLER_291_124 ();
 b15zdnd11an1n64x5 FILLER_291_150 ();
 b15zdnd11an1n64x5 FILLER_291_214 ();
 b15zdnd11an1n64x5 FILLER_291_278 ();
 b15zdnd11an1n64x5 FILLER_291_342 ();
 b15zdnd11an1n64x5 FILLER_291_406 ();
 b15zdnd11an1n32x5 FILLER_291_470 ();
 b15zdnd11an1n08x5 FILLER_291_502 ();
 b15zdnd11an1n04x5 FILLER_291_510 ();
 b15zdnd11an1n64x5 FILLER_291_517 ();
 b15zdnd11an1n64x5 FILLER_291_581 ();
 b15zdnd11an1n08x5 FILLER_291_645 ();
 b15zdnd11an1n08x5 FILLER_291_656 ();
 b15zdnd00an1n02x5 FILLER_291_664 ();
 b15zdnd00an1n01x5 FILLER_291_666 ();
 b15zdnd11an1n32x5 FILLER_291_709 ();
 b15zdnd11an1n16x5 FILLER_291_741 ();
 b15zdnd11an1n08x5 FILLER_291_757 ();
 b15zdnd11an1n04x5 FILLER_291_765 ();
 b15zdnd00an1n02x5 FILLER_291_769 ();
 b15zdnd11an1n04x5 FILLER_291_811 ();
 b15zdnd11an1n64x5 FILLER_291_818 ();
 b15zdnd11an1n64x5 FILLER_291_882 ();
 b15zdnd11an1n64x5 FILLER_291_946 ();
 b15zdnd11an1n64x5 FILLER_291_1010 ();
 b15zdnd11an1n64x5 FILLER_291_1074 ();
 b15zdnd11an1n64x5 FILLER_291_1138 ();
 b15zdnd11an1n64x5 FILLER_291_1202 ();
 b15zdnd11an1n64x5 FILLER_291_1266 ();
 b15zdnd11an1n64x5 FILLER_291_1330 ();
 b15zdnd11an1n16x5 FILLER_291_1394 ();
 b15zdnd11an1n04x5 FILLER_291_1410 ();
 b15zdnd00an1n02x5 FILLER_291_1414 ();
 b15zdnd11an1n64x5 FILLER_291_1468 ();
 b15zdnd11an1n16x5 FILLER_291_1532 ();
 b15zdnd11an1n08x5 FILLER_291_1548 ();
 b15zdnd00an1n01x5 FILLER_291_1556 ();
 b15zdnd11an1n04x5 FILLER_291_1560 ();
 b15zdnd11an1n64x5 FILLER_291_1567 ();
 b15zdnd11an1n64x5 FILLER_291_1631 ();
 b15zdnd11an1n04x5 FILLER_291_1695 ();
 b15zdnd00an1n02x5 FILLER_291_1699 ();
 b15zdnd00an1n01x5 FILLER_291_1701 ();
 b15zdnd11an1n04x5 FILLER_291_1705 ();
 b15zdnd11an1n04x5 FILLER_291_1712 ();
 b15zdnd11an1n32x5 FILLER_291_1719 ();
 b15zdnd11an1n08x5 FILLER_291_1751 ();
 b15zdnd00an1n02x5 FILLER_291_1759 ();
 b15zdnd00an1n01x5 FILLER_291_1761 ();
 b15zdnd11an1n64x5 FILLER_291_1814 ();
 b15zdnd11an1n32x5 FILLER_291_1878 ();
 b15zdnd00an1n02x5 FILLER_291_1910 ();
 b15zdnd11an1n04x5 FILLER_291_1926 ();
 b15zdnd11an1n64x5 FILLER_291_1933 ();
 b15zdnd11an1n64x5 FILLER_291_1997 ();
 b15zdnd11an1n16x5 FILLER_291_2061 ();
 b15zdnd11an1n08x5 FILLER_291_2077 ();
 b15zdnd00an1n02x5 FILLER_291_2085 ();
 b15zdnd00an1n01x5 FILLER_291_2087 ();
 b15zdnd11an1n64x5 FILLER_291_2091 ();
 b15zdnd11an1n64x5 FILLER_291_2155 ();
 b15zdnd11an1n64x5 FILLER_291_2219 ();
 b15zdnd00an1n01x5 FILLER_291_2283 ();
 b15zdnd11an1n32x5 FILLER_292_8 ();
 b15zdnd11an1n08x5 FILLER_292_40 ();
 b15zdnd11an1n64x5 FILLER_292_90 ();
 b15zdnd11an1n64x5 FILLER_292_154 ();
 b15zdnd11an1n64x5 FILLER_292_218 ();
 b15zdnd11an1n64x5 FILLER_292_282 ();
 b15zdnd11an1n64x5 FILLER_292_346 ();
 b15zdnd11an1n64x5 FILLER_292_410 ();
 b15zdnd11an1n32x5 FILLER_292_474 ();
 b15zdnd11an1n04x5 FILLER_292_506 ();
 b15zdnd11an1n64x5 FILLER_292_515 ();
 b15zdnd11an1n64x5 FILLER_292_579 ();
 b15zdnd11an1n08x5 FILLER_292_643 ();
 b15zdnd00an1n02x5 FILLER_292_651 ();
 b15zdnd11an1n32x5 FILLER_292_680 ();
 b15zdnd11an1n04x5 FILLER_292_712 ();
 b15zdnd00an1n02x5 FILLER_292_716 ();
 b15zdnd11an1n64x5 FILLER_292_726 ();
 b15zdnd11an1n64x5 FILLER_292_790 ();
 b15zdnd00an1n02x5 FILLER_292_854 ();
 b15zdnd11an1n64x5 FILLER_292_860 ();
 b15zdnd11an1n64x5 FILLER_292_924 ();
 b15zdnd11an1n64x5 FILLER_292_988 ();
 b15zdnd11an1n16x5 FILLER_292_1052 ();
 b15zdnd11an1n08x5 FILLER_292_1068 ();
 b15zdnd00an1n01x5 FILLER_292_1076 ();
 b15zdnd11an1n64x5 FILLER_292_1083 ();
 b15zdnd11an1n64x5 FILLER_292_1147 ();
 b15zdnd11an1n16x5 FILLER_292_1211 ();
 b15zdnd00an1n02x5 FILLER_292_1227 ();
 b15zdnd00an1n01x5 FILLER_292_1229 ();
 b15zdnd11an1n64x5 FILLER_292_1250 ();
 b15zdnd11an1n64x5 FILLER_292_1314 ();
 b15zdnd11an1n32x5 FILLER_292_1378 ();
 b15zdnd11an1n04x5 FILLER_292_1410 ();
 b15zdnd00an1n01x5 FILLER_292_1414 ();
 b15zdnd11an1n64x5 FILLER_292_1467 ();
 b15zdnd00an1n01x5 FILLER_292_1531 ();
 b15zdnd11an1n64x5 FILLER_292_1584 ();
 b15zdnd11an1n64x5 FILLER_292_1648 ();
 b15zdnd11an1n16x5 FILLER_292_1712 ();
 b15zdnd11an1n08x5 FILLER_292_1728 ();
 b15zdnd00an1n02x5 FILLER_292_1736 ();
 b15zdnd11an1n32x5 FILLER_292_1747 ();
 b15zdnd00an1n01x5 FILLER_292_1779 ();
 b15zdnd11an1n04x5 FILLER_292_1783 ();
 b15zdnd11an1n64x5 FILLER_292_1790 ();
 b15zdnd11an1n64x5 FILLER_292_1854 ();
 b15zdnd11an1n64x5 FILLER_292_1918 ();
 b15zdnd11an1n64x5 FILLER_292_1982 ();
 b15zdnd11an1n32x5 FILLER_292_2046 ();
 b15zdnd11an1n08x5 FILLER_292_2078 ();
 b15zdnd00an1n02x5 FILLER_292_2086 ();
 b15zdnd00an1n01x5 FILLER_292_2088 ();
 b15zdnd11an1n16x5 FILLER_292_2092 ();
 b15zdnd11an1n08x5 FILLER_292_2108 ();
 b15zdnd11an1n04x5 FILLER_292_2116 ();
 b15zdnd11an1n08x5 FILLER_292_2145 ();
 b15zdnd00an1n01x5 FILLER_292_2153 ();
 b15zdnd11an1n64x5 FILLER_292_2162 ();
 b15zdnd11an1n32x5 FILLER_292_2226 ();
 b15zdnd11an1n16x5 FILLER_292_2258 ();
 b15zdnd00an1n02x5 FILLER_292_2274 ();
 b15zdnd11an1n32x5 FILLER_293_0 ();
 b15zdnd11an1n16x5 FILLER_293_32 ();
 b15zdnd11an1n08x5 FILLER_293_48 ();
 b15zdnd00an1n02x5 FILLER_293_56 ();
 b15zdnd11an1n32x5 FILLER_293_83 ();
 b15zdnd11an1n08x5 FILLER_293_115 ();
 b15zdnd11an1n04x5 FILLER_293_123 ();
 b15zdnd00an1n01x5 FILLER_293_127 ();
 b15zdnd11an1n04x5 FILLER_293_153 ();
 b15zdnd11an1n64x5 FILLER_293_197 ();
 b15zdnd11an1n64x5 FILLER_293_261 ();
 b15zdnd11an1n64x5 FILLER_293_325 ();
 b15zdnd11an1n64x5 FILLER_293_389 ();
 b15zdnd11an1n32x5 FILLER_293_453 ();
 b15zdnd11an1n16x5 FILLER_293_485 ();
 b15zdnd11an1n04x5 FILLER_293_512 ();
 b15zdnd11an1n64x5 FILLER_293_522 ();
 b15zdnd11an1n64x5 FILLER_293_586 ();
 b15zdnd11an1n64x5 FILLER_293_650 ();
 b15zdnd11an1n64x5 FILLER_293_714 ();
 b15zdnd11an1n64x5 FILLER_293_778 ();
 b15zdnd11an1n64x5 FILLER_293_842 ();
 b15zdnd11an1n64x5 FILLER_293_906 ();
 b15zdnd11an1n64x5 FILLER_293_970 ();
 b15zdnd00an1n02x5 FILLER_293_1034 ();
 b15zdnd00an1n01x5 FILLER_293_1036 ();
 b15zdnd11an1n32x5 FILLER_293_1041 ();
 b15zdnd11an1n16x5 FILLER_293_1073 ();
 b15zdnd11an1n04x5 FILLER_293_1089 ();
 b15zdnd00an1n01x5 FILLER_293_1093 ();
 b15zdnd11an1n64x5 FILLER_293_1101 ();
 b15zdnd11an1n64x5 FILLER_293_1165 ();
 b15zdnd11an1n64x5 FILLER_293_1229 ();
 b15zdnd11an1n04x5 FILLER_293_1293 ();
 b15zdnd00an1n02x5 FILLER_293_1297 ();
 b15zdnd00an1n01x5 FILLER_293_1299 ();
 b15zdnd11an1n64x5 FILLER_293_1314 ();
 b15zdnd11an1n32x5 FILLER_293_1378 ();
 b15zdnd11an1n16x5 FILLER_293_1410 ();
 b15zdnd11an1n04x5 FILLER_293_1426 ();
 b15zdnd00an1n02x5 FILLER_293_1430 ();
 b15zdnd00an1n01x5 FILLER_293_1432 ();
 b15zdnd11an1n04x5 FILLER_293_1436 ();
 b15zdnd11an1n04x5 FILLER_293_1443 ();
 b15zdnd11an1n04x5 FILLER_293_1450 ();
 b15zdnd11an1n64x5 FILLER_293_1457 ();
 b15zdnd11an1n32x5 FILLER_293_1521 ();
 b15zdnd11an1n04x5 FILLER_293_1553 ();
 b15zdnd00an1n01x5 FILLER_293_1557 ();
 b15zdnd11an1n64x5 FILLER_293_1561 ();
 b15zdnd11an1n64x5 FILLER_293_1625 ();
 b15zdnd11an1n16x5 FILLER_293_1689 ();
 b15zdnd00an1n02x5 FILLER_293_1705 ();
 b15zdnd00an1n01x5 FILLER_293_1707 ();
 b15zdnd11an1n64x5 FILLER_293_1718 ();
 b15zdnd11an1n64x5 FILLER_293_1782 ();
 b15zdnd11an1n64x5 FILLER_293_1846 ();
 b15zdnd11an1n64x5 FILLER_293_1910 ();
 b15zdnd11an1n64x5 FILLER_293_1974 ();
 b15zdnd11an1n16x5 FILLER_293_2038 ();
 b15zdnd11an1n08x5 FILLER_293_2054 ();
 b15zdnd00an1n02x5 FILLER_293_2062 ();
 b15zdnd11an1n04x5 FILLER_293_2116 ();
 b15zdnd11an1n64x5 FILLER_293_2162 ();
 b15zdnd11an1n32x5 FILLER_293_2226 ();
 b15zdnd11an1n16x5 FILLER_293_2258 ();
 b15zdnd11an1n08x5 FILLER_293_2274 ();
 b15zdnd00an1n02x5 FILLER_293_2282 ();
 b15zdnd11an1n32x5 FILLER_294_8 ();
 b15zdnd11an1n16x5 FILLER_294_40 ();
 b15zdnd11an1n08x5 FILLER_294_56 ();
 b15zdnd00an1n02x5 FILLER_294_64 ();
 b15zdnd00an1n01x5 FILLER_294_66 ();
 b15zdnd11an1n04x5 FILLER_294_109 ();
 b15zdnd00an1n02x5 FILLER_294_113 ();
 b15zdnd11an1n64x5 FILLER_294_118 ();
 b15zdnd11an1n64x5 FILLER_294_182 ();
 b15zdnd11an1n64x5 FILLER_294_246 ();
 b15zdnd11an1n64x5 FILLER_294_310 ();
 b15zdnd11an1n64x5 FILLER_294_374 ();
 b15zdnd11an1n32x5 FILLER_294_438 ();
 b15zdnd11an1n16x5 FILLER_294_470 ();
 b15zdnd11an1n04x5 FILLER_294_486 ();
 b15zdnd11an1n04x5 FILLER_294_494 ();
 b15zdnd11an1n04x5 FILLER_294_507 ();
 b15zdnd11an1n64x5 FILLER_294_524 ();
 b15zdnd11an1n64x5 FILLER_294_588 ();
 b15zdnd11an1n64x5 FILLER_294_652 ();
 b15zdnd00an1n02x5 FILLER_294_716 ();
 b15zdnd11an1n64x5 FILLER_294_726 ();
 b15zdnd11an1n64x5 FILLER_294_790 ();
 b15zdnd11an1n64x5 FILLER_294_854 ();
 b15zdnd11an1n16x5 FILLER_294_918 ();
 b15zdnd00an1n02x5 FILLER_294_934 ();
 b15zdnd00an1n01x5 FILLER_294_936 ();
 b15zdnd11an1n16x5 FILLER_294_940 ();
 b15zdnd11an1n08x5 FILLER_294_956 ();
 b15zdnd11an1n04x5 FILLER_294_964 ();
 b15zdnd11an1n08x5 FILLER_294_971 ();
 b15zdnd11an1n04x5 FILLER_294_979 ();
 b15zdnd00an1n01x5 FILLER_294_983 ();
 b15zdnd11an1n64x5 FILLER_294_987 ();
 b15zdnd11an1n16x5 FILLER_294_1051 ();
 b15zdnd11an1n04x5 FILLER_294_1067 ();
 b15zdnd00an1n02x5 FILLER_294_1071 ();
 b15zdnd11an1n64x5 FILLER_294_1100 ();
 b15zdnd11an1n32x5 FILLER_294_1164 ();
 b15zdnd11an1n16x5 FILLER_294_1196 ();
 b15zdnd00an1n01x5 FILLER_294_1212 ();
 b15zdnd11an1n64x5 FILLER_294_1227 ();
 b15zdnd11an1n64x5 FILLER_294_1291 ();
 b15zdnd11an1n64x5 FILLER_294_1355 ();
 b15zdnd11an1n16x5 FILLER_294_1419 ();
 b15zdnd11an1n04x5 FILLER_294_1438 ();
 b15zdnd11an1n64x5 FILLER_294_1445 ();
 b15zdnd11an1n64x5 FILLER_294_1509 ();
 b15zdnd11an1n64x5 FILLER_294_1573 ();
 b15zdnd11an1n64x5 FILLER_294_1637 ();
 b15zdnd11an1n64x5 FILLER_294_1701 ();
 b15zdnd11an1n64x5 FILLER_294_1765 ();
 b15zdnd11an1n64x5 FILLER_294_1829 ();
 b15zdnd11an1n64x5 FILLER_294_1893 ();
 b15zdnd11an1n64x5 FILLER_294_1957 ();
 b15zdnd11an1n64x5 FILLER_294_2021 ();
 b15zdnd11an1n04x5 FILLER_294_2085 ();
 b15zdnd11an1n32x5 FILLER_294_2092 ();
 b15zdnd11an1n16x5 FILLER_294_2124 ();
 b15zdnd11an1n08x5 FILLER_294_2140 ();
 b15zdnd11an1n04x5 FILLER_294_2148 ();
 b15zdnd00an1n02x5 FILLER_294_2152 ();
 b15zdnd11an1n64x5 FILLER_294_2162 ();
 b15zdnd11an1n32x5 FILLER_294_2226 ();
 b15zdnd11an1n16x5 FILLER_294_2258 ();
 b15zdnd00an1n02x5 FILLER_294_2274 ();
 b15zdnd00an1n02x5 FILLER_295_0 ();
 b15zdnd11an1n08x5 FILLER_295_7 ();
 b15zdnd11an1n04x5 FILLER_295_15 ();
 b15zdnd00an1n02x5 FILLER_295_19 ();
 b15zdnd11an1n32x5 FILLER_295_25 ();
 b15zdnd11an1n16x5 FILLER_295_57 ();
 b15zdnd11an1n08x5 FILLER_295_73 ();
 b15zdnd00an1n01x5 FILLER_295_81 ();
 b15zdnd11an1n04x5 FILLER_295_122 ();
 b15zdnd11an1n08x5 FILLER_295_129 ();
 b15zdnd00an1n02x5 FILLER_295_137 ();
 b15zdnd00an1n01x5 FILLER_295_139 ();
 b15zdnd11an1n64x5 FILLER_295_158 ();
 b15zdnd11an1n64x5 FILLER_295_222 ();
 b15zdnd11an1n64x5 FILLER_295_286 ();
 b15zdnd11an1n64x5 FILLER_295_350 ();
 b15zdnd11an1n64x5 FILLER_295_414 ();
 b15zdnd11an1n08x5 FILLER_295_478 ();
 b15zdnd11an1n04x5 FILLER_295_486 ();
 b15zdnd00an1n02x5 FILLER_295_490 ();
 b15zdnd11an1n04x5 FILLER_295_499 ();
 b15zdnd00an1n02x5 FILLER_295_503 ();
 b15zdnd11an1n64x5 FILLER_295_547 ();
 b15zdnd11an1n64x5 FILLER_295_611 ();
 b15zdnd11an1n64x5 FILLER_295_675 ();
 b15zdnd11an1n64x5 FILLER_295_739 ();
 b15zdnd11an1n64x5 FILLER_295_803 ();
 b15zdnd11an1n32x5 FILLER_295_867 ();
 b15zdnd11an1n08x5 FILLER_295_899 ();
 b15zdnd11an1n04x5 FILLER_295_907 ();
 b15zdnd11an1n04x5 FILLER_295_963 ();
 b15zdnd11an1n16x5 FILLER_295_1019 ();
 b15zdnd11an1n08x5 FILLER_295_1043 ();
 b15zdnd11an1n08x5 FILLER_295_1055 ();
 b15zdnd11an1n04x5 FILLER_295_1063 ();
 b15zdnd11an1n32x5 FILLER_295_1071 ();
 b15zdnd11an1n08x5 FILLER_295_1103 ();
 b15zdnd11an1n64x5 FILLER_295_1114 ();
 b15zdnd11an1n32x5 FILLER_295_1178 ();
 b15zdnd11an1n16x5 FILLER_295_1210 ();
 b15zdnd00an1n02x5 FILLER_295_1226 ();
 b15zdnd00an1n01x5 FILLER_295_1228 ();
 b15zdnd11an1n32x5 FILLER_295_1271 ();
 b15zdnd11an1n04x5 FILLER_295_1303 ();
 b15zdnd00an1n02x5 FILLER_295_1307 ();
 b15zdnd00an1n01x5 FILLER_295_1309 ();
 b15zdnd11an1n04x5 FILLER_295_1324 ();
 b15zdnd00an1n02x5 FILLER_295_1328 ();
 b15zdnd00an1n01x5 FILLER_295_1330 ();
 b15zdnd11an1n64x5 FILLER_295_1345 ();
 b15zdnd11an1n64x5 FILLER_295_1409 ();
 b15zdnd11an1n64x5 FILLER_295_1473 ();
 b15zdnd11an1n64x5 FILLER_295_1537 ();
 b15zdnd11an1n64x5 FILLER_295_1601 ();
 b15zdnd11an1n64x5 FILLER_295_1665 ();
 b15zdnd11an1n64x5 FILLER_295_1729 ();
 b15zdnd11an1n64x5 FILLER_295_1793 ();
 b15zdnd11an1n64x5 FILLER_295_1857 ();
 b15zdnd11an1n64x5 FILLER_295_1921 ();
 b15zdnd11an1n64x5 FILLER_295_1985 ();
 b15zdnd11an1n64x5 FILLER_295_2049 ();
 b15zdnd11an1n64x5 FILLER_295_2113 ();
 b15zdnd11an1n64x5 FILLER_295_2177 ();
 b15zdnd11an1n32x5 FILLER_295_2241 ();
 b15zdnd11an1n08x5 FILLER_295_2273 ();
 b15zdnd00an1n02x5 FILLER_295_2281 ();
 b15zdnd00an1n01x5 FILLER_295_2283 ();
 b15zdnd00an1n02x5 FILLER_296_8 ();
 b15zdnd11an1n08x5 FILLER_296_17 ();
 b15zdnd00an1n02x5 FILLER_296_25 ();
 b15zdnd00an1n01x5 FILLER_296_27 ();
 b15zdnd11an1n64x5 FILLER_296_36 ();
 b15zdnd11an1n04x5 FILLER_296_100 ();
 b15zdnd00an1n02x5 FILLER_296_104 ();
 b15zdnd11an1n04x5 FILLER_296_148 ();
 b15zdnd00an1n02x5 FILLER_296_152 ();
 b15zdnd00an1n01x5 FILLER_296_154 ();
 b15zdnd11an1n64x5 FILLER_296_180 ();
 b15zdnd11an1n64x5 FILLER_296_244 ();
 b15zdnd11an1n64x5 FILLER_296_308 ();
 b15zdnd11an1n64x5 FILLER_296_372 ();
 b15zdnd11an1n64x5 FILLER_296_436 ();
 b15zdnd11an1n08x5 FILLER_296_500 ();
 b15zdnd11an1n04x5 FILLER_296_511 ();
 b15zdnd11an1n64x5 FILLER_296_557 ();
 b15zdnd11an1n64x5 FILLER_296_621 ();
 b15zdnd11an1n32x5 FILLER_296_685 ();
 b15zdnd00an1n01x5 FILLER_296_717 ();
 b15zdnd11an1n64x5 FILLER_296_726 ();
 b15zdnd11an1n64x5 FILLER_296_790 ();
 b15zdnd11an1n64x5 FILLER_296_854 ();
 b15zdnd11an1n08x5 FILLER_296_918 ();
 b15zdnd00an1n02x5 FILLER_296_926 ();
 b15zdnd00an1n01x5 FILLER_296_928 ();
 b15zdnd11an1n04x5 FILLER_296_932 ();
 b15zdnd00an1n02x5 FILLER_296_936 ();
 b15zdnd11an1n16x5 FILLER_296_941 ();
 b15zdnd11an1n04x5 FILLER_296_957 ();
 b15zdnd00an1n02x5 FILLER_296_961 ();
 b15zdnd00an1n01x5 FILLER_296_963 ();
 b15zdnd11an1n64x5 FILLER_296_1016 ();
 b15zdnd11an1n08x5 FILLER_296_1080 ();
 b15zdnd00an1n01x5 FILLER_296_1088 ();
 b15zdnd11an1n64x5 FILLER_296_1141 ();
 b15zdnd11an1n04x5 FILLER_296_1205 ();
 b15zdnd00an1n01x5 FILLER_296_1209 ();
 b15zdnd11an1n08x5 FILLER_296_1227 ();
 b15zdnd00an1n02x5 FILLER_296_1235 ();
 b15zdnd00an1n01x5 FILLER_296_1237 ();
 b15zdnd11an1n64x5 FILLER_296_1244 ();
 b15zdnd11an1n64x5 FILLER_296_1308 ();
 b15zdnd11an1n08x5 FILLER_296_1372 ();
 b15zdnd11an1n04x5 FILLER_296_1380 ();
 b15zdnd00an1n02x5 FILLER_296_1384 ();
 b15zdnd11an1n64x5 FILLER_296_1390 ();
 b15zdnd11an1n64x5 FILLER_296_1454 ();
 b15zdnd11an1n64x5 FILLER_296_1518 ();
 b15zdnd11an1n64x5 FILLER_296_1582 ();
 b15zdnd11an1n64x5 FILLER_296_1646 ();
 b15zdnd11an1n64x5 FILLER_296_1710 ();
 b15zdnd11an1n64x5 FILLER_296_1774 ();
 b15zdnd11an1n64x5 FILLER_296_1838 ();
 b15zdnd11an1n64x5 FILLER_296_1902 ();
 b15zdnd11an1n64x5 FILLER_296_1966 ();
 b15zdnd11an1n32x5 FILLER_296_2030 ();
 b15zdnd11an1n16x5 FILLER_296_2062 ();
 b15zdnd11an1n32x5 FILLER_296_2120 ();
 b15zdnd00an1n02x5 FILLER_296_2152 ();
 b15zdnd11an1n64x5 FILLER_296_2162 ();
 b15zdnd11an1n32x5 FILLER_296_2226 ();
 b15zdnd11an1n16x5 FILLER_296_2258 ();
 b15zdnd00an1n02x5 FILLER_296_2274 ();
 b15zdnd11an1n16x5 FILLER_297_0 ();
 b15zdnd00an1n01x5 FILLER_297_16 ();
 b15zdnd11an1n32x5 FILLER_297_21 ();
 b15zdnd11an1n16x5 FILLER_297_53 ();
 b15zdnd11an1n04x5 FILLER_297_69 ();
 b15zdnd00an1n02x5 FILLER_297_73 ();
 b15zdnd00an1n01x5 FILLER_297_75 ();
 b15zdnd11an1n08x5 FILLER_297_121 ();
 b15zdnd00an1n01x5 FILLER_297_129 ();
 b15zdnd11an1n64x5 FILLER_297_161 ();
 b15zdnd11an1n64x5 FILLER_297_225 ();
 b15zdnd11an1n64x5 FILLER_297_289 ();
 b15zdnd11an1n64x5 FILLER_297_353 ();
 b15zdnd11an1n64x5 FILLER_297_417 ();
 b15zdnd11an1n08x5 FILLER_297_481 ();
 b15zdnd11an1n04x5 FILLER_297_489 ();
 b15zdnd00an1n02x5 FILLER_297_493 ();
 b15zdnd11an1n64x5 FILLER_297_547 ();
 b15zdnd11an1n64x5 FILLER_297_611 ();
 b15zdnd11an1n64x5 FILLER_297_675 ();
 b15zdnd11an1n64x5 FILLER_297_739 ();
 b15zdnd11an1n64x5 FILLER_297_803 ();
 b15zdnd11an1n64x5 FILLER_297_867 ();
 b15zdnd11an1n08x5 FILLER_297_931 ();
 b15zdnd11an1n16x5 FILLER_297_942 ();
 b15zdnd11an1n08x5 FILLER_297_958 ();
 b15zdnd11an1n04x5 FILLER_297_966 ();
 b15zdnd00an1n01x5 FILLER_297_970 ();
 b15zdnd11an1n08x5 FILLER_297_974 ();
 b15zdnd00an1n02x5 FILLER_297_982 ();
 b15zdnd11an1n64x5 FILLER_297_987 ();
 b15zdnd11an1n32x5 FILLER_297_1051 ();
 b15zdnd11an1n16x5 FILLER_297_1083 ();
 b15zdnd11an1n08x5 FILLER_297_1099 ();
 b15zdnd11an1n04x5 FILLER_297_1107 ();
 b15zdnd11an1n04x5 FILLER_297_1114 ();
 b15zdnd11an1n16x5 FILLER_297_1121 ();
 b15zdnd11an1n08x5 FILLER_297_1137 ();
 b15zdnd00an1n02x5 FILLER_297_1145 ();
 b15zdnd00an1n01x5 FILLER_297_1147 ();
 b15zdnd11an1n08x5 FILLER_297_1190 ();
 b15zdnd11an1n04x5 FILLER_297_1198 ();
 b15zdnd00an1n02x5 FILLER_297_1202 ();
 b15zdnd00an1n01x5 FILLER_297_1204 ();
 b15zdnd11an1n64x5 FILLER_297_1219 ();
 b15zdnd11an1n04x5 FILLER_297_1283 ();
 b15zdnd00an1n02x5 FILLER_297_1287 ();
 b15zdnd11an1n64x5 FILLER_297_1303 ();
 b15zdnd11an1n64x5 FILLER_297_1367 ();
 b15zdnd11an1n64x5 FILLER_297_1431 ();
 b15zdnd11an1n64x5 FILLER_297_1495 ();
 b15zdnd11an1n64x5 FILLER_297_1559 ();
 b15zdnd11an1n64x5 FILLER_297_1623 ();
 b15zdnd11an1n64x5 FILLER_297_1687 ();
 b15zdnd11an1n64x5 FILLER_297_1751 ();
 b15zdnd11an1n64x5 FILLER_297_1815 ();
 b15zdnd11an1n32x5 FILLER_297_1879 ();
 b15zdnd00an1n02x5 FILLER_297_1911 ();
 b15zdnd11an1n64x5 FILLER_297_1919 ();
 b15zdnd11an1n64x5 FILLER_297_1983 ();
 b15zdnd11an1n64x5 FILLER_297_2047 ();
 b15zdnd11an1n64x5 FILLER_297_2111 ();
 b15zdnd11an1n64x5 FILLER_297_2175 ();
 b15zdnd11an1n32x5 FILLER_297_2239 ();
 b15zdnd11an1n08x5 FILLER_297_2271 ();
 b15zdnd11an1n04x5 FILLER_297_2279 ();
 b15zdnd00an1n01x5 FILLER_297_2283 ();
 b15zdnd11an1n64x5 FILLER_298_8 ();
 b15zdnd11an1n64x5 FILLER_298_72 ();
 b15zdnd11an1n16x5 FILLER_298_136 ();
 b15zdnd11an1n04x5 FILLER_298_152 ();
 b15zdnd11an1n16x5 FILLER_298_198 ();
 b15zdnd00an1n02x5 FILLER_298_214 ();
 b15zdnd00an1n01x5 FILLER_298_216 ();
 b15zdnd11an1n64x5 FILLER_298_257 ();
 b15zdnd11an1n64x5 FILLER_298_321 ();
 b15zdnd11an1n64x5 FILLER_298_385 ();
 b15zdnd11an1n64x5 FILLER_298_449 ();
 b15zdnd00an1n02x5 FILLER_298_513 ();
 b15zdnd11an1n04x5 FILLER_298_518 ();
 b15zdnd11an1n64x5 FILLER_298_525 ();
 b15zdnd11an1n32x5 FILLER_298_589 ();
 b15zdnd11an1n04x5 FILLER_298_621 ();
 b15zdnd00an1n02x5 FILLER_298_625 ();
 b15zdnd00an1n01x5 FILLER_298_627 ();
 b15zdnd11an1n32x5 FILLER_298_670 ();
 b15zdnd11an1n16x5 FILLER_298_702 ();
 b15zdnd11an1n64x5 FILLER_298_726 ();
 b15zdnd11an1n64x5 FILLER_298_790 ();
 b15zdnd11an1n32x5 FILLER_298_854 ();
 b15zdnd11an1n08x5 FILLER_298_886 ();
 b15zdnd11an1n04x5 FILLER_298_894 ();
 b15zdnd00an1n01x5 FILLER_298_898 ();
 b15zdnd11an1n08x5 FILLER_298_904 ();
 b15zdnd11an1n04x5 FILLER_298_912 ();
 b15zdnd11an1n08x5 FILLER_298_968 ();
 b15zdnd00an1n02x5 FILLER_298_976 ();
 b15zdnd00an1n01x5 FILLER_298_978 ();
 b15zdnd11an1n08x5 FILLER_298_982 ();
 b15zdnd11an1n64x5 FILLER_298_993 ();
 b15zdnd11an1n32x5 FILLER_298_1057 ();
 b15zdnd11an1n04x5 FILLER_298_1089 ();
 b15zdnd11an1n16x5 FILLER_298_1114 ();
 b15zdnd11an1n08x5 FILLER_298_1130 ();
 b15zdnd11an1n04x5 FILLER_298_1180 ();
 b15zdnd00an1n01x5 FILLER_298_1184 ();
 b15zdnd11an1n16x5 FILLER_298_1188 ();
 b15zdnd11an1n04x5 FILLER_298_1204 ();
 b15zdnd00an1n02x5 FILLER_298_1208 ();
 b15zdnd00an1n01x5 FILLER_298_1210 ();
 b15zdnd11an1n16x5 FILLER_298_1253 ();
 b15zdnd11an1n08x5 FILLER_298_1269 ();
 b15zdnd00an1n02x5 FILLER_298_1277 ();
 b15zdnd00an1n01x5 FILLER_298_1279 ();
 b15zdnd11an1n64x5 FILLER_298_1283 ();
 b15zdnd11an1n64x5 FILLER_298_1347 ();
 b15zdnd11an1n32x5 FILLER_298_1411 ();
 b15zdnd11an1n04x5 FILLER_298_1443 ();
 b15zdnd00an1n02x5 FILLER_298_1447 ();
 b15zdnd11an1n64x5 FILLER_298_1460 ();
 b15zdnd11an1n64x5 FILLER_298_1524 ();
 b15zdnd11an1n64x5 FILLER_298_1588 ();
 b15zdnd11an1n64x5 FILLER_298_1652 ();
 b15zdnd11an1n32x5 FILLER_298_1716 ();
 b15zdnd11an1n04x5 FILLER_298_1748 ();
 b15zdnd00an1n01x5 FILLER_298_1752 ();
 b15zdnd11an1n64x5 FILLER_298_1762 ();
 b15zdnd11an1n32x5 FILLER_298_1826 ();
 b15zdnd11an1n16x5 FILLER_298_1858 ();
 b15zdnd11an1n08x5 FILLER_298_1874 ();
 b15zdnd11an1n04x5 FILLER_298_1882 ();
 b15zdnd00an1n01x5 FILLER_298_1886 ();
 b15zdnd11an1n64x5 FILLER_298_1929 ();
 b15zdnd11an1n64x5 FILLER_298_1993 ();
 b15zdnd11an1n32x5 FILLER_298_2057 ();
 b15zdnd11an1n32x5 FILLER_298_2093 ();
 b15zdnd11an1n16x5 FILLER_298_2125 ();
 b15zdnd11an1n08x5 FILLER_298_2141 ();
 b15zdnd11an1n04x5 FILLER_298_2149 ();
 b15zdnd00an1n01x5 FILLER_298_2153 ();
 b15zdnd11an1n64x5 FILLER_298_2162 ();
 b15zdnd11an1n32x5 FILLER_298_2226 ();
 b15zdnd11an1n16x5 FILLER_298_2258 ();
 b15zdnd00an1n02x5 FILLER_298_2274 ();
 b15zdnd11an1n64x5 FILLER_299_0 ();
 b15zdnd11an1n08x5 FILLER_299_64 ();
 b15zdnd11an1n04x5 FILLER_299_72 ();
 b15zdnd00an1n01x5 FILLER_299_76 ();
 b15zdnd11an1n64x5 FILLER_299_85 ();
 b15zdnd11an1n32x5 FILLER_299_149 ();
 b15zdnd11an1n08x5 FILLER_299_181 ();
 b15zdnd11an1n16x5 FILLER_299_231 ();
 b15zdnd11an1n08x5 FILLER_299_247 ();
 b15zdnd11an1n04x5 FILLER_299_255 ();
 b15zdnd00an1n02x5 FILLER_299_259 ();
 b15zdnd11an1n64x5 FILLER_299_264 ();
 b15zdnd11an1n64x5 FILLER_299_328 ();
 b15zdnd11an1n64x5 FILLER_299_392 ();
 b15zdnd11an1n64x5 FILLER_299_456 ();
 b15zdnd11an1n64x5 FILLER_299_520 ();
 b15zdnd11an1n64x5 FILLER_299_584 ();
 b15zdnd11an1n64x5 FILLER_299_648 ();
 b15zdnd11an1n64x5 FILLER_299_712 ();
 b15zdnd11an1n32x5 FILLER_299_776 ();
 b15zdnd11an1n04x5 FILLER_299_808 ();
 b15zdnd00an1n01x5 FILLER_299_812 ();
 b15zdnd11an1n64x5 FILLER_299_816 ();
 b15zdnd11an1n32x5 FILLER_299_880 ();
 b15zdnd11an1n16x5 FILLER_299_912 ();
 b15zdnd11an1n08x5 FILLER_299_928 ();
 b15zdnd11an1n04x5 FILLER_299_939 ();
 b15zdnd11an1n64x5 FILLER_299_946 ();
 b15zdnd11an1n64x5 FILLER_299_1010 ();
 b15zdnd11an1n32x5 FILLER_299_1074 ();
 b15zdnd11an1n16x5 FILLER_299_1106 ();
 b15zdnd11an1n08x5 FILLER_299_1122 ();
 b15zdnd00an1n01x5 FILLER_299_1130 ();
 b15zdnd11an1n04x5 FILLER_299_1138 ();
 b15zdnd11an1n32x5 FILLER_299_1149 ();
 b15zdnd11an1n04x5 FILLER_299_1181 ();
 b15zdnd00an1n01x5 FILLER_299_1185 ();
 b15zdnd11an1n16x5 FILLER_299_1189 ();
 b15zdnd11an1n08x5 FILLER_299_1205 ();
 b15zdnd00an1n01x5 FILLER_299_1213 ();
 b15zdnd11an1n16x5 FILLER_299_1256 ();
 b15zdnd11an1n08x5 FILLER_299_1272 ();
 b15zdnd11an1n04x5 FILLER_299_1280 ();
 b15zdnd00an1n01x5 FILLER_299_1284 ();
 b15zdnd11an1n64x5 FILLER_299_1299 ();
 b15zdnd11an1n64x5 FILLER_299_1363 ();
 b15zdnd11an1n64x5 FILLER_299_1427 ();
 b15zdnd11an1n64x5 FILLER_299_1491 ();
 b15zdnd11an1n64x5 FILLER_299_1555 ();
 b15zdnd11an1n64x5 FILLER_299_1619 ();
 b15zdnd11an1n64x5 FILLER_299_1683 ();
 b15zdnd11an1n64x5 FILLER_299_1747 ();
 b15zdnd11an1n64x5 FILLER_299_1811 ();
 b15zdnd11an1n16x5 FILLER_299_1875 ();
 b15zdnd11an1n08x5 FILLER_299_1891 ();
 b15zdnd11an1n04x5 FILLER_299_1899 ();
 b15zdnd00an1n01x5 FILLER_299_1903 ();
 b15zdnd11an1n64x5 FILLER_299_1925 ();
 b15zdnd11an1n64x5 FILLER_299_1989 ();
 b15zdnd11an1n64x5 FILLER_299_2053 ();
 b15zdnd11an1n64x5 FILLER_299_2117 ();
 b15zdnd11an1n64x5 FILLER_299_2181 ();
 b15zdnd11an1n32x5 FILLER_299_2245 ();
 b15zdnd11an1n04x5 FILLER_299_2277 ();
 b15zdnd00an1n02x5 FILLER_299_2281 ();
 b15zdnd00an1n01x5 FILLER_299_2283 ();
 b15zdnd00an1n02x5 FILLER_300_8 ();
 b15zdnd11an1n32x5 FILLER_300_17 ();
 b15zdnd11an1n16x5 FILLER_300_49 ();
 b15zdnd11an1n08x5 FILLER_300_65 ();
 b15zdnd11an1n04x5 FILLER_300_73 ();
 b15zdnd00an1n02x5 FILLER_300_77 ();
 b15zdnd00an1n01x5 FILLER_300_79 ();
 b15zdnd11an1n64x5 FILLER_300_94 ();
 b15zdnd11an1n64x5 FILLER_300_158 ();
 b15zdnd11an1n32x5 FILLER_300_222 ();
 b15zdnd11an1n16x5 FILLER_300_254 ();
 b15zdnd11an1n04x5 FILLER_300_270 ();
 b15zdnd00an1n01x5 FILLER_300_274 ();
 b15zdnd11an1n64x5 FILLER_300_286 ();
 b15zdnd11an1n64x5 FILLER_300_350 ();
 b15zdnd11an1n64x5 FILLER_300_414 ();
 b15zdnd11an1n64x5 FILLER_300_478 ();
 b15zdnd11an1n64x5 FILLER_300_542 ();
 b15zdnd11an1n64x5 FILLER_300_606 ();
 b15zdnd11an1n32x5 FILLER_300_670 ();
 b15zdnd11an1n16x5 FILLER_300_702 ();
 b15zdnd11an1n32x5 FILLER_300_726 ();
 b15zdnd11an1n16x5 FILLER_300_758 ();
 b15zdnd11an1n08x5 FILLER_300_774 ();
 b15zdnd11an1n04x5 FILLER_300_782 ();
 b15zdnd11an1n64x5 FILLER_300_838 ();
 b15zdnd11an1n64x5 FILLER_300_902 ();
 b15zdnd11an1n64x5 FILLER_300_966 ();
 b15zdnd11an1n64x5 FILLER_300_1030 ();
 b15zdnd11an1n64x5 FILLER_300_1094 ();
 b15zdnd00an1n02x5 FILLER_300_1158 ();
 b15zdnd00an1n01x5 FILLER_300_1160 ();
 b15zdnd11an1n64x5 FILLER_300_1213 ();
 b15zdnd11an1n64x5 FILLER_300_1277 ();
 b15zdnd00an1n01x5 FILLER_300_1341 ();
 b15zdnd11an1n64x5 FILLER_300_1345 ();
 b15zdnd11an1n64x5 FILLER_300_1409 ();
 b15zdnd11an1n64x5 FILLER_300_1473 ();
 b15zdnd11an1n16x5 FILLER_300_1537 ();
 b15zdnd11an1n04x5 FILLER_300_1553 ();
 b15zdnd00an1n01x5 FILLER_300_1557 ();
 b15zdnd11an1n04x5 FILLER_300_1562 ();
 b15zdnd11an1n64x5 FILLER_300_1586 ();
 b15zdnd11an1n64x5 FILLER_300_1650 ();
 b15zdnd11an1n64x5 FILLER_300_1714 ();
 b15zdnd11an1n64x5 FILLER_300_1778 ();
 b15zdnd11an1n64x5 FILLER_300_1842 ();
 b15zdnd11an1n64x5 FILLER_300_1906 ();
 b15zdnd11an1n64x5 FILLER_300_1970 ();
 b15zdnd11an1n64x5 FILLER_300_2034 ();
 b15zdnd11an1n08x5 FILLER_300_2098 ();
 b15zdnd11an1n04x5 FILLER_300_2106 ();
 b15zdnd00an1n02x5 FILLER_300_2110 ();
 b15zdnd00an1n01x5 FILLER_300_2112 ();
 b15zdnd11an1n32x5 FILLER_300_2118 ();
 b15zdnd11an1n04x5 FILLER_300_2150 ();
 b15zdnd11an1n64x5 FILLER_300_2162 ();
 b15zdnd11an1n32x5 FILLER_300_2226 ();
 b15zdnd11an1n16x5 FILLER_300_2258 ();
 b15zdnd00an1n02x5 FILLER_300_2274 ();
 b15zdnd11an1n64x5 FILLER_301_0 ();
 b15zdnd11an1n64x5 FILLER_301_64 ();
 b15zdnd11an1n64x5 FILLER_301_128 ();
 b15zdnd11an1n64x5 FILLER_301_192 ();
 b15zdnd11an1n64x5 FILLER_301_256 ();
 b15zdnd11an1n64x5 FILLER_301_320 ();
 b15zdnd11an1n64x5 FILLER_301_384 ();
 b15zdnd11an1n64x5 FILLER_301_448 ();
 b15zdnd11an1n08x5 FILLER_301_512 ();
 b15zdnd11an1n04x5 FILLER_301_520 ();
 b15zdnd00an1n01x5 FILLER_301_524 ();
 b15zdnd11an1n64x5 FILLER_301_530 ();
 b15zdnd11an1n64x5 FILLER_301_594 ();
 b15zdnd11an1n64x5 FILLER_301_658 ();
 b15zdnd11an1n64x5 FILLER_301_722 ();
 b15zdnd11an1n16x5 FILLER_301_786 ();
 b15zdnd00an1n02x5 FILLER_301_802 ();
 b15zdnd11an1n04x5 FILLER_301_807 ();
 b15zdnd11an1n64x5 FILLER_301_814 ();
 b15zdnd11an1n64x5 FILLER_301_878 ();
 b15zdnd11an1n64x5 FILLER_301_942 ();
 b15zdnd11an1n64x5 FILLER_301_1006 ();
 b15zdnd11an1n32x5 FILLER_301_1070 ();
 b15zdnd11an1n08x5 FILLER_301_1102 ();
 b15zdnd00an1n02x5 FILLER_301_1110 ();
 b15zdnd00an1n01x5 FILLER_301_1112 ();
 b15zdnd11an1n64x5 FILLER_301_1121 ();
 b15zdnd00an1n01x5 FILLER_301_1185 ();
 b15zdnd11an1n64x5 FILLER_301_1189 ();
 b15zdnd00an1n02x5 FILLER_301_1253 ();
 b15zdnd00an1n01x5 FILLER_301_1255 ();
 b15zdnd11an1n64x5 FILLER_301_1263 ();
 b15zdnd11an1n08x5 FILLER_301_1327 ();
 b15zdnd00an1n02x5 FILLER_301_1335 ();
 b15zdnd11an1n04x5 FILLER_301_1340 ();
 b15zdnd11an1n64x5 FILLER_301_1358 ();
 b15zdnd11an1n64x5 FILLER_301_1422 ();
 b15zdnd11an1n64x5 FILLER_301_1486 ();
 b15zdnd11an1n64x5 FILLER_301_1550 ();
 b15zdnd11an1n64x5 FILLER_301_1614 ();
 b15zdnd11an1n64x5 FILLER_301_1678 ();
 b15zdnd11an1n64x5 FILLER_301_1742 ();
 b15zdnd11an1n64x5 FILLER_301_1806 ();
 b15zdnd11an1n64x5 FILLER_301_1870 ();
 b15zdnd11an1n64x5 FILLER_301_1934 ();
 b15zdnd11an1n64x5 FILLER_301_1998 ();
 b15zdnd11an1n64x5 FILLER_301_2062 ();
 b15zdnd11an1n64x5 FILLER_301_2126 ();
 b15zdnd11an1n64x5 FILLER_301_2190 ();
 b15zdnd11an1n16x5 FILLER_301_2254 ();
 b15zdnd11an1n08x5 FILLER_301_2270 ();
 b15zdnd11an1n04x5 FILLER_301_2278 ();
 b15zdnd00an1n02x5 FILLER_301_2282 ();
 b15zdnd11an1n16x5 FILLER_302_8 ();
 b15zdnd00an1n01x5 FILLER_302_24 ();
 b15zdnd11an1n64x5 FILLER_302_43 ();
 b15zdnd11an1n64x5 FILLER_302_107 ();
 b15zdnd11an1n64x5 FILLER_302_171 ();
 b15zdnd11an1n16x5 FILLER_302_235 ();
 b15zdnd00an1n01x5 FILLER_302_251 ();
 b15zdnd11an1n64x5 FILLER_302_255 ();
 b15zdnd11an1n64x5 FILLER_302_319 ();
 b15zdnd11an1n64x5 FILLER_302_383 ();
 b15zdnd11an1n64x5 FILLER_302_447 ();
 b15zdnd11an1n64x5 FILLER_302_511 ();
 b15zdnd11an1n64x5 FILLER_302_575 ();
 b15zdnd11an1n64x5 FILLER_302_639 ();
 b15zdnd11an1n08x5 FILLER_302_703 ();
 b15zdnd11an1n04x5 FILLER_302_711 ();
 b15zdnd00an1n02x5 FILLER_302_715 ();
 b15zdnd00an1n01x5 FILLER_302_717 ();
 b15zdnd11an1n64x5 FILLER_302_726 ();
 b15zdnd11an1n64x5 FILLER_302_790 ();
 b15zdnd11an1n64x5 FILLER_302_854 ();
 b15zdnd11an1n64x5 FILLER_302_918 ();
 b15zdnd11an1n64x5 FILLER_302_982 ();
 b15zdnd11an1n64x5 FILLER_302_1046 ();
 b15zdnd11an1n64x5 FILLER_302_1110 ();
 b15zdnd11an1n64x5 FILLER_302_1174 ();
 b15zdnd11an1n64x5 FILLER_302_1238 ();
 b15zdnd11an1n64x5 FILLER_302_1302 ();
 b15zdnd11an1n64x5 FILLER_302_1366 ();
 b15zdnd11an1n64x5 FILLER_302_1430 ();
 b15zdnd11an1n64x5 FILLER_302_1494 ();
 b15zdnd11an1n32x5 FILLER_302_1558 ();
 b15zdnd00an1n02x5 FILLER_302_1590 ();
 b15zdnd00an1n01x5 FILLER_302_1592 ();
 b15zdnd11an1n64x5 FILLER_302_1601 ();
 b15zdnd11an1n64x5 FILLER_302_1665 ();
 b15zdnd11an1n08x5 FILLER_302_1729 ();
 b15zdnd00an1n01x5 FILLER_302_1737 ();
 b15zdnd11an1n64x5 FILLER_302_1747 ();
 b15zdnd11an1n64x5 FILLER_302_1811 ();
 b15zdnd11an1n32x5 FILLER_302_1875 ();
 b15zdnd11an1n04x5 FILLER_302_1907 ();
 b15zdnd00an1n02x5 FILLER_302_1911 ();
 b15zdnd00an1n01x5 FILLER_302_1913 ();
 b15zdnd11an1n08x5 FILLER_302_1921 ();
 b15zdnd11an1n04x5 FILLER_302_1929 ();
 b15zdnd00an1n01x5 FILLER_302_1933 ();
 b15zdnd11an1n04x5 FILLER_302_1937 ();
 b15zdnd11an1n64x5 FILLER_302_1944 ();
 b15zdnd11an1n64x5 FILLER_302_2008 ();
 b15zdnd11an1n64x5 FILLER_302_2072 ();
 b15zdnd11an1n16x5 FILLER_302_2136 ();
 b15zdnd00an1n02x5 FILLER_302_2152 ();
 b15zdnd11an1n64x5 FILLER_302_2162 ();
 b15zdnd11an1n32x5 FILLER_302_2226 ();
 b15zdnd11an1n16x5 FILLER_302_2258 ();
 b15zdnd00an1n02x5 FILLER_302_2274 ();
 b15zdnd11an1n04x5 FILLER_303_0 ();
 b15zdnd00an1n02x5 FILLER_303_4 ();
 b15zdnd00an1n01x5 FILLER_303_6 ();
 b15zdnd11an1n64x5 FILLER_303_13 ();
 b15zdnd11an1n64x5 FILLER_303_77 ();
 b15zdnd11an1n64x5 FILLER_303_141 ();
 b15zdnd11an1n64x5 FILLER_303_205 ();
 b15zdnd11an1n64x5 FILLER_303_269 ();
 b15zdnd11an1n32x5 FILLER_303_333 ();
 b15zdnd00an1n02x5 FILLER_303_365 ();
 b15zdnd11an1n04x5 FILLER_303_385 ();
 b15zdnd11an1n64x5 FILLER_303_393 ();
 b15zdnd11an1n64x5 FILLER_303_457 ();
 b15zdnd11an1n64x5 FILLER_303_521 ();
 b15zdnd11an1n64x5 FILLER_303_585 ();
 b15zdnd11an1n64x5 FILLER_303_649 ();
 b15zdnd11an1n64x5 FILLER_303_713 ();
 b15zdnd11an1n64x5 FILLER_303_777 ();
 b15zdnd11an1n64x5 FILLER_303_841 ();
 b15zdnd11an1n64x5 FILLER_303_905 ();
 b15zdnd11an1n64x5 FILLER_303_969 ();
 b15zdnd11an1n64x5 FILLER_303_1033 ();
 b15zdnd11an1n64x5 FILLER_303_1097 ();
 b15zdnd11an1n32x5 FILLER_303_1161 ();
 b15zdnd11an1n04x5 FILLER_303_1193 ();
 b15zdnd00an1n02x5 FILLER_303_1197 ();
 b15zdnd00an1n01x5 FILLER_303_1199 ();
 b15zdnd11an1n64x5 FILLER_303_1220 ();
 b15zdnd11an1n04x5 FILLER_303_1284 ();
 b15zdnd00an1n02x5 FILLER_303_1288 ();
 b15zdnd00an1n01x5 FILLER_303_1290 ();
 b15zdnd11an1n16x5 FILLER_303_1299 ();
 b15zdnd11an1n04x5 FILLER_303_1315 ();
 b15zdnd00an1n02x5 FILLER_303_1319 ();
 b15zdnd00an1n01x5 FILLER_303_1321 ();
 b15zdnd11an1n08x5 FILLER_303_1343 ();
 b15zdnd11an1n64x5 FILLER_303_1369 ();
 b15zdnd11an1n64x5 FILLER_303_1433 ();
 b15zdnd11an1n64x5 FILLER_303_1497 ();
 b15zdnd11an1n64x5 FILLER_303_1561 ();
 b15zdnd11an1n64x5 FILLER_303_1625 ();
 b15zdnd11an1n64x5 FILLER_303_1689 ();
 b15zdnd11an1n64x5 FILLER_303_1753 ();
 b15zdnd11an1n64x5 FILLER_303_1817 ();
 b15zdnd11an1n32x5 FILLER_303_1881 ();
 b15zdnd11an1n04x5 FILLER_303_1913 ();
 b15zdnd00an1n02x5 FILLER_303_1917 ();
 b15zdnd11an1n64x5 FILLER_303_1963 ();
 b15zdnd11an1n64x5 FILLER_303_2027 ();
 b15zdnd11an1n32x5 FILLER_303_2091 ();
 b15zdnd11an1n08x5 FILLER_303_2123 ();
 b15zdnd00an1n02x5 FILLER_303_2131 ();
 b15zdnd00an1n01x5 FILLER_303_2133 ();
 b15zdnd11an1n64x5 FILLER_303_2176 ();
 b15zdnd11an1n32x5 FILLER_303_2240 ();
 b15zdnd11an1n08x5 FILLER_303_2272 ();
 b15zdnd11an1n04x5 FILLER_303_2280 ();
 b15zdnd11an1n16x5 FILLER_304_8 ();
 b15zdnd11an1n04x5 FILLER_304_24 ();
 b15zdnd00an1n02x5 FILLER_304_28 ();
 b15zdnd11an1n64x5 FILLER_304_36 ();
 b15zdnd11an1n64x5 FILLER_304_100 ();
 b15zdnd11an1n64x5 FILLER_304_164 ();
 b15zdnd11an1n64x5 FILLER_304_228 ();
 b15zdnd11an1n64x5 FILLER_304_292 ();
 b15zdnd11an1n32x5 FILLER_304_356 ();
 b15zdnd11an1n16x5 FILLER_304_407 ();
 b15zdnd11an1n08x5 FILLER_304_423 ();
 b15zdnd11an1n04x5 FILLER_304_431 ();
 b15zdnd00an1n02x5 FILLER_304_435 ();
 b15zdnd11an1n32x5 FILLER_304_445 ();
 b15zdnd11an1n16x5 FILLER_304_477 ();
 b15zdnd11an1n04x5 FILLER_304_493 ();
 b15zdnd00an1n02x5 FILLER_304_497 ();
 b15zdnd11an1n04x5 FILLER_304_515 ();
 b15zdnd11an1n32x5 FILLER_304_533 ();
 b15zdnd00an1n02x5 FILLER_304_565 ();
 b15zdnd11an1n04x5 FILLER_304_572 ();
 b15zdnd00an1n01x5 FILLER_304_576 ();
 b15zdnd11an1n64x5 FILLER_304_619 ();
 b15zdnd11an1n32x5 FILLER_304_683 ();
 b15zdnd00an1n02x5 FILLER_304_715 ();
 b15zdnd00an1n01x5 FILLER_304_717 ();
 b15zdnd11an1n64x5 FILLER_304_726 ();
 b15zdnd11an1n64x5 FILLER_304_790 ();
 b15zdnd11an1n08x5 FILLER_304_854 ();
 b15zdnd00an1n02x5 FILLER_304_862 ();
 b15zdnd11an1n64x5 FILLER_304_906 ();
 b15zdnd11an1n64x5 FILLER_304_970 ();
 b15zdnd11an1n64x5 FILLER_304_1034 ();
 b15zdnd11an1n64x5 FILLER_304_1098 ();
 b15zdnd11an1n64x5 FILLER_304_1162 ();
 b15zdnd11an1n04x5 FILLER_304_1226 ();
 b15zdnd00an1n02x5 FILLER_304_1230 ();
 b15zdnd11an1n04x5 FILLER_304_1235 ();
 b15zdnd11an1n64x5 FILLER_304_1242 ();
 b15zdnd11an1n08x5 FILLER_304_1306 ();
 b15zdnd00an1n02x5 FILLER_304_1314 ();
 b15zdnd00an1n01x5 FILLER_304_1316 ();
 b15zdnd11an1n64x5 FILLER_304_1328 ();
 b15zdnd11an1n64x5 FILLER_304_1392 ();
 b15zdnd11an1n64x5 FILLER_304_1456 ();
 b15zdnd11an1n64x5 FILLER_304_1520 ();
 b15zdnd11an1n64x5 FILLER_304_1584 ();
 b15zdnd11an1n32x5 FILLER_304_1648 ();
 b15zdnd11an1n16x5 FILLER_304_1680 ();
 b15zdnd11an1n08x5 FILLER_304_1696 ();
 b15zdnd00an1n02x5 FILLER_304_1704 ();
 b15zdnd00an1n01x5 FILLER_304_1706 ();
 b15zdnd11an1n08x5 FILLER_304_1710 ();
 b15zdnd11an1n64x5 FILLER_304_1745 ();
 b15zdnd11an1n64x5 FILLER_304_1809 ();
 b15zdnd11an1n64x5 FILLER_304_1873 ();
 b15zdnd11an1n04x5 FILLER_304_1937 ();
 b15zdnd00an1n01x5 FILLER_304_1941 ();
 b15zdnd11an1n04x5 FILLER_304_1945 ();
 b15zdnd00an1n01x5 FILLER_304_1949 ();
 b15zdnd11an1n64x5 FILLER_304_1977 ();
 b15zdnd11an1n64x5 FILLER_304_2041 ();
 b15zdnd11an1n32x5 FILLER_304_2105 ();
 b15zdnd11an1n16x5 FILLER_304_2137 ();
 b15zdnd00an1n01x5 FILLER_304_2153 ();
 b15zdnd11an1n64x5 FILLER_304_2162 ();
 b15zdnd11an1n32x5 FILLER_304_2226 ();
 b15zdnd11an1n16x5 FILLER_304_2258 ();
 b15zdnd00an1n02x5 FILLER_304_2274 ();
 b15zdnd11an1n04x5 FILLER_305_0 ();
 b15zdnd11an1n08x5 FILLER_305_10 ();
 b15zdnd11an1n04x5 FILLER_305_18 ();
 b15zdnd00an1n02x5 FILLER_305_22 ();
 b15zdnd00an1n01x5 FILLER_305_24 ();
 b15zdnd11an1n64x5 FILLER_305_30 ();
 b15zdnd11an1n64x5 FILLER_305_94 ();
 b15zdnd11an1n64x5 FILLER_305_158 ();
 b15zdnd11an1n64x5 FILLER_305_222 ();
 b15zdnd11an1n64x5 FILLER_305_286 ();
 b15zdnd11an1n64x5 FILLER_305_350 ();
 b15zdnd11an1n64x5 FILLER_305_427 ();
 b15zdnd11an1n64x5 FILLER_305_491 ();
 b15zdnd11an1n16x5 FILLER_305_555 ();
 b15zdnd11an1n08x5 FILLER_305_571 ();
 b15zdnd11an1n04x5 FILLER_305_579 ();
 b15zdnd00an1n01x5 FILLER_305_583 ();
 b15zdnd11an1n64x5 FILLER_305_636 ();
 b15zdnd11an1n32x5 FILLER_305_700 ();
 b15zdnd11an1n16x5 FILLER_305_732 ();
 b15zdnd11an1n08x5 FILLER_305_748 ();
 b15zdnd00an1n02x5 FILLER_305_756 ();
 b15zdnd11an1n64x5 FILLER_305_762 ();
 b15zdnd11an1n64x5 FILLER_305_826 ();
 b15zdnd11an1n64x5 FILLER_305_890 ();
 b15zdnd11an1n64x5 FILLER_305_954 ();
 b15zdnd11an1n64x5 FILLER_305_1018 ();
 b15zdnd11an1n64x5 FILLER_305_1082 ();
 b15zdnd11an1n64x5 FILLER_305_1146 ();
 b15zdnd11an1n04x5 FILLER_305_1210 ();
 b15zdnd00an1n02x5 FILLER_305_1214 ();
 b15zdnd00an1n01x5 FILLER_305_1216 ();
 b15zdnd11an1n64x5 FILLER_305_1261 ();
 b15zdnd11an1n64x5 FILLER_305_1325 ();
 b15zdnd11an1n64x5 FILLER_305_1389 ();
 b15zdnd11an1n64x5 FILLER_305_1453 ();
 b15zdnd11an1n64x5 FILLER_305_1517 ();
 b15zdnd11an1n64x5 FILLER_305_1581 ();
 b15zdnd11an1n32x5 FILLER_305_1645 ();
 b15zdnd11an1n04x5 FILLER_305_1677 ();
 b15zdnd00an1n01x5 FILLER_305_1681 ();
 b15zdnd11an1n64x5 FILLER_305_1734 ();
 b15zdnd11an1n64x5 FILLER_305_1798 ();
 b15zdnd11an1n64x5 FILLER_305_1862 ();
 b15zdnd11an1n16x5 FILLER_305_1926 ();
 b15zdnd11an1n08x5 FILLER_305_1942 ();
 b15zdnd11an1n04x5 FILLER_305_1950 ();
 b15zdnd11an1n64x5 FILLER_305_1962 ();
 b15zdnd11an1n64x5 FILLER_305_2026 ();
 b15zdnd11an1n04x5 FILLER_305_2090 ();
 b15zdnd11an1n64x5 FILLER_305_2100 ();
 b15zdnd11an1n64x5 FILLER_305_2164 ();
 b15zdnd11an1n32x5 FILLER_305_2228 ();
 b15zdnd11an1n16x5 FILLER_305_2260 ();
 b15zdnd11an1n08x5 FILLER_305_2276 ();
 b15zdnd11an1n08x5 FILLER_306_8 ();
 b15zdnd00an1n02x5 FILLER_306_16 ();
 b15zdnd00an1n01x5 FILLER_306_18 ();
 b15zdnd11an1n32x5 FILLER_306_24 ();
 b15zdnd11an1n08x5 FILLER_306_56 ();
 b15zdnd11an1n64x5 FILLER_306_76 ();
 b15zdnd11an1n64x5 FILLER_306_140 ();
 b15zdnd11an1n64x5 FILLER_306_204 ();
 b15zdnd11an1n64x5 FILLER_306_268 ();
 b15zdnd11an1n64x5 FILLER_306_332 ();
 b15zdnd11an1n64x5 FILLER_306_396 ();
 b15zdnd11an1n64x5 FILLER_306_460 ();
 b15zdnd11an1n64x5 FILLER_306_524 ();
 b15zdnd11an1n16x5 FILLER_306_588 ();
 b15zdnd11an1n04x5 FILLER_306_607 ();
 b15zdnd11an1n64x5 FILLER_306_614 ();
 b15zdnd11an1n32x5 FILLER_306_678 ();
 b15zdnd11an1n08x5 FILLER_306_710 ();
 b15zdnd11an1n64x5 FILLER_306_726 ();
 b15zdnd11an1n64x5 FILLER_306_790 ();
 b15zdnd11an1n64x5 FILLER_306_854 ();
 b15zdnd11an1n64x5 FILLER_306_918 ();
 b15zdnd11an1n64x5 FILLER_306_982 ();
 b15zdnd11an1n64x5 FILLER_306_1046 ();
 b15zdnd11an1n64x5 FILLER_306_1110 ();
 b15zdnd11an1n64x5 FILLER_306_1174 ();
 b15zdnd00an1n02x5 FILLER_306_1238 ();
 b15zdnd11an1n32x5 FILLER_306_1243 ();
 b15zdnd11an1n08x5 FILLER_306_1275 ();
 b15zdnd11an1n04x5 FILLER_306_1283 ();
 b15zdnd00an1n01x5 FILLER_306_1287 ();
 b15zdnd11an1n64x5 FILLER_306_1291 ();
 b15zdnd11an1n64x5 FILLER_306_1355 ();
 b15zdnd11an1n64x5 FILLER_306_1419 ();
 b15zdnd11an1n64x5 FILLER_306_1483 ();
 b15zdnd11an1n64x5 FILLER_306_1547 ();
 b15zdnd11an1n64x5 FILLER_306_1611 ();
 b15zdnd11an1n04x5 FILLER_306_1675 ();
 b15zdnd00an1n01x5 FILLER_306_1679 ();
 b15zdnd11an1n32x5 FILLER_306_1732 ();
 b15zdnd11an1n08x5 FILLER_306_1764 ();
 b15zdnd11an1n04x5 FILLER_306_1772 ();
 b15zdnd00an1n01x5 FILLER_306_1776 ();
 b15zdnd11an1n04x5 FILLER_306_1780 ();
 b15zdnd11an1n64x5 FILLER_306_1787 ();
 b15zdnd11an1n64x5 FILLER_306_1851 ();
 b15zdnd11an1n64x5 FILLER_306_1915 ();
 b15zdnd11an1n64x5 FILLER_306_1979 ();
 b15zdnd11an1n64x5 FILLER_306_2043 ();
 b15zdnd11an1n32x5 FILLER_306_2107 ();
 b15zdnd11an1n08x5 FILLER_306_2139 ();
 b15zdnd11an1n04x5 FILLER_306_2147 ();
 b15zdnd00an1n02x5 FILLER_306_2151 ();
 b15zdnd00an1n01x5 FILLER_306_2153 ();
 b15zdnd11an1n64x5 FILLER_306_2162 ();
 b15zdnd11an1n32x5 FILLER_306_2226 ();
 b15zdnd11an1n16x5 FILLER_306_2258 ();
 b15zdnd00an1n02x5 FILLER_306_2274 ();
 b15zdnd11an1n08x5 FILLER_307_0 ();
 b15zdnd11an1n04x5 FILLER_307_8 ();
 b15zdnd00an1n01x5 FILLER_307_12 ();
 b15zdnd11an1n08x5 FILLER_307_20 ();
 b15zdnd11an1n04x5 FILLER_307_28 ();
 b15zdnd00an1n02x5 FILLER_307_32 ();
 b15zdnd00an1n01x5 FILLER_307_34 ();
 b15zdnd11an1n04x5 FILLER_307_60 ();
 b15zdnd11an1n32x5 FILLER_307_74 ();
 b15zdnd11an1n64x5 FILLER_307_131 ();
 b15zdnd11an1n16x5 FILLER_307_195 ();
 b15zdnd11an1n08x5 FILLER_307_211 ();
 b15zdnd00an1n02x5 FILLER_307_219 ();
 b15zdnd11an1n08x5 FILLER_307_238 ();
 b15zdnd11an1n04x5 FILLER_307_246 ();
 b15zdnd00an1n01x5 FILLER_307_250 ();
 b15zdnd11an1n08x5 FILLER_307_255 ();
 b15zdnd11an1n04x5 FILLER_307_263 ();
 b15zdnd11an1n32x5 FILLER_307_287 ();
 b15zdnd11an1n16x5 FILLER_307_319 ();
 b15zdnd11an1n08x5 FILLER_307_335 ();
 b15zdnd00an1n02x5 FILLER_307_343 ();
 b15zdnd00an1n01x5 FILLER_307_345 ();
 b15zdnd11an1n04x5 FILLER_307_363 ();
 b15zdnd11an1n04x5 FILLER_307_379 ();
 b15zdnd11an1n64x5 FILLER_307_388 ();
 b15zdnd11an1n64x5 FILLER_307_452 ();
 b15zdnd11an1n64x5 FILLER_307_516 ();
 b15zdnd11an1n16x5 FILLER_307_580 ();
 b15zdnd11an1n08x5 FILLER_307_596 ();
 b15zdnd11an1n64x5 FILLER_307_607 ();
 b15zdnd11an1n64x5 FILLER_307_671 ();
 b15zdnd11an1n64x5 FILLER_307_735 ();
 b15zdnd11an1n64x5 FILLER_307_799 ();
 b15zdnd11an1n16x5 FILLER_307_863 ();
 b15zdnd11an1n04x5 FILLER_307_879 ();
 b15zdnd00an1n01x5 FILLER_307_883 ();
 b15zdnd11an1n64x5 FILLER_307_895 ();
 b15zdnd11an1n64x5 FILLER_307_959 ();
 b15zdnd11an1n64x5 FILLER_307_1023 ();
 b15zdnd11an1n64x5 FILLER_307_1087 ();
 b15zdnd11an1n64x5 FILLER_307_1151 ();
 b15zdnd11an1n64x5 FILLER_307_1215 ();
 b15zdnd11an1n32x5 FILLER_307_1279 ();
 b15zdnd00an1n02x5 FILLER_307_1311 ();
 b15zdnd00an1n01x5 FILLER_307_1313 ();
 b15zdnd11an1n64x5 FILLER_307_1323 ();
 b15zdnd11an1n64x5 FILLER_307_1387 ();
 b15zdnd11an1n64x5 FILLER_307_1451 ();
 b15zdnd11an1n64x5 FILLER_307_1515 ();
 b15zdnd11an1n32x5 FILLER_307_1579 ();
 b15zdnd11an1n16x5 FILLER_307_1611 ();
 b15zdnd11an1n04x5 FILLER_307_1627 ();
 b15zdnd00an1n02x5 FILLER_307_1631 ();
 b15zdnd11an1n32x5 FILLER_307_1637 ();
 b15zdnd11an1n16x5 FILLER_307_1669 ();
 b15zdnd11an1n08x5 FILLER_307_1685 ();
 b15zdnd11an1n04x5 FILLER_307_1693 ();
 b15zdnd00an1n01x5 FILLER_307_1697 ();
 b15zdnd11an1n04x5 FILLER_307_1701 ();
 b15zdnd11an1n04x5 FILLER_307_1708 ();
 b15zdnd11an1n04x5 FILLER_307_1715 ();
 b15zdnd11an1n32x5 FILLER_307_1722 ();
 b15zdnd11an1n04x5 FILLER_307_1754 ();
 b15zdnd00an1n01x5 FILLER_307_1758 ();
 b15zdnd11an1n64x5 FILLER_307_1811 ();
 b15zdnd11an1n32x5 FILLER_307_1875 ();
 b15zdnd11an1n08x5 FILLER_307_1907 ();
 b15zdnd11an1n04x5 FILLER_307_1915 ();
 b15zdnd00an1n02x5 FILLER_307_1919 ();
 b15zdnd11an1n64x5 FILLER_307_1963 ();
 b15zdnd11an1n64x5 FILLER_307_2027 ();
 b15zdnd11an1n64x5 FILLER_307_2091 ();
 b15zdnd11an1n64x5 FILLER_307_2155 ();
 b15zdnd11an1n64x5 FILLER_307_2219 ();
 b15zdnd00an1n01x5 FILLER_307_2283 ();
 b15zdnd00an1n02x5 FILLER_308_8 ();
 b15zdnd11an1n04x5 FILLER_308_17 ();
 b15zdnd00an1n02x5 FILLER_308_21 ();
 b15zdnd11an1n16x5 FILLER_308_31 ();
 b15zdnd11an1n08x5 FILLER_308_47 ();
 b15zdnd00an1n01x5 FILLER_308_55 ();
 b15zdnd11an1n64x5 FILLER_308_81 ();
 b15zdnd11an1n64x5 FILLER_308_145 ();
 b15zdnd11an1n08x5 FILLER_308_209 ();
 b15zdnd11an1n04x5 FILLER_308_217 ();
 b15zdnd00an1n01x5 FILLER_308_221 ();
 b15zdnd11an1n04x5 FILLER_308_225 ();
 b15zdnd11an1n32x5 FILLER_308_246 ();
 b15zdnd11an1n08x5 FILLER_308_278 ();
 b15zdnd00an1n01x5 FILLER_308_286 ();
 b15zdnd11an1n32x5 FILLER_308_307 ();
 b15zdnd11an1n08x5 FILLER_308_339 ();
 b15zdnd00an1n02x5 FILLER_308_347 ();
 b15zdnd11an1n04x5 FILLER_308_358 ();
 b15zdnd11an1n04x5 FILLER_308_372 ();
 b15zdnd11an1n64x5 FILLER_308_391 ();
 b15zdnd11an1n64x5 FILLER_308_455 ();
 b15zdnd11an1n64x5 FILLER_308_535 ();
 b15zdnd11an1n64x5 FILLER_308_599 ();
 b15zdnd11an1n32x5 FILLER_308_663 ();
 b15zdnd11an1n16x5 FILLER_308_695 ();
 b15zdnd11an1n04x5 FILLER_308_711 ();
 b15zdnd00an1n02x5 FILLER_308_715 ();
 b15zdnd00an1n01x5 FILLER_308_717 ();
 b15zdnd11an1n64x5 FILLER_308_726 ();
 b15zdnd11an1n64x5 FILLER_308_790 ();
 b15zdnd11an1n64x5 FILLER_308_854 ();
 b15zdnd11an1n64x5 FILLER_308_918 ();
 b15zdnd11an1n64x5 FILLER_308_982 ();
 b15zdnd11an1n64x5 FILLER_308_1046 ();
 b15zdnd11an1n64x5 FILLER_308_1110 ();
 b15zdnd11an1n64x5 FILLER_308_1174 ();
 b15zdnd11an1n64x5 FILLER_308_1238 ();
 b15zdnd11an1n04x5 FILLER_308_1302 ();
 b15zdnd00an1n02x5 FILLER_308_1306 ();
 b15zdnd11an1n64x5 FILLER_308_1320 ();
 b15zdnd11an1n32x5 FILLER_308_1384 ();
 b15zdnd11an1n16x5 FILLER_308_1416 ();
 b15zdnd11an1n04x5 FILLER_308_1432 ();
 b15zdnd00an1n02x5 FILLER_308_1436 ();
 b15zdnd00an1n01x5 FILLER_308_1438 ();
 b15zdnd11an1n64x5 FILLER_308_1453 ();
 b15zdnd11an1n64x5 FILLER_308_1517 ();
 b15zdnd11an1n64x5 FILLER_308_1581 ();
 b15zdnd11an1n32x5 FILLER_308_1645 ();
 b15zdnd11an1n16x5 FILLER_308_1677 ();
 b15zdnd11an1n08x5 FILLER_308_1693 ();
 b15zdnd00an1n02x5 FILLER_308_1701 ();
 b15zdnd00an1n01x5 FILLER_308_1703 ();
 b15zdnd11an1n04x5 FILLER_308_1707 ();
 b15zdnd11an1n64x5 FILLER_308_1714 ();
 b15zdnd11an1n04x5 FILLER_308_1778 ();
 b15zdnd00an1n02x5 FILLER_308_1782 ();
 b15zdnd11an1n08x5 FILLER_308_1787 ();
 b15zdnd00an1n02x5 FILLER_308_1795 ();
 b15zdnd00an1n01x5 FILLER_308_1797 ();
 b15zdnd11an1n64x5 FILLER_308_1802 ();
 b15zdnd11an1n04x5 FILLER_308_1866 ();
 b15zdnd00an1n02x5 FILLER_308_1870 ();
 b15zdnd11an1n64x5 FILLER_308_1889 ();
 b15zdnd11an1n32x5 FILLER_308_1953 ();
 b15zdnd11an1n08x5 FILLER_308_1985 ();
 b15zdnd11an1n04x5 FILLER_308_1993 ();
 b15zdnd00an1n02x5 FILLER_308_1997 ();
 b15zdnd00an1n01x5 FILLER_308_1999 ();
 b15zdnd11an1n32x5 FILLER_308_2006 ();
 b15zdnd11an1n16x5 FILLER_308_2038 ();
 b15zdnd00an1n02x5 FILLER_308_2054 ();
 b15zdnd11an1n64x5 FILLER_308_2059 ();
 b15zdnd11an1n16x5 FILLER_308_2123 ();
 b15zdnd11an1n08x5 FILLER_308_2139 ();
 b15zdnd11an1n04x5 FILLER_308_2147 ();
 b15zdnd00an1n02x5 FILLER_308_2151 ();
 b15zdnd00an1n01x5 FILLER_308_2153 ();
 b15zdnd11an1n64x5 FILLER_308_2162 ();
 b15zdnd11an1n32x5 FILLER_308_2226 ();
 b15zdnd11an1n16x5 FILLER_308_2258 ();
 b15zdnd00an1n02x5 FILLER_308_2274 ();
 b15zdnd11an1n08x5 FILLER_309_0 ();
 b15zdnd11an1n04x5 FILLER_309_8 ();
 b15zdnd00an1n02x5 FILLER_309_12 ();
 b15zdnd11an1n16x5 FILLER_309_21 ();
 b15zdnd11an1n16x5 FILLER_309_45 ();
 b15zdnd11an1n08x5 FILLER_309_61 ();
 b15zdnd11an1n04x5 FILLER_309_69 ();
 b15zdnd00an1n02x5 FILLER_309_73 ();
 b15zdnd11an1n64x5 FILLER_309_85 ();
 b15zdnd11an1n64x5 FILLER_309_149 ();
 b15zdnd11an1n32x5 FILLER_309_213 ();
 b15zdnd11an1n08x5 FILLER_309_245 ();
 b15zdnd00an1n01x5 FILLER_309_253 ();
 b15zdnd11an1n16x5 FILLER_309_259 ();
 b15zdnd11an1n08x5 FILLER_309_275 ();
 b15zdnd11an1n04x5 FILLER_309_283 ();
 b15zdnd00an1n01x5 FILLER_309_287 ();
 b15zdnd11an1n08x5 FILLER_309_319 ();
 b15zdnd11an1n04x5 FILLER_309_327 ();
 b15zdnd00an1n02x5 FILLER_309_331 ();
 b15zdnd11an1n16x5 FILLER_309_337 ();
 b15zdnd00an1n02x5 FILLER_309_353 ();
 b15zdnd11an1n04x5 FILLER_309_369 ();
 b15zdnd11an1n16x5 FILLER_309_376 ();
 b15zdnd00an1n01x5 FILLER_309_392 ();
 b15zdnd11an1n64x5 FILLER_309_407 ();
 b15zdnd11an1n64x5 FILLER_309_471 ();
 b15zdnd11an1n64x5 FILLER_309_535 ();
 b15zdnd11an1n64x5 FILLER_309_599 ();
 b15zdnd11an1n64x5 FILLER_309_663 ();
 b15zdnd11an1n64x5 FILLER_309_727 ();
 b15zdnd11an1n64x5 FILLER_309_791 ();
 b15zdnd11an1n64x5 FILLER_309_855 ();
 b15zdnd11an1n64x5 FILLER_309_919 ();
 b15zdnd11an1n64x5 FILLER_309_983 ();
 b15zdnd11an1n64x5 FILLER_309_1047 ();
 b15zdnd11an1n64x5 FILLER_309_1111 ();
 b15zdnd11an1n08x5 FILLER_309_1175 ();
 b15zdnd00an1n02x5 FILLER_309_1183 ();
 b15zdnd00an1n01x5 FILLER_309_1185 ();
 b15zdnd11an1n64x5 FILLER_309_1228 ();
 b15zdnd11an1n16x5 FILLER_309_1292 ();
 b15zdnd11an1n04x5 FILLER_309_1308 ();
 b15zdnd11an1n64x5 FILLER_309_1332 ();
 b15zdnd11an1n64x5 FILLER_309_1396 ();
 b15zdnd11an1n04x5 FILLER_309_1460 ();
 b15zdnd00an1n02x5 FILLER_309_1464 ();
 b15zdnd00an1n01x5 FILLER_309_1466 ();
 b15zdnd11an1n16x5 FILLER_309_1471 ();
 b15zdnd11an1n08x5 FILLER_309_1487 ();
 b15zdnd00an1n02x5 FILLER_309_1495 ();
 b15zdnd11an1n32x5 FILLER_309_1506 ();
 b15zdnd11an1n08x5 FILLER_309_1538 ();
 b15zdnd11an1n04x5 FILLER_309_1546 ();
 b15zdnd00an1n02x5 FILLER_309_1550 ();
 b15zdnd11an1n64x5 FILLER_309_1594 ();
 b15zdnd11an1n64x5 FILLER_309_1658 ();
 b15zdnd11an1n64x5 FILLER_309_1722 ();
 b15zdnd11an1n64x5 FILLER_309_1786 ();
 b15zdnd11an1n64x5 FILLER_309_1850 ();
 b15zdnd11an1n64x5 FILLER_309_1914 ();
 b15zdnd11an1n64x5 FILLER_309_1978 ();
 b15zdnd11an1n08x5 FILLER_309_2042 ();
 b15zdnd11an1n04x5 FILLER_309_2050 ();
 b15zdnd00an1n01x5 FILLER_309_2054 ();
 b15zdnd11an1n64x5 FILLER_309_2058 ();
 b15zdnd11an1n64x5 FILLER_309_2122 ();
 b15zdnd11an1n64x5 FILLER_309_2186 ();
 b15zdnd11an1n32x5 FILLER_309_2250 ();
 b15zdnd00an1n02x5 FILLER_309_2282 ();
 b15zdnd00an1n02x5 FILLER_310_8 ();
 b15zdnd00an1n01x5 FILLER_310_10 ();
 b15zdnd11an1n16x5 FILLER_310_19 ();
 b15zdnd11an1n64x5 FILLER_310_42 ();
 b15zdnd11an1n64x5 FILLER_310_106 ();
 b15zdnd11an1n64x5 FILLER_310_170 ();
 b15zdnd11an1n64x5 FILLER_310_234 ();
 b15zdnd00an1n01x5 FILLER_310_298 ();
 b15zdnd11an1n32x5 FILLER_310_309 ();
 b15zdnd11an1n16x5 FILLER_310_341 ();
 b15zdnd00an1n02x5 FILLER_310_357 ();
 b15zdnd00an1n01x5 FILLER_310_359 ();
 b15zdnd11an1n04x5 FILLER_310_370 ();
 b15zdnd11an1n64x5 FILLER_310_382 ();
 b15zdnd11an1n64x5 FILLER_310_446 ();
 b15zdnd11an1n64x5 FILLER_310_510 ();
 b15zdnd11an1n64x5 FILLER_310_574 ();
 b15zdnd11an1n32x5 FILLER_310_638 ();
 b15zdnd11an1n16x5 FILLER_310_670 ();
 b15zdnd00an1n02x5 FILLER_310_686 ();
 b15zdnd11an1n08x5 FILLER_310_696 ();
 b15zdnd11an1n04x5 FILLER_310_704 ();
 b15zdnd00an1n02x5 FILLER_310_716 ();
 b15zdnd11an1n32x5 FILLER_310_726 ();
 b15zdnd11an1n08x5 FILLER_310_758 ();
 b15zdnd11an1n64x5 FILLER_310_775 ();
 b15zdnd11an1n64x5 FILLER_310_839 ();
 b15zdnd11an1n64x5 FILLER_310_903 ();
 b15zdnd11an1n64x5 FILLER_310_967 ();
 b15zdnd11an1n64x5 FILLER_310_1031 ();
 b15zdnd11an1n64x5 FILLER_310_1095 ();
 b15zdnd11an1n64x5 FILLER_310_1159 ();
 b15zdnd00an1n02x5 FILLER_310_1223 ();
 b15zdnd11an1n64x5 FILLER_310_1233 ();
 b15zdnd11an1n32x5 FILLER_310_1297 ();
 b15zdnd00an1n02x5 FILLER_310_1329 ();
 b15zdnd11an1n64x5 FILLER_310_1345 ();
 b15zdnd11an1n16x5 FILLER_310_1409 ();
 b15zdnd11an1n08x5 FILLER_310_1425 ();
 b15zdnd11an1n04x5 FILLER_310_1433 ();
 b15zdnd00an1n02x5 FILLER_310_1437 ();
 b15zdnd11an1n32x5 FILLER_310_1453 ();
 b15zdnd11an1n04x5 FILLER_310_1485 ();
 b15zdnd00an1n01x5 FILLER_310_1489 ();
 b15zdnd11an1n64x5 FILLER_310_1498 ();
 b15zdnd11an1n64x5 FILLER_310_1562 ();
 b15zdnd11an1n64x5 FILLER_310_1626 ();
 b15zdnd11an1n64x5 FILLER_310_1690 ();
 b15zdnd11an1n64x5 FILLER_310_1754 ();
 b15zdnd11an1n32x5 FILLER_310_1818 ();
 b15zdnd11an1n16x5 FILLER_310_1850 ();
 b15zdnd11an1n08x5 FILLER_310_1866 ();
 b15zdnd00an1n02x5 FILLER_310_1874 ();
 b15zdnd11an1n64x5 FILLER_310_1918 ();
 b15zdnd11an1n08x5 FILLER_310_1982 ();
 b15zdnd11an1n04x5 FILLER_310_1990 ();
 b15zdnd00an1n01x5 FILLER_310_1994 ();
 b15zdnd11an1n04x5 FILLER_310_2026 ();
 b15zdnd11an1n32x5 FILLER_310_2082 ();
 b15zdnd11an1n16x5 FILLER_310_2114 ();
 b15zdnd11an1n08x5 FILLER_310_2130 ();
 b15zdnd11an1n04x5 FILLER_310_2138 ();
 b15zdnd11an1n08x5 FILLER_310_2145 ();
 b15zdnd00an1n01x5 FILLER_310_2153 ();
 b15zdnd11an1n16x5 FILLER_310_2162 ();
 b15zdnd00an1n02x5 FILLER_310_2178 ();
 b15zdnd11an1n04x5 FILLER_310_2183 ();
 b15zdnd11an1n64x5 FILLER_310_2190 ();
 b15zdnd11an1n16x5 FILLER_310_2254 ();
 b15zdnd11an1n04x5 FILLER_310_2270 ();
 b15zdnd00an1n02x5 FILLER_310_2274 ();
 b15zdnd11an1n64x5 FILLER_311_0 ();
 b15zdnd11an1n32x5 FILLER_311_64 ();
 b15zdnd11an1n08x5 FILLER_311_96 ();
 b15zdnd00an1n02x5 FILLER_311_104 ();
 b15zdnd00an1n01x5 FILLER_311_106 ();
 b15zdnd11an1n64x5 FILLER_311_138 ();
 b15zdnd11an1n64x5 FILLER_311_202 ();
 b15zdnd11an1n32x5 FILLER_311_266 ();
 b15zdnd11an1n16x5 FILLER_311_298 ();
 b15zdnd11an1n08x5 FILLER_311_314 ();
 b15zdnd00an1n02x5 FILLER_311_322 ();
 b15zdnd00an1n01x5 FILLER_311_324 ();
 b15zdnd11an1n16x5 FILLER_311_331 ();
 b15zdnd11an1n04x5 FILLER_311_347 ();
 b15zdnd00an1n02x5 FILLER_311_351 ();
 b15zdnd00an1n01x5 FILLER_311_353 ();
 b15zdnd11an1n04x5 FILLER_311_359 ();
 b15zdnd11an1n04x5 FILLER_311_369 ();
 b15zdnd11an1n64x5 FILLER_311_380 ();
 b15zdnd11an1n64x5 FILLER_311_444 ();
 b15zdnd11an1n64x5 FILLER_311_508 ();
 b15zdnd11an1n64x5 FILLER_311_572 ();
 b15zdnd11an1n64x5 FILLER_311_636 ();
 b15zdnd11an1n64x5 FILLER_311_700 ();
 b15zdnd11an1n64x5 FILLER_311_764 ();
 b15zdnd11an1n64x5 FILLER_311_828 ();
 b15zdnd11an1n64x5 FILLER_311_892 ();
 b15zdnd11an1n64x5 FILLER_311_956 ();
 b15zdnd11an1n64x5 FILLER_311_1020 ();
 b15zdnd11an1n64x5 FILLER_311_1084 ();
 b15zdnd11an1n64x5 FILLER_311_1148 ();
 b15zdnd11an1n64x5 FILLER_311_1212 ();
 b15zdnd11an1n32x5 FILLER_311_1276 ();
 b15zdnd11an1n16x5 FILLER_311_1308 ();
 b15zdnd11an1n08x5 FILLER_311_1324 ();
 b15zdnd11an1n64x5 FILLER_311_1374 ();
 b15zdnd11an1n64x5 FILLER_311_1441 ();
 b15zdnd11an1n64x5 FILLER_311_1505 ();
 b15zdnd11an1n64x5 FILLER_311_1569 ();
 b15zdnd11an1n64x5 FILLER_311_1633 ();
 b15zdnd11an1n64x5 FILLER_311_1697 ();
 b15zdnd11an1n64x5 FILLER_311_1761 ();
 b15zdnd11an1n32x5 FILLER_311_1825 ();
 b15zdnd11an1n16x5 FILLER_311_1857 ();
 b15zdnd00an1n02x5 FILLER_311_1873 ();
 b15zdnd00an1n01x5 FILLER_311_1875 ();
 b15zdnd11an1n64x5 FILLER_311_1928 ();
 b15zdnd11an1n32x5 FILLER_311_1992 ();
 b15zdnd11an1n16x5 FILLER_311_2024 ();
 b15zdnd11an1n08x5 FILLER_311_2040 ();
 b15zdnd11an1n04x5 FILLER_311_2048 ();
 b15zdnd00an1n02x5 FILLER_311_2052 ();
 b15zdnd00an1n01x5 FILLER_311_2054 ();
 b15zdnd11an1n32x5 FILLER_311_2058 ();
 b15zdnd11an1n16x5 FILLER_311_2090 ();
 b15zdnd11an1n08x5 FILLER_311_2106 ();
 b15zdnd11an1n16x5 FILLER_311_2120 ();
 b15zdnd11an1n04x5 FILLER_311_2136 ();
 b15zdnd00an1n02x5 FILLER_311_2140 ();
 b15zdnd11an1n08x5 FILLER_311_2149 ();
 b15zdnd11an1n04x5 FILLER_311_2157 ();
 b15zdnd00an1n01x5 FILLER_311_2161 ();
 b15zdnd11an1n64x5 FILLER_311_2214 ();
 b15zdnd11an1n04x5 FILLER_311_2278 ();
 b15zdnd00an1n02x5 FILLER_311_2282 ();
 b15zdnd11an1n64x5 FILLER_312_8 ();
 b15zdnd11an1n64x5 FILLER_312_72 ();
 b15zdnd11an1n64x5 FILLER_312_136 ();
 b15zdnd11an1n64x5 FILLER_312_200 ();
 b15zdnd11an1n16x5 FILLER_312_264 ();
 b15zdnd11an1n04x5 FILLER_312_280 ();
 b15zdnd00an1n01x5 FILLER_312_284 ();
 b15zdnd11an1n64x5 FILLER_312_289 ();
 b15zdnd11an1n64x5 FILLER_312_353 ();
 b15zdnd11an1n64x5 FILLER_312_417 ();
 b15zdnd11an1n64x5 FILLER_312_481 ();
 b15zdnd11an1n64x5 FILLER_312_545 ();
 b15zdnd11an1n16x5 FILLER_312_609 ();
 b15zdnd00an1n01x5 FILLER_312_625 ();
 b15zdnd11an1n64x5 FILLER_312_637 ();
 b15zdnd11an1n16x5 FILLER_312_701 ();
 b15zdnd00an1n01x5 FILLER_312_717 ();
 b15zdnd11an1n64x5 FILLER_312_726 ();
 b15zdnd11an1n64x5 FILLER_312_790 ();
 b15zdnd11an1n64x5 FILLER_312_854 ();
 b15zdnd11an1n64x5 FILLER_312_918 ();
 b15zdnd11an1n64x5 FILLER_312_982 ();
 b15zdnd11an1n64x5 FILLER_312_1046 ();
 b15zdnd11an1n64x5 FILLER_312_1110 ();
 b15zdnd11an1n64x5 FILLER_312_1174 ();
 b15zdnd11an1n16x5 FILLER_312_1238 ();
 b15zdnd11an1n08x5 FILLER_312_1254 ();
 b15zdnd11an1n04x5 FILLER_312_1262 ();
 b15zdnd00an1n02x5 FILLER_312_1266 ();
 b15zdnd00an1n01x5 FILLER_312_1268 ();
 b15zdnd11an1n32x5 FILLER_312_1286 ();
 b15zdnd11an1n08x5 FILLER_312_1318 ();
 b15zdnd11an1n04x5 FILLER_312_1326 ();
 b15zdnd00an1n02x5 FILLER_312_1330 ();
 b15zdnd11an1n64x5 FILLER_312_1339 ();
 b15zdnd11an1n32x5 FILLER_312_1403 ();
 b15zdnd11an1n16x5 FILLER_312_1435 ();
 b15zdnd11an1n64x5 FILLER_312_1454 ();
 b15zdnd11an1n64x5 FILLER_312_1518 ();
 b15zdnd11an1n64x5 FILLER_312_1582 ();
 b15zdnd11an1n64x5 FILLER_312_1646 ();
 b15zdnd11an1n64x5 FILLER_312_1710 ();
 b15zdnd11an1n64x5 FILLER_312_1774 ();
 b15zdnd11an1n32x5 FILLER_312_1838 ();
 b15zdnd11an1n16x5 FILLER_312_1870 ();
 b15zdnd11an1n08x5 FILLER_312_1886 ();
 b15zdnd11an1n04x5 FILLER_312_1897 ();
 b15zdnd11an1n64x5 FILLER_312_1904 ();
 b15zdnd11an1n64x5 FILLER_312_1968 ();
 b15zdnd11an1n64x5 FILLER_312_2032 ();
 b15zdnd11an1n08x5 FILLER_312_2096 ();
 b15zdnd11an1n04x5 FILLER_312_2104 ();
 b15zdnd00an1n02x5 FILLER_312_2108 ();
 b15zdnd00an1n01x5 FILLER_312_2110 ();
 b15zdnd11an1n04x5 FILLER_312_2124 ();
 b15zdnd00an1n02x5 FILLER_312_2128 ();
 b15zdnd11an1n08x5 FILLER_312_2143 ();
 b15zdnd00an1n02x5 FILLER_312_2151 ();
 b15zdnd00an1n01x5 FILLER_312_2153 ();
 b15zdnd00an1n02x5 FILLER_312_2162 ();
 b15zdnd11an1n64x5 FILLER_312_2206 ();
 b15zdnd11an1n04x5 FILLER_312_2270 ();
 b15zdnd00an1n02x5 FILLER_312_2274 ();
 b15zdnd11an1n64x5 FILLER_313_0 ();
 b15zdnd11an1n64x5 FILLER_313_64 ();
 b15zdnd11an1n64x5 FILLER_313_128 ();
 b15zdnd11an1n64x5 FILLER_313_192 ();
 b15zdnd11an1n16x5 FILLER_313_256 ();
 b15zdnd11an1n08x5 FILLER_313_272 ();
 b15zdnd00an1n02x5 FILLER_313_280 ();
 b15zdnd11an1n64x5 FILLER_313_294 ();
 b15zdnd11an1n64x5 FILLER_313_358 ();
 b15zdnd11an1n64x5 FILLER_313_422 ();
 b15zdnd11an1n64x5 FILLER_313_486 ();
 b15zdnd11an1n64x5 FILLER_313_550 ();
 b15zdnd11an1n64x5 FILLER_313_614 ();
 b15zdnd11an1n64x5 FILLER_313_678 ();
 b15zdnd11an1n64x5 FILLER_313_742 ();
 b15zdnd11an1n64x5 FILLER_313_806 ();
 b15zdnd11an1n64x5 FILLER_313_870 ();
 b15zdnd11an1n64x5 FILLER_313_934 ();
 b15zdnd11an1n64x5 FILLER_313_998 ();
 b15zdnd11an1n64x5 FILLER_313_1062 ();
 b15zdnd11an1n64x5 FILLER_313_1126 ();
 b15zdnd11an1n64x5 FILLER_313_1190 ();
 b15zdnd11an1n64x5 FILLER_313_1254 ();
 b15zdnd00an1n02x5 FILLER_313_1318 ();
 b15zdnd00an1n01x5 FILLER_313_1320 ();
 b15zdnd11an1n08x5 FILLER_313_1341 ();
 b15zdnd11an1n04x5 FILLER_313_1349 ();
 b15zdnd00an1n02x5 FILLER_313_1353 ();
 b15zdnd00an1n01x5 FILLER_313_1355 ();
 b15zdnd11an1n64x5 FILLER_313_1373 ();
 b15zdnd11an1n64x5 FILLER_313_1437 ();
 b15zdnd11an1n64x5 FILLER_313_1501 ();
 b15zdnd11an1n64x5 FILLER_313_1565 ();
 b15zdnd11an1n64x5 FILLER_313_1629 ();
 b15zdnd11an1n64x5 FILLER_313_1693 ();
 b15zdnd11an1n64x5 FILLER_313_1757 ();
 b15zdnd11an1n64x5 FILLER_313_1821 ();
 b15zdnd11an1n16x5 FILLER_313_1885 ();
 b15zdnd11an1n32x5 FILLER_313_1904 ();
 b15zdnd11an1n16x5 FILLER_313_1936 ();
 b15zdnd11an1n04x5 FILLER_313_1952 ();
 b15zdnd00an1n02x5 FILLER_313_1956 ();
 b15zdnd00an1n01x5 FILLER_313_1958 ();
 b15zdnd11an1n64x5 FILLER_313_2001 ();
 b15zdnd11an1n64x5 FILLER_313_2065 ();
 b15zdnd11an1n04x5 FILLER_313_2140 ();
 b15zdnd11an1n32x5 FILLER_313_2149 ();
 b15zdnd11an1n04x5 FILLER_313_2181 ();
 b15zdnd00an1n02x5 FILLER_313_2185 ();
 b15zdnd00an1n01x5 FILLER_313_2187 ();
 b15zdnd11an1n64x5 FILLER_313_2191 ();
 b15zdnd11an1n16x5 FILLER_313_2255 ();
 b15zdnd11an1n08x5 FILLER_313_2271 ();
 b15zdnd11an1n04x5 FILLER_313_2279 ();
 b15zdnd00an1n01x5 FILLER_313_2283 ();
 b15zdnd11an1n08x5 FILLER_314_8 ();
 b15zdnd00an1n02x5 FILLER_314_16 ();
 b15zdnd11an1n04x5 FILLER_314_24 ();
 b15zdnd11an1n64x5 FILLER_314_33 ();
 b15zdnd11an1n64x5 FILLER_314_97 ();
 b15zdnd11an1n16x5 FILLER_314_161 ();
 b15zdnd11an1n08x5 FILLER_314_177 ();
 b15zdnd11an1n04x5 FILLER_314_185 ();
 b15zdnd00an1n02x5 FILLER_314_189 ();
 b15zdnd00an1n01x5 FILLER_314_191 ();
 b15zdnd11an1n64x5 FILLER_314_197 ();
 b15zdnd11an1n16x5 FILLER_314_261 ();
 b15zdnd11an1n08x5 FILLER_314_277 ();
 b15zdnd11an1n04x5 FILLER_314_285 ();
 b15zdnd00an1n02x5 FILLER_314_289 ();
 b15zdnd11an1n64x5 FILLER_314_296 ();
 b15zdnd11an1n64x5 FILLER_314_360 ();
 b15zdnd11an1n64x5 FILLER_314_424 ();
 b15zdnd11an1n64x5 FILLER_314_488 ();
 b15zdnd11an1n64x5 FILLER_314_552 ();
 b15zdnd11an1n64x5 FILLER_314_616 ();
 b15zdnd11an1n32x5 FILLER_314_680 ();
 b15zdnd11an1n04x5 FILLER_314_712 ();
 b15zdnd00an1n02x5 FILLER_314_716 ();
 b15zdnd11an1n04x5 FILLER_314_726 ();
 b15zdnd00an1n02x5 FILLER_314_730 ();
 b15zdnd00an1n01x5 FILLER_314_732 ();
 b15zdnd11an1n32x5 FILLER_314_738 ();
 b15zdnd11an1n16x5 FILLER_314_770 ();
 b15zdnd11an1n04x5 FILLER_314_786 ();
 b15zdnd11an1n64x5 FILLER_314_832 ();
 b15zdnd11an1n64x5 FILLER_314_896 ();
 b15zdnd11an1n64x5 FILLER_314_960 ();
 b15zdnd11an1n64x5 FILLER_314_1024 ();
 b15zdnd11an1n64x5 FILLER_314_1088 ();
 b15zdnd11an1n64x5 FILLER_314_1152 ();
 b15zdnd11an1n64x5 FILLER_314_1216 ();
 b15zdnd11an1n64x5 FILLER_314_1280 ();
 b15zdnd00an1n02x5 FILLER_314_1344 ();
 b15zdnd00an1n01x5 FILLER_314_1346 ();
 b15zdnd11an1n64x5 FILLER_314_1389 ();
 b15zdnd11an1n64x5 FILLER_314_1453 ();
 b15zdnd11an1n64x5 FILLER_314_1517 ();
 b15zdnd11an1n64x5 FILLER_314_1581 ();
 b15zdnd11an1n64x5 FILLER_314_1645 ();
 b15zdnd11an1n64x5 FILLER_314_1709 ();
 b15zdnd11an1n64x5 FILLER_314_1773 ();
 b15zdnd11an1n64x5 FILLER_314_1837 ();
 b15zdnd11an1n64x5 FILLER_314_1901 ();
 b15zdnd11an1n64x5 FILLER_314_1965 ();
 b15zdnd11an1n32x5 FILLER_314_2029 ();
 b15zdnd11an1n16x5 FILLER_314_2061 ();
 b15zdnd11an1n04x5 FILLER_314_2077 ();
 b15zdnd00an1n01x5 FILLER_314_2081 ();
 b15zdnd11an1n16x5 FILLER_314_2124 ();
 b15zdnd11an1n08x5 FILLER_314_2140 ();
 b15zdnd11an1n04x5 FILLER_314_2148 ();
 b15zdnd00an1n02x5 FILLER_314_2152 ();
 b15zdnd11an1n64x5 FILLER_314_2162 ();
 b15zdnd11an1n32x5 FILLER_314_2226 ();
 b15zdnd11an1n16x5 FILLER_314_2258 ();
 b15zdnd00an1n02x5 FILLER_314_2274 ();
 b15zdnd11an1n32x5 FILLER_315_0 ();
 b15zdnd11an1n08x5 FILLER_315_32 ();
 b15zdnd11an1n64x5 FILLER_315_58 ();
 b15zdnd00an1n02x5 FILLER_315_122 ();
 b15zdnd11an1n64x5 FILLER_315_139 ();
 b15zdnd11an1n64x5 FILLER_315_203 ();
 b15zdnd11an1n64x5 FILLER_315_267 ();
 b15zdnd11an1n64x5 FILLER_315_331 ();
 b15zdnd11an1n64x5 FILLER_315_395 ();
 b15zdnd11an1n64x5 FILLER_315_459 ();
 b15zdnd11an1n64x5 FILLER_315_523 ();
 b15zdnd11an1n64x5 FILLER_315_587 ();
 b15zdnd11an1n32x5 FILLER_315_651 ();
 b15zdnd11an1n16x5 FILLER_315_683 ();
 b15zdnd11an1n04x5 FILLER_315_699 ();
 b15zdnd11an1n64x5 FILLER_315_716 ();
 b15zdnd11an1n64x5 FILLER_315_780 ();
 b15zdnd11an1n32x5 FILLER_315_844 ();
 b15zdnd11an1n16x5 FILLER_315_876 ();
 b15zdnd11an1n08x5 FILLER_315_892 ();
 b15zdnd11an1n04x5 FILLER_315_900 ();
 b15zdnd00an1n01x5 FILLER_315_904 ();
 b15zdnd11an1n64x5 FILLER_315_926 ();
 b15zdnd11an1n64x5 FILLER_315_990 ();
 b15zdnd00an1n02x5 FILLER_315_1054 ();
 b15zdnd00an1n01x5 FILLER_315_1056 ();
 b15zdnd11an1n04x5 FILLER_315_1060 ();
 b15zdnd11an1n64x5 FILLER_315_1067 ();
 b15zdnd11an1n64x5 FILLER_315_1131 ();
 b15zdnd11an1n64x5 FILLER_315_1195 ();
 b15zdnd11an1n64x5 FILLER_315_1259 ();
 b15zdnd11an1n32x5 FILLER_315_1323 ();
 b15zdnd11an1n04x5 FILLER_315_1355 ();
 b15zdnd00an1n02x5 FILLER_315_1359 ();
 b15zdnd11an1n32x5 FILLER_315_1369 ();
 b15zdnd11an1n64x5 FILLER_315_1415 ();
 b15zdnd11an1n64x5 FILLER_315_1479 ();
 b15zdnd11an1n16x5 FILLER_315_1543 ();
 b15zdnd11an1n08x5 FILLER_315_1559 ();
 b15zdnd00an1n02x5 FILLER_315_1567 ();
 b15zdnd00an1n01x5 FILLER_315_1569 ();
 b15zdnd11an1n04x5 FILLER_315_1577 ();
 b15zdnd11an1n16x5 FILLER_315_1588 ();
 b15zdnd11an1n04x5 FILLER_315_1604 ();
 b15zdnd00an1n02x5 FILLER_315_1608 ();
 b15zdnd11an1n32x5 FILLER_315_1652 ();
 b15zdnd00an1n02x5 FILLER_315_1684 ();
 b15zdnd11an1n64x5 FILLER_315_1728 ();
 b15zdnd11an1n64x5 FILLER_315_1792 ();
 b15zdnd11an1n64x5 FILLER_315_1856 ();
 b15zdnd11an1n64x5 FILLER_315_1920 ();
 b15zdnd11an1n64x5 FILLER_315_1984 ();
 b15zdnd11an1n08x5 FILLER_315_2048 ();
 b15zdnd00an1n02x5 FILLER_315_2056 ();
 b15zdnd11an1n32x5 FILLER_315_2100 ();
 b15zdnd00an1n02x5 FILLER_315_2132 ();
 b15zdnd11an1n64x5 FILLER_315_2141 ();
 b15zdnd11an1n64x5 FILLER_315_2205 ();
 b15zdnd11an1n08x5 FILLER_315_2269 ();
 b15zdnd11an1n04x5 FILLER_315_2277 ();
 b15zdnd00an1n02x5 FILLER_315_2281 ();
 b15zdnd00an1n01x5 FILLER_315_2283 ();
 b15zdnd11an1n64x5 FILLER_316_8 ();
 b15zdnd11an1n64x5 FILLER_316_72 ();
 b15zdnd11an1n64x5 FILLER_316_136 ();
 b15zdnd11an1n32x5 FILLER_316_200 ();
 b15zdnd00an1n02x5 FILLER_316_232 ();
 b15zdnd00an1n01x5 FILLER_316_234 ();
 b15zdnd11an1n64x5 FILLER_316_247 ();
 b15zdnd11an1n64x5 FILLER_316_311 ();
 b15zdnd11an1n64x5 FILLER_316_375 ();
 b15zdnd11an1n64x5 FILLER_316_439 ();
 b15zdnd11an1n64x5 FILLER_316_503 ();
 b15zdnd11an1n64x5 FILLER_316_567 ();
 b15zdnd11an1n64x5 FILLER_316_631 ();
 b15zdnd11an1n04x5 FILLER_316_695 ();
 b15zdnd00an1n01x5 FILLER_316_699 ();
 b15zdnd00an1n02x5 FILLER_316_715 ();
 b15zdnd00an1n01x5 FILLER_316_717 ();
 b15zdnd00an1n02x5 FILLER_316_726 ();
 b15zdnd11an1n32x5 FILLER_316_731 ();
 b15zdnd11an1n16x5 FILLER_316_763 ();
 b15zdnd11an1n64x5 FILLER_316_804 ();
 b15zdnd11an1n32x5 FILLER_316_868 ();
 b15zdnd11an1n16x5 FILLER_316_900 ();
 b15zdnd11an1n04x5 FILLER_316_916 ();
 b15zdnd11an1n64x5 FILLER_316_926 ();
 b15zdnd11an1n32x5 FILLER_316_990 ();
 b15zdnd11an1n08x5 FILLER_316_1022 ();
 b15zdnd11an1n04x5 FILLER_316_1030 ();
 b15zdnd00an1n02x5 FILLER_316_1034 ();
 b15zdnd11an1n64x5 FILLER_316_1088 ();
 b15zdnd11an1n64x5 FILLER_316_1152 ();
 b15zdnd11an1n64x5 FILLER_316_1216 ();
 b15zdnd11an1n64x5 FILLER_316_1280 ();
 b15zdnd11an1n64x5 FILLER_316_1344 ();
 b15zdnd11an1n64x5 FILLER_316_1408 ();
 b15zdnd11an1n64x5 FILLER_316_1472 ();
 b15zdnd11an1n08x5 FILLER_316_1536 ();
 b15zdnd00an1n02x5 FILLER_316_1544 ();
 b15zdnd00an1n01x5 FILLER_316_1546 ();
 b15zdnd11an1n04x5 FILLER_316_1589 ();
 b15zdnd11an1n64x5 FILLER_316_1596 ();
 b15zdnd11an1n64x5 FILLER_316_1660 ();
 b15zdnd11an1n64x5 FILLER_316_1724 ();
 b15zdnd11an1n64x5 FILLER_316_1788 ();
 b15zdnd11an1n64x5 FILLER_316_1852 ();
 b15zdnd11an1n64x5 FILLER_316_1916 ();
 b15zdnd11an1n64x5 FILLER_316_1980 ();
 b15zdnd11an1n32x5 FILLER_316_2044 ();
 b15zdnd11an1n16x5 FILLER_316_2076 ();
 b15zdnd11an1n08x5 FILLER_316_2092 ();
 b15zdnd00an1n02x5 FILLER_316_2100 ();
 b15zdnd00an1n01x5 FILLER_316_2102 ();
 b15zdnd11an1n08x5 FILLER_316_2145 ();
 b15zdnd00an1n01x5 FILLER_316_2153 ();
 b15zdnd11an1n64x5 FILLER_316_2162 ();
 b15zdnd11an1n32x5 FILLER_316_2226 ();
 b15zdnd11an1n16x5 FILLER_316_2258 ();
 b15zdnd00an1n02x5 FILLER_316_2274 ();
 b15zdnd11an1n16x5 FILLER_317_0 ();
 b15zdnd11an1n08x5 FILLER_317_16 ();
 b15zdnd11an1n64x5 FILLER_317_28 ();
 b15zdnd11an1n64x5 FILLER_317_92 ();
 b15zdnd11an1n32x5 FILLER_317_156 ();
 b15zdnd11an1n04x5 FILLER_317_188 ();
 b15zdnd00an1n01x5 FILLER_317_192 ();
 b15zdnd11an1n64x5 FILLER_317_224 ();
 b15zdnd11an1n64x5 FILLER_317_288 ();
 b15zdnd11an1n64x5 FILLER_317_352 ();
 b15zdnd11an1n64x5 FILLER_317_416 ();
 b15zdnd11an1n64x5 FILLER_317_480 ();
 b15zdnd11an1n64x5 FILLER_317_544 ();
 b15zdnd11an1n64x5 FILLER_317_608 ();
 b15zdnd11an1n16x5 FILLER_317_672 ();
 b15zdnd11an1n08x5 FILLER_317_688 ();
 b15zdnd11an1n04x5 FILLER_317_696 ();
 b15zdnd00an1n02x5 FILLER_317_700 ();
 b15zdnd11an1n16x5 FILLER_317_744 ();
 b15zdnd11an1n04x5 FILLER_317_760 ();
 b15zdnd11an1n64x5 FILLER_317_806 ();
 b15zdnd11an1n16x5 FILLER_317_870 ();
 b15zdnd11an1n04x5 FILLER_317_886 ();
 b15zdnd00an1n02x5 FILLER_317_890 ();
 b15zdnd00an1n01x5 FILLER_317_892 ();
 b15zdnd11an1n64x5 FILLER_317_896 ();
 b15zdnd11an1n64x5 FILLER_317_960 ();
 b15zdnd11an1n16x5 FILLER_317_1024 ();
 b15zdnd11an1n08x5 FILLER_317_1040 ();
 b15zdnd11an1n04x5 FILLER_317_1048 ();
 b15zdnd00an1n02x5 FILLER_317_1052 ();
 b15zdnd00an1n01x5 FILLER_317_1054 ();
 b15zdnd11an1n64x5 FILLER_317_1058 ();
 b15zdnd11an1n64x5 FILLER_317_1122 ();
 b15zdnd11an1n64x5 FILLER_317_1186 ();
 b15zdnd11an1n64x5 FILLER_317_1250 ();
 b15zdnd11an1n32x5 FILLER_317_1314 ();
 b15zdnd00an1n02x5 FILLER_317_1346 ();
 b15zdnd00an1n01x5 FILLER_317_1348 ();
 b15zdnd11an1n64x5 FILLER_317_1391 ();
 b15zdnd11an1n32x5 FILLER_317_1455 ();
 b15zdnd11an1n16x5 FILLER_317_1487 ();
 b15zdnd11an1n04x5 FILLER_317_1503 ();
 b15zdnd00an1n01x5 FILLER_317_1507 ();
 b15zdnd11an1n04x5 FILLER_317_1560 ();
 b15zdnd11an1n64x5 FILLER_317_1606 ();
 b15zdnd11an1n04x5 FILLER_317_1670 ();
 b15zdnd00an1n01x5 FILLER_317_1674 ();
 b15zdnd11an1n32x5 FILLER_317_1687 ();
 b15zdnd11an1n08x5 FILLER_317_1719 ();
 b15zdnd11an1n04x5 FILLER_317_1727 ();
 b15zdnd00an1n02x5 FILLER_317_1731 ();
 b15zdnd11an1n64x5 FILLER_317_1775 ();
 b15zdnd11an1n64x5 FILLER_317_1839 ();
 b15zdnd11an1n64x5 FILLER_317_1903 ();
 b15zdnd11an1n64x5 FILLER_317_1967 ();
 b15zdnd11an1n64x5 FILLER_317_2031 ();
 b15zdnd11an1n64x5 FILLER_317_2095 ();
 b15zdnd11an1n64x5 FILLER_317_2159 ();
 b15zdnd11an1n32x5 FILLER_317_2223 ();
 b15zdnd11an1n16x5 FILLER_317_2255 ();
 b15zdnd11an1n08x5 FILLER_317_2271 ();
 b15zdnd11an1n04x5 FILLER_317_2279 ();
 b15zdnd00an1n01x5 FILLER_317_2283 ();
 b15zdnd11an1n08x5 FILLER_318_8 ();
 b15zdnd00an1n02x5 FILLER_318_16 ();
 b15zdnd11an1n64x5 FILLER_318_36 ();
 b15zdnd11an1n16x5 FILLER_318_100 ();
 b15zdnd11an1n04x5 FILLER_318_116 ();
 b15zdnd00an1n02x5 FILLER_318_120 ();
 b15zdnd11an1n64x5 FILLER_318_153 ();
 b15zdnd11an1n64x5 FILLER_318_217 ();
 b15zdnd11an1n64x5 FILLER_318_281 ();
 b15zdnd11an1n64x5 FILLER_318_345 ();
 b15zdnd11an1n64x5 FILLER_318_409 ();
 b15zdnd11an1n64x5 FILLER_318_473 ();
 b15zdnd11an1n64x5 FILLER_318_537 ();
 b15zdnd11an1n64x5 FILLER_318_601 ();
 b15zdnd11an1n08x5 FILLER_318_665 ();
 b15zdnd11an1n04x5 FILLER_318_673 ();
 b15zdnd11an1n08x5 FILLER_318_680 ();
 b15zdnd11an1n04x5 FILLER_318_688 ();
 b15zdnd00an1n02x5 FILLER_318_692 ();
 b15zdnd00an1n01x5 FILLER_318_694 ();
 b15zdnd11an1n04x5 FILLER_318_700 ();
 b15zdnd00an1n02x5 FILLER_318_715 ();
 b15zdnd00an1n01x5 FILLER_318_717 ();
 b15zdnd11an1n08x5 FILLER_318_726 ();
 b15zdnd11an1n04x5 FILLER_318_750 ();
 b15zdnd11an1n04x5 FILLER_318_759 ();
 b15zdnd11an1n16x5 FILLER_318_767 ();
 b15zdnd11an1n08x5 FILLER_318_783 ();
 b15zdnd11an1n04x5 FILLER_318_791 ();
 b15zdnd00an1n01x5 FILLER_318_795 ();
 b15zdnd11an1n32x5 FILLER_318_838 ();
 b15zdnd11an1n16x5 FILLER_318_870 ();
 b15zdnd11an1n04x5 FILLER_318_886 ();
 b15zdnd00an1n02x5 FILLER_318_890 ();
 b15zdnd11an1n64x5 FILLER_318_934 ();
 b15zdnd11an1n64x5 FILLER_318_998 ();
 b15zdnd11an1n32x5 FILLER_318_1062 ();
 b15zdnd11an1n04x5 FILLER_318_1094 ();
 b15zdnd00an1n02x5 FILLER_318_1098 ();
 b15zdnd11an1n04x5 FILLER_318_1103 ();
 b15zdnd11an1n64x5 FILLER_318_1110 ();
 b15zdnd11an1n64x5 FILLER_318_1174 ();
 b15zdnd11an1n64x5 FILLER_318_1238 ();
 b15zdnd11an1n32x5 FILLER_318_1302 ();
 b15zdnd11an1n16x5 FILLER_318_1334 ();
 b15zdnd11an1n04x5 FILLER_318_1350 ();
 b15zdnd00an1n02x5 FILLER_318_1354 ();
 b15zdnd11an1n16x5 FILLER_318_1359 ();
 b15zdnd11an1n08x5 FILLER_318_1375 ();
 b15zdnd00an1n02x5 FILLER_318_1383 ();
 b15zdnd11an1n64x5 FILLER_318_1427 ();
 b15zdnd11an1n32x5 FILLER_318_1491 ();
 b15zdnd11an1n04x5 FILLER_318_1523 ();
 b15zdnd11an1n04x5 FILLER_318_1530 ();
 b15zdnd11an1n16x5 FILLER_318_1537 ();
 b15zdnd00an1n02x5 FILLER_318_1553 ();
 b15zdnd00an1n01x5 FILLER_318_1555 ();
 b15zdnd11an1n04x5 FILLER_318_1598 ();
 b15zdnd11an1n64x5 FILLER_318_1608 ();
 b15zdnd11an1n64x5 FILLER_318_1672 ();
 b15zdnd11an1n64x5 FILLER_318_1736 ();
 b15zdnd11an1n32x5 FILLER_318_1800 ();
 b15zdnd11an1n16x5 FILLER_318_1832 ();
 b15zdnd11an1n16x5 FILLER_318_1852 ();
 b15zdnd11an1n04x5 FILLER_318_1868 ();
 b15zdnd00an1n02x5 FILLER_318_1872 ();
 b15zdnd00an1n01x5 FILLER_318_1874 ();
 b15zdnd11an1n64x5 FILLER_318_1886 ();
 b15zdnd11an1n32x5 FILLER_318_1950 ();
 b15zdnd11an1n04x5 FILLER_318_1982 ();
 b15zdnd11an1n04x5 FILLER_318_1989 ();
 b15zdnd11an1n64x5 FILLER_318_1996 ();
 b15zdnd11an1n64x5 FILLER_318_2060 ();
 b15zdnd11an1n08x5 FILLER_318_2124 ();
 b15zdnd11an1n04x5 FILLER_318_2132 ();
 b15zdnd00an1n01x5 FILLER_318_2136 ();
 b15zdnd11an1n08x5 FILLER_318_2141 ();
 b15zdnd11an1n04x5 FILLER_318_2149 ();
 b15zdnd00an1n01x5 FILLER_318_2153 ();
 b15zdnd11an1n64x5 FILLER_318_2162 ();
 b15zdnd11an1n32x5 FILLER_318_2226 ();
 b15zdnd11an1n16x5 FILLER_318_2258 ();
 b15zdnd00an1n02x5 FILLER_318_2274 ();
 b15zdnd11an1n64x5 FILLER_319_0 ();
 b15zdnd11an1n32x5 FILLER_319_64 ();
 b15zdnd11an1n08x5 FILLER_319_96 ();
 b15zdnd11an1n04x5 FILLER_319_104 ();
 b15zdnd00an1n02x5 FILLER_319_108 ();
 b15zdnd00an1n01x5 FILLER_319_110 ();
 b15zdnd11an1n32x5 FILLER_319_129 ();
 b15zdnd11an1n04x5 FILLER_319_161 ();
 b15zdnd00an1n02x5 FILLER_319_165 ();
 b15zdnd00an1n01x5 FILLER_319_167 ();
 b15zdnd11an1n08x5 FILLER_319_199 ();
 b15zdnd11an1n64x5 FILLER_319_225 ();
 b15zdnd11an1n64x5 FILLER_319_289 ();
 b15zdnd11an1n64x5 FILLER_319_353 ();
 b15zdnd11an1n64x5 FILLER_319_417 ();
 b15zdnd11an1n64x5 FILLER_319_481 ();
 b15zdnd11an1n64x5 FILLER_319_545 ();
 b15zdnd11an1n32x5 FILLER_319_609 ();
 b15zdnd11an1n08x5 FILLER_319_641 ();
 b15zdnd11an1n04x5 FILLER_319_649 ();
 b15zdnd00an1n01x5 FILLER_319_653 ();
 b15zdnd11an1n04x5 FILLER_319_706 ();
 b15zdnd11an1n08x5 FILLER_319_752 ();
 b15zdnd00an1n02x5 FILLER_319_760 ();
 b15zdnd11an1n32x5 FILLER_319_814 ();
 b15zdnd11an1n08x5 FILLER_319_846 ();
 b15zdnd00an1n02x5 FILLER_319_854 ();
 b15zdnd11an1n04x5 FILLER_319_896 ();
 b15zdnd11an1n04x5 FILLER_319_903 ();
 b15zdnd11an1n64x5 FILLER_319_911 ();
 b15zdnd11an1n64x5 FILLER_319_975 ();
 b15zdnd11an1n32x5 FILLER_319_1039 ();
 b15zdnd11an1n08x5 FILLER_319_1071 ();
 b15zdnd00an1n01x5 FILLER_319_1079 ();
 b15zdnd11an1n04x5 FILLER_319_1132 ();
 b15zdnd11an1n04x5 FILLER_319_1146 ();
 b15zdnd00an1n01x5 FILLER_319_1150 ();
 b15zdnd11an1n64x5 FILLER_319_1165 ();
 b15zdnd11an1n64x5 FILLER_319_1229 ();
 b15zdnd11an1n32x5 FILLER_319_1293 ();
 b15zdnd11an1n16x5 FILLER_319_1325 ();
 b15zdnd11an1n08x5 FILLER_319_1341 ();
 b15zdnd11an1n04x5 FILLER_319_1349 ();
 b15zdnd00an1n02x5 FILLER_319_1353 ();
 b15zdnd00an1n01x5 FILLER_319_1355 ();
 b15zdnd11an1n64x5 FILLER_319_1359 ();
 b15zdnd11an1n64x5 FILLER_319_1423 ();
 b15zdnd11an1n32x5 FILLER_319_1487 ();
 b15zdnd11an1n08x5 FILLER_319_1519 ();
 b15zdnd11an1n04x5 FILLER_319_1527 ();
 b15zdnd11an1n16x5 FILLER_319_1534 ();
 b15zdnd11an1n08x5 FILLER_319_1550 ();
 b15zdnd11an1n04x5 FILLER_319_1558 ();
 b15zdnd00an1n02x5 FILLER_319_1562 ();
 b15zdnd11an1n04x5 FILLER_319_1577 ();
 b15zdnd11an1n04x5 FILLER_319_1590 ();
 b15zdnd11an1n04x5 FILLER_319_1599 ();
 b15zdnd11an1n64x5 FILLER_319_1607 ();
 b15zdnd11an1n64x5 FILLER_319_1671 ();
 b15zdnd11an1n04x5 FILLER_319_1735 ();
 b15zdnd00an1n02x5 FILLER_319_1739 ();
 b15zdnd00an1n01x5 FILLER_319_1741 ();
 b15zdnd11an1n64x5 FILLER_319_1784 ();
 b15zdnd11an1n64x5 FILLER_319_1848 ();
 b15zdnd11an1n32x5 FILLER_319_1912 ();
 b15zdnd11an1n08x5 FILLER_319_1944 ();
 b15zdnd00an1n02x5 FILLER_319_1952 ();
 b15zdnd00an1n01x5 FILLER_319_1954 ();
 b15zdnd11an1n64x5 FILLER_319_1995 ();
 b15zdnd11an1n04x5 FILLER_319_2059 ();
 b15zdnd11an1n64x5 FILLER_319_2115 ();
 b15zdnd11an1n64x5 FILLER_319_2179 ();
 b15zdnd11an1n32x5 FILLER_319_2243 ();
 b15zdnd11an1n08x5 FILLER_319_2275 ();
 b15zdnd00an1n01x5 FILLER_319_2283 ();
 b15zdnd11an1n64x5 FILLER_320_8 ();
 b15zdnd11an1n64x5 FILLER_320_72 ();
 b15zdnd11an1n64x5 FILLER_320_136 ();
 b15zdnd11an1n64x5 FILLER_320_200 ();
 b15zdnd11an1n64x5 FILLER_320_264 ();
 b15zdnd11an1n64x5 FILLER_320_328 ();
 b15zdnd11an1n64x5 FILLER_320_392 ();
 b15zdnd11an1n64x5 FILLER_320_456 ();
 b15zdnd11an1n64x5 FILLER_320_520 ();
 b15zdnd11an1n64x5 FILLER_320_584 ();
 b15zdnd11an1n16x5 FILLER_320_648 ();
 b15zdnd11an1n08x5 FILLER_320_664 ();
 b15zdnd00an1n01x5 FILLER_320_672 ();
 b15zdnd11an1n04x5 FILLER_320_676 ();
 b15zdnd11an1n16x5 FILLER_320_683 ();
 b15zdnd11an1n04x5 FILLER_320_703 ();
 b15zdnd11an1n04x5 FILLER_320_714 ();
 b15zdnd11an1n08x5 FILLER_320_726 ();
 b15zdnd11an1n04x5 FILLER_320_734 ();
 b15zdnd00an1n01x5 FILLER_320_738 ();
 b15zdnd11an1n16x5 FILLER_320_747 ();
 b15zdnd11an1n04x5 FILLER_320_763 ();
 b15zdnd00an1n02x5 FILLER_320_767 ();
 b15zdnd00an1n01x5 FILLER_320_769 ();
 b15zdnd11an1n64x5 FILLER_320_812 ();
 b15zdnd11an1n08x5 FILLER_320_876 ();
 b15zdnd00an1n02x5 FILLER_320_884 ();
 b15zdnd00an1n01x5 FILLER_320_886 ();
 b15zdnd11an1n64x5 FILLER_320_896 ();
 b15zdnd11an1n64x5 FILLER_320_960 ();
 b15zdnd11an1n64x5 FILLER_320_1024 ();
 b15zdnd11an1n08x5 FILLER_320_1088 ();
 b15zdnd11an1n04x5 FILLER_320_1096 ();
 b15zdnd00an1n02x5 FILLER_320_1100 ();
 b15zdnd11an1n08x5 FILLER_320_1105 ();
 b15zdnd00an1n02x5 FILLER_320_1113 ();
 b15zdnd00an1n01x5 FILLER_320_1115 ();
 b15zdnd11an1n32x5 FILLER_320_1158 ();
 b15zdnd11an1n64x5 FILLER_320_1203 ();
 b15zdnd11an1n64x5 FILLER_320_1267 ();
 b15zdnd00an1n02x5 FILLER_320_1331 ();
 b15zdnd00an1n01x5 FILLER_320_1333 ();
 b15zdnd11an1n64x5 FILLER_320_1378 ();
 b15zdnd11an1n64x5 FILLER_320_1442 ();
 b15zdnd11an1n64x5 FILLER_320_1506 ();
 b15zdnd11an1n08x5 FILLER_320_1570 ();
 b15zdnd00an1n02x5 FILLER_320_1578 ();
 b15zdnd11an1n64x5 FILLER_320_1622 ();
 b15zdnd11an1n64x5 FILLER_320_1686 ();
 b15zdnd11an1n64x5 FILLER_320_1750 ();
 b15zdnd11an1n64x5 FILLER_320_1814 ();
 b15zdnd11an1n64x5 FILLER_320_1878 ();
 b15zdnd11an1n64x5 FILLER_320_1942 ();
 b15zdnd11an1n64x5 FILLER_320_2006 ();
 b15zdnd11an1n16x5 FILLER_320_2070 ();
 b15zdnd11an1n64x5 FILLER_320_2089 ();
 b15zdnd00an1n01x5 FILLER_320_2153 ();
 b15zdnd11an1n64x5 FILLER_320_2162 ();
 b15zdnd11an1n32x5 FILLER_320_2226 ();
 b15zdnd11an1n16x5 FILLER_320_2258 ();
 b15zdnd00an1n02x5 FILLER_320_2274 ();
 b15zdnd11an1n64x5 FILLER_321_0 ();
 b15zdnd11an1n64x5 FILLER_321_64 ();
 b15zdnd11an1n64x5 FILLER_321_128 ();
 b15zdnd11an1n64x5 FILLER_321_192 ();
 b15zdnd11an1n64x5 FILLER_321_256 ();
 b15zdnd11an1n64x5 FILLER_321_320 ();
 b15zdnd11an1n64x5 FILLER_321_384 ();
 b15zdnd11an1n08x5 FILLER_321_448 ();
 b15zdnd11an1n04x5 FILLER_321_456 ();
 b15zdnd11an1n16x5 FILLER_321_471 ();
 b15zdnd11an1n08x5 FILLER_321_487 ();
 b15zdnd11an1n64x5 FILLER_321_547 ();
 b15zdnd11an1n64x5 FILLER_321_611 ();
 b15zdnd11an1n64x5 FILLER_321_675 ();
 b15zdnd11an1n32x5 FILLER_321_739 ();
 b15zdnd11an1n08x5 FILLER_321_771 ();
 b15zdnd00an1n02x5 FILLER_321_779 ();
 b15zdnd00an1n01x5 FILLER_321_781 ();
 b15zdnd11an1n04x5 FILLER_321_785 ();
 b15zdnd11an1n32x5 FILLER_321_792 ();
 b15zdnd11an1n16x5 FILLER_321_824 ();
 b15zdnd11an1n08x5 FILLER_321_840 ();
 b15zdnd00an1n01x5 FILLER_321_848 ();
 b15zdnd11an1n08x5 FILLER_321_858 ();
 b15zdnd11an1n04x5 FILLER_321_866 ();
 b15zdnd00an1n02x5 FILLER_321_870 ();
 b15zdnd00an1n01x5 FILLER_321_872 ();
 b15zdnd11an1n64x5 FILLER_321_925 ();
 b15zdnd11an1n64x5 FILLER_321_989 ();
 b15zdnd11an1n32x5 FILLER_321_1053 ();
 b15zdnd11an1n16x5 FILLER_321_1085 ();
 b15zdnd11an1n04x5 FILLER_321_1101 ();
 b15zdnd00an1n02x5 FILLER_321_1105 ();
 b15zdnd00an1n01x5 FILLER_321_1107 ();
 b15zdnd11an1n04x5 FILLER_321_1150 ();
 b15zdnd11an1n04x5 FILLER_321_1164 ();
 b15zdnd11an1n16x5 FILLER_321_1171 ();
 b15zdnd11an1n08x5 FILLER_321_1187 ();
 b15zdnd11an1n04x5 FILLER_321_1195 ();
 b15zdnd00an1n01x5 FILLER_321_1199 ();
 b15zdnd11an1n64x5 FILLER_321_1214 ();
 b15zdnd11an1n08x5 FILLER_321_1278 ();
 b15zdnd11an1n04x5 FILLER_321_1286 ();
 b15zdnd00an1n02x5 FILLER_321_1290 ();
 b15zdnd11an1n32x5 FILLER_321_1323 ();
 b15zdnd00an1n02x5 FILLER_321_1355 ();
 b15zdnd11an1n16x5 FILLER_321_1360 ();
 b15zdnd11an1n04x5 FILLER_321_1376 ();
 b15zdnd11an1n04x5 FILLER_321_1383 ();
 b15zdnd11an1n64x5 FILLER_321_1390 ();
 b15zdnd11an1n64x5 FILLER_321_1454 ();
 b15zdnd11an1n32x5 FILLER_321_1518 ();
 b15zdnd11an1n16x5 FILLER_321_1550 ();
 b15zdnd00an1n01x5 FILLER_321_1566 ();
 b15zdnd11an1n04x5 FILLER_321_1576 ();
 b15zdnd11an1n04x5 FILLER_321_1590 ();
 b15zdnd11an1n04x5 FILLER_321_1599 ();
 b15zdnd11an1n64x5 FILLER_321_1606 ();
 b15zdnd11an1n64x5 FILLER_321_1670 ();
 b15zdnd11an1n32x5 FILLER_321_1734 ();
 b15zdnd11an1n04x5 FILLER_321_1766 ();
 b15zdnd00an1n02x5 FILLER_321_1770 ();
 b15zdnd00an1n01x5 FILLER_321_1772 ();
 b15zdnd11an1n16x5 FILLER_321_1815 ();
 b15zdnd11an1n64x5 FILLER_321_1873 ();
 b15zdnd11an1n64x5 FILLER_321_1937 ();
 b15zdnd11an1n64x5 FILLER_321_2001 ();
 b15zdnd11an1n16x5 FILLER_321_2065 ();
 b15zdnd11an1n04x5 FILLER_321_2081 ();
 b15zdnd00an1n01x5 FILLER_321_2085 ();
 b15zdnd11an1n04x5 FILLER_321_2089 ();
 b15zdnd11an1n64x5 FILLER_321_2096 ();
 b15zdnd11an1n64x5 FILLER_321_2160 ();
 b15zdnd11an1n32x5 FILLER_321_2224 ();
 b15zdnd11an1n16x5 FILLER_321_2256 ();
 b15zdnd11an1n08x5 FILLER_321_2272 ();
 b15zdnd11an1n04x5 FILLER_321_2280 ();
 b15zdnd11an1n64x5 FILLER_322_8 ();
 b15zdnd11an1n64x5 FILLER_322_72 ();
 b15zdnd11an1n64x5 FILLER_322_136 ();
 b15zdnd11an1n64x5 FILLER_322_200 ();
 b15zdnd11an1n64x5 FILLER_322_264 ();
 b15zdnd11an1n64x5 FILLER_322_328 ();
 b15zdnd11an1n64x5 FILLER_322_392 ();
 b15zdnd11an1n32x5 FILLER_322_456 ();
 b15zdnd11an1n16x5 FILLER_322_488 ();
 b15zdnd11an1n08x5 FILLER_322_504 ();
 b15zdnd00an1n02x5 FILLER_322_512 ();
 b15zdnd00an1n01x5 FILLER_322_514 ();
 b15zdnd11an1n04x5 FILLER_322_518 ();
 b15zdnd11an1n04x5 FILLER_322_525 ();
 b15zdnd11an1n64x5 FILLER_322_532 ();
 b15zdnd11an1n64x5 FILLER_322_596 ();
 b15zdnd11an1n32x5 FILLER_322_660 ();
 b15zdnd11an1n16x5 FILLER_322_692 ();
 b15zdnd11an1n08x5 FILLER_322_708 ();
 b15zdnd00an1n02x5 FILLER_322_716 ();
 b15zdnd11an1n32x5 FILLER_322_726 ();
 b15zdnd11an1n16x5 FILLER_322_758 ();
 b15zdnd11an1n08x5 FILLER_322_774 ();
 b15zdnd00an1n01x5 FILLER_322_782 ();
 b15zdnd11an1n64x5 FILLER_322_786 ();
 b15zdnd11an1n32x5 FILLER_322_850 ();
 b15zdnd11an1n04x5 FILLER_322_882 ();
 b15zdnd00an1n02x5 FILLER_322_886 ();
 b15zdnd00an1n01x5 FILLER_322_888 ();
 b15zdnd11an1n64x5 FILLER_322_931 ();
 b15zdnd11an1n64x5 FILLER_322_995 ();
 b15zdnd11an1n64x5 FILLER_322_1059 ();
 b15zdnd11an1n08x5 FILLER_322_1123 ();
 b15zdnd11an1n04x5 FILLER_322_1131 ();
 b15zdnd00an1n02x5 FILLER_322_1135 ();
 b15zdnd00an1n01x5 FILLER_322_1137 ();
 b15zdnd11an1n16x5 FILLER_322_1143 ();
 b15zdnd11an1n08x5 FILLER_322_1159 ();
 b15zdnd11an1n04x5 FILLER_322_1167 ();
 b15zdnd00an1n02x5 FILLER_322_1171 ();
 b15zdnd11an1n64x5 FILLER_322_1215 ();
 b15zdnd11an1n64x5 FILLER_322_1279 ();
 b15zdnd11an1n16x5 FILLER_322_1343 ();
 b15zdnd00an1n02x5 FILLER_322_1359 ();
 b15zdnd00an1n01x5 FILLER_322_1361 ();
 b15zdnd11an1n64x5 FILLER_322_1414 ();
 b15zdnd11an1n32x5 FILLER_322_1478 ();
 b15zdnd11an1n16x5 FILLER_322_1510 ();
 b15zdnd11an1n08x5 FILLER_322_1526 ();
 b15zdnd11an1n04x5 FILLER_322_1534 ();
 b15zdnd00an1n02x5 FILLER_322_1538 ();
 b15zdnd11an1n32x5 FILLER_322_1548 ();
 b15zdnd11an1n04x5 FILLER_322_1580 ();
 b15zdnd00an1n02x5 FILLER_322_1584 ();
 b15zdnd11an1n64x5 FILLER_322_1592 ();
 b15zdnd11an1n64x5 FILLER_322_1656 ();
 b15zdnd11an1n64x5 FILLER_322_1720 ();
 b15zdnd11an1n64x5 FILLER_322_1784 ();
 b15zdnd11an1n64x5 FILLER_322_1848 ();
 b15zdnd11an1n64x5 FILLER_322_1912 ();
 b15zdnd11an1n64x5 FILLER_322_1976 ();
 b15zdnd11an1n64x5 FILLER_322_2040 ();
 b15zdnd11an1n32x5 FILLER_322_2104 ();
 b15zdnd11an1n16x5 FILLER_322_2136 ();
 b15zdnd00an1n02x5 FILLER_322_2152 ();
 b15zdnd11an1n64x5 FILLER_322_2162 ();
 b15zdnd11an1n32x5 FILLER_322_2226 ();
 b15zdnd11an1n08x5 FILLER_322_2262 ();
 b15zdnd11an1n04x5 FILLER_322_2270 ();
 b15zdnd00an1n02x5 FILLER_322_2274 ();
 b15zdnd11an1n64x5 FILLER_323_0 ();
 b15zdnd11an1n32x5 FILLER_323_64 ();
 b15zdnd11an1n16x5 FILLER_323_96 ();
 b15zdnd11an1n04x5 FILLER_323_112 ();
 b15zdnd11an1n64x5 FILLER_323_140 ();
 b15zdnd11an1n64x5 FILLER_323_204 ();
 b15zdnd11an1n64x5 FILLER_323_268 ();
 b15zdnd11an1n64x5 FILLER_323_332 ();
 b15zdnd11an1n64x5 FILLER_323_396 ();
 b15zdnd11an1n64x5 FILLER_323_460 ();
 b15zdnd11an1n16x5 FILLER_323_524 ();
 b15zdnd11an1n04x5 FILLER_323_540 ();
 b15zdnd00an1n01x5 FILLER_323_544 ();
 b15zdnd11an1n16x5 FILLER_323_587 ();
 b15zdnd11an1n64x5 FILLER_323_606 ();
 b15zdnd11an1n64x5 FILLER_323_670 ();
 b15zdnd11an1n32x5 FILLER_323_734 ();
 b15zdnd11an1n16x5 FILLER_323_766 ();
 b15zdnd00an1n02x5 FILLER_323_782 ();
 b15zdnd11an1n04x5 FILLER_323_826 ();
 b15zdnd11an1n16x5 FILLER_323_872 ();
 b15zdnd11an1n04x5 FILLER_323_888 ();
 b15zdnd00an1n01x5 FILLER_323_892 ();
 b15zdnd11an1n04x5 FILLER_323_896 ();
 b15zdnd11an1n04x5 FILLER_323_903 ();
 b15zdnd11an1n64x5 FILLER_323_910 ();
 b15zdnd11an1n64x5 FILLER_323_974 ();
 b15zdnd11an1n64x5 FILLER_323_1038 ();
 b15zdnd11an1n64x5 FILLER_323_1102 ();
 b15zdnd11an1n16x5 FILLER_323_1166 ();
 b15zdnd11an1n08x5 FILLER_323_1182 ();
 b15zdnd00an1n02x5 FILLER_323_1190 ();
 b15zdnd11an1n04x5 FILLER_323_1198 ();
 b15zdnd11an1n64x5 FILLER_323_1206 ();
 b15zdnd11an1n64x5 FILLER_323_1270 ();
 b15zdnd11an1n32x5 FILLER_323_1334 ();
 b15zdnd11an1n16x5 FILLER_323_1366 ();
 b15zdnd11an1n04x5 FILLER_323_1382 ();
 b15zdnd00an1n01x5 FILLER_323_1386 ();
 b15zdnd11an1n64x5 FILLER_323_1390 ();
 b15zdnd11an1n32x5 FILLER_323_1454 ();
 b15zdnd11an1n16x5 FILLER_323_1486 ();
 b15zdnd11an1n04x5 FILLER_323_1502 ();
 b15zdnd00an1n02x5 FILLER_323_1506 ();
 b15zdnd00an1n01x5 FILLER_323_1508 ();
 b15zdnd11an1n64x5 FILLER_323_1548 ();
 b15zdnd11an1n64x5 FILLER_323_1612 ();
 b15zdnd11an1n64x5 FILLER_323_1676 ();
 b15zdnd11an1n64x5 FILLER_323_1740 ();
 b15zdnd11an1n64x5 FILLER_323_1804 ();
 b15zdnd11an1n64x5 FILLER_323_1868 ();
 b15zdnd11an1n64x5 FILLER_323_1932 ();
 b15zdnd11an1n64x5 FILLER_323_1996 ();
 b15zdnd11an1n64x5 FILLER_323_2060 ();
 b15zdnd11an1n64x5 FILLER_323_2124 ();
 b15zdnd11an1n64x5 FILLER_323_2188 ();
 b15zdnd11an1n16x5 FILLER_323_2252 ();
 b15zdnd11an1n08x5 FILLER_323_2268 ();
 b15zdnd00an1n02x5 FILLER_323_2276 ();
 b15zdnd00an1n02x5 FILLER_323_2282 ();
 b15zdnd11an1n16x5 FILLER_324_8 ();
 b15zdnd11an1n08x5 FILLER_324_24 ();
 b15zdnd11an1n04x5 FILLER_324_32 ();
 b15zdnd00an1n02x5 FILLER_324_36 ();
 b15zdnd11an1n16x5 FILLER_324_63 ();
 b15zdnd11an1n64x5 FILLER_324_97 ();
 b15zdnd11an1n64x5 FILLER_324_161 ();
 b15zdnd11an1n64x5 FILLER_324_225 ();
 b15zdnd11an1n64x5 FILLER_324_289 ();
 b15zdnd11an1n64x5 FILLER_324_353 ();
 b15zdnd11an1n64x5 FILLER_324_417 ();
 b15zdnd11an1n08x5 FILLER_324_481 ();
 b15zdnd11an1n04x5 FILLER_324_489 ();
 b15zdnd00an1n02x5 FILLER_324_493 ();
 b15zdnd00an1n01x5 FILLER_324_495 ();
 b15zdnd11an1n04x5 FILLER_324_538 ();
 b15zdnd00an1n02x5 FILLER_324_542 ();
 b15zdnd11an1n04x5 FILLER_324_569 ();
 b15zdnd00an1n02x5 FILLER_324_573 ();
 b15zdnd00an1n01x5 FILLER_324_575 ();
 b15zdnd11an1n64x5 FILLER_324_628 ();
 b15zdnd11an1n16x5 FILLER_324_692 ();
 b15zdnd11an1n08x5 FILLER_324_708 ();
 b15zdnd00an1n02x5 FILLER_324_716 ();
 b15zdnd11an1n64x5 FILLER_324_726 ();
 b15zdnd11an1n64x5 FILLER_324_790 ();
 b15zdnd11an1n64x5 FILLER_324_854 ();
 b15zdnd11an1n64x5 FILLER_324_918 ();
 b15zdnd11an1n64x5 FILLER_324_982 ();
 b15zdnd11an1n64x5 FILLER_324_1046 ();
 b15zdnd11an1n64x5 FILLER_324_1110 ();
 b15zdnd11an1n32x5 FILLER_324_1174 ();
 b15zdnd00an1n01x5 FILLER_324_1206 ();
 b15zdnd11an1n32x5 FILLER_324_1212 ();
 b15zdnd11an1n16x5 FILLER_324_1244 ();
 b15zdnd11an1n08x5 FILLER_324_1260 ();
 b15zdnd00an1n01x5 FILLER_324_1268 ();
 b15zdnd11an1n08x5 FILLER_324_1300 ();
 b15zdnd11an1n04x5 FILLER_324_1308 ();
 b15zdnd00an1n02x5 FILLER_324_1312 ();
 b15zdnd00an1n01x5 FILLER_324_1314 ();
 b15zdnd11an1n08x5 FILLER_324_1322 ();
 b15zdnd00an1n02x5 FILLER_324_1330 ();
 b15zdnd11an1n64x5 FILLER_324_1339 ();
 b15zdnd11an1n64x5 FILLER_324_1403 ();
 b15zdnd11an1n32x5 FILLER_324_1467 ();
 b15zdnd11an1n16x5 FILLER_324_1499 ();
 b15zdnd11an1n04x5 FILLER_324_1515 ();
 b15zdnd11an1n64x5 FILLER_324_1526 ();
 b15zdnd11an1n08x5 FILLER_324_1590 ();
 b15zdnd11an1n04x5 FILLER_324_1598 ();
 b15zdnd00an1n02x5 FILLER_324_1602 ();
 b15zdnd00an1n01x5 FILLER_324_1604 ();
 b15zdnd11an1n16x5 FILLER_324_1647 ();
 b15zdnd11an1n08x5 FILLER_324_1663 ();
 b15zdnd00an1n02x5 FILLER_324_1671 ();
 b15zdnd00an1n01x5 FILLER_324_1673 ();
 b15zdnd11an1n04x5 FILLER_324_1699 ();
 b15zdnd11an1n64x5 FILLER_324_1706 ();
 b15zdnd11an1n32x5 FILLER_324_1770 ();
 b15zdnd11an1n04x5 FILLER_324_1802 ();
 b15zdnd00an1n02x5 FILLER_324_1806 ();
 b15zdnd00an1n01x5 FILLER_324_1808 ();
 b15zdnd11an1n04x5 FILLER_324_1849 ();
 b15zdnd11an1n16x5 FILLER_324_1856 ();
 b15zdnd00an1n02x5 FILLER_324_1872 ();
 b15zdnd11an1n64x5 FILLER_324_1877 ();
 b15zdnd11an1n64x5 FILLER_324_1941 ();
 b15zdnd11an1n64x5 FILLER_324_2005 ();
 b15zdnd11an1n64x5 FILLER_324_2069 ();
 b15zdnd11an1n16x5 FILLER_324_2133 ();
 b15zdnd11an1n04x5 FILLER_324_2149 ();
 b15zdnd00an1n01x5 FILLER_324_2153 ();
 b15zdnd11an1n64x5 FILLER_324_2162 ();
 b15zdnd11an1n32x5 FILLER_324_2226 ();
 b15zdnd11an1n16x5 FILLER_324_2258 ();
 b15zdnd00an1n02x5 FILLER_324_2274 ();
 b15zdnd11an1n64x5 FILLER_325_0 ();
 b15zdnd11an1n32x5 FILLER_325_64 ();
 b15zdnd11an1n16x5 FILLER_325_96 ();
 b15zdnd11an1n08x5 FILLER_325_112 ();
 b15zdnd11an1n04x5 FILLER_325_120 ();
 b15zdnd00an1n01x5 FILLER_325_124 ();
 b15zdnd11an1n64x5 FILLER_325_156 ();
 b15zdnd11an1n64x5 FILLER_325_220 ();
 b15zdnd11an1n64x5 FILLER_325_284 ();
 b15zdnd11an1n64x5 FILLER_325_348 ();
 b15zdnd11an1n64x5 FILLER_325_412 ();
 b15zdnd11an1n64x5 FILLER_325_476 ();
 b15zdnd11an1n32x5 FILLER_325_540 ();
 b15zdnd11an1n16x5 FILLER_325_572 ();
 b15zdnd11an1n04x5 FILLER_325_588 ();
 b15zdnd00an1n02x5 FILLER_325_592 ();
 b15zdnd11an1n04x5 FILLER_325_597 ();
 b15zdnd11an1n64x5 FILLER_325_604 ();
 b15zdnd11an1n64x5 FILLER_325_668 ();
 b15zdnd11an1n64x5 FILLER_325_732 ();
 b15zdnd11an1n64x5 FILLER_325_796 ();
 b15zdnd11an1n64x5 FILLER_325_860 ();
 b15zdnd11an1n64x5 FILLER_325_924 ();
 b15zdnd11an1n04x5 FILLER_325_988 ();
 b15zdnd00an1n01x5 FILLER_325_992 ();
 b15zdnd11an1n64x5 FILLER_325_1001 ();
 b15zdnd11an1n64x5 FILLER_325_1065 ();
 b15zdnd11an1n64x5 FILLER_325_1129 ();
 b15zdnd11an1n16x5 FILLER_325_1193 ();
 b15zdnd00an1n01x5 FILLER_325_1209 ();
 b15zdnd11an1n04x5 FILLER_325_1216 ();
 b15zdnd11an1n16x5 FILLER_325_1223 ();
 b15zdnd11an1n32x5 FILLER_325_1281 ();
 b15zdnd11an1n04x5 FILLER_325_1313 ();
 b15zdnd00an1n02x5 FILLER_325_1317 ();
 b15zdnd11an1n64x5 FILLER_325_1330 ();
 b15zdnd11an1n64x5 FILLER_325_1394 ();
 b15zdnd11an1n64x5 FILLER_325_1458 ();
 b15zdnd11an1n32x5 FILLER_325_1522 ();
 b15zdnd11an1n16x5 FILLER_325_1554 ();
 b15zdnd11an1n08x5 FILLER_325_1570 ();
 b15zdnd00an1n02x5 FILLER_325_1578 ();
 b15zdnd11an1n32x5 FILLER_325_1622 ();
 b15zdnd11an1n08x5 FILLER_325_1654 ();
 b15zdnd11an1n04x5 FILLER_325_1662 ();
 b15zdnd11an1n64x5 FILLER_325_1706 ();
 b15zdnd11an1n64x5 FILLER_325_1770 ();
 b15zdnd11an1n08x5 FILLER_325_1834 ();
 b15zdnd00an1n02x5 FILLER_325_1842 ();
 b15zdnd00an1n01x5 FILLER_325_1844 ();
 b15zdnd11an1n64x5 FILLER_325_1848 ();
 b15zdnd11an1n64x5 FILLER_325_1912 ();
 b15zdnd11an1n64x5 FILLER_325_1976 ();
 b15zdnd11an1n64x5 FILLER_325_2040 ();
 b15zdnd11an1n64x5 FILLER_325_2104 ();
 b15zdnd11an1n64x5 FILLER_325_2168 ();
 b15zdnd11an1n32x5 FILLER_325_2232 ();
 b15zdnd11an1n16x5 FILLER_325_2264 ();
 b15zdnd11an1n04x5 FILLER_325_2280 ();
 b15zdnd11an1n64x5 FILLER_326_8 ();
 b15zdnd11an1n16x5 FILLER_326_72 ();
 b15zdnd11an1n04x5 FILLER_326_88 ();
 b15zdnd11an1n04x5 FILLER_326_110 ();
 b15zdnd11an1n64x5 FILLER_326_139 ();
 b15zdnd11an1n64x5 FILLER_326_203 ();
 b15zdnd11an1n64x5 FILLER_326_267 ();
 b15zdnd11an1n64x5 FILLER_326_331 ();
 b15zdnd11an1n64x5 FILLER_326_395 ();
 b15zdnd11an1n32x5 FILLER_326_459 ();
 b15zdnd00an1n01x5 FILLER_326_491 ();
 b15zdnd11an1n64x5 FILLER_326_534 ();
 b15zdnd11an1n64x5 FILLER_326_598 ();
 b15zdnd11an1n32x5 FILLER_326_662 ();
 b15zdnd11an1n16x5 FILLER_326_694 ();
 b15zdnd11an1n08x5 FILLER_326_710 ();
 b15zdnd11an1n64x5 FILLER_326_726 ();
 b15zdnd11an1n64x5 FILLER_326_790 ();
 b15zdnd11an1n64x5 FILLER_326_854 ();
 b15zdnd11an1n64x5 FILLER_326_918 ();
 b15zdnd11an1n64x5 FILLER_326_982 ();
 b15zdnd11an1n64x5 FILLER_326_1046 ();
 b15zdnd11an1n64x5 FILLER_326_1110 ();
 b15zdnd00an1n02x5 FILLER_326_1174 ();
 b15zdnd11an1n16x5 FILLER_326_1218 ();
 b15zdnd00an1n02x5 FILLER_326_1234 ();
 b15zdnd11an1n64x5 FILLER_326_1278 ();
 b15zdnd11an1n64x5 FILLER_326_1342 ();
 b15zdnd11an1n16x5 FILLER_326_1406 ();
 b15zdnd11an1n08x5 FILLER_326_1422 ();
 b15zdnd00an1n02x5 FILLER_326_1430 ();
 b15zdnd11an1n64x5 FILLER_326_1441 ();
 b15zdnd11an1n64x5 FILLER_326_1505 ();
 b15zdnd11an1n64x5 FILLER_326_1569 ();
 b15zdnd11an1n32x5 FILLER_326_1633 ();
 b15zdnd11an1n16x5 FILLER_326_1665 ();
 b15zdnd11an1n04x5 FILLER_326_1681 ();
 b15zdnd00an1n02x5 FILLER_326_1685 ();
 b15zdnd11an1n04x5 FILLER_326_1693 ();
 b15zdnd11an1n64x5 FILLER_326_1700 ();
 b15zdnd11an1n64x5 FILLER_326_1764 ();
 b15zdnd11an1n64x5 FILLER_326_1828 ();
 b15zdnd11an1n64x5 FILLER_326_1892 ();
 b15zdnd11an1n64x5 FILLER_326_1956 ();
 b15zdnd11an1n64x5 FILLER_326_2020 ();
 b15zdnd11an1n64x5 FILLER_326_2084 ();
 b15zdnd11an1n04x5 FILLER_326_2148 ();
 b15zdnd00an1n02x5 FILLER_326_2152 ();
 b15zdnd11an1n64x5 FILLER_326_2162 ();
 b15zdnd11an1n32x5 FILLER_326_2226 ();
 b15zdnd11an1n16x5 FILLER_326_2258 ();
 b15zdnd00an1n02x5 FILLER_326_2274 ();
 b15zdnd11an1n64x5 FILLER_327_0 ();
 b15zdnd11an1n64x5 FILLER_327_64 ();
 b15zdnd11an1n64x5 FILLER_327_128 ();
 b15zdnd11an1n64x5 FILLER_327_192 ();
 b15zdnd11an1n64x5 FILLER_327_256 ();
 b15zdnd11an1n64x5 FILLER_327_320 ();
 b15zdnd11an1n64x5 FILLER_327_384 ();
 b15zdnd11an1n32x5 FILLER_327_448 ();
 b15zdnd11an1n08x5 FILLER_327_480 ();
 b15zdnd11an1n04x5 FILLER_327_488 ();
 b15zdnd00an1n01x5 FILLER_327_492 ();
 b15zdnd11an1n64x5 FILLER_327_499 ();
 b15zdnd11an1n64x5 FILLER_327_563 ();
 b15zdnd11an1n64x5 FILLER_327_627 ();
 b15zdnd11an1n64x5 FILLER_327_691 ();
 b15zdnd11an1n64x5 FILLER_327_755 ();
 b15zdnd11an1n64x5 FILLER_327_819 ();
 b15zdnd11an1n64x5 FILLER_327_883 ();
 b15zdnd11an1n64x5 FILLER_327_947 ();
 b15zdnd11an1n64x5 FILLER_327_1011 ();
 b15zdnd11an1n64x5 FILLER_327_1075 ();
 b15zdnd11an1n64x5 FILLER_327_1139 ();
 b15zdnd11an1n16x5 FILLER_327_1203 ();
 b15zdnd11an1n08x5 FILLER_327_1219 ();
 b15zdnd11an1n04x5 FILLER_327_1227 ();
 b15zdnd00an1n02x5 FILLER_327_1231 ();
 b15zdnd00an1n01x5 FILLER_327_1233 ();
 b15zdnd11an1n64x5 FILLER_327_1276 ();
 b15zdnd11an1n64x5 FILLER_327_1340 ();
 b15zdnd11an1n64x5 FILLER_327_1404 ();
 b15zdnd11an1n64x5 FILLER_327_1468 ();
 b15zdnd11an1n32x5 FILLER_327_1532 ();
 b15zdnd11an1n16x5 FILLER_327_1564 ();
 b15zdnd11an1n08x5 FILLER_327_1580 ();
 b15zdnd00an1n02x5 FILLER_327_1588 ();
 b15zdnd11an1n04x5 FILLER_327_1593 ();
 b15zdnd11an1n64x5 FILLER_327_1600 ();
 b15zdnd11an1n64x5 FILLER_327_1664 ();
 b15zdnd11an1n64x5 FILLER_327_1728 ();
 b15zdnd11an1n64x5 FILLER_327_1792 ();
 b15zdnd11an1n64x5 FILLER_327_1856 ();
 b15zdnd11an1n08x5 FILLER_327_1920 ();
 b15zdnd11an1n04x5 FILLER_327_1928 ();
 b15zdnd00an1n02x5 FILLER_327_1932 ();
 b15zdnd00an1n01x5 FILLER_327_1934 ();
 b15zdnd11an1n04x5 FILLER_327_1938 ();
 b15zdnd11an1n64x5 FILLER_327_1945 ();
 b15zdnd11an1n64x5 FILLER_327_2009 ();
 b15zdnd11an1n64x5 FILLER_327_2073 ();
 b15zdnd11an1n64x5 FILLER_327_2137 ();
 b15zdnd11an1n04x5 FILLER_327_2201 ();
 b15zdnd00an1n02x5 FILLER_327_2205 ();
 b15zdnd11an1n64x5 FILLER_327_2210 ();
 b15zdnd11an1n08x5 FILLER_327_2274 ();
 b15zdnd00an1n02x5 FILLER_327_2282 ();
 b15zdnd11an1n64x5 FILLER_328_8 ();
 b15zdnd11an1n64x5 FILLER_328_72 ();
 b15zdnd11an1n64x5 FILLER_328_136 ();
 b15zdnd11an1n64x5 FILLER_328_200 ();
 b15zdnd11an1n64x5 FILLER_328_264 ();
 b15zdnd11an1n64x5 FILLER_328_328 ();
 b15zdnd11an1n08x5 FILLER_328_392 ();
 b15zdnd00an1n02x5 FILLER_328_400 ();
 b15zdnd11an1n16x5 FILLER_328_441 ();
 b15zdnd00an1n01x5 FILLER_328_457 ();
 b15zdnd11an1n64x5 FILLER_328_479 ();
 b15zdnd11an1n64x5 FILLER_328_543 ();
 b15zdnd11an1n64x5 FILLER_328_607 ();
 b15zdnd11an1n32x5 FILLER_328_671 ();
 b15zdnd11an1n08x5 FILLER_328_703 ();
 b15zdnd11an1n04x5 FILLER_328_711 ();
 b15zdnd00an1n02x5 FILLER_328_715 ();
 b15zdnd00an1n01x5 FILLER_328_717 ();
 b15zdnd11an1n64x5 FILLER_328_726 ();
 b15zdnd11an1n64x5 FILLER_328_790 ();
 b15zdnd11an1n64x5 FILLER_328_854 ();
 b15zdnd11an1n64x5 FILLER_328_918 ();
 b15zdnd11an1n08x5 FILLER_328_982 ();
 b15zdnd11an1n04x5 FILLER_328_990 ();
 b15zdnd00an1n02x5 FILLER_328_994 ();
 b15zdnd00an1n01x5 FILLER_328_996 ();
 b15zdnd11an1n64x5 FILLER_328_1039 ();
 b15zdnd11an1n64x5 FILLER_328_1103 ();
 b15zdnd11an1n32x5 FILLER_328_1167 ();
 b15zdnd11an1n16x5 FILLER_328_1199 ();
 b15zdnd00an1n02x5 FILLER_328_1215 ();
 b15zdnd11an1n64x5 FILLER_328_1269 ();
 b15zdnd11an1n64x5 FILLER_328_1333 ();
 b15zdnd11an1n64x5 FILLER_328_1397 ();
 b15zdnd11an1n64x5 FILLER_328_1461 ();
 b15zdnd11an1n32x5 FILLER_328_1525 ();
 b15zdnd11an1n08x5 FILLER_328_1557 ();
 b15zdnd11an1n04x5 FILLER_328_1565 ();
 b15zdnd00an1n02x5 FILLER_328_1569 ();
 b15zdnd00an1n01x5 FILLER_328_1571 ();
 b15zdnd11an1n64x5 FILLER_328_1624 ();
 b15zdnd11an1n16x5 FILLER_328_1688 ();
 b15zdnd11an1n08x5 FILLER_328_1704 ();
 b15zdnd00an1n01x5 FILLER_328_1712 ();
 b15zdnd11an1n04x5 FILLER_328_1716 ();
 b15zdnd11an1n64x5 FILLER_328_1723 ();
 b15zdnd11an1n64x5 FILLER_328_1787 ();
 b15zdnd11an1n32x5 FILLER_328_1851 ();
 b15zdnd11an1n16x5 FILLER_328_1883 ();
 b15zdnd11an1n08x5 FILLER_328_1899 ();
 b15zdnd00an1n02x5 FILLER_328_1907 ();
 b15zdnd00an1n01x5 FILLER_328_1909 ();
 b15zdnd11an1n64x5 FILLER_328_1962 ();
 b15zdnd11an1n64x5 FILLER_328_2026 ();
 b15zdnd11an1n64x5 FILLER_328_2090 ();
 b15zdnd11an1n32x5 FILLER_328_2162 ();
 b15zdnd11an1n08x5 FILLER_328_2194 ();
 b15zdnd11an1n04x5 FILLER_328_2202 ();
 b15zdnd11an1n64x5 FILLER_328_2209 ();
 b15zdnd00an1n02x5 FILLER_328_2273 ();
 b15zdnd00an1n01x5 FILLER_328_2275 ();
 b15zdnd11an1n64x5 FILLER_329_0 ();
 b15zdnd11an1n64x5 FILLER_329_64 ();
 b15zdnd11an1n64x5 FILLER_329_128 ();
 b15zdnd11an1n64x5 FILLER_329_192 ();
 b15zdnd11an1n64x5 FILLER_329_256 ();
 b15zdnd11an1n32x5 FILLER_329_320 ();
 b15zdnd11an1n16x5 FILLER_329_352 ();
 b15zdnd11an1n08x5 FILLER_329_368 ();
 b15zdnd11an1n04x5 FILLER_329_376 ();
 b15zdnd11an1n08x5 FILLER_329_383 ();
 b15zdnd00an1n01x5 FILLER_329_391 ();
 b15zdnd11an1n32x5 FILLER_329_395 ();
 b15zdnd11an1n04x5 FILLER_329_427 ();
 b15zdnd00an1n01x5 FILLER_329_431 ();
 b15zdnd11an1n08x5 FILLER_329_474 ();
 b15zdnd00an1n01x5 FILLER_329_482 ();
 b15zdnd11an1n64x5 FILLER_329_491 ();
 b15zdnd11an1n64x5 FILLER_329_555 ();
 b15zdnd11an1n64x5 FILLER_329_619 ();
 b15zdnd11an1n64x5 FILLER_329_683 ();
 b15zdnd11an1n64x5 FILLER_329_747 ();
 b15zdnd11an1n64x5 FILLER_329_811 ();
 b15zdnd11an1n64x5 FILLER_329_875 ();
 b15zdnd11an1n64x5 FILLER_329_939 ();
 b15zdnd11an1n16x5 FILLER_329_1003 ();
 b15zdnd11an1n08x5 FILLER_329_1019 ();
 b15zdnd00an1n01x5 FILLER_329_1027 ();
 b15zdnd11an1n64x5 FILLER_329_1031 ();
 b15zdnd11an1n64x5 FILLER_329_1095 ();
 b15zdnd11an1n64x5 FILLER_329_1159 ();
 b15zdnd11an1n16x5 FILLER_329_1223 ();
 b15zdnd11an1n04x5 FILLER_329_1239 ();
 b15zdnd11an1n08x5 FILLER_329_1246 ();
 b15zdnd00an1n02x5 FILLER_329_1254 ();
 b15zdnd00an1n01x5 FILLER_329_1256 ();
 b15zdnd11an1n64x5 FILLER_329_1260 ();
 b15zdnd11an1n64x5 FILLER_329_1324 ();
 b15zdnd11an1n64x5 FILLER_329_1388 ();
 b15zdnd11an1n64x5 FILLER_329_1452 ();
 b15zdnd11an1n64x5 FILLER_329_1516 ();
 b15zdnd11an1n16x5 FILLER_329_1580 ();
 b15zdnd00an1n02x5 FILLER_329_1596 ();
 b15zdnd11an1n64x5 FILLER_329_1601 ();
 b15zdnd11an1n16x5 FILLER_329_1665 ();
 b15zdnd11an1n08x5 FILLER_329_1681 ();
 b15zdnd11an1n04x5 FILLER_329_1689 ();
 b15zdnd00an1n02x5 FILLER_329_1693 ();
 b15zdnd11an1n64x5 FILLER_329_1747 ();
 b15zdnd11an1n64x5 FILLER_329_1811 ();
 b15zdnd11an1n32x5 FILLER_329_1875 ();
 b15zdnd11an1n16x5 FILLER_329_1907 ();
 b15zdnd11an1n08x5 FILLER_329_1923 ();
 b15zdnd11an1n04x5 FILLER_329_1931 ();
 b15zdnd00an1n01x5 FILLER_329_1935 ();
 b15zdnd11an1n04x5 FILLER_329_1939 ();
 b15zdnd00an1n02x5 FILLER_329_1943 ();
 b15zdnd11an1n64x5 FILLER_329_1987 ();
 b15zdnd11an1n32x5 FILLER_329_2051 ();
 b15zdnd00an1n02x5 FILLER_329_2083 ();
 b15zdnd00an1n01x5 FILLER_329_2085 ();
 b15zdnd11an1n32x5 FILLER_329_2128 ();
 b15zdnd11an1n16x5 FILLER_329_2160 ();
 b15zdnd11an1n04x5 FILLER_329_2176 ();
 b15zdnd00an1n01x5 FILLER_329_2180 ();
 b15zdnd11an1n32x5 FILLER_329_2233 ();
 b15zdnd11an1n16x5 FILLER_329_2265 ();
 b15zdnd00an1n02x5 FILLER_329_2281 ();
 b15zdnd00an1n01x5 FILLER_329_2283 ();
 b15zdnd11an1n64x5 FILLER_330_8 ();
 b15zdnd11an1n64x5 FILLER_330_72 ();
 b15zdnd11an1n64x5 FILLER_330_136 ();
 b15zdnd11an1n64x5 FILLER_330_200 ();
 b15zdnd11an1n64x5 FILLER_330_264 ();
 b15zdnd11an1n32x5 FILLER_330_328 ();
 b15zdnd00an1n02x5 FILLER_330_360 ();
 b15zdnd11an1n04x5 FILLER_330_366 ();
 b15zdnd11an1n04x5 FILLER_330_422 ();
 b15zdnd11an1n04x5 FILLER_330_434 ();
 b15zdnd11an1n04x5 FILLER_330_480 ();
 b15zdnd11an1n64x5 FILLER_330_489 ();
 b15zdnd11an1n32x5 FILLER_330_553 ();
 b15zdnd11an1n16x5 FILLER_330_585 ();
 b15zdnd00an1n02x5 FILLER_330_601 ();
 b15zdnd00an1n01x5 FILLER_330_603 ();
 b15zdnd11an1n08x5 FILLER_330_610 ();
 b15zdnd00an1n01x5 FILLER_330_618 ();
 b15zdnd11an1n64x5 FILLER_330_628 ();
 b15zdnd11an1n16x5 FILLER_330_692 ();
 b15zdnd11an1n08x5 FILLER_330_708 ();
 b15zdnd00an1n02x5 FILLER_330_716 ();
 b15zdnd11an1n64x5 FILLER_330_726 ();
 b15zdnd11an1n64x5 FILLER_330_790 ();
 b15zdnd11an1n64x5 FILLER_330_854 ();
 b15zdnd11an1n32x5 FILLER_330_918 ();
 b15zdnd11an1n16x5 FILLER_330_950 ();
 b15zdnd00an1n02x5 FILLER_330_966 ();
 b15zdnd00an1n01x5 FILLER_330_968 ();
 b15zdnd11an1n04x5 FILLER_330_972 ();
 b15zdnd00an1n02x5 FILLER_330_976 ();
 b15zdnd11an1n08x5 FILLER_330_981 ();
 b15zdnd00an1n02x5 FILLER_330_989 ();
 b15zdnd00an1n01x5 FILLER_330_991 ();
 b15zdnd11an1n04x5 FILLER_330_1032 ();
 b15zdnd11an1n64x5 FILLER_330_1039 ();
 b15zdnd11an1n64x5 FILLER_330_1103 ();
 b15zdnd11an1n64x5 FILLER_330_1167 ();
 b15zdnd11an1n08x5 FILLER_330_1231 ();
 b15zdnd00an1n02x5 FILLER_330_1239 ();
 b15zdnd00an1n01x5 FILLER_330_1241 ();
 b15zdnd11an1n64x5 FILLER_330_1245 ();
 b15zdnd11an1n64x5 FILLER_330_1309 ();
 b15zdnd11an1n64x5 FILLER_330_1373 ();
 b15zdnd11an1n64x5 FILLER_330_1437 ();
 b15zdnd11an1n64x5 FILLER_330_1501 ();
 b15zdnd11an1n64x5 FILLER_330_1565 ();
 b15zdnd11an1n64x5 FILLER_330_1629 ();
 b15zdnd11an1n16x5 FILLER_330_1693 ();
 b15zdnd11an1n08x5 FILLER_330_1709 ();
 b15zdnd00an1n02x5 FILLER_330_1717 ();
 b15zdnd00an1n01x5 FILLER_330_1719 ();
 b15zdnd11an1n64x5 FILLER_330_1723 ();
 b15zdnd11an1n64x5 FILLER_330_1787 ();
 b15zdnd11an1n64x5 FILLER_330_1851 ();
 b15zdnd11an1n32x5 FILLER_330_1915 ();
 b15zdnd11an1n04x5 FILLER_330_1947 ();
 b15zdnd00an1n01x5 FILLER_330_1951 ();
 b15zdnd11an1n04x5 FILLER_330_1967 ();
 b15zdnd11an1n16x5 FILLER_330_1975 ();
 b15zdnd11an1n08x5 FILLER_330_1991 ();
 b15zdnd11an1n04x5 FILLER_330_1999 ();
 b15zdnd11an1n64x5 FILLER_330_2006 ();
 b15zdnd11an1n64x5 FILLER_330_2070 ();
 b15zdnd11an1n16x5 FILLER_330_2134 ();
 b15zdnd11an1n04x5 FILLER_330_2150 ();
 b15zdnd11an1n32x5 FILLER_330_2162 ();
 b15zdnd11an1n08x5 FILLER_330_2194 ();
 b15zdnd11an1n04x5 FILLER_330_2202 ();
 b15zdnd11an1n64x5 FILLER_330_2209 ();
 b15zdnd00an1n02x5 FILLER_330_2273 ();
 b15zdnd00an1n01x5 FILLER_330_2275 ();
 b15zdnd11an1n64x5 FILLER_331_0 ();
 b15zdnd11an1n64x5 FILLER_331_64 ();
 b15zdnd11an1n64x5 FILLER_331_128 ();
 b15zdnd11an1n64x5 FILLER_331_192 ();
 b15zdnd11an1n64x5 FILLER_331_256 ();
 b15zdnd11an1n64x5 FILLER_331_320 ();
 b15zdnd11an1n08x5 FILLER_331_384 ();
 b15zdnd00an1n01x5 FILLER_331_392 ();
 b15zdnd11an1n32x5 FILLER_331_396 ();
 b15zdnd11an1n16x5 FILLER_331_428 ();
 b15zdnd00an1n02x5 FILLER_331_444 ();
 b15zdnd11an1n04x5 FILLER_331_453 ();
 b15zdnd11an1n64x5 FILLER_331_499 ();
 b15zdnd11an1n64x5 FILLER_331_563 ();
 b15zdnd11an1n64x5 FILLER_331_627 ();
 b15zdnd11an1n64x5 FILLER_331_691 ();
 b15zdnd11an1n64x5 FILLER_331_755 ();
 b15zdnd11an1n64x5 FILLER_331_819 ();
 b15zdnd11an1n64x5 FILLER_331_883 ();
 b15zdnd11an1n04x5 FILLER_331_947 ();
 b15zdnd11an1n64x5 FILLER_331_1003 ();
 b15zdnd11an1n64x5 FILLER_331_1067 ();
 b15zdnd11an1n64x5 FILLER_331_1131 ();
 b15zdnd11an1n64x5 FILLER_331_1195 ();
 b15zdnd11an1n64x5 FILLER_331_1259 ();
 b15zdnd11an1n64x5 FILLER_331_1323 ();
 b15zdnd11an1n64x5 FILLER_331_1387 ();
 b15zdnd11an1n64x5 FILLER_331_1451 ();
 b15zdnd11an1n64x5 FILLER_331_1515 ();
 b15zdnd11an1n64x5 FILLER_331_1579 ();
 b15zdnd11an1n64x5 FILLER_331_1643 ();
 b15zdnd11an1n64x5 FILLER_331_1707 ();
 b15zdnd11an1n64x5 FILLER_331_1771 ();
 b15zdnd11an1n64x5 FILLER_331_1835 ();
 b15zdnd11an1n64x5 FILLER_331_1899 ();
 b15zdnd11an1n04x5 FILLER_331_1963 ();
 b15zdnd00an1n01x5 FILLER_331_1967 ();
 b15zdnd11an1n64x5 FILLER_331_2010 ();
 b15zdnd11an1n64x5 FILLER_331_2074 ();
 b15zdnd11an1n64x5 FILLER_331_2138 ();
 b15zdnd11an1n64x5 FILLER_331_2202 ();
 b15zdnd11an1n16x5 FILLER_331_2266 ();
 b15zdnd00an1n02x5 FILLER_331_2282 ();
 b15zdnd11an1n64x5 FILLER_332_8 ();
 b15zdnd11an1n64x5 FILLER_332_72 ();
 b15zdnd11an1n64x5 FILLER_332_136 ();
 b15zdnd11an1n64x5 FILLER_332_200 ();
 b15zdnd00an1n02x5 FILLER_332_264 ();
 b15zdnd00an1n01x5 FILLER_332_266 ();
 b15zdnd11an1n64x5 FILLER_332_270 ();
 b15zdnd11an1n64x5 FILLER_332_334 ();
 b15zdnd11an1n16x5 FILLER_332_398 ();
 b15zdnd11an1n08x5 FILLER_332_414 ();
 b15zdnd11an1n04x5 FILLER_332_422 ();
 b15zdnd00an1n01x5 FILLER_332_426 ();
 b15zdnd11an1n04x5 FILLER_332_469 ();
 b15zdnd11an1n04x5 FILLER_332_477 ();
 b15zdnd11an1n64x5 FILLER_332_484 ();
 b15zdnd11an1n64x5 FILLER_332_548 ();
 b15zdnd11an1n64x5 FILLER_332_612 ();
 b15zdnd11an1n32x5 FILLER_332_676 ();
 b15zdnd11an1n08x5 FILLER_332_708 ();
 b15zdnd00an1n02x5 FILLER_332_716 ();
 b15zdnd11an1n64x5 FILLER_332_726 ();
 b15zdnd11an1n64x5 FILLER_332_790 ();
 b15zdnd11an1n64x5 FILLER_332_854 ();
 b15zdnd11an1n32x5 FILLER_332_918 ();
 b15zdnd11an1n04x5 FILLER_332_950 ();
 b15zdnd00an1n02x5 FILLER_332_954 ();
 b15zdnd00an1n01x5 FILLER_332_956 ();
 b15zdnd11an1n08x5 FILLER_332_999 ();
 b15zdnd11an1n04x5 FILLER_332_1007 ();
 b15zdnd00an1n02x5 FILLER_332_1011 ();
 b15zdnd11an1n32x5 FILLER_332_1055 ();
 b15zdnd11an1n16x5 FILLER_332_1087 ();
 b15zdnd11an1n04x5 FILLER_332_1103 ();
 b15zdnd00an1n01x5 FILLER_332_1107 ();
 b15zdnd11an1n64x5 FILLER_332_1111 ();
 b15zdnd11an1n32x5 FILLER_332_1175 ();
 b15zdnd11an1n08x5 FILLER_332_1207 ();
 b15zdnd00an1n01x5 FILLER_332_1215 ();
 b15zdnd11an1n64x5 FILLER_332_1226 ();
 b15zdnd11an1n64x5 FILLER_332_1290 ();
 b15zdnd11an1n64x5 FILLER_332_1354 ();
 b15zdnd11an1n64x5 FILLER_332_1418 ();
 b15zdnd11an1n64x5 FILLER_332_1482 ();
 b15zdnd11an1n64x5 FILLER_332_1546 ();
 b15zdnd11an1n64x5 FILLER_332_1610 ();
 b15zdnd11an1n64x5 FILLER_332_1674 ();
 b15zdnd11an1n64x5 FILLER_332_1738 ();
 b15zdnd11an1n64x5 FILLER_332_1802 ();
 b15zdnd11an1n64x5 FILLER_332_1866 ();
 b15zdnd11an1n32x5 FILLER_332_1930 ();
 b15zdnd11an1n04x5 FILLER_332_1962 ();
 b15zdnd11an1n64x5 FILLER_332_2006 ();
 b15zdnd11an1n64x5 FILLER_332_2070 ();
 b15zdnd11an1n16x5 FILLER_332_2134 ();
 b15zdnd11an1n04x5 FILLER_332_2150 ();
 b15zdnd11an1n64x5 FILLER_332_2162 ();
 b15zdnd11an1n32x5 FILLER_332_2226 ();
 b15zdnd11an1n16x5 FILLER_332_2258 ();
 b15zdnd00an1n02x5 FILLER_332_2274 ();
 b15zdnd11an1n64x5 FILLER_333_0 ();
 b15zdnd11an1n64x5 FILLER_333_64 ();
 b15zdnd11an1n64x5 FILLER_333_128 ();
 b15zdnd11an1n32x5 FILLER_333_192 ();
 b15zdnd11an1n08x5 FILLER_333_224 ();
 b15zdnd00an1n01x5 FILLER_333_232 ();
 b15zdnd11an1n04x5 FILLER_333_273 ();
 b15zdnd11an1n64x5 FILLER_333_280 ();
 b15zdnd11an1n64x5 FILLER_333_344 ();
 b15zdnd11an1n32x5 FILLER_333_408 ();
 b15zdnd11an1n08x5 FILLER_333_440 ();
 b15zdnd11an1n04x5 FILLER_333_452 ();
 b15zdnd00an1n02x5 FILLER_333_456 ();
 b15zdnd00an1n01x5 FILLER_333_458 ();
 b15zdnd11an1n04x5 FILLER_333_468 ();
 b15zdnd11an1n64x5 FILLER_333_477 ();
 b15zdnd11an1n64x5 FILLER_333_541 ();
 b15zdnd11an1n64x5 FILLER_333_605 ();
 b15zdnd11an1n64x5 FILLER_333_669 ();
 b15zdnd11an1n16x5 FILLER_333_733 ();
 b15zdnd11an1n04x5 FILLER_333_749 ();
 b15zdnd00an1n01x5 FILLER_333_753 ();
 b15zdnd11an1n64x5 FILLER_333_757 ();
 b15zdnd11an1n64x5 FILLER_333_821 ();
 b15zdnd11an1n64x5 FILLER_333_885 ();
 b15zdnd11an1n08x5 FILLER_333_949 ();
 b15zdnd00an1n02x5 FILLER_333_957 ();
 b15zdnd00an1n01x5 FILLER_333_959 ();
 b15zdnd11an1n08x5 FILLER_333_967 ();
 b15zdnd00an1n01x5 FILLER_333_975 ();
 b15zdnd11an1n32x5 FILLER_333_979 ();
 b15zdnd11an1n08x5 FILLER_333_1011 ();
 b15zdnd11an1n04x5 FILLER_333_1019 ();
 b15zdnd11an1n64x5 FILLER_333_1030 ();
 b15zdnd11an1n08x5 FILLER_333_1094 ();
 b15zdnd11an1n04x5 FILLER_333_1102 ();
 b15zdnd00an1n02x5 FILLER_333_1106 ();
 b15zdnd00an1n01x5 FILLER_333_1108 ();
 b15zdnd11an1n64x5 FILLER_333_1116 ();
 b15zdnd11an1n32x5 FILLER_333_1180 ();
 b15zdnd11an1n08x5 FILLER_333_1212 ();
 b15zdnd00an1n02x5 FILLER_333_1220 ();
 b15zdnd11an1n64x5 FILLER_333_1229 ();
 b15zdnd11an1n32x5 FILLER_333_1293 ();
 b15zdnd11an1n16x5 FILLER_333_1325 ();
 b15zdnd11an1n04x5 FILLER_333_1341 ();
 b15zdnd00an1n02x5 FILLER_333_1345 ();
 b15zdnd00an1n01x5 FILLER_333_1347 ();
 b15zdnd11an1n64x5 FILLER_333_1353 ();
 b15zdnd11an1n16x5 FILLER_333_1417 ();
 b15zdnd11an1n08x5 FILLER_333_1433 ();
 b15zdnd11an1n04x5 FILLER_333_1441 ();
 b15zdnd00an1n02x5 FILLER_333_1445 ();
 b15zdnd11an1n04x5 FILLER_333_1450 ();
 b15zdnd11an1n64x5 FILLER_333_1481 ();
 b15zdnd11an1n64x5 FILLER_333_1545 ();
 b15zdnd11an1n64x5 FILLER_333_1609 ();
 b15zdnd11an1n64x5 FILLER_333_1673 ();
 b15zdnd11an1n64x5 FILLER_333_1737 ();
 b15zdnd11an1n64x5 FILLER_333_1801 ();
 b15zdnd11an1n64x5 FILLER_333_1865 ();
 b15zdnd11an1n64x5 FILLER_333_1929 ();
 b15zdnd11an1n08x5 FILLER_333_1993 ();
 b15zdnd00an1n01x5 FILLER_333_2001 ();
 b15zdnd11an1n64x5 FILLER_333_2005 ();
 b15zdnd11an1n16x5 FILLER_333_2069 ();
 b15zdnd11an1n04x5 FILLER_333_2085 ();
 b15zdnd00an1n01x5 FILLER_333_2089 ();
 b15zdnd11an1n64x5 FILLER_333_2093 ();
 b15zdnd11an1n64x5 FILLER_333_2157 ();
 b15zdnd11an1n32x5 FILLER_333_2221 ();
 b15zdnd11an1n16x5 FILLER_333_2253 ();
 b15zdnd11an1n08x5 FILLER_333_2269 ();
 b15zdnd11an1n04x5 FILLER_333_2277 ();
 b15zdnd00an1n02x5 FILLER_333_2281 ();
 b15zdnd00an1n01x5 FILLER_333_2283 ();
 b15zdnd11an1n64x5 FILLER_334_8 ();
 b15zdnd11an1n64x5 FILLER_334_72 ();
 b15zdnd11an1n64x5 FILLER_334_136 ();
 b15zdnd11an1n64x5 FILLER_334_200 ();
 b15zdnd11an1n64x5 FILLER_334_264 ();
 b15zdnd11an1n64x5 FILLER_334_328 ();
 b15zdnd11an1n64x5 FILLER_334_392 ();
 b15zdnd11an1n04x5 FILLER_334_461 ();
 b15zdnd11an1n64x5 FILLER_334_468 ();
 b15zdnd11an1n64x5 FILLER_334_532 ();
 b15zdnd11an1n16x5 FILLER_334_596 ();
 b15zdnd11an1n08x5 FILLER_334_612 ();
 b15zdnd00an1n01x5 FILLER_334_620 ();
 b15zdnd11an1n64x5 FILLER_334_627 ();
 b15zdnd11an1n16x5 FILLER_334_691 ();
 b15zdnd11an1n08x5 FILLER_334_707 ();
 b15zdnd00an1n02x5 FILLER_334_715 ();
 b15zdnd00an1n01x5 FILLER_334_717 ();
 b15zdnd00an1n02x5 FILLER_334_726 ();
 b15zdnd11an1n64x5 FILLER_334_780 ();
 b15zdnd11an1n64x5 FILLER_334_844 ();
 b15zdnd11an1n64x5 FILLER_334_908 ();
 b15zdnd11an1n64x5 FILLER_334_972 ();
 b15zdnd11an1n32x5 FILLER_334_1036 ();
 b15zdnd11an1n04x5 FILLER_334_1068 ();
 b15zdnd00an1n02x5 FILLER_334_1072 ();
 b15zdnd00an1n01x5 FILLER_334_1074 ();
 b15zdnd11an1n16x5 FILLER_334_1080 ();
 b15zdnd00an1n01x5 FILLER_334_1096 ();
 b15zdnd11an1n64x5 FILLER_334_1139 ();
 b15zdnd11an1n16x5 FILLER_334_1203 ();
 b15zdnd11an1n08x5 FILLER_334_1219 ();
 b15zdnd11an1n04x5 FILLER_334_1227 ();
 b15zdnd00an1n02x5 FILLER_334_1231 ();
 b15zdnd00an1n01x5 FILLER_334_1233 ();
 b15zdnd11an1n08x5 FILLER_334_1276 ();
 b15zdnd00an1n01x5 FILLER_334_1284 ();
 b15zdnd11an1n08x5 FILLER_334_1327 ();
 b15zdnd11an1n64x5 FILLER_334_1377 ();
 b15zdnd11an1n64x5 FILLER_334_1441 ();
 b15zdnd11an1n64x5 FILLER_334_1505 ();
 b15zdnd11an1n64x5 FILLER_334_1569 ();
 b15zdnd11an1n64x5 FILLER_334_1633 ();
 b15zdnd11an1n64x5 FILLER_334_1697 ();
 b15zdnd11an1n64x5 FILLER_334_1761 ();
 b15zdnd11an1n16x5 FILLER_334_1825 ();
 b15zdnd00an1n01x5 FILLER_334_1841 ();
 b15zdnd11an1n04x5 FILLER_334_1845 ();
 b15zdnd00an1n01x5 FILLER_334_1849 ();
 b15zdnd11an1n64x5 FILLER_334_1853 ();
 b15zdnd11an1n64x5 FILLER_334_1917 ();
 b15zdnd11an1n64x5 FILLER_334_1981 ();
 b15zdnd11an1n16x5 FILLER_334_2045 ();
 b15zdnd11an1n08x5 FILLER_334_2061 ();
 b15zdnd11an1n04x5 FILLER_334_2069 ();
 b15zdnd11an1n04x5 FILLER_334_2101 ();
 b15zdnd11an1n04x5 FILLER_334_2108 ();
 b15zdnd11an1n32x5 FILLER_334_2115 ();
 b15zdnd11an1n04x5 FILLER_334_2147 ();
 b15zdnd00an1n02x5 FILLER_334_2151 ();
 b15zdnd00an1n01x5 FILLER_334_2153 ();
 b15zdnd11an1n64x5 FILLER_334_2162 ();
 b15zdnd11an1n32x5 FILLER_334_2226 ();
 b15zdnd11an1n16x5 FILLER_334_2258 ();
 b15zdnd00an1n02x5 FILLER_334_2274 ();
 b15zdnd11an1n64x5 FILLER_335_0 ();
 b15zdnd11an1n64x5 FILLER_335_64 ();
 b15zdnd11an1n64x5 FILLER_335_128 ();
 b15zdnd11an1n64x5 FILLER_335_192 ();
 b15zdnd11an1n64x5 FILLER_335_256 ();
 b15zdnd11an1n16x5 FILLER_335_320 ();
 b15zdnd11an1n04x5 FILLER_335_336 ();
 b15zdnd00an1n01x5 FILLER_335_340 ();
 b15zdnd11an1n64x5 FILLER_335_352 ();
 b15zdnd11an1n32x5 FILLER_335_416 ();
 b15zdnd11an1n08x5 FILLER_335_448 ();
 b15zdnd11an1n64x5 FILLER_335_459 ();
 b15zdnd11an1n64x5 FILLER_335_523 ();
 b15zdnd11an1n16x5 FILLER_335_587 ();
 b15zdnd00an1n01x5 FILLER_335_603 ();
 b15zdnd11an1n04x5 FILLER_335_609 ();
 b15zdnd11an1n64x5 FILLER_335_627 ();
 b15zdnd11an1n32x5 FILLER_335_691 ();
 b15zdnd11an1n16x5 FILLER_335_723 ();
 b15zdnd11an1n08x5 FILLER_335_739 ();
 b15zdnd11an1n04x5 FILLER_335_747 ();
 b15zdnd00an1n01x5 FILLER_335_751 ();
 b15zdnd11an1n64x5 FILLER_335_755 ();
 b15zdnd11an1n64x5 FILLER_335_819 ();
 b15zdnd11an1n64x5 FILLER_335_883 ();
 b15zdnd11an1n64x5 FILLER_335_947 ();
 b15zdnd11an1n32x5 FILLER_335_1011 ();
 b15zdnd11an1n16x5 FILLER_335_1043 ();
 b15zdnd11an1n04x5 FILLER_335_1059 ();
 b15zdnd00an1n02x5 FILLER_335_1063 ();
 b15zdnd00an1n01x5 FILLER_335_1065 ();
 b15zdnd11an1n08x5 FILLER_335_1108 ();
 b15zdnd11an1n04x5 FILLER_335_1158 ();
 b15zdnd11an1n64x5 FILLER_335_1165 ();
 b15zdnd11an1n04x5 FILLER_335_1229 ();
 b15zdnd00an1n02x5 FILLER_335_1233 ();
 b15zdnd00an1n01x5 FILLER_335_1235 ();
 b15zdnd11an1n64x5 FILLER_335_1243 ();
 b15zdnd11an1n32x5 FILLER_335_1307 ();
 b15zdnd11an1n08x5 FILLER_335_1339 ();
 b15zdnd00an1n01x5 FILLER_335_1347 ();
 b15zdnd11an1n64x5 FILLER_335_1379 ();
 b15zdnd11an1n64x5 FILLER_335_1443 ();
 b15zdnd11an1n64x5 FILLER_335_1507 ();
 b15zdnd11an1n64x5 FILLER_335_1571 ();
 b15zdnd11an1n64x5 FILLER_335_1635 ();
 b15zdnd11an1n64x5 FILLER_335_1699 ();
 b15zdnd11an1n64x5 FILLER_335_1763 ();
 b15zdnd11an1n08x5 FILLER_335_1827 ();
 b15zdnd00an1n02x5 FILLER_335_1835 ();
 b15zdnd00an1n01x5 FILLER_335_1837 ();
 b15zdnd11an1n04x5 FILLER_335_1841 ();
 b15zdnd11an1n08x5 FILLER_335_1854 ();
 b15zdnd11an1n64x5 FILLER_335_1893 ();
 b15zdnd11an1n32x5 FILLER_335_1957 ();
 b15zdnd11an1n08x5 FILLER_335_1989 ();
 b15zdnd11an1n64x5 FILLER_335_2001 ();
 b15zdnd11an1n08x5 FILLER_335_2065 ();
 b15zdnd11an1n04x5 FILLER_335_2073 ();
 b15zdnd00an1n02x5 FILLER_335_2077 ();
 b15zdnd11an1n64x5 FILLER_335_2121 ();
 b15zdnd11an1n64x5 FILLER_335_2185 ();
 b15zdnd11an1n08x5 FILLER_335_2249 ();
 b15zdnd00an1n02x5 FILLER_335_2257 ();
 b15zdnd11an1n16x5 FILLER_335_2263 ();
 b15zdnd11an1n04x5 FILLER_335_2279 ();
 b15zdnd00an1n01x5 FILLER_335_2283 ();
 b15zdnd11an1n64x5 FILLER_336_8 ();
 b15zdnd11an1n64x5 FILLER_336_72 ();
 b15zdnd11an1n64x5 FILLER_336_136 ();
 b15zdnd11an1n64x5 FILLER_336_200 ();
 b15zdnd11an1n64x5 FILLER_336_264 ();
 b15zdnd11an1n64x5 FILLER_336_328 ();
 b15zdnd11an1n64x5 FILLER_336_392 ();
 b15zdnd11an1n04x5 FILLER_336_456 ();
 b15zdnd11an1n16x5 FILLER_336_470 ();
 b15zdnd11an1n04x5 FILLER_336_486 ();
 b15zdnd00an1n02x5 FILLER_336_490 ();
 b15zdnd00an1n01x5 FILLER_336_492 ();
 b15zdnd11an1n64x5 FILLER_336_502 ();
 b15zdnd11an1n32x5 FILLER_336_566 ();
 b15zdnd11an1n04x5 FILLER_336_598 ();
 b15zdnd00an1n02x5 FILLER_336_602 ();
 b15zdnd00an1n01x5 FILLER_336_604 ();
 b15zdnd11an1n08x5 FILLER_336_608 ();
 b15zdnd11an1n04x5 FILLER_336_616 ();
 b15zdnd00an1n02x5 FILLER_336_620 ();
 b15zdnd11an1n64x5 FILLER_336_625 ();
 b15zdnd11an1n16x5 FILLER_336_689 ();
 b15zdnd11an1n08x5 FILLER_336_705 ();
 b15zdnd11an1n04x5 FILLER_336_713 ();
 b15zdnd00an1n01x5 FILLER_336_717 ();
 b15zdnd11an1n16x5 FILLER_336_726 ();
 b15zdnd11an1n08x5 FILLER_336_742 ();
 b15zdnd00an1n01x5 FILLER_336_750 ();
 b15zdnd11an1n64x5 FILLER_336_754 ();
 b15zdnd11an1n64x5 FILLER_336_818 ();
 b15zdnd11an1n64x5 FILLER_336_882 ();
 b15zdnd11an1n64x5 FILLER_336_946 ();
 b15zdnd11an1n64x5 FILLER_336_1010 ();
 b15zdnd11an1n04x5 FILLER_336_1074 ();
 b15zdnd00an1n02x5 FILLER_336_1078 ();
 b15zdnd00an1n01x5 FILLER_336_1080 ();
 b15zdnd11an1n16x5 FILLER_336_1133 ();
 b15zdnd11an1n08x5 FILLER_336_1149 ();
 b15zdnd11an1n04x5 FILLER_336_1157 ();
 b15zdnd00an1n01x5 FILLER_336_1161 ();
 b15zdnd11an1n64x5 FILLER_336_1165 ();
 b15zdnd11an1n64x5 FILLER_336_1229 ();
 b15zdnd11an1n64x5 FILLER_336_1293 ();
 b15zdnd11an1n64x5 FILLER_336_1357 ();
 b15zdnd11an1n32x5 FILLER_336_1421 ();
 b15zdnd11an1n04x5 FILLER_336_1453 ();
 b15zdnd00an1n02x5 FILLER_336_1457 ();
 b15zdnd00an1n01x5 FILLER_336_1459 ();
 b15zdnd11an1n64x5 FILLER_336_1463 ();
 b15zdnd11an1n64x5 FILLER_336_1527 ();
 b15zdnd11an1n64x5 FILLER_336_1591 ();
 b15zdnd11an1n64x5 FILLER_336_1655 ();
 b15zdnd11an1n64x5 FILLER_336_1719 ();
 b15zdnd11an1n32x5 FILLER_336_1783 ();
 b15zdnd11an1n04x5 FILLER_336_1815 ();
 b15zdnd00an1n01x5 FILLER_336_1819 ();
 b15zdnd11an1n64x5 FILLER_336_1872 ();
 b15zdnd11an1n64x5 FILLER_336_1936 ();
 b15zdnd11an1n32x5 FILLER_336_2000 ();
 b15zdnd11an1n16x5 FILLER_336_2032 ();
 b15zdnd11an1n08x5 FILLER_336_2048 ();
 b15zdnd11an1n04x5 FILLER_336_2056 ();
 b15zdnd00an1n02x5 FILLER_336_2060 ();
 b15zdnd00an1n01x5 FILLER_336_2062 ();
 b15zdnd11an1n32x5 FILLER_336_2115 ();
 b15zdnd11an1n04x5 FILLER_336_2147 ();
 b15zdnd00an1n02x5 FILLER_336_2151 ();
 b15zdnd00an1n01x5 FILLER_336_2153 ();
 b15zdnd11an1n64x5 FILLER_336_2162 ();
 b15zdnd11an1n32x5 FILLER_336_2226 ();
 b15zdnd11an1n16x5 FILLER_336_2258 ();
 b15zdnd00an1n02x5 FILLER_336_2274 ();
 b15zdnd11an1n64x5 FILLER_337_0 ();
 b15zdnd11an1n64x5 FILLER_337_64 ();
 b15zdnd11an1n64x5 FILLER_337_128 ();
 b15zdnd11an1n64x5 FILLER_337_192 ();
 b15zdnd11an1n64x5 FILLER_337_256 ();
 b15zdnd11an1n64x5 FILLER_337_320 ();
 b15zdnd11an1n64x5 FILLER_337_384 ();
 b15zdnd11an1n64x5 FILLER_337_448 ();
 b15zdnd11an1n64x5 FILLER_337_512 ();
 b15zdnd11an1n16x5 FILLER_337_576 ();
 b15zdnd11an1n08x5 FILLER_337_592 ();
 b15zdnd11an1n04x5 FILLER_337_600 ();
 b15zdnd00an1n01x5 FILLER_337_604 ();
 b15zdnd11an1n64x5 FILLER_337_610 ();
 b15zdnd11an1n64x5 FILLER_337_674 ();
 b15zdnd11an1n64x5 FILLER_337_738 ();
 b15zdnd11an1n64x5 FILLER_337_802 ();
 b15zdnd11an1n64x5 FILLER_337_866 ();
 b15zdnd11an1n64x5 FILLER_337_930 ();
 b15zdnd11an1n64x5 FILLER_337_994 ();
 b15zdnd11an1n32x5 FILLER_337_1058 ();
 b15zdnd00an1n01x5 FILLER_337_1090 ();
 b15zdnd11an1n04x5 FILLER_337_1133 ();
 b15zdnd11an1n64x5 FILLER_337_1189 ();
 b15zdnd11an1n64x5 FILLER_337_1253 ();
 b15zdnd11an1n16x5 FILLER_337_1317 ();
 b15zdnd11an1n08x5 FILLER_337_1333 ();
 b15zdnd00an1n01x5 FILLER_337_1341 ();
 b15zdnd11an1n32x5 FILLER_337_1353 ();
 b15zdnd11an1n16x5 FILLER_337_1385 ();
 b15zdnd11an1n16x5 FILLER_337_1443 ();
 b15zdnd11an1n64x5 FILLER_337_1462 ();
 b15zdnd11an1n64x5 FILLER_337_1526 ();
 b15zdnd11an1n64x5 FILLER_337_1590 ();
 b15zdnd11an1n64x5 FILLER_337_1654 ();
 b15zdnd11an1n64x5 FILLER_337_1718 ();
 b15zdnd11an1n64x5 FILLER_337_1782 ();
 b15zdnd11an1n64x5 FILLER_337_1846 ();
 b15zdnd11an1n64x5 FILLER_337_1910 ();
 b15zdnd11an1n16x5 FILLER_337_1974 ();
 b15zdnd11an1n04x5 FILLER_337_1990 ();
 b15zdnd00an1n01x5 FILLER_337_1994 ();
 b15zdnd11an1n32x5 FILLER_337_2020 ();
 b15zdnd11an1n16x5 FILLER_337_2052 ();
 b15zdnd11an1n08x5 FILLER_337_2068 ();
 b15zdnd11an1n04x5 FILLER_337_2076 ();
 b15zdnd00an1n01x5 FILLER_337_2080 ();
 b15zdnd11an1n04x5 FILLER_337_2084 ();
 b15zdnd11an1n08x5 FILLER_337_2091 ();
 b15zdnd11an1n04x5 FILLER_337_2099 ();
 b15zdnd00an1n01x5 FILLER_337_2103 ();
 b15zdnd11an1n64x5 FILLER_337_2146 ();
 b15zdnd11an1n64x5 FILLER_337_2210 ();
 b15zdnd11an1n08x5 FILLER_337_2274 ();
 b15zdnd00an1n02x5 FILLER_337_2282 ();
 b15zdnd11an1n64x5 FILLER_338_8 ();
 b15zdnd11an1n64x5 FILLER_338_72 ();
 b15zdnd11an1n64x5 FILLER_338_136 ();
 b15zdnd11an1n64x5 FILLER_338_200 ();
 b15zdnd11an1n64x5 FILLER_338_264 ();
 b15zdnd11an1n64x5 FILLER_338_328 ();
 b15zdnd11an1n64x5 FILLER_338_392 ();
 b15zdnd11an1n64x5 FILLER_338_456 ();
 b15zdnd11an1n64x5 FILLER_338_520 ();
 b15zdnd11an1n64x5 FILLER_338_584 ();
 b15zdnd11an1n64x5 FILLER_338_648 ();
 b15zdnd11an1n04x5 FILLER_338_712 ();
 b15zdnd00an1n02x5 FILLER_338_716 ();
 b15zdnd11an1n64x5 FILLER_338_726 ();
 b15zdnd11an1n64x5 FILLER_338_790 ();
 b15zdnd11an1n64x5 FILLER_338_854 ();
 b15zdnd11an1n64x5 FILLER_338_918 ();
 b15zdnd11an1n64x5 FILLER_338_982 ();
 b15zdnd11an1n32x5 FILLER_338_1046 ();
 b15zdnd11an1n16x5 FILLER_338_1078 ();
 b15zdnd11an1n04x5 FILLER_338_1094 ();
 b15zdnd00an1n01x5 FILLER_338_1098 ();
 b15zdnd11an1n04x5 FILLER_338_1102 ();
 b15zdnd11an1n32x5 FILLER_338_1109 ();
 b15zdnd11an1n16x5 FILLER_338_1141 ();
 b15zdnd11an1n04x5 FILLER_338_1157 ();
 b15zdnd00an1n02x5 FILLER_338_1161 ();
 b15zdnd11an1n64x5 FILLER_338_1166 ();
 b15zdnd11an1n64x5 FILLER_338_1230 ();
 b15zdnd11an1n64x5 FILLER_338_1294 ();
 b15zdnd11an1n64x5 FILLER_338_1358 ();
 b15zdnd11an1n08x5 FILLER_338_1422 ();
 b15zdnd11an1n04x5 FILLER_338_1430 ();
 b15zdnd11an1n64x5 FILLER_338_1486 ();
 b15zdnd11an1n64x5 FILLER_338_1550 ();
 b15zdnd11an1n64x5 FILLER_338_1614 ();
 b15zdnd11an1n64x5 FILLER_338_1678 ();
 b15zdnd11an1n64x5 FILLER_338_1742 ();
 b15zdnd11an1n64x5 FILLER_338_1806 ();
 b15zdnd11an1n64x5 FILLER_338_1870 ();
 b15zdnd11an1n64x5 FILLER_338_1934 ();
 b15zdnd11an1n64x5 FILLER_338_1998 ();
 b15zdnd11an1n64x5 FILLER_338_2062 ();
 b15zdnd11an1n16x5 FILLER_338_2126 ();
 b15zdnd11an1n08x5 FILLER_338_2142 ();
 b15zdnd11an1n04x5 FILLER_338_2150 ();
 b15zdnd11an1n64x5 FILLER_338_2162 ();
 b15zdnd11an1n32x5 FILLER_338_2226 ();
 b15zdnd11an1n16x5 FILLER_338_2258 ();
 b15zdnd00an1n02x5 FILLER_338_2274 ();
 b15zdnd11an1n64x5 FILLER_339_0 ();
 b15zdnd11an1n64x5 FILLER_339_64 ();
 b15zdnd11an1n64x5 FILLER_339_128 ();
 b15zdnd11an1n64x5 FILLER_339_192 ();
 b15zdnd11an1n64x5 FILLER_339_256 ();
 b15zdnd11an1n08x5 FILLER_339_320 ();
 b15zdnd11an1n04x5 FILLER_339_328 ();
 b15zdnd00an1n02x5 FILLER_339_332 ();
 b15zdnd11an1n64x5 FILLER_339_376 ();
 b15zdnd11an1n64x5 FILLER_339_440 ();
 b15zdnd11an1n64x5 FILLER_339_504 ();
 b15zdnd11an1n32x5 FILLER_339_568 ();
 b15zdnd11an1n04x5 FILLER_339_600 ();
 b15zdnd00an1n01x5 FILLER_339_604 ();
 b15zdnd11an1n64x5 FILLER_339_609 ();
 b15zdnd11an1n64x5 FILLER_339_673 ();
 b15zdnd11an1n64x5 FILLER_339_737 ();
 b15zdnd11an1n64x5 FILLER_339_801 ();
 b15zdnd11an1n64x5 FILLER_339_865 ();
 b15zdnd11an1n64x5 FILLER_339_929 ();
 b15zdnd11an1n64x5 FILLER_339_993 ();
 b15zdnd11an1n08x5 FILLER_339_1057 ();
 b15zdnd11an1n04x5 FILLER_339_1065 ();
 b15zdnd11an1n04x5 FILLER_339_1114 ();
 b15zdnd11an1n64x5 FILLER_339_1125 ();
 b15zdnd11an1n16x5 FILLER_339_1189 ();
 b15zdnd11an1n08x5 FILLER_339_1205 ();
 b15zdnd00an1n01x5 FILLER_339_1213 ();
 b15zdnd11an1n64x5 FILLER_339_1256 ();
 b15zdnd11an1n64x5 FILLER_339_1320 ();
 b15zdnd11an1n64x5 FILLER_339_1384 ();
 b15zdnd11an1n08x5 FILLER_339_1448 ();
 b15zdnd00an1n02x5 FILLER_339_1456 ();
 b15zdnd00an1n01x5 FILLER_339_1458 ();
 b15zdnd11an1n64x5 FILLER_339_1462 ();
 b15zdnd11an1n64x5 FILLER_339_1526 ();
 b15zdnd11an1n64x5 FILLER_339_1590 ();
 b15zdnd11an1n64x5 FILLER_339_1654 ();
 b15zdnd11an1n64x5 FILLER_339_1718 ();
 b15zdnd11an1n64x5 FILLER_339_1782 ();
 b15zdnd11an1n64x5 FILLER_339_1846 ();
 b15zdnd11an1n64x5 FILLER_339_1910 ();
 b15zdnd11an1n64x5 FILLER_339_1974 ();
 b15zdnd11an1n64x5 FILLER_339_2038 ();
 b15zdnd11an1n64x5 FILLER_339_2102 ();
 b15zdnd11an1n64x5 FILLER_339_2166 ();
 b15zdnd11an1n32x5 FILLER_339_2230 ();
 b15zdnd11an1n16x5 FILLER_339_2262 ();
 b15zdnd11an1n04x5 FILLER_339_2278 ();
 b15zdnd00an1n02x5 FILLER_339_2282 ();
 b15zdnd11an1n64x5 FILLER_340_8 ();
 b15zdnd11an1n64x5 FILLER_340_72 ();
 b15zdnd11an1n64x5 FILLER_340_136 ();
 b15zdnd11an1n64x5 FILLER_340_200 ();
 b15zdnd11an1n64x5 FILLER_340_264 ();
 b15zdnd11an1n64x5 FILLER_340_328 ();
 b15zdnd11an1n64x5 FILLER_340_392 ();
 b15zdnd11an1n64x5 FILLER_340_456 ();
 b15zdnd11an1n64x5 FILLER_340_520 ();
 b15zdnd11an1n64x5 FILLER_340_584 ();
 b15zdnd11an1n64x5 FILLER_340_648 ();
 b15zdnd11an1n04x5 FILLER_340_712 ();
 b15zdnd00an1n02x5 FILLER_340_716 ();
 b15zdnd11an1n32x5 FILLER_340_726 ();
 b15zdnd11an1n16x5 FILLER_340_758 ();
 b15zdnd11an1n32x5 FILLER_340_816 ();
 b15zdnd11an1n16x5 FILLER_340_848 ();
 b15zdnd11an1n04x5 FILLER_340_864 ();
 b15zdnd00an1n02x5 FILLER_340_868 ();
 b15zdnd00an1n01x5 FILLER_340_870 ();
 b15zdnd11an1n64x5 FILLER_340_874 ();
 b15zdnd11an1n64x5 FILLER_340_938 ();
 b15zdnd11an1n64x5 FILLER_340_1002 ();
 b15zdnd11an1n64x5 FILLER_340_1066 ();
 b15zdnd11an1n64x5 FILLER_340_1130 ();
 b15zdnd11an1n64x5 FILLER_340_1194 ();
 b15zdnd11an1n64x5 FILLER_340_1258 ();
 b15zdnd11an1n64x5 FILLER_340_1322 ();
 b15zdnd11an1n64x5 FILLER_340_1386 ();
 b15zdnd11an1n64x5 FILLER_340_1450 ();
 b15zdnd11an1n64x5 FILLER_340_1514 ();
 b15zdnd11an1n64x5 FILLER_340_1578 ();
 b15zdnd11an1n64x5 FILLER_340_1642 ();
 b15zdnd11an1n64x5 FILLER_340_1706 ();
 b15zdnd11an1n16x5 FILLER_340_1770 ();
 b15zdnd11an1n08x5 FILLER_340_1786 ();
 b15zdnd00an1n01x5 FILLER_340_1794 ();
 b15zdnd11an1n64x5 FILLER_340_1804 ();
 b15zdnd11an1n64x5 FILLER_340_1868 ();
 b15zdnd11an1n64x5 FILLER_340_1932 ();
 b15zdnd11an1n64x5 FILLER_340_1996 ();
 b15zdnd11an1n64x5 FILLER_340_2060 ();
 b15zdnd11an1n16x5 FILLER_340_2124 ();
 b15zdnd11an1n08x5 FILLER_340_2140 ();
 b15zdnd11an1n04x5 FILLER_340_2148 ();
 b15zdnd00an1n02x5 FILLER_340_2152 ();
 b15zdnd11an1n64x5 FILLER_340_2162 ();
 b15zdnd11an1n32x5 FILLER_340_2226 ();
 b15zdnd11an1n16x5 FILLER_340_2258 ();
 b15zdnd00an1n02x5 FILLER_340_2274 ();
 b15zdnd11an1n64x5 FILLER_341_0 ();
 b15zdnd11an1n64x5 FILLER_341_64 ();
 b15zdnd11an1n64x5 FILLER_341_128 ();
 b15zdnd11an1n64x5 FILLER_341_192 ();
 b15zdnd11an1n64x5 FILLER_341_256 ();
 b15zdnd11an1n64x5 FILLER_341_320 ();
 b15zdnd11an1n64x5 FILLER_341_384 ();
 b15zdnd11an1n64x5 FILLER_341_448 ();
 b15zdnd11an1n64x5 FILLER_341_512 ();
 b15zdnd11an1n64x5 FILLER_341_576 ();
 b15zdnd11an1n64x5 FILLER_341_640 ();
 b15zdnd11an1n64x5 FILLER_341_704 ();
 b15zdnd11an1n64x5 FILLER_341_768 ();
 b15zdnd11an1n04x5 FILLER_341_832 ();
 b15zdnd00an1n01x5 FILLER_341_836 ();
 b15zdnd11an1n04x5 FILLER_341_877 ();
 b15zdnd11an1n64x5 FILLER_341_884 ();
 b15zdnd11an1n64x5 FILLER_341_948 ();
 b15zdnd11an1n64x5 FILLER_341_1012 ();
 b15zdnd11an1n64x5 FILLER_341_1076 ();
 b15zdnd11an1n64x5 FILLER_341_1140 ();
 b15zdnd11an1n64x5 FILLER_341_1204 ();
 b15zdnd11an1n64x5 FILLER_341_1268 ();
 b15zdnd11an1n64x5 FILLER_341_1332 ();
 b15zdnd11an1n64x5 FILLER_341_1396 ();
 b15zdnd11an1n64x5 FILLER_341_1460 ();
 b15zdnd11an1n64x5 FILLER_341_1524 ();
 b15zdnd11an1n64x5 FILLER_341_1588 ();
 b15zdnd11an1n64x5 FILLER_341_1652 ();
 b15zdnd11an1n64x5 FILLER_341_1716 ();
 b15zdnd11an1n16x5 FILLER_341_1780 ();
 b15zdnd11an1n08x5 FILLER_341_1796 ();
 b15zdnd00an1n02x5 FILLER_341_1804 ();
 b15zdnd00an1n01x5 FILLER_341_1806 ();
 b15zdnd11an1n64x5 FILLER_341_1813 ();
 b15zdnd11an1n64x5 FILLER_341_1877 ();
 b15zdnd11an1n64x5 FILLER_341_1941 ();
 b15zdnd11an1n64x5 FILLER_341_2005 ();
 b15zdnd11an1n64x5 FILLER_341_2069 ();
 b15zdnd11an1n64x5 FILLER_341_2133 ();
 b15zdnd11an1n64x5 FILLER_341_2197 ();
 b15zdnd11an1n16x5 FILLER_341_2261 ();
 b15zdnd11an1n04x5 FILLER_341_2277 ();
 b15zdnd00an1n02x5 FILLER_341_2281 ();
 b15zdnd00an1n01x5 FILLER_341_2283 ();
 b15zdnd11an1n64x5 FILLER_342_8 ();
 b15zdnd11an1n64x5 FILLER_342_72 ();
 b15zdnd11an1n64x5 FILLER_342_136 ();
 b15zdnd11an1n64x5 FILLER_342_200 ();
 b15zdnd11an1n64x5 FILLER_342_264 ();
 b15zdnd11an1n64x5 FILLER_342_328 ();
 b15zdnd11an1n64x5 FILLER_342_392 ();
 b15zdnd11an1n64x5 FILLER_342_456 ();
 b15zdnd11an1n64x5 FILLER_342_520 ();
 b15zdnd11an1n64x5 FILLER_342_584 ();
 b15zdnd11an1n64x5 FILLER_342_648 ();
 b15zdnd11an1n04x5 FILLER_342_712 ();
 b15zdnd00an1n02x5 FILLER_342_716 ();
 b15zdnd11an1n64x5 FILLER_342_726 ();
 b15zdnd11an1n64x5 FILLER_342_790 ();
 b15zdnd11an1n64x5 FILLER_342_854 ();
 b15zdnd11an1n64x5 FILLER_342_918 ();
 b15zdnd11an1n64x5 FILLER_342_982 ();
 b15zdnd11an1n64x5 FILLER_342_1046 ();
 b15zdnd11an1n64x5 FILLER_342_1110 ();
 b15zdnd11an1n64x5 FILLER_342_1174 ();
 b15zdnd11an1n64x5 FILLER_342_1238 ();
 b15zdnd11an1n08x5 FILLER_342_1302 ();
 b15zdnd11an1n04x5 FILLER_342_1310 ();
 b15zdnd00an1n02x5 FILLER_342_1314 ();
 b15zdnd00an1n01x5 FILLER_342_1316 ();
 b15zdnd11an1n64x5 FILLER_342_1359 ();
 b15zdnd11an1n64x5 FILLER_342_1423 ();
 b15zdnd11an1n64x5 FILLER_342_1487 ();
 b15zdnd11an1n64x5 FILLER_342_1551 ();
 b15zdnd11an1n64x5 FILLER_342_1615 ();
 b15zdnd11an1n64x5 FILLER_342_1679 ();
 b15zdnd11an1n32x5 FILLER_342_1743 ();
 b15zdnd11an1n08x5 FILLER_342_1775 ();
 b15zdnd00an1n02x5 FILLER_342_1783 ();
 b15zdnd11an1n04x5 FILLER_342_1788 ();
 b15zdnd11an1n08x5 FILLER_342_1795 ();
 b15zdnd11an1n04x5 FILLER_342_1803 ();
 b15zdnd00an1n01x5 FILLER_342_1807 ();
 b15zdnd11an1n64x5 FILLER_342_1850 ();
 b15zdnd11an1n64x5 FILLER_342_1914 ();
 b15zdnd11an1n64x5 FILLER_342_1978 ();
 b15zdnd11an1n64x5 FILLER_342_2042 ();
 b15zdnd11an1n32x5 FILLER_342_2106 ();
 b15zdnd11an1n16x5 FILLER_342_2138 ();
 b15zdnd11an1n64x5 FILLER_342_2162 ();
 b15zdnd11an1n32x5 FILLER_342_2226 ();
 b15zdnd11an1n16x5 FILLER_342_2258 ();
 b15zdnd00an1n02x5 FILLER_342_2274 ();
 b15zdnd11an1n64x5 FILLER_343_0 ();
 b15zdnd11an1n64x5 FILLER_343_64 ();
 b15zdnd11an1n64x5 FILLER_343_128 ();
 b15zdnd11an1n64x5 FILLER_343_192 ();
 b15zdnd11an1n64x5 FILLER_343_256 ();
 b15zdnd11an1n64x5 FILLER_343_320 ();
 b15zdnd11an1n64x5 FILLER_343_384 ();
 b15zdnd11an1n64x5 FILLER_343_448 ();
 b15zdnd11an1n04x5 FILLER_343_512 ();
 b15zdnd00an1n02x5 FILLER_343_516 ();
 b15zdnd11an1n08x5 FILLER_343_521 ();
 b15zdnd11an1n04x5 FILLER_343_529 ();
 b15zdnd00an1n02x5 FILLER_343_533 ();
 b15zdnd00an1n01x5 FILLER_343_535 ();
 b15zdnd11an1n32x5 FILLER_343_547 ();
 b15zdnd11an1n16x5 FILLER_343_579 ();
 b15zdnd11an1n08x5 FILLER_343_595 ();
 b15zdnd11an1n04x5 FILLER_343_603 ();
 b15zdnd00an1n01x5 FILLER_343_607 ();
 b15zdnd11an1n64x5 FILLER_343_614 ();
 b15zdnd11an1n64x5 FILLER_343_678 ();
 b15zdnd11an1n64x5 FILLER_343_742 ();
 b15zdnd11an1n16x5 FILLER_343_806 ();
 b15zdnd00an1n02x5 FILLER_343_822 ();
 b15zdnd11an1n64x5 FILLER_343_827 ();
 b15zdnd11an1n64x5 FILLER_343_891 ();
 b15zdnd11an1n64x5 FILLER_343_955 ();
 b15zdnd11an1n64x5 FILLER_343_1019 ();
 b15zdnd11an1n08x5 FILLER_343_1083 ();
 b15zdnd11an1n64x5 FILLER_343_1133 ();
 b15zdnd11an1n64x5 FILLER_343_1197 ();
 b15zdnd11an1n64x5 FILLER_343_1261 ();
 b15zdnd11an1n64x5 FILLER_343_1325 ();
 b15zdnd11an1n64x5 FILLER_343_1389 ();
 b15zdnd11an1n64x5 FILLER_343_1453 ();
 b15zdnd11an1n64x5 FILLER_343_1517 ();
 b15zdnd11an1n64x5 FILLER_343_1581 ();
 b15zdnd11an1n64x5 FILLER_343_1645 ();
 b15zdnd11an1n32x5 FILLER_343_1709 ();
 b15zdnd11an1n16x5 FILLER_343_1741 ();
 b15zdnd11an1n08x5 FILLER_343_1757 ();
 b15zdnd00an1n02x5 FILLER_343_1765 ();
 b15zdnd11an1n64x5 FILLER_343_1819 ();
 b15zdnd11an1n64x5 FILLER_343_1883 ();
 b15zdnd11an1n64x5 FILLER_343_1947 ();
 b15zdnd11an1n64x5 FILLER_343_2011 ();
 b15zdnd11an1n64x5 FILLER_343_2075 ();
 b15zdnd11an1n64x5 FILLER_343_2139 ();
 b15zdnd11an1n64x5 FILLER_343_2203 ();
 b15zdnd11an1n16x5 FILLER_343_2267 ();
 b15zdnd00an1n01x5 FILLER_343_2283 ();
 b15zdnd11an1n64x5 FILLER_344_8 ();
 b15zdnd11an1n64x5 FILLER_344_72 ();
 b15zdnd11an1n64x5 FILLER_344_136 ();
 b15zdnd11an1n64x5 FILLER_344_200 ();
 b15zdnd11an1n64x5 FILLER_344_264 ();
 b15zdnd11an1n64x5 FILLER_344_328 ();
 b15zdnd11an1n64x5 FILLER_344_392 ();
 b15zdnd11an1n16x5 FILLER_344_456 ();
 b15zdnd11an1n08x5 FILLER_344_472 ();
 b15zdnd11an1n04x5 FILLER_344_480 ();
 b15zdnd11an1n64x5 FILLER_344_524 ();
 b15zdnd11an1n16x5 FILLER_344_588 ();
 b15zdnd11an1n04x5 FILLER_344_604 ();
 b15zdnd00an1n02x5 FILLER_344_608 ();
 b15zdnd00an1n01x5 FILLER_344_610 ();
 b15zdnd11an1n64x5 FILLER_344_614 ();
 b15zdnd11an1n32x5 FILLER_344_678 ();
 b15zdnd11an1n08x5 FILLER_344_710 ();
 b15zdnd11an1n64x5 FILLER_344_726 ();
 b15zdnd11an1n16x5 FILLER_344_790 ();
 b15zdnd11an1n08x5 FILLER_344_806 ();
 b15zdnd11an1n04x5 FILLER_344_814 ();
 b15zdnd00an1n02x5 FILLER_344_818 ();
 b15zdnd00an1n01x5 FILLER_344_820 ();
 b15zdnd11an1n64x5 FILLER_344_863 ();
 b15zdnd11an1n64x5 FILLER_344_927 ();
 b15zdnd11an1n64x5 FILLER_344_991 ();
 b15zdnd11an1n64x5 FILLER_344_1055 ();
 b15zdnd11an1n64x5 FILLER_344_1119 ();
 b15zdnd11an1n32x5 FILLER_344_1183 ();
 b15zdnd11an1n16x5 FILLER_344_1215 ();
 b15zdnd11an1n08x5 FILLER_344_1231 ();
 b15zdnd00an1n01x5 FILLER_344_1239 ();
 b15zdnd11an1n32x5 FILLER_344_1292 ();
 b15zdnd00an1n02x5 FILLER_344_1324 ();
 b15zdnd11an1n16x5 FILLER_344_1368 ();
 b15zdnd00an1n02x5 FILLER_344_1384 ();
 b15zdnd11an1n64x5 FILLER_344_1396 ();
 b15zdnd11an1n32x5 FILLER_344_1460 ();
 b15zdnd11an1n04x5 FILLER_344_1492 ();
 b15zdnd00an1n01x5 FILLER_344_1496 ();
 b15zdnd11an1n32x5 FILLER_344_1522 ();
 b15zdnd11an1n16x5 FILLER_344_1554 ();
 b15zdnd11an1n04x5 FILLER_344_1570 ();
 b15zdnd00an1n01x5 FILLER_344_1574 ();
 b15zdnd11an1n64x5 FILLER_344_1586 ();
 b15zdnd11an1n64x5 FILLER_344_1650 ();
 b15zdnd11an1n64x5 FILLER_344_1714 ();
 b15zdnd11an1n08x5 FILLER_344_1778 ();
 b15zdnd11an1n04x5 FILLER_344_1786 ();
 b15zdnd00an1n02x5 FILLER_344_1790 ();
 b15zdnd11an1n04x5 FILLER_344_1795 ();
 b15zdnd11an1n04x5 FILLER_344_1805 ();
 b15zdnd00an1n01x5 FILLER_344_1809 ();
 b15zdnd11an1n64x5 FILLER_344_1852 ();
 b15zdnd11an1n64x5 FILLER_344_1916 ();
 b15zdnd11an1n64x5 FILLER_344_1980 ();
 b15zdnd11an1n64x5 FILLER_344_2044 ();
 b15zdnd11an1n32x5 FILLER_344_2108 ();
 b15zdnd11an1n08x5 FILLER_344_2140 ();
 b15zdnd11an1n04x5 FILLER_344_2148 ();
 b15zdnd00an1n02x5 FILLER_344_2152 ();
 b15zdnd11an1n64x5 FILLER_344_2162 ();
 b15zdnd11an1n32x5 FILLER_344_2226 ();
 b15zdnd11an1n16x5 FILLER_344_2258 ();
 b15zdnd00an1n02x5 FILLER_344_2274 ();
 b15zdnd11an1n64x5 FILLER_345_0 ();
 b15zdnd11an1n64x5 FILLER_345_64 ();
 b15zdnd11an1n64x5 FILLER_345_128 ();
 b15zdnd11an1n64x5 FILLER_345_192 ();
 b15zdnd11an1n64x5 FILLER_345_256 ();
 b15zdnd11an1n16x5 FILLER_345_320 ();
 b15zdnd11an1n08x5 FILLER_345_336 ();
 b15zdnd00an1n02x5 FILLER_345_344 ();
 b15zdnd11an1n64x5 FILLER_345_349 ();
 b15zdnd11an1n64x5 FILLER_345_413 ();
 b15zdnd11an1n32x5 FILLER_345_477 ();
 b15zdnd11an1n08x5 FILLER_345_509 ();
 b15zdnd00an1n02x5 FILLER_345_517 ();
 b15zdnd00an1n01x5 FILLER_345_519 ();
 b15zdnd11an1n64x5 FILLER_345_523 ();
 b15zdnd11an1n64x5 FILLER_345_587 ();
 b15zdnd11an1n32x5 FILLER_345_651 ();
 b15zdnd11an1n16x5 FILLER_345_683 ();
 b15zdnd00an1n01x5 FILLER_345_699 ();
 b15zdnd11an1n04x5 FILLER_345_752 ();
 b15zdnd11an1n04x5 FILLER_345_760 ();
 b15zdnd11an1n16x5 FILLER_345_768 ();
 b15zdnd11an1n08x5 FILLER_345_784 ();
 b15zdnd11an1n04x5 FILLER_345_792 ();
 b15zdnd00an1n01x5 FILLER_345_796 ();
 b15zdnd11an1n64x5 FILLER_345_849 ();
 b15zdnd11an1n64x5 FILLER_345_913 ();
 b15zdnd11an1n64x5 FILLER_345_977 ();
 b15zdnd11an1n64x5 FILLER_345_1041 ();
 b15zdnd11an1n16x5 FILLER_345_1105 ();
 b15zdnd11an1n04x5 FILLER_345_1121 ();
 b15zdnd00an1n02x5 FILLER_345_1125 ();
 b15zdnd00an1n01x5 FILLER_345_1127 ();
 b15zdnd11an1n64x5 FILLER_345_1142 ();
 b15zdnd11an1n32x5 FILLER_345_1206 ();
 b15zdnd11an1n08x5 FILLER_345_1238 ();
 b15zdnd00an1n01x5 FILLER_345_1246 ();
 b15zdnd11an1n04x5 FILLER_345_1254 ();
 b15zdnd11an1n04x5 FILLER_345_1261 ();
 b15zdnd11an1n32x5 FILLER_345_1268 ();
 b15zdnd11an1n04x5 FILLER_345_1300 ();
 b15zdnd00an1n02x5 FILLER_345_1304 ();
 b15zdnd00an1n01x5 FILLER_345_1306 ();
 b15zdnd11an1n64x5 FILLER_345_1317 ();
 b15zdnd11an1n32x5 FILLER_345_1381 ();
 b15zdnd11an1n08x5 FILLER_345_1413 ();
 b15zdnd11an1n04x5 FILLER_345_1421 ();
 b15zdnd00an1n01x5 FILLER_345_1425 ();
 b15zdnd11an1n64x5 FILLER_345_1444 ();
 b15zdnd11an1n64x5 FILLER_345_1508 ();
 b15zdnd11an1n64x5 FILLER_345_1572 ();
 b15zdnd11an1n32x5 FILLER_345_1636 ();
 b15zdnd11an1n16x5 FILLER_345_1668 ();
 b15zdnd11an1n08x5 FILLER_345_1684 ();
 b15zdnd11an1n04x5 FILLER_345_1692 ();
 b15zdnd00an1n01x5 FILLER_345_1696 ();
 b15zdnd11an1n04x5 FILLER_345_1739 ();
 b15zdnd11an1n64x5 FILLER_345_1785 ();
 b15zdnd11an1n64x5 FILLER_345_1849 ();
 b15zdnd11an1n64x5 FILLER_345_1913 ();
 b15zdnd11an1n64x5 FILLER_345_1977 ();
 b15zdnd11an1n64x5 FILLER_345_2041 ();
 b15zdnd11an1n64x5 FILLER_345_2105 ();
 b15zdnd11an1n64x5 FILLER_345_2169 ();
 b15zdnd11an1n32x5 FILLER_345_2233 ();
 b15zdnd11an1n16x5 FILLER_345_2265 ();
 b15zdnd00an1n02x5 FILLER_345_2281 ();
 b15zdnd00an1n01x5 FILLER_345_2283 ();
 b15zdnd11an1n64x5 FILLER_346_8 ();
 b15zdnd11an1n64x5 FILLER_346_72 ();
 b15zdnd11an1n64x5 FILLER_346_136 ();
 b15zdnd11an1n64x5 FILLER_346_200 ();
 b15zdnd11an1n32x5 FILLER_346_264 ();
 b15zdnd11an1n16x5 FILLER_346_296 ();
 b15zdnd11an1n04x5 FILLER_346_312 ();
 b15zdnd00an1n02x5 FILLER_346_316 ();
 b15zdnd00an1n01x5 FILLER_346_318 ();
 b15zdnd11an1n64x5 FILLER_346_371 ();
 b15zdnd11an1n64x5 FILLER_346_435 ();
 b15zdnd11an1n64x5 FILLER_346_499 ();
 b15zdnd11an1n64x5 FILLER_346_563 ();
 b15zdnd11an1n64x5 FILLER_346_627 ();
 b15zdnd11an1n16x5 FILLER_346_691 ();
 b15zdnd11an1n08x5 FILLER_346_707 ();
 b15zdnd00an1n02x5 FILLER_346_715 ();
 b15zdnd00an1n01x5 FILLER_346_717 ();
 b15zdnd11an1n04x5 FILLER_346_726 ();
 b15zdnd11an1n08x5 FILLER_346_772 ();
 b15zdnd11an1n04x5 FILLER_346_822 ();
 b15zdnd11an1n64x5 FILLER_346_829 ();
 b15zdnd11an1n64x5 FILLER_346_893 ();
 b15zdnd11an1n64x5 FILLER_346_957 ();
 b15zdnd11an1n64x5 FILLER_346_1021 ();
 b15zdnd11an1n64x5 FILLER_346_1085 ();
 b15zdnd11an1n64x5 FILLER_346_1149 ();
 b15zdnd11an1n32x5 FILLER_346_1213 ();
 b15zdnd11an1n16x5 FILLER_346_1245 ();
 b15zdnd00an1n02x5 FILLER_346_1261 ();
 b15zdnd11an1n16x5 FILLER_346_1266 ();
 b15zdnd11an1n08x5 FILLER_346_1282 ();
 b15zdnd11an1n04x5 FILLER_346_1290 ();
 b15zdnd00an1n02x5 FILLER_346_1294 ();
 b15zdnd00an1n01x5 FILLER_346_1296 ();
 b15zdnd11an1n32x5 FILLER_346_1302 ();
 b15zdnd11an1n16x5 FILLER_346_1334 ();
 b15zdnd00an1n02x5 FILLER_346_1350 ();
 b15zdnd11an1n04x5 FILLER_346_1370 ();
 b15zdnd11an1n64x5 FILLER_346_1389 ();
 b15zdnd11an1n64x5 FILLER_346_1453 ();
 b15zdnd11an1n64x5 FILLER_346_1517 ();
 b15zdnd00an1n02x5 FILLER_346_1581 ();
 b15zdnd11an1n64x5 FILLER_346_1608 ();
 b15zdnd11an1n64x5 FILLER_346_1672 ();
 b15zdnd11an1n32x5 FILLER_346_1736 ();
 b15zdnd11an1n16x5 FILLER_346_1768 ();
 b15zdnd11an1n08x5 FILLER_346_1784 ();
 b15zdnd11an1n04x5 FILLER_346_1792 ();
 b15zdnd00an1n01x5 FILLER_346_1796 ();
 b15zdnd11an1n64x5 FILLER_346_1839 ();
 b15zdnd11an1n64x5 FILLER_346_1903 ();
 b15zdnd11an1n64x5 FILLER_346_1967 ();
 b15zdnd11an1n64x5 FILLER_346_2031 ();
 b15zdnd11an1n32x5 FILLER_346_2095 ();
 b15zdnd11an1n16x5 FILLER_346_2127 ();
 b15zdnd11an1n08x5 FILLER_346_2143 ();
 b15zdnd00an1n02x5 FILLER_346_2151 ();
 b15zdnd00an1n01x5 FILLER_346_2153 ();
 b15zdnd11an1n64x5 FILLER_346_2162 ();
 b15zdnd11an1n32x5 FILLER_346_2226 ();
 b15zdnd11an1n16x5 FILLER_346_2258 ();
 b15zdnd00an1n02x5 FILLER_346_2274 ();
 b15zdnd11an1n64x5 FILLER_347_0 ();
 b15zdnd11an1n64x5 FILLER_347_64 ();
 b15zdnd11an1n64x5 FILLER_347_128 ();
 b15zdnd11an1n64x5 FILLER_347_192 ();
 b15zdnd11an1n32x5 FILLER_347_256 ();
 b15zdnd11an1n16x5 FILLER_347_288 ();
 b15zdnd11an1n08x5 FILLER_347_304 ();
 b15zdnd11an1n16x5 FILLER_347_327 ();
 b15zdnd00an1n01x5 FILLER_347_343 ();
 b15zdnd11an1n64x5 FILLER_347_347 ();
 b15zdnd11an1n64x5 FILLER_347_411 ();
 b15zdnd11an1n64x5 FILLER_347_475 ();
 b15zdnd11an1n64x5 FILLER_347_539 ();
 b15zdnd11an1n08x5 FILLER_347_603 ();
 b15zdnd00an1n02x5 FILLER_347_611 ();
 b15zdnd00an1n01x5 FILLER_347_613 ();
 b15zdnd11an1n64x5 FILLER_347_618 ();
 b15zdnd11an1n32x5 FILLER_347_682 ();
 b15zdnd00an1n02x5 FILLER_347_714 ();
 b15zdnd00an1n01x5 FILLER_347_716 ();
 b15zdnd11an1n04x5 FILLER_347_720 ();
 b15zdnd11an1n04x5 FILLER_347_727 ();
 b15zdnd11an1n04x5 FILLER_347_734 ();
 b15zdnd11an1n04x5 FILLER_347_745 ();
 b15zdnd00an1n01x5 FILLER_347_749 ();
 b15zdnd11an1n16x5 FILLER_347_792 ();
 b15zdnd11an1n04x5 FILLER_347_808 ();
 b15zdnd00an1n02x5 FILLER_347_812 ();
 b15zdnd00an1n01x5 FILLER_347_814 ();
 b15zdnd11an1n64x5 FILLER_347_818 ();
 b15zdnd11an1n64x5 FILLER_347_882 ();
 b15zdnd11an1n64x5 FILLER_347_946 ();
 b15zdnd11an1n64x5 FILLER_347_1010 ();
 b15zdnd11an1n64x5 FILLER_347_1074 ();
 b15zdnd11an1n64x5 FILLER_347_1138 ();
 b15zdnd11an1n64x5 FILLER_347_1202 ();
 b15zdnd11an1n64x5 FILLER_347_1266 ();
 b15zdnd11an1n32x5 FILLER_347_1330 ();
 b15zdnd11an1n16x5 FILLER_347_1362 ();
 b15zdnd11an1n04x5 FILLER_347_1378 ();
 b15zdnd00an1n01x5 FILLER_347_1382 ();
 b15zdnd11an1n64x5 FILLER_347_1398 ();
 b15zdnd11an1n64x5 FILLER_347_1462 ();
 b15zdnd11an1n64x5 FILLER_347_1526 ();
 b15zdnd11an1n64x5 FILLER_347_1590 ();
 b15zdnd11an1n64x5 FILLER_347_1654 ();
 b15zdnd11an1n64x5 FILLER_347_1718 ();
 b15zdnd11an1n04x5 FILLER_347_1782 ();
 b15zdnd00an1n02x5 FILLER_347_1786 ();
 b15zdnd00an1n01x5 FILLER_347_1788 ();
 b15zdnd11an1n04x5 FILLER_347_1792 ();
 b15zdnd11an1n04x5 FILLER_347_1803 ();
 b15zdnd00an1n01x5 FILLER_347_1807 ();
 b15zdnd11an1n64x5 FILLER_347_1850 ();
 b15zdnd11an1n64x5 FILLER_347_1914 ();
 b15zdnd11an1n64x5 FILLER_347_1978 ();
 b15zdnd11an1n64x5 FILLER_347_2042 ();
 b15zdnd11an1n64x5 FILLER_347_2106 ();
 b15zdnd11an1n64x5 FILLER_347_2170 ();
 b15zdnd11an1n32x5 FILLER_347_2234 ();
 b15zdnd11an1n16x5 FILLER_347_2266 ();
 b15zdnd00an1n02x5 FILLER_347_2282 ();
 b15zdnd11an1n64x5 FILLER_348_8 ();
 b15zdnd11an1n64x5 FILLER_348_72 ();
 b15zdnd11an1n64x5 FILLER_348_136 ();
 b15zdnd11an1n64x5 FILLER_348_200 ();
 b15zdnd11an1n32x5 FILLER_348_264 ();
 b15zdnd11an1n16x5 FILLER_348_296 ();
 b15zdnd11an1n04x5 FILLER_348_312 ();
 b15zdnd00an1n02x5 FILLER_348_316 ();
 b15zdnd11an1n64x5 FILLER_348_360 ();
 b15zdnd11an1n64x5 FILLER_348_424 ();
 b15zdnd11an1n64x5 FILLER_348_488 ();
 b15zdnd11an1n64x5 FILLER_348_552 ();
 b15zdnd11an1n64x5 FILLER_348_616 ();
 b15zdnd11an1n32x5 FILLER_348_680 ();
 b15zdnd11an1n04x5 FILLER_348_712 ();
 b15zdnd00an1n02x5 FILLER_348_716 ();
 b15zdnd11an1n08x5 FILLER_348_726 ();
 b15zdnd11an1n04x5 FILLER_348_734 ();
 b15zdnd00an1n02x5 FILLER_348_738 ();
 b15zdnd00an1n01x5 FILLER_348_740 ();
 b15zdnd11an1n64x5 FILLER_348_783 ();
 b15zdnd11an1n64x5 FILLER_348_847 ();
 b15zdnd11an1n64x5 FILLER_348_911 ();
 b15zdnd11an1n16x5 FILLER_348_975 ();
 b15zdnd11an1n08x5 FILLER_348_991 ();
 b15zdnd00an1n02x5 FILLER_348_999 ();
 b15zdnd11an1n64x5 FILLER_348_1004 ();
 b15zdnd11an1n64x5 FILLER_348_1068 ();
 b15zdnd11an1n64x5 FILLER_348_1132 ();
 b15zdnd11an1n64x5 FILLER_348_1196 ();
 b15zdnd11an1n64x5 FILLER_348_1260 ();
 b15zdnd11an1n64x5 FILLER_348_1324 ();
 b15zdnd11an1n64x5 FILLER_348_1388 ();
 b15zdnd11an1n16x5 FILLER_348_1452 ();
 b15zdnd00an1n02x5 FILLER_348_1468 ();
 b15zdnd00an1n01x5 FILLER_348_1470 ();
 b15zdnd11an1n04x5 FILLER_348_1477 ();
 b15zdnd11an1n64x5 FILLER_348_1487 ();
 b15zdnd11an1n32x5 FILLER_348_1551 ();
 b15zdnd11an1n16x5 FILLER_348_1583 ();
 b15zdnd00an1n02x5 FILLER_348_1599 ();
 b15zdnd00an1n01x5 FILLER_348_1601 ();
 b15zdnd11an1n64x5 FILLER_348_1605 ();
 b15zdnd11an1n04x5 FILLER_348_1669 ();
 b15zdnd00an1n02x5 FILLER_348_1673 ();
 b15zdnd00an1n01x5 FILLER_348_1675 ();
 b15zdnd11an1n04x5 FILLER_348_1679 ();
 b15zdnd11an1n64x5 FILLER_348_1686 ();
 b15zdnd11an1n32x5 FILLER_348_1750 ();
 b15zdnd11an1n64x5 FILLER_348_1824 ();
 b15zdnd11an1n64x5 FILLER_348_1888 ();
 b15zdnd11an1n64x5 FILLER_348_1952 ();
 b15zdnd11an1n64x5 FILLER_348_2016 ();
 b15zdnd11an1n64x5 FILLER_348_2080 ();
 b15zdnd11an1n08x5 FILLER_348_2144 ();
 b15zdnd00an1n02x5 FILLER_348_2152 ();
 b15zdnd11an1n64x5 FILLER_348_2162 ();
 b15zdnd11an1n32x5 FILLER_348_2226 ();
 b15zdnd11an1n16x5 FILLER_348_2258 ();
 b15zdnd00an1n02x5 FILLER_348_2274 ();
 b15zdnd11an1n64x5 FILLER_349_0 ();
 b15zdnd11an1n64x5 FILLER_349_64 ();
 b15zdnd11an1n64x5 FILLER_349_128 ();
 b15zdnd11an1n64x5 FILLER_349_192 ();
 b15zdnd11an1n64x5 FILLER_349_256 ();
 b15zdnd11an1n16x5 FILLER_349_320 ();
 b15zdnd11an1n08x5 FILLER_349_336 ();
 b15zdnd11an1n16x5 FILLER_349_347 ();
 b15zdnd11an1n08x5 FILLER_349_363 ();
 b15zdnd11an1n04x5 FILLER_349_371 ();
 b15zdnd11an1n64x5 FILLER_349_417 ();
 b15zdnd11an1n64x5 FILLER_349_481 ();
 b15zdnd11an1n32x5 FILLER_349_545 ();
 b15zdnd11an1n16x5 FILLER_349_577 ();
 b15zdnd11an1n08x5 FILLER_349_593 ();
 b15zdnd11an1n04x5 FILLER_349_601 ();
 b15zdnd00an1n02x5 FILLER_349_605 ();
 b15zdnd11an1n04x5 FILLER_349_613 ();
 b15zdnd11an1n64x5 FILLER_349_621 ();
 b15zdnd11an1n32x5 FILLER_349_685 ();
 b15zdnd11an1n16x5 FILLER_349_717 ();
 b15zdnd11an1n08x5 FILLER_349_733 ();
 b15zdnd00an1n01x5 FILLER_349_741 ();
 b15zdnd11an1n04x5 FILLER_349_745 ();
 b15zdnd11an1n64x5 FILLER_349_754 ();
 b15zdnd11an1n64x5 FILLER_349_818 ();
 b15zdnd11an1n16x5 FILLER_349_882 ();
 b15zdnd11an1n04x5 FILLER_349_898 ();
 b15zdnd11an1n16x5 FILLER_349_920 ();
 b15zdnd11an1n08x5 FILLER_349_936 ();
 b15zdnd00an1n02x5 FILLER_349_944 ();
 b15zdnd00an1n01x5 FILLER_349_946 ();
 b15zdnd11an1n16x5 FILLER_349_954 ();
 b15zdnd11an1n04x5 FILLER_349_970 ();
 b15zdnd11an1n64x5 FILLER_349_1026 ();
 b15zdnd11an1n04x5 FILLER_349_1090 ();
 b15zdnd11an1n16x5 FILLER_349_1102 ();
 b15zdnd00an1n01x5 FILLER_349_1118 ();
 b15zdnd11an1n64x5 FILLER_349_1122 ();
 b15zdnd11an1n64x5 FILLER_349_1186 ();
 b15zdnd11an1n64x5 FILLER_349_1250 ();
 b15zdnd11an1n32x5 FILLER_349_1314 ();
 b15zdnd00an1n02x5 FILLER_349_1346 ();
 b15zdnd11an1n04x5 FILLER_349_1363 ();
 b15zdnd11an1n64x5 FILLER_349_1370 ();
 b15zdnd11an1n32x5 FILLER_349_1434 ();
 b15zdnd11an1n16x5 FILLER_349_1466 ();
 b15zdnd11an1n04x5 FILLER_349_1482 ();
 b15zdnd11an1n64x5 FILLER_349_1503 ();
 b15zdnd11an1n16x5 FILLER_349_1567 ();
 b15zdnd11an1n04x5 FILLER_349_1583 ();
 b15zdnd11an1n04x5 FILLER_349_1590 ();
 b15zdnd11an1n08x5 FILLER_349_1597 ();
 b15zdnd00an1n01x5 FILLER_349_1605 ();
 b15zdnd11an1n08x5 FILLER_349_1648 ();
 b15zdnd00an1n02x5 FILLER_349_1656 ();
 b15zdnd11an1n32x5 FILLER_349_1710 ();
 b15zdnd00an1n01x5 FILLER_349_1742 ();
 b15zdnd11an1n08x5 FILLER_349_1785 ();
 b15zdnd11an1n64x5 FILLER_349_1797 ();
 b15zdnd11an1n64x5 FILLER_349_1861 ();
 b15zdnd11an1n64x5 FILLER_349_1925 ();
 b15zdnd11an1n64x5 FILLER_349_1989 ();
 b15zdnd11an1n64x5 FILLER_349_2053 ();
 b15zdnd11an1n64x5 FILLER_349_2117 ();
 b15zdnd11an1n64x5 FILLER_349_2181 ();
 b15zdnd11an1n32x5 FILLER_349_2245 ();
 b15zdnd11an1n04x5 FILLER_349_2277 ();
 b15zdnd00an1n02x5 FILLER_349_2281 ();
 b15zdnd00an1n01x5 FILLER_349_2283 ();
 b15zdnd11an1n64x5 FILLER_350_8 ();
 b15zdnd11an1n64x5 FILLER_350_72 ();
 b15zdnd11an1n64x5 FILLER_350_136 ();
 b15zdnd11an1n64x5 FILLER_350_200 ();
 b15zdnd11an1n64x5 FILLER_350_264 ();
 b15zdnd11an1n32x5 FILLER_350_328 ();
 b15zdnd11an1n16x5 FILLER_350_360 ();
 b15zdnd11an1n08x5 FILLER_350_376 ();
 b15zdnd11an1n04x5 FILLER_350_384 ();
 b15zdnd11an1n64x5 FILLER_350_391 ();
 b15zdnd11an1n64x5 FILLER_350_455 ();
 b15zdnd11an1n64x5 FILLER_350_519 ();
 b15zdnd11an1n16x5 FILLER_350_583 ();
 b15zdnd11an1n08x5 FILLER_350_599 ();
 b15zdnd00an1n01x5 FILLER_350_607 ();
 b15zdnd11an1n08x5 FILLER_350_612 ();
 b15zdnd11an1n04x5 FILLER_350_620 ();
 b15zdnd11an1n16x5 FILLER_350_627 ();
 b15zdnd11an1n08x5 FILLER_350_643 ();
 b15zdnd11an1n04x5 FILLER_350_651 ();
 b15zdnd00an1n01x5 FILLER_350_655 ();
 b15zdnd11an1n32x5 FILLER_350_676 ();
 b15zdnd11an1n08x5 FILLER_350_708 ();
 b15zdnd00an1n02x5 FILLER_350_716 ();
 b15zdnd11an1n16x5 FILLER_350_726 ();
 b15zdnd11an1n04x5 FILLER_350_742 ();
 b15zdnd00an1n02x5 FILLER_350_746 ();
 b15zdnd00an1n01x5 FILLER_350_748 ();
 b15zdnd11an1n64x5 FILLER_350_755 ();
 b15zdnd11an1n64x5 FILLER_350_819 ();
 b15zdnd11an1n08x5 FILLER_350_883 ();
 b15zdnd00an1n02x5 FILLER_350_891 ();
 b15zdnd00an1n01x5 FILLER_350_893 ();
 b15zdnd11an1n32x5 FILLER_350_897 ();
 b15zdnd11an1n08x5 FILLER_350_929 ();
 b15zdnd00an1n02x5 FILLER_350_937 ();
 b15zdnd00an1n01x5 FILLER_350_939 ();
 b15zdnd11an1n08x5 FILLER_350_982 ();
 b15zdnd00an1n02x5 FILLER_350_990 ();
 b15zdnd11an1n04x5 FILLER_350_995 ();
 b15zdnd11an1n64x5 FILLER_350_1002 ();
 b15zdnd11an1n16x5 FILLER_350_1066 ();
 b15zdnd11an1n08x5 FILLER_350_1082 ();
 b15zdnd11an1n04x5 FILLER_350_1090 ();
 b15zdnd00an1n01x5 FILLER_350_1094 ();
 b15zdnd11an1n64x5 FILLER_350_1137 ();
 b15zdnd11an1n64x5 FILLER_350_1201 ();
 b15zdnd11an1n64x5 FILLER_350_1265 ();
 b15zdnd11an1n64x5 FILLER_350_1329 ();
 b15zdnd11an1n64x5 FILLER_350_1393 ();
 b15zdnd11an1n16x5 FILLER_350_1457 ();
 b15zdnd11an1n08x5 FILLER_350_1473 ();
 b15zdnd00an1n02x5 FILLER_350_1481 ();
 b15zdnd00an1n01x5 FILLER_350_1483 ();
 b15zdnd11an1n32x5 FILLER_350_1536 ();
 b15zdnd11an1n04x5 FILLER_350_1568 ();
 b15zdnd11an1n32x5 FILLER_350_1624 ();
 b15zdnd11an1n16x5 FILLER_350_1656 ();
 b15zdnd11an1n08x5 FILLER_350_1672 ();
 b15zdnd00an1n02x5 FILLER_350_1680 ();
 b15zdnd00an1n01x5 FILLER_350_1682 ();
 b15zdnd11an1n32x5 FILLER_350_1686 ();
 b15zdnd11an1n16x5 FILLER_350_1718 ();
 b15zdnd11an1n04x5 FILLER_350_1776 ();
 b15zdnd11an1n08x5 FILLER_350_1785 ();
 b15zdnd00an1n01x5 FILLER_350_1793 ();
 b15zdnd11an1n64x5 FILLER_350_1799 ();
 b15zdnd11an1n64x5 FILLER_350_1863 ();
 b15zdnd11an1n32x5 FILLER_350_1927 ();
 b15zdnd00an1n01x5 FILLER_350_1959 ();
 b15zdnd11an1n16x5 FILLER_350_1964 ();
 b15zdnd11an1n08x5 FILLER_350_1980 ();
 b15zdnd11an1n04x5 FILLER_350_1988 ();
 b15zdnd00an1n02x5 FILLER_350_1992 ();
 b15zdnd11an1n64x5 FILLER_350_2036 ();
 b15zdnd11an1n32x5 FILLER_350_2100 ();
 b15zdnd11an1n16x5 FILLER_350_2132 ();
 b15zdnd11an1n04x5 FILLER_350_2148 ();
 b15zdnd00an1n02x5 FILLER_350_2152 ();
 b15zdnd11an1n64x5 FILLER_350_2162 ();
 b15zdnd11an1n32x5 FILLER_350_2226 ();
 b15zdnd11an1n16x5 FILLER_350_2258 ();
 b15zdnd00an1n02x5 FILLER_350_2274 ();
 b15zdnd11an1n64x5 FILLER_351_0 ();
 b15zdnd11an1n64x5 FILLER_351_64 ();
 b15zdnd11an1n64x5 FILLER_351_128 ();
 b15zdnd11an1n32x5 FILLER_351_192 ();
 b15zdnd11an1n16x5 FILLER_351_224 ();
 b15zdnd11an1n04x5 FILLER_351_240 ();
 b15zdnd11an1n64x5 FILLER_351_253 ();
 b15zdnd11an1n32x5 FILLER_351_317 ();
 b15zdnd11an1n08x5 FILLER_351_349 ();
 b15zdnd11an1n04x5 FILLER_351_357 ();
 b15zdnd11an1n64x5 FILLER_351_413 ();
 b15zdnd11an1n64x5 FILLER_351_477 ();
 b15zdnd11an1n32x5 FILLER_351_541 ();
 b15zdnd11an1n16x5 FILLER_351_573 ();
 b15zdnd11an1n08x5 FILLER_351_589 ();
 b15zdnd11an1n04x5 FILLER_351_597 ();
 b15zdnd11an1n64x5 FILLER_351_653 ();
 b15zdnd11an1n16x5 FILLER_351_717 ();
 b15zdnd00an1n02x5 FILLER_351_733 ();
 b15zdnd00an1n01x5 FILLER_351_735 ();
 b15zdnd11an1n04x5 FILLER_351_741 ();
 b15zdnd11an1n64x5 FILLER_351_755 ();
 b15zdnd11an1n32x5 FILLER_351_819 ();
 b15zdnd11an1n08x5 FILLER_351_851 ();
 b15zdnd00an1n02x5 FILLER_351_859 ();
 b15zdnd11an1n04x5 FILLER_351_867 ();
 b15zdnd11an1n08x5 FILLER_351_923 ();
 b15zdnd11an1n04x5 FILLER_351_931 ();
 b15zdnd11an1n32x5 FILLER_351_977 ();
 b15zdnd00an1n01x5 FILLER_351_1009 ();
 b15zdnd11an1n64x5 FILLER_351_1018 ();
 b15zdnd11an1n08x5 FILLER_351_1082 ();
 b15zdnd00an1n02x5 FILLER_351_1090 ();
 b15zdnd11an1n32x5 FILLER_351_1144 ();
 b15zdnd11an1n04x5 FILLER_351_1176 ();
 b15zdnd00an1n01x5 FILLER_351_1180 ();
 b15zdnd11an1n04x5 FILLER_351_1223 ();
 b15zdnd11an1n64x5 FILLER_351_1269 ();
 b15zdnd11an1n32x5 FILLER_351_1333 ();
 b15zdnd11an1n16x5 FILLER_351_1365 ();
 b15zdnd00an1n02x5 FILLER_351_1381 ();
 b15zdnd11an1n64x5 FILLER_351_1401 ();
 b15zdnd11an1n32x5 FILLER_351_1465 ();
 b15zdnd11an1n04x5 FILLER_351_1497 ();
 b15zdnd00an1n01x5 FILLER_351_1501 ();
 b15zdnd11an1n04x5 FILLER_351_1505 ();
 b15zdnd11an1n64x5 FILLER_351_1512 ();
 b15zdnd11an1n64x5 FILLER_351_1576 ();
 b15zdnd11an1n64x5 FILLER_351_1640 ();
 b15zdnd11an1n64x5 FILLER_351_1704 ();
 b15zdnd11an1n04x5 FILLER_351_1768 ();
 b15zdnd11an1n08x5 FILLER_351_1781 ();
 b15zdnd11an1n04x5 FILLER_351_1789 ();
 b15zdnd00an1n01x5 FILLER_351_1793 ();
 b15zdnd11an1n64x5 FILLER_351_1801 ();
 b15zdnd11an1n64x5 FILLER_351_1865 ();
 b15zdnd11an1n16x5 FILLER_351_1929 ();
 b15zdnd11an1n08x5 FILLER_351_1948 ();
 b15zdnd11an1n04x5 FILLER_351_1956 ();
 b15zdnd11an1n08x5 FILLER_351_1966 ();
 b15zdnd00an1n01x5 FILLER_351_1974 ();
 b15zdnd11an1n64x5 FILLER_351_2017 ();
 b15zdnd11an1n64x5 FILLER_351_2081 ();
 b15zdnd11an1n64x5 FILLER_351_2145 ();
 b15zdnd11an1n64x5 FILLER_351_2209 ();
 b15zdnd11an1n08x5 FILLER_351_2273 ();
 b15zdnd00an1n02x5 FILLER_351_2281 ();
 b15zdnd00an1n01x5 FILLER_351_2283 ();
 b15zdnd11an1n64x5 FILLER_352_8 ();
 b15zdnd11an1n64x5 FILLER_352_72 ();
 b15zdnd11an1n64x5 FILLER_352_136 ();
 b15zdnd11an1n32x5 FILLER_352_200 ();
 b15zdnd11an1n16x5 FILLER_352_232 ();
 b15zdnd11an1n04x5 FILLER_352_248 ();
 b15zdnd11an1n64x5 FILLER_352_255 ();
 b15zdnd11an1n64x5 FILLER_352_319 ();
 b15zdnd00an1n02x5 FILLER_352_383 ();
 b15zdnd00an1n01x5 FILLER_352_385 ();
 b15zdnd11an1n64x5 FILLER_352_389 ();
 b15zdnd11an1n64x5 FILLER_352_453 ();
 b15zdnd11an1n64x5 FILLER_352_517 ();
 b15zdnd11an1n32x5 FILLER_352_581 ();
 b15zdnd11an1n08x5 FILLER_352_613 ();
 b15zdnd00an1n02x5 FILLER_352_621 ();
 b15zdnd11an1n04x5 FILLER_352_626 ();
 b15zdnd11an1n64x5 FILLER_352_650 ();
 b15zdnd11an1n04x5 FILLER_352_714 ();
 b15zdnd11an1n16x5 FILLER_352_726 ();
 b15zdnd11an1n08x5 FILLER_352_742 ();
 b15zdnd11an1n64x5 FILLER_352_766 ();
 b15zdnd11an1n32x5 FILLER_352_830 ();
 b15zdnd11an1n08x5 FILLER_352_862 ();
 b15zdnd11an1n04x5 FILLER_352_870 ();
 b15zdnd11an1n64x5 FILLER_352_916 ();
 b15zdnd11an1n64x5 FILLER_352_980 ();
 b15zdnd11an1n32x5 FILLER_352_1044 ();
 b15zdnd11an1n16x5 FILLER_352_1076 ();
 b15zdnd11an1n64x5 FILLER_352_1134 ();
 b15zdnd11an1n64x5 FILLER_352_1198 ();
 b15zdnd11an1n64x5 FILLER_352_1262 ();
 b15zdnd11an1n32x5 FILLER_352_1326 ();
 b15zdnd11an1n08x5 FILLER_352_1358 ();
 b15zdnd11an1n04x5 FILLER_352_1366 ();
 b15zdnd11an1n64x5 FILLER_352_1410 ();
 b15zdnd11an1n32x5 FILLER_352_1474 ();
 b15zdnd11an1n04x5 FILLER_352_1506 ();
 b15zdnd11an1n16x5 FILLER_352_1513 ();
 b15zdnd11an1n08x5 FILLER_352_1529 ();
 b15zdnd00an1n02x5 FILLER_352_1537 ();
 b15zdnd00an1n01x5 FILLER_352_1539 ();
 b15zdnd11an1n64x5 FILLER_352_1547 ();
 b15zdnd11an1n64x5 FILLER_352_1611 ();
 b15zdnd11an1n64x5 FILLER_352_1675 ();
 b15zdnd11an1n64x5 FILLER_352_1739 ();
 b15zdnd11an1n64x5 FILLER_352_1803 ();
 b15zdnd11an1n64x5 FILLER_352_1867 ();
 b15zdnd11an1n04x5 FILLER_352_1931 ();
 b15zdnd00an1n02x5 FILLER_352_1935 ();
 b15zdnd11an1n04x5 FILLER_352_1942 ();
 b15zdnd11an1n08x5 FILLER_352_1951 ();
 b15zdnd11an1n04x5 FILLER_352_1969 ();
 b15zdnd00an1n02x5 FILLER_352_1973 ();
 b15zdnd00an1n01x5 FILLER_352_1975 ();
 b15zdnd11an1n64x5 FILLER_352_2028 ();
 b15zdnd11an1n32x5 FILLER_352_2092 ();
 b15zdnd11an1n16x5 FILLER_352_2124 ();
 b15zdnd11an1n08x5 FILLER_352_2140 ();
 b15zdnd11an1n04x5 FILLER_352_2148 ();
 b15zdnd00an1n02x5 FILLER_352_2152 ();
 b15zdnd11an1n64x5 FILLER_352_2162 ();
 b15zdnd11an1n32x5 FILLER_352_2226 ();
 b15zdnd11an1n16x5 FILLER_352_2258 ();
 b15zdnd00an1n02x5 FILLER_352_2274 ();
 b15zdnd11an1n64x5 FILLER_353_0 ();
 b15zdnd11an1n64x5 FILLER_353_64 ();
 b15zdnd11an1n64x5 FILLER_353_128 ();
 b15zdnd11an1n32x5 FILLER_353_192 ();
 b15zdnd00an1n01x5 FILLER_353_224 ();
 b15zdnd11an1n64x5 FILLER_353_277 ();
 b15zdnd11an1n32x5 FILLER_353_341 ();
 b15zdnd11an1n08x5 FILLER_353_373 ();
 b15zdnd00an1n02x5 FILLER_353_381 ();
 b15zdnd00an1n01x5 FILLER_353_383 ();
 b15zdnd11an1n64x5 FILLER_353_387 ();
 b15zdnd11an1n64x5 FILLER_353_451 ();
 b15zdnd11an1n64x5 FILLER_353_515 ();
 b15zdnd11an1n32x5 FILLER_353_579 ();
 b15zdnd11an1n16x5 FILLER_353_611 ();
 b15zdnd11an1n64x5 FILLER_353_630 ();
 b15zdnd11an1n32x5 FILLER_353_694 ();
 b15zdnd11an1n16x5 FILLER_353_726 ();
 b15zdnd11an1n08x5 FILLER_353_742 ();
 b15zdnd00an1n01x5 FILLER_353_750 ();
 b15zdnd11an1n64x5 FILLER_353_764 ();
 b15zdnd11an1n32x5 FILLER_353_828 ();
 b15zdnd11an1n08x5 FILLER_353_860 ();
 b15zdnd11an1n04x5 FILLER_353_868 ();
 b15zdnd00an1n01x5 FILLER_353_872 ();
 b15zdnd11an1n08x5 FILLER_353_880 ();
 b15zdnd00an1n02x5 FILLER_353_888 ();
 b15zdnd00an1n01x5 FILLER_353_890 ();
 b15zdnd11an1n04x5 FILLER_353_894 ();
 b15zdnd11an1n64x5 FILLER_353_901 ();
 b15zdnd11an1n64x5 FILLER_353_965 ();
 b15zdnd11an1n32x5 FILLER_353_1029 ();
 b15zdnd11an1n08x5 FILLER_353_1061 ();
 b15zdnd11an1n04x5 FILLER_353_1121 ();
 b15zdnd11an1n16x5 FILLER_353_1128 ();
 b15zdnd11an1n64x5 FILLER_353_1186 ();
 b15zdnd11an1n64x5 FILLER_353_1250 ();
 b15zdnd11an1n08x5 FILLER_353_1314 ();
 b15zdnd11an1n04x5 FILLER_353_1322 ();
 b15zdnd11an1n64x5 FILLER_353_1336 ();
 b15zdnd11an1n64x5 FILLER_353_1400 ();
 b15zdnd11an1n16x5 FILLER_353_1464 ();
 b15zdnd11an1n08x5 FILLER_353_1480 ();
 b15zdnd11an1n04x5 FILLER_353_1488 ();
 b15zdnd00an1n01x5 FILLER_353_1492 ();
 b15zdnd11an1n32x5 FILLER_353_1524 ();
 b15zdnd11an1n16x5 FILLER_353_1556 ();
 b15zdnd11an1n08x5 FILLER_353_1572 ();
 b15zdnd00an1n02x5 FILLER_353_1580 ();
 b15zdnd00an1n01x5 FILLER_353_1582 ();
 b15zdnd11an1n64x5 FILLER_353_1608 ();
 b15zdnd11an1n64x5 FILLER_353_1672 ();
 b15zdnd11an1n64x5 FILLER_353_1736 ();
 b15zdnd11an1n64x5 FILLER_353_1800 ();
 b15zdnd11an1n64x5 FILLER_353_1864 ();
 b15zdnd00an1n02x5 FILLER_353_1928 ();
 b15zdnd00an1n01x5 FILLER_353_1930 ();
 b15zdnd11an1n04x5 FILLER_353_1937 ();
 b15zdnd11an1n04x5 FILLER_353_1945 ();
 b15zdnd11an1n08x5 FILLER_353_1956 ();
 b15zdnd11an1n04x5 FILLER_353_2006 ();
 b15zdnd11an1n04x5 FILLER_353_2013 ();
 b15zdnd11an1n64x5 FILLER_353_2020 ();
 b15zdnd11an1n64x5 FILLER_353_2084 ();
 b15zdnd11an1n64x5 FILLER_353_2148 ();
 b15zdnd11an1n64x5 FILLER_353_2212 ();
 b15zdnd11an1n08x5 FILLER_353_2276 ();
 b15zdnd11an1n64x5 FILLER_354_8 ();
 b15zdnd11an1n64x5 FILLER_354_72 ();
 b15zdnd11an1n64x5 FILLER_354_136 ();
 b15zdnd11an1n32x5 FILLER_354_200 ();
 b15zdnd11an1n08x5 FILLER_354_232 ();
 b15zdnd00an1n02x5 FILLER_354_240 ();
 b15zdnd00an1n01x5 FILLER_354_242 ();
 b15zdnd11an1n04x5 FILLER_354_246 ();
 b15zdnd11an1n64x5 FILLER_354_253 ();
 b15zdnd11an1n64x5 FILLER_354_317 ();
 b15zdnd11an1n64x5 FILLER_354_381 ();
 b15zdnd11an1n64x5 FILLER_354_445 ();
 b15zdnd11an1n08x5 FILLER_354_509 ();
 b15zdnd11an1n04x5 FILLER_354_517 ();
 b15zdnd11an1n64x5 FILLER_354_563 ();
 b15zdnd11an1n64x5 FILLER_354_627 ();
 b15zdnd11an1n16x5 FILLER_354_691 ();
 b15zdnd11an1n08x5 FILLER_354_707 ();
 b15zdnd00an1n02x5 FILLER_354_715 ();
 b15zdnd00an1n01x5 FILLER_354_717 ();
 b15zdnd11an1n64x5 FILLER_354_726 ();
 b15zdnd11an1n64x5 FILLER_354_790 ();
 b15zdnd11an1n64x5 FILLER_354_854 ();
 b15zdnd11an1n64x5 FILLER_354_918 ();
 b15zdnd11an1n64x5 FILLER_354_982 ();
 b15zdnd11an1n32x5 FILLER_354_1046 ();
 b15zdnd11an1n08x5 FILLER_354_1078 ();
 b15zdnd00an1n01x5 FILLER_354_1086 ();
 b15zdnd11an1n04x5 FILLER_354_1090 ();
 b15zdnd11an1n08x5 FILLER_354_1101 ();
 b15zdnd00an1n01x5 FILLER_354_1109 ();
 b15zdnd11an1n08x5 FILLER_354_1113 ();
 b15zdnd11an1n64x5 FILLER_354_1163 ();
 b15zdnd11an1n16x5 FILLER_354_1227 ();
 b15zdnd11an1n08x5 FILLER_354_1243 ();
 b15zdnd00an1n01x5 FILLER_354_1251 ();
 b15zdnd11an1n64x5 FILLER_354_1263 ();
 b15zdnd11an1n64x5 FILLER_354_1334 ();
 b15zdnd11an1n64x5 FILLER_354_1398 ();
 b15zdnd11an1n64x5 FILLER_354_1462 ();
 b15zdnd11an1n64x5 FILLER_354_1526 ();
 b15zdnd11an1n64x5 FILLER_354_1590 ();
 b15zdnd11an1n64x5 FILLER_354_1654 ();
 b15zdnd11an1n32x5 FILLER_354_1718 ();
 b15zdnd11an1n16x5 FILLER_354_1750 ();
 b15zdnd11an1n04x5 FILLER_354_1766 ();
 b15zdnd00an1n01x5 FILLER_354_1770 ();
 b15zdnd11an1n64x5 FILLER_354_1776 ();
 b15zdnd11an1n64x5 FILLER_354_1840 ();
 b15zdnd11an1n16x5 FILLER_354_1904 ();
 b15zdnd00an1n02x5 FILLER_354_1920 ();
 b15zdnd00an1n01x5 FILLER_354_1922 ();
 b15zdnd11an1n04x5 FILLER_354_1933 ();
 b15zdnd11an1n08x5 FILLER_354_1944 ();
 b15zdnd11an1n04x5 FILLER_354_1994 ();
 b15zdnd11an1n64x5 FILLER_354_2001 ();
 b15zdnd11an1n64x5 FILLER_354_2065 ();
 b15zdnd11an1n16x5 FILLER_354_2129 ();
 b15zdnd11an1n08x5 FILLER_354_2145 ();
 b15zdnd00an1n01x5 FILLER_354_2153 ();
 b15zdnd11an1n64x5 FILLER_354_2162 ();
 b15zdnd11an1n32x5 FILLER_354_2226 ();
 b15zdnd11an1n16x5 FILLER_354_2258 ();
 b15zdnd00an1n02x5 FILLER_354_2274 ();
 b15zdnd11an1n64x5 FILLER_355_0 ();
 b15zdnd11an1n64x5 FILLER_355_64 ();
 b15zdnd11an1n64x5 FILLER_355_128 ();
 b15zdnd11an1n32x5 FILLER_355_192 ();
 b15zdnd11an1n16x5 FILLER_355_224 ();
 b15zdnd11an1n08x5 FILLER_355_240 ();
 b15zdnd00an1n01x5 FILLER_355_248 ();
 b15zdnd11an1n64x5 FILLER_355_291 ();
 b15zdnd11an1n64x5 FILLER_355_355 ();
 b15zdnd11an1n64x5 FILLER_355_419 ();
 b15zdnd11an1n64x5 FILLER_355_483 ();
 b15zdnd11an1n64x5 FILLER_355_547 ();
 b15zdnd11an1n64x5 FILLER_355_611 ();
 b15zdnd11an1n64x5 FILLER_355_675 ();
 b15zdnd11an1n64x5 FILLER_355_739 ();
 b15zdnd11an1n64x5 FILLER_355_803 ();
 b15zdnd11an1n64x5 FILLER_355_867 ();
 b15zdnd11an1n64x5 FILLER_355_931 ();
 b15zdnd11an1n64x5 FILLER_355_995 ();
 b15zdnd00an1n01x5 FILLER_355_1059 ();
 b15zdnd11an1n08x5 FILLER_355_1091 ();
 b15zdnd11an1n16x5 FILLER_355_1102 ();
 b15zdnd11an1n04x5 FILLER_355_1118 ();
 b15zdnd11an1n64x5 FILLER_355_1129 ();
 b15zdnd11an1n64x5 FILLER_355_1193 ();
 b15zdnd11an1n64x5 FILLER_355_1257 ();
 b15zdnd00an1n02x5 FILLER_355_1321 ();
 b15zdnd00an1n01x5 FILLER_355_1323 ();
 b15zdnd11an1n64x5 FILLER_355_1328 ();
 b15zdnd11an1n64x5 FILLER_355_1392 ();
 b15zdnd11an1n64x5 FILLER_355_1456 ();
 b15zdnd11an1n64x5 FILLER_355_1520 ();
 b15zdnd11an1n64x5 FILLER_355_1584 ();
 b15zdnd11an1n64x5 FILLER_355_1648 ();
 b15zdnd11an1n64x5 FILLER_355_1712 ();
 b15zdnd11an1n64x5 FILLER_355_1780 ();
 b15zdnd11an1n64x5 FILLER_355_1844 ();
 b15zdnd11an1n16x5 FILLER_355_1908 ();
 b15zdnd11an1n04x5 FILLER_355_1966 ();
 b15zdnd11an1n64x5 FILLER_355_1976 ();
 b15zdnd11an1n64x5 FILLER_355_2040 ();
 b15zdnd11an1n64x5 FILLER_355_2104 ();
 b15zdnd11an1n64x5 FILLER_355_2168 ();
 b15zdnd11an1n32x5 FILLER_355_2232 ();
 b15zdnd11an1n16x5 FILLER_355_2264 ();
 b15zdnd11an1n04x5 FILLER_355_2280 ();
 b15zdnd11an1n64x5 FILLER_356_8 ();
 b15zdnd11an1n64x5 FILLER_356_72 ();
 b15zdnd11an1n64x5 FILLER_356_136 ();
 b15zdnd11an1n32x5 FILLER_356_200 ();
 b15zdnd11an1n16x5 FILLER_356_232 ();
 b15zdnd00an1n02x5 FILLER_356_248 ();
 b15zdnd11an1n64x5 FILLER_356_255 ();
 b15zdnd11an1n64x5 FILLER_356_319 ();
 b15zdnd11an1n64x5 FILLER_356_383 ();
 b15zdnd11an1n64x5 FILLER_356_447 ();
 b15zdnd11an1n64x5 FILLER_356_511 ();
 b15zdnd11an1n64x5 FILLER_356_575 ();
 b15zdnd11an1n64x5 FILLER_356_639 ();
 b15zdnd11an1n08x5 FILLER_356_703 ();
 b15zdnd11an1n04x5 FILLER_356_711 ();
 b15zdnd00an1n02x5 FILLER_356_715 ();
 b15zdnd00an1n01x5 FILLER_356_717 ();
 b15zdnd11an1n64x5 FILLER_356_726 ();
 b15zdnd11an1n64x5 FILLER_356_790 ();
 b15zdnd11an1n64x5 FILLER_356_854 ();
 b15zdnd11an1n64x5 FILLER_356_918 ();
 b15zdnd11an1n64x5 FILLER_356_982 ();
 b15zdnd11an1n32x5 FILLER_356_1046 ();
 b15zdnd11an1n16x5 FILLER_356_1078 ();
 b15zdnd00an1n01x5 FILLER_356_1094 ();
 b15zdnd11an1n64x5 FILLER_356_1098 ();
 b15zdnd11an1n64x5 FILLER_356_1162 ();
 b15zdnd11an1n64x5 FILLER_356_1226 ();
 b15zdnd00an1n02x5 FILLER_356_1290 ();
 b15zdnd00an1n01x5 FILLER_356_1292 ();
 b15zdnd11an1n64x5 FILLER_356_1335 ();
 b15zdnd11an1n64x5 FILLER_356_1399 ();
 b15zdnd11an1n64x5 FILLER_356_1463 ();
 b15zdnd11an1n64x5 FILLER_356_1527 ();
 b15zdnd11an1n64x5 FILLER_356_1591 ();
 b15zdnd11an1n64x5 FILLER_356_1655 ();
 b15zdnd11an1n64x5 FILLER_356_1719 ();
 b15zdnd11an1n64x5 FILLER_356_1783 ();
 b15zdnd11an1n64x5 FILLER_356_1847 ();
 b15zdnd11an1n08x5 FILLER_356_1911 ();
 b15zdnd11an1n04x5 FILLER_356_1922 ();
 b15zdnd00an1n02x5 FILLER_356_1926 ();
 b15zdnd11an1n64x5 FILLER_356_1970 ();
 b15zdnd11an1n64x5 FILLER_356_2034 ();
 b15zdnd11an1n32x5 FILLER_356_2098 ();
 b15zdnd11an1n16x5 FILLER_356_2130 ();
 b15zdnd11an1n08x5 FILLER_356_2146 ();
 b15zdnd11an1n64x5 FILLER_356_2162 ();
 b15zdnd11an1n32x5 FILLER_356_2226 ();
 b15zdnd11an1n16x5 FILLER_356_2258 ();
 b15zdnd00an1n02x5 FILLER_356_2274 ();
 b15zdnd11an1n64x5 FILLER_357_0 ();
 b15zdnd11an1n64x5 FILLER_357_64 ();
 b15zdnd11an1n64x5 FILLER_357_128 ();
 b15zdnd11an1n32x5 FILLER_357_192 ();
 b15zdnd11an1n16x5 FILLER_357_224 ();
 b15zdnd11an1n08x5 FILLER_357_240 ();
 b15zdnd11an1n04x5 FILLER_357_248 ();
 b15zdnd00an1n02x5 FILLER_357_252 ();
 b15zdnd00an1n01x5 FILLER_357_254 ();
 b15zdnd11an1n64x5 FILLER_357_259 ();
 b15zdnd11an1n64x5 FILLER_357_323 ();
 b15zdnd11an1n64x5 FILLER_357_387 ();
 b15zdnd11an1n64x5 FILLER_357_451 ();
 b15zdnd11an1n64x5 FILLER_357_515 ();
 b15zdnd11an1n64x5 FILLER_357_579 ();
 b15zdnd11an1n64x5 FILLER_357_643 ();
 b15zdnd11an1n64x5 FILLER_357_707 ();
 b15zdnd11an1n64x5 FILLER_357_771 ();
 b15zdnd11an1n08x5 FILLER_357_835 ();
 b15zdnd11an1n04x5 FILLER_357_843 ();
 b15zdnd00an1n02x5 FILLER_357_847 ();
 b15zdnd00an1n01x5 FILLER_357_849 ();
 b15zdnd11an1n64x5 FILLER_357_892 ();
 b15zdnd11an1n64x5 FILLER_357_956 ();
 b15zdnd11an1n64x5 FILLER_357_1020 ();
 b15zdnd11an1n64x5 FILLER_357_1084 ();
 b15zdnd11an1n64x5 FILLER_357_1148 ();
 b15zdnd11an1n64x5 FILLER_357_1212 ();
 b15zdnd11an1n32x5 FILLER_357_1276 ();
 b15zdnd11an1n16x5 FILLER_357_1308 ();
 b15zdnd11an1n08x5 FILLER_357_1324 ();
 b15zdnd11an1n04x5 FILLER_357_1332 ();
 b15zdnd00an1n01x5 FILLER_357_1336 ();
 b15zdnd11an1n04x5 FILLER_357_1379 ();
 b15zdnd11an1n64x5 FILLER_357_1386 ();
 b15zdnd11an1n64x5 FILLER_357_1450 ();
 b15zdnd11an1n64x5 FILLER_357_1514 ();
 b15zdnd11an1n64x5 FILLER_357_1578 ();
 b15zdnd11an1n64x5 FILLER_357_1642 ();
 b15zdnd11an1n64x5 FILLER_357_1706 ();
 b15zdnd11an1n64x5 FILLER_357_1770 ();
 b15zdnd11an1n64x5 FILLER_357_1834 ();
 b15zdnd11an1n16x5 FILLER_357_1898 ();
 b15zdnd11an1n64x5 FILLER_357_1956 ();
 b15zdnd11an1n64x5 FILLER_357_2020 ();
 b15zdnd11an1n64x5 FILLER_357_2084 ();
 b15zdnd11an1n64x5 FILLER_357_2148 ();
 b15zdnd11an1n64x5 FILLER_357_2212 ();
 b15zdnd11an1n08x5 FILLER_357_2276 ();
 b15zdnd11an1n64x5 FILLER_358_8 ();
 b15zdnd11an1n64x5 FILLER_358_72 ();
 b15zdnd11an1n64x5 FILLER_358_136 ();
 b15zdnd11an1n64x5 FILLER_358_200 ();
 b15zdnd11an1n64x5 FILLER_358_264 ();
 b15zdnd11an1n64x5 FILLER_358_328 ();
 b15zdnd11an1n64x5 FILLER_358_392 ();
 b15zdnd11an1n64x5 FILLER_358_456 ();
 b15zdnd11an1n64x5 FILLER_358_520 ();
 b15zdnd11an1n64x5 FILLER_358_584 ();
 b15zdnd11an1n64x5 FILLER_358_648 ();
 b15zdnd11an1n04x5 FILLER_358_712 ();
 b15zdnd00an1n02x5 FILLER_358_716 ();
 b15zdnd11an1n64x5 FILLER_358_726 ();
 b15zdnd11an1n64x5 FILLER_358_790 ();
 b15zdnd11an1n64x5 FILLER_358_854 ();
 b15zdnd11an1n64x5 FILLER_358_918 ();
 b15zdnd11an1n64x5 FILLER_358_982 ();
 b15zdnd11an1n16x5 FILLER_358_1046 ();
 b15zdnd11an1n16x5 FILLER_358_1107 ();
 b15zdnd11an1n08x5 FILLER_358_1123 ();
 b15zdnd00an1n02x5 FILLER_358_1131 ();
 b15zdnd00an1n01x5 FILLER_358_1133 ();
 b15zdnd11an1n16x5 FILLER_358_1144 ();
 b15zdnd11an1n08x5 FILLER_358_1160 ();
 b15zdnd00an1n02x5 FILLER_358_1168 ();
 b15zdnd00an1n01x5 FILLER_358_1170 ();
 b15zdnd11an1n64x5 FILLER_358_1189 ();
 b15zdnd11an1n64x5 FILLER_358_1253 ();
 b15zdnd11an1n16x5 FILLER_358_1317 ();
 b15zdnd00an1n01x5 FILLER_358_1333 ();
 b15zdnd11an1n64x5 FILLER_358_1374 ();
 b15zdnd11an1n64x5 FILLER_358_1438 ();
 b15zdnd11an1n64x5 FILLER_358_1502 ();
 b15zdnd11an1n64x5 FILLER_358_1566 ();
 b15zdnd11an1n64x5 FILLER_358_1630 ();
 b15zdnd11an1n32x5 FILLER_358_1694 ();
 b15zdnd00an1n02x5 FILLER_358_1726 ();
 b15zdnd11an1n64x5 FILLER_358_1770 ();
 b15zdnd11an1n32x5 FILLER_358_1834 ();
 b15zdnd11an1n16x5 FILLER_358_1866 ();
 b15zdnd11an1n08x5 FILLER_358_1882 ();
 b15zdnd11an1n04x5 FILLER_358_1890 ();
 b15zdnd11an1n64x5 FILLER_358_1946 ();
 b15zdnd11an1n64x5 FILLER_358_2010 ();
 b15zdnd11an1n64x5 FILLER_358_2074 ();
 b15zdnd11an1n16x5 FILLER_358_2138 ();
 b15zdnd11an1n64x5 FILLER_358_2162 ();
 b15zdnd11an1n32x5 FILLER_358_2226 ();
 b15zdnd11an1n16x5 FILLER_358_2258 ();
 b15zdnd00an1n02x5 FILLER_358_2274 ();
 b15zdnd11an1n64x5 FILLER_359_0 ();
 b15zdnd11an1n64x5 FILLER_359_64 ();
 b15zdnd11an1n64x5 FILLER_359_128 ();
 b15zdnd11an1n32x5 FILLER_359_192 ();
 b15zdnd11an1n16x5 FILLER_359_224 ();
 b15zdnd11an1n08x5 FILLER_359_240 ();
 b15zdnd00an1n01x5 FILLER_359_248 ();
 b15zdnd11an1n08x5 FILLER_359_256 ();
 b15zdnd11an1n64x5 FILLER_359_267 ();
 b15zdnd11an1n64x5 FILLER_359_331 ();
 b15zdnd11an1n64x5 FILLER_359_395 ();
 b15zdnd11an1n64x5 FILLER_359_459 ();
 b15zdnd11an1n64x5 FILLER_359_523 ();
 b15zdnd11an1n64x5 FILLER_359_587 ();
 b15zdnd11an1n64x5 FILLER_359_651 ();
 b15zdnd11an1n64x5 FILLER_359_715 ();
 b15zdnd11an1n64x5 FILLER_359_779 ();
 b15zdnd11an1n64x5 FILLER_359_843 ();
 b15zdnd11an1n64x5 FILLER_359_907 ();
 b15zdnd11an1n64x5 FILLER_359_971 ();
 b15zdnd11an1n64x5 FILLER_359_1035 ();
 b15zdnd11an1n64x5 FILLER_359_1099 ();
 b15zdnd11an1n64x5 FILLER_359_1163 ();
 b15zdnd11an1n64x5 FILLER_359_1227 ();
 b15zdnd11an1n32x5 FILLER_359_1291 ();
 b15zdnd11an1n16x5 FILLER_359_1323 ();
 b15zdnd11an1n04x5 FILLER_359_1339 ();
 b15zdnd00an1n01x5 FILLER_359_1343 ();
 b15zdnd11an1n04x5 FILLER_359_1384 ();
 b15zdnd11an1n64x5 FILLER_359_1391 ();
 b15zdnd11an1n64x5 FILLER_359_1455 ();
 b15zdnd11an1n64x5 FILLER_359_1519 ();
 b15zdnd11an1n64x5 FILLER_359_1583 ();
 b15zdnd11an1n32x5 FILLER_359_1647 ();
 b15zdnd11an1n16x5 FILLER_359_1679 ();
 b15zdnd11an1n64x5 FILLER_359_1737 ();
 b15zdnd11an1n64x5 FILLER_359_1801 ();
 b15zdnd11an1n32x5 FILLER_359_1865 ();
 b15zdnd11an1n16x5 FILLER_359_1897 ();
 b15zdnd00an1n02x5 FILLER_359_1913 ();
 b15zdnd00an1n01x5 FILLER_359_1915 ();
 b15zdnd11an1n04x5 FILLER_359_1919 ();
 b15zdnd00an1n02x5 FILLER_359_1923 ();
 b15zdnd00an1n01x5 FILLER_359_1925 ();
 b15zdnd11an1n04x5 FILLER_359_1929 ();
 b15zdnd00an1n02x5 FILLER_359_1933 ();
 b15zdnd00an1n01x5 FILLER_359_1935 ();
 b15zdnd11an1n64x5 FILLER_359_1978 ();
 b15zdnd11an1n64x5 FILLER_359_2042 ();
 b15zdnd11an1n64x5 FILLER_359_2106 ();
 b15zdnd11an1n64x5 FILLER_359_2170 ();
 b15zdnd11an1n32x5 FILLER_359_2234 ();
 b15zdnd11an1n16x5 FILLER_359_2266 ();
 b15zdnd00an1n02x5 FILLER_359_2282 ();
 b15zdnd11an1n64x5 FILLER_360_8 ();
 b15zdnd11an1n64x5 FILLER_360_72 ();
 b15zdnd11an1n64x5 FILLER_360_136 ();
 b15zdnd11an1n32x5 FILLER_360_200 ();
 b15zdnd11an1n08x5 FILLER_360_232 ();
 b15zdnd11an1n04x5 FILLER_360_240 ();
 b15zdnd00an1n01x5 FILLER_360_244 ();
 b15zdnd11an1n04x5 FILLER_360_250 ();
 b15zdnd11an1n64x5 FILLER_360_258 ();
 b15zdnd11an1n64x5 FILLER_360_322 ();
 b15zdnd11an1n64x5 FILLER_360_386 ();
 b15zdnd11an1n64x5 FILLER_360_450 ();
 b15zdnd11an1n64x5 FILLER_360_514 ();
 b15zdnd11an1n64x5 FILLER_360_578 ();
 b15zdnd11an1n64x5 FILLER_360_642 ();
 b15zdnd11an1n08x5 FILLER_360_706 ();
 b15zdnd11an1n04x5 FILLER_360_714 ();
 b15zdnd11an1n16x5 FILLER_360_726 ();
 b15zdnd11an1n08x5 FILLER_360_742 ();
 b15zdnd00an1n02x5 FILLER_360_750 ();
 b15zdnd11an1n64x5 FILLER_360_757 ();
 b15zdnd11an1n64x5 FILLER_360_821 ();
 b15zdnd11an1n64x5 FILLER_360_885 ();
 b15zdnd11an1n64x5 FILLER_360_949 ();
 b15zdnd11an1n64x5 FILLER_360_1013 ();
 b15zdnd11an1n64x5 FILLER_360_1077 ();
 b15zdnd11an1n64x5 FILLER_360_1141 ();
 b15zdnd11an1n64x5 FILLER_360_1205 ();
 b15zdnd11an1n64x5 FILLER_360_1269 ();
 b15zdnd11an1n64x5 FILLER_360_1333 ();
 b15zdnd11an1n32x5 FILLER_360_1397 ();
 b15zdnd00an1n01x5 FILLER_360_1429 ();
 b15zdnd11an1n64x5 FILLER_360_1455 ();
 b15zdnd11an1n64x5 FILLER_360_1519 ();
 b15zdnd11an1n64x5 FILLER_360_1583 ();
 b15zdnd11an1n64x5 FILLER_360_1647 ();
 b15zdnd11an1n64x5 FILLER_360_1711 ();
 b15zdnd11an1n64x5 FILLER_360_1775 ();
 b15zdnd11an1n64x5 FILLER_360_1839 ();
 b15zdnd11an1n64x5 FILLER_360_1903 ();
 b15zdnd11an1n64x5 FILLER_360_1967 ();
 b15zdnd11an1n64x5 FILLER_360_2031 ();
 b15zdnd11an1n32x5 FILLER_360_2095 ();
 b15zdnd11an1n16x5 FILLER_360_2127 ();
 b15zdnd11an1n08x5 FILLER_360_2143 ();
 b15zdnd00an1n02x5 FILLER_360_2151 ();
 b15zdnd00an1n01x5 FILLER_360_2153 ();
 b15zdnd11an1n64x5 FILLER_360_2162 ();
 b15zdnd11an1n32x5 FILLER_360_2226 ();
 b15zdnd11an1n16x5 FILLER_360_2258 ();
 b15zdnd00an1n02x5 FILLER_360_2274 ();
 b15zdnd11an1n64x5 FILLER_361_0 ();
 b15zdnd11an1n64x5 FILLER_361_64 ();
 b15zdnd11an1n64x5 FILLER_361_128 ();
 b15zdnd11an1n64x5 FILLER_361_192 ();
 b15zdnd11an1n64x5 FILLER_361_256 ();
 b15zdnd11an1n64x5 FILLER_361_320 ();
 b15zdnd11an1n64x5 FILLER_361_384 ();
 b15zdnd11an1n64x5 FILLER_361_448 ();
 b15zdnd11an1n64x5 FILLER_361_512 ();
 b15zdnd11an1n64x5 FILLER_361_576 ();
 b15zdnd11an1n64x5 FILLER_361_640 ();
 b15zdnd11an1n64x5 FILLER_361_704 ();
 b15zdnd11an1n64x5 FILLER_361_768 ();
 b15zdnd11an1n64x5 FILLER_361_832 ();
 b15zdnd11an1n64x5 FILLER_361_896 ();
 b15zdnd11an1n64x5 FILLER_361_960 ();
 b15zdnd11an1n64x5 FILLER_361_1024 ();
 b15zdnd00an1n02x5 FILLER_361_1088 ();
 b15zdnd11an1n32x5 FILLER_361_1132 ();
 b15zdnd11an1n16x5 FILLER_361_1164 ();
 b15zdnd11an1n08x5 FILLER_361_1180 ();
 b15zdnd00an1n01x5 FILLER_361_1188 ();
 b15zdnd11an1n64x5 FILLER_361_1207 ();
 b15zdnd11an1n64x5 FILLER_361_1271 ();
 b15zdnd11an1n32x5 FILLER_361_1335 ();
 b15zdnd11an1n16x5 FILLER_361_1367 ();
 b15zdnd11an1n08x5 FILLER_361_1383 ();
 b15zdnd11an1n64x5 FILLER_361_1409 ();
 b15zdnd11an1n64x5 FILLER_361_1473 ();
 b15zdnd11an1n32x5 FILLER_361_1537 ();
 b15zdnd11an1n08x5 FILLER_361_1569 ();
 b15zdnd11an1n04x5 FILLER_361_1577 ();
 b15zdnd00an1n02x5 FILLER_361_1581 ();
 b15zdnd11an1n04x5 FILLER_361_1625 ();
 b15zdnd11an1n64x5 FILLER_361_1671 ();
 b15zdnd11an1n64x5 FILLER_361_1735 ();
 b15zdnd11an1n64x5 FILLER_361_1799 ();
 b15zdnd11an1n64x5 FILLER_361_1863 ();
 b15zdnd11an1n64x5 FILLER_361_1927 ();
 b15zdnd11an1n64x5 FILLER_361_1991 ();
 b15zdnd11an1n64x5 FILLER_361_2055 ();
 b15zdnd11an1n64x5 FILLER_361_2119 ();
 b15zdnd11an1n64x5 FILLER_361_2183 ();
 b15zdnd11an1n32x5 FILLER_361_2247 ();
 b15zdnd11an1n04x5 FILLER_361_2279 ();
 b15zdnd00an1n01x5 FILLER_361_2283 ();
 b15zdnd11an1n64x5 FILLER_362_8 ();
 b15zdnd11an1n64x5 FILLER_362_72 ();
 b15zdnd11an1n64x5 FILLER_362_136 ();
 b15zdnd11an1n32x5 FILLER_362_200 ();
 b15zdnd11an1n16x5 FILLER_362_232 ();
 b15zdnd11an1n04x5 FILLER_362_254 ();
 b15zdnd11an1n64x5 FILLER_362_262 ();
 b15zdnd11an1n64x5 FILLER_362_326 ();
 b15zdnd11an1n64x5 FILLER_362_390 ();
 b15zdnd11an1n64x5 FILLER_362_454 ();
 b15zdnd11an1n64x5 FILLER_362_518 ();
 b15zdnd11an1n64x5 FILLER_362_582 ();
 b15zdnd11an1n64x5 FILLER_362_646 ();
 b15zdnd11an1n08x5 FILLER_362_710 ();
 b15zdnd11an1n16x5 FILLER_362_726 ();
 b15zdnd11an1n08x5 FILLER_362_742 ();
 b15zdnd11an1n04x5 FILLER_362_750 ();
 b15zdnd00an1n01x5 FILLER_362_754 ();
 b15zdnd11an1n64x5 FILLER_362_759 ();
 b15zdnd11an1n64x5 FILLER_362_823 ();
 b15zdnd11an1n64x5 FILLER_362_887 ();
 b15zdnd11an1n64x5 FILLER_362_951 ();
 b15zdnd11an1n64x5 FILLER_362_1015 ();
 b15zdnd11an1n64x5 FILLER_362_1079 ();
 b15zdnd11an1n32x5 FILLER_362_1143 ();
 b15zdnd11an1n08x5 FILLER_362_1175 ();
 b15zdnd11an1n04x5 FILLER_362_1183 ();
 b15zdnd00an1n02x5 FILLER_362_1187 ();
 b15zdnd00an1n01x5 FILLER_362_1189 ();
 b15zdnd11an1n64x5 FILLER_362_1232 ();
 b15zdnd11an1n64x5 FILLER_362_1296 ();
 b15zdnd11an1n64x5 FILLER_362_1360 ();
 b15zdnd11an1n04x5 FILLER_362_1424 ();
 b15zdnd00an1n01x5 FILLER_362_1428 ();
 b15zdnd11an1n64x5 FILLER_362_1454 ();
 b15zdnd11an1n64x5 FILLER_362_1518 ();
 b15zdnd11an1n64x5 FILLER_362_1582 ();
 b15zdnd11an1n64x5 FILLER_362_1646 ();
 b15zdnd11an1n64x5 FILLER_362_1710 ();
 b15zdnd11an1n64x5 FILLER_362_1774 ();
 b15zdnd11an1n64x5 FILLER_362_1838 ();
 b15zdnd11an1n64x5 FILLER_362_1902 ();
 b15zdnd11an1n64x5 FILLER_362_1966 ();
 b15zdnd11an1n64x5 FILLER_362_2030 ();
 b15zdnd11an1n32x5 FILLER_362_2094 ();
 b15zdnd11an1n16x5 FILLER_362_2126 ();
 b15zdnd11an1n08x5 FILLER_362_2142 ();
 b15zdnd11an1n04x5 FILLER_362_2150 ();
 b15zdnd11an1n64x5 FILLER_362_2162 ();
 b15zdnd11an1n32x5 FILLER_362_2226 ();
 b15zdnd11an1n16x5 FILLER_362_2258 ();
 b15zdnd00an1n02x5 FILLER_362_2274 ();
 b15zdnd11an1n08x5 FILLER_363_0 ();
 b15zdnd11an1n04x5 FILLER_363_8 ();
 b15zdnd11an1n64x5 FILLER_363_32 ();
 b15zdnd11an1n64x5 FILLER_363_96 ();
 b15zdnd11an1n64x5 FILLER_363_160 ();
 b15zdnd11an1n16x5 FILLER_363_224 ();
 b15zdnd11an1n08x5 FILLER_363_240 ();
 b15zdnd00an1n02x5 FILLER_363_248 ();
 b15zdnd00an1n01x5 FILLER_363_250 ();
 b15zdnd11an1n64x5 FILLER_363_256 ();
 b15zdnd11an1n64x5 FILLER_363_320 ();
 b15zdnd11an1n64x5 FILLER_363_384 ();
 b15zdnd11an1n64x5 FILLER_363_448 ();
 b15zdnd11an1n32x5 FILLER_363_512 ();
 b15zdnd11an1n08x5 FILLER_363_544 ();
 b15zdnd00an1n02x5 FILLER_363_552 ();
 b15zdnd11an1n64x5 FILLER_363_596 ();
 b15zdnd11an1n64x5 FILLER_363_660 ();
 b15zdnd11an1n64x5 FILLER_363_724 ();
 b15zdnd11an1n32x5 FILLER_363_788 ();
 b15zdnd11an1n16x5 FILLER_363_820 ();
 b15zdnd11an1n04x5 FILLER_363_836 ();
 b15zdnd00an1n02x5 FILLER_363_840 ();
 b15zdnd11an1n64x5 FILLER_363_853 ();
 b15zdnd11an1n64x5 FILLER_363_917 ();
 b15zdnd11an1n64x5 FILLER_363_981 ();
 b15zdnd11an1n64x5 FILLER_363_1045 ();
 b15zdnd11an1n08x5 FILLER_363_1109 ();
 b15zdnd00an1n01x5 FILLER_363_1117 ();
 b15zdnd11an1n64x5 FILLER_363_1160 ();
 b15zdnd11an1n32x5 FILLER_363_1224 ();
 b15zdnd00an1n02x5 FILLER_363_1256 ();
 b15zdnd11an1n64x5 FILLER_363_1300 ();
 b15zdnd11an1n16x5 FILLER_363_1364 ();
 b15zdnd11an1n08x5 FILLER_363_1380 ();
 b15zdnd11an1n64x5 FILLER_363_1419 ();
 b15zdnd11an1n64x5 FILLER_363_1483 ();
 b15zdnd11an1n64x5 FILLER_363_1547 ();
 b15zdnd11an1n64x5 FILLER_363_1611 ();
 b15zdnd11an1n64x5 FILLER_363_1675 ();
 b15zdnd11an1n64x5 FILLER_363_1739 ();
 b15zdnd11an1n64x5 FILLER_363_1803 ();
 b15zdnd11an1n64x5 FILLER_363_1867 ();
 b15zdnd11an1n64x5 FILLER_363_1931 ();
 b15zdnd11an1n64x5 FILLER_363_1995 ();
 b15zdnd11an1n64x5 FILLER_363_2059 ();
 b15zdnd11an1n64x5 FILLER_363_2123 ();
 b15zdnd11an1n64x5 FILLER_363_2187 ();
 b15zdnd11an1n32x5 FILLER_363_2251 ();
 b15zdnd00an1n01x5 FILLER_363_2283 ();
 b15zdnd00an1n02x5 FILLER_364_8 ();
 b15zdnd11an1n04x5 FILLER_364_52 ();
 b15zdnd11an1n64x5 FILLER_364_70 ();
 b15zdnd11an1n64x5 FILLER_364_134 ();
 b15zdnd11an1n32x5 FILLER_364_198 ();
 b15zdnd11an1n16x5 FILLER_364_230 ();
 b15zdnd11an1n08x5 FILLER_364_246 ();
 b15zdnd00an1n01x5 FILLER_364_254 ();
 b15zdnd11an1n64x5 FILLER_364_297 ();
 b15zdnd11an1n64x5 FILLER_364_361 ();
 b15zdnd11an1n64x5 FILLER_364_425 ();
 b15zdnd11an1n64x5 FILLER_364_489 ();
 b15zdnd11an1n64x5 FILLER_364_553 ();
 b15zdnd11an1n64x5 FILLER_364_617 ();
 b15zdnd11an1n32x5 FILLER_364_681 ();
 b15zdnd11an1n04x5 FILLER_364_713 ();
 b15zdnd00an1n01x5 FILLER_364_717 ();
 b15zdnd11an1n64x5 FILLER_364_726 ();
 b15zdnd11an1n64x5 FILLER_364_790 ();
 b15zdnd11an1n64x5 FILLER_364_854 ();
 b15zdnd11an1n64x5 FILLER_364_918 ();
 b15zdnd11an1n64x5 FILLER_364_982 ();
 b15zdnd11an1n64x5 FILLER_364_1046 ();
 b15zdnd11an1n64x5 FILLER_364_1110 ();
 b15zdnd11an1n64x5 FILLER_364_1174 ();
 b15zdnd11an1n16x5 FILLER_364_1238 ();
 b15zdnd11an1n04x5 FILLER_364_1254 ();
 b15zdnd00an1n01x5 FILLER_364_1258 ();
 b15zdnd11an1n64x5 FILLER_364_1277 ();
 b15zdnd11an1n64x5 FILLER_364_1341 ();
 b15zdnd11an1n64x5 FILLER_364_1405 ();
 b15zdnd11an1n64x5 FILLER_364_1469 ();
 b15zdnd11an1n64x5 FILLER_364_1533 ();
 b15zdnd11an1n64x5 FILLER_364_1597 ();
 b15zdnd11an1n64x5 FILLER_364_1661 ();
 b15zdnd11an1n64x5 FILLER_364_1725 ();
 b15zdnd11an1n64x5 FILLER_364_1789 ();
 b15zdnd11an1n64x5 FILLER_364_1853 ();
 b15zdnd11an1n64x5 FILLER_364_1917 ();
 b15zdnd11an1n64x5 FILLER_364_1981 ();
 b15zdnd11an1n64x5 FILLER_364_2045 ();
 b15zdnd11an1n32x5 FILLER_364_2109 ();
 b15zdnd11an1n08x5 FILLER_364_2141 ();
 b15zdnd11an1n04x5 FILLER_364_2149 ();
 b15zdnd00an1n01x5 FILLER_364_2153 ();
 b15zdnd11an1n64x5 FILLER_364_2162 ();
 b15zdnd11an1n32x5 FILLER_364_2226 ();
 b15zdnd11an1n16x5 FILLER_364_2258 ();
 b15zdnd00an1n02x5 FILLER_364_2274 ();
 b15zdnd11an1n64x5 FILLER_365_0 ();
 b15zdnd11an1n64x5 FILLER_365_64 ();
 b15zdnd11an1n64x5 FILLER_365_128 ();
 b15zdnd11an1n32x5 FILLER_365_192 ();
 b15zdnd11an1n08x5 FILLER_365_224 ();
 b15zdnd11an1n04x5 FILLER_365_274 ();
 b15zdnd11an1n64x5 FILLER_365_281 ();
 b15zdnd11an1n64x5 FILLER_365_345 ();
 b15zdnd11an1n64x5 FILLER_365_409 ();
 b15zdnd11an1n64x5 FILLER_365_473 ();
 b15zdnd11an1n64x5 FILLER_365_537 ();
 b15zdnd11an1n64x5 FILLER_365_601 ();
 b15zdnd11an1n64x5 FILLER_365_665 ();
 b15zdnd11an1n64x5 FILLER_365_729 ();
 b15zdnd11an1n64x5 FILLER_365_793 ();
 b15zdnd11an1n08x5 FILLER_365_857 ();
 b15zdnd11an1n04x5 FILLER_365_865 ();
 b15zdnd11an1n16x5 FILLER_365_872 ();
 b15zdnd11an1n04x5 FILLER_365_888 ();
 b15zdnd11an1n64x5 FILLER_365_899 ();
 b15zdnd11an1n64x5 FILLER_365_963 ();
 b15zdnd11an1n64x5 FILLER_365_1027 ();
 b15zdnd11an1n64x5 FILLER_365_1091 ();
 b15zdnd11an1n16x5 FILLER_365_1155 ();
 b15zdnd11an1n08x5 FILLER_365_1171 ();
 b15zdnd11an1n64x5 FILLER_365_1191 ();
 b15zdnd11an1n64x5 FILLER_365_1255 ();
 b15zdnd11an1n64x5 FILLER_365_1319 ();
 b15zdnd11an1n64x5 FILLER_365_1383 ();
 b15zdnd11an1n64x5 FILLER_365_1447 ();
 b15zdnd11an1n64x5 FILLER_365_1511 ();
 b15zdnd11an1n64x5 FILLER_365_1575 ();
 b15zdnd11an1n32x5 FILLER_365_1639 ();
 b15zdnd11an1n16x5 FILLER_365_1671 ();
 b15zdnd11an1n04x5 FILLER_365_1687 ();
 b15zdnd00an1n02x5 FILLER_365_1691 ();
 b15zdnd11an1n64x5 FILLER_365_1696 ();
 b15zdnd11an1n64x5 FILLER_365_1760 ();
 b15zdnd11an1n64x5 FILLER_365_1824 ();
 b15zdnd11an1n64x5 FILLER_365_1888 ();
 b15zdnd11an1n64x5 FILLER_365_1952 ();
 b15zdnd11an1n64x5 FILLER_365_2016 ();
 b15zdnd11an1n64x5 FILLER_365_2080 ();
 b15zdnd11an1n64x5 FILLER_365_2144 ();
 b15zdnd11an1n64x5 FILLER_365_2208 ();
 b15zdnd11an1n08x5 FILLER_365_2272 ();
 b15zdnd11an1n04x5 FILLER_365_2280 ();
 b15zdnd11an1n64x5 FILLER_366_8 ();
 b15zdnd11an1n64x5 FILLER_366_72 ();
 b15zdnd11an1n64x5 FILLER_366_136 ();
 b15zdnd11an1n32x5 FILLER_366_200 ();
 b15zdnd00an1n02x5 FILLER_366_232 ();
 b15zdnd11an1n64x5 FILLER_366_276 ();
 b15zdnd11an1n64x5 FILLER_366_340 ();
 b15zdnd11an1n64x5 FILLER_366_404 ();
 b15zdnd11an1n64x5 FILLER_366_468 ();
 b15zdnd11an1n64x5 FILLER_366_532 ();
 b15zdnd11an1n64x5 FILLER_366_596 ();
 b15zdnd11an1n32x5 FILLER_366_660 ();
 b15zdnd11an1n16x5 FILLER_366_692 ();
 b15zdnd11an1n08x5 FILLER_366_708 ();
 b15zdnd00an1n02x5 FILLER_366_716 ();
 b15zdnd11an1n64x5 FILLER_366_726 ();
 b15zdnd11an1n32x5 FILLER_366_790 ();
 b15zdnd11an1n16x5 FILLER_366_822 ();
 b15zdnd11an1n04x5 FILLER_366_838 ();
 b15zdnd11an1n04x5 FILLER_366_894 ();
 b15zdnd11an1n64x5 FILLER_366_940 ();
 b15zdnd11an1n64x5 FILLER_366_1004 ();
 b15zdnd11an1n64x5 FILLER_366_1068 ();
 b15zdnd11an1n16x5 FILLER_366_1132 ();
 b15zdnd11an1n08x5 FILLER_366_1148 ();
 b15zdnd00an1n01x5 FILLER_366_1156 ();
 b15zdnd11an1n04x5 FILLER_366_1199 ();
 b15zdnd00an1n01x5 FILLER_366_1203 ();
 b15zdnd11an1n64x5 FILLER_366_1216 ();
 b15zdnd11an1n64x5 FILLER_366_1280 ();
 b15zdnd11an1n64x5 FILLER_366_1344 ();
 b15zdnd11an1n64x5 FILLER_366_1408 ();
 b15zdnd11an1n64x5 FILLER_366_1472 ();
 b15zdnd11an1n64x5 FILLER_366_1536 ();
 b15zdnd11an1n16x5 FILLER_366_1600 ();
 b15zdnd11an1n64x5 FILLER_366_1619 ();
 b15zdnd00an1n02x5 FILLER_366_1683 ();
 b15zdnd11an1n04x5 FILLER_366_1688 ();
 b15zdnd11an1n64x5 FILLER_366_1695 ();
 b15zdnd11an1n04x5 FILLER_366_1759 ();
 b15zdnd00an1n02x5 FILLER_366_1763 ();
 b15zdnd11an1n04x5 FILLER_366_1768 ();
 b15zdnd11an1n64x5 FILLER_366_1775 ();
 b15zdnd11an1n64x5 FILLER_366_1839 ();
 b15zdnd11an1n64x5 FILLER_366_1903 ();
 b15zdnd11an1n64x5 FILLER_366_1967 ();
 b15zdnd11an1n64x5 FILLER_366_2031 ();
 b15zdnd11an1n32x5 FILLER_366_2095 ();
 b15zdnd11an1n16x5 FILLER_366_2127 ();
 b15zdnd11an1n08x5 FILLER_366_2143 ();
 b15zdnd00an1n02x5 FILLER_366_2151 ();
 b15zdnd00an1n01x5 FILLER_366_2153 ();
 b15zdnd11an1n64x5 FILLER_366_2162 ();
 b15zdnd11an1n32x5 FILLER_366_2226 ();
 b15zdnd11an1n16x5 FILLER_366_2258 ();
 b15zdnd00an1n02x5 FILLER_366_2274 ();
 b15zdnd11an1n64x5 FILLER_367_0 ();
 b15zdnd11an1n64x5 FILLER_367_64 ();
 b15zdnd11an1n64x5 FILLER_367_128 ();
 b15zdnd11an1n32x5 FILLER_367_192 ();
 b15zdnd11an1n16x5 FILLER_367_224 ();
 b15zdnd00an1n02x5 FILLER_367_240 ();
 b15zdnd00an1n01x5 FILLER_367_242 ();
 b15zdnd11an1n04x5 FILLER_367_249 ();
 b15zdnd11an1n64x5 FILLER_367_260 ();
 b15zdnd11an1n64x5 FILLER_367_324 ();
 b15zdnd11an1n32x5 FILLER_367_388 ();
 b15zdnd11an1n04x5 FILLER_367_420 ();
 b15zdnd00an1n02x5 FILLER_367_424 ();
 b15zdnd11an1n64x5 FILLER_367_429 ();
 b15zdnd11an1n64x5 FILLER_367_493 ();
 b15zdnd00an1n02x5 FILLER_367_557 ();
 b15zdnd00an1n01x5 FILLER_367_559 ();
 b15zdnd11an1n04x5 FILLER_367_600 ();
 b15zdnd00an1n02x5 FILLER_367_604 ();
 b15zdnd00an1n01x5 FILLER_367_606 ();
 b15zdnd11an1n64x5 FILLER_367_610 ();
 b15zdnd11an1n64x5 FILLER_367_674 ();
 b15zdnd11an1n64x5 FILLER_367_738 ();
 b15zdnd11an1n32x5 FILLER_367_802 ();
 b15zdnd11an1n08x5 FILLER_367_834 ();
 b15zdnd11an1n04x5 FILLER_367_842 ();
 b15zdnd00an1n01x5 FILLER_367_846 ();
 b15zdnd11an1n04x5 FILLER_367_889 ();
 b15zdnd11an1n64x5 FILLER_367_935 ();
 b15zdnd11an1n64x5 FILLER_367_999 ();
 b15zdnd11an1n64x5 FILLER_367_1063 ();
 b15zdnd11an1n16x5 FILLER_367_1127 ();
 b15zdnd11an1n08x5 FILLER_367_1143 ();
 b15zdnd11an1n04x5 FILLER_367_1151 ();
 b15zdnd11an1n32x5 FILLER_367_1175 ();
 b15zdnd11an1n16x5 FILLER_367_1219 ();
 b15zdnd11an1n08x5 FILLER_367_1235 ();
 b15zdnd11an1n08x5 FILLER_367_1285 ();
 b15zdnd00an1n02x5 FILLER_367_1293 ();
 b15zdnd11an1n04x5 FILLER_367_1337 ();
 b15zdnd11an1n64x5 FILLER_367_1383 ();
 b15zdnd11an1n64x5 FILLER_367_1447 ();
 b15zdnd11an1n64x5 FILLER_367_1511 ();
 b15zdnd11an1n32x5 FILLER_367_1575 ();
 b15zdnd11an1n04x5 FILLER_367_1607 ();
 b15zdnd00an1n02x5 FILLER_367_1611 ();
 b15zdnd00an1n01x5 FILLER_367_1613 ();
 b15zdnd11an1n04x5 FILLER_367_1617 ();
 b15zdnd11an1n32x5 FILLER_367_1624 ();
 b15zdnd11an1n08x5 FILLER_367_1656 ();
 b15zdnd00an1n02x5 FILLER_367_1664 ();
 b15zdnd00an1n01x5 FILLER_367_1666 ();
 b15zdnd11an1n32x5 FILLER_367_1719 ();
 b15zdnd00an1n02x5 FILLER_367_1751 ();
 b15zdnd00an1n01x5 FILLER_367_1753 ();
 b15zdnd11an1n04x5 FILLER_367_1757 ();
 b15zdnd11an1n64x5 FILLER_367_1803 ();
 b15zdnd11an1n64x5 FILLER_367_1867 ();
 b15zdnd11an1n64x5 FILLER_367_1931 ();
 b15zdnd11an1n64x5 FILLER_367_1995 ();
 b15zdnd11an1n64x5 FILLER_367_2059 ();
 b15zdnd11an1n64x5 FILLER_367_2123 ();
 b15zdnd11an1n64x5 FILLER_367_2187 ();
 b15zdnd11an1n32x5 FILLER_367_2251 ();
 b15zdnd00an1n01x5 FILLER_367_2283 ();
 b15zdnd11an1n64x5 FILLER_368_8 ();
 b15zdnd11an1n64x5 FILLER_368_72 ();
 b15zdnd11an1n64x5 FILLER_368_136 ();
 b15zdnd11an1n32x5 FILLER_368_200 ();
 b15zdnd11an1n04x5 FILLER_368_232 ();
 b15zdnd00an1n01x5 FILLER_368_236 ();
 b15zdnd11an1n04x5 FILLER_368_240 ();
 b15zdnd11an1n64x5 FILLER_368_286 ();
 b15zdnd11an1n32x5 FILLER_368_350 ();
 b15zdnd11an1n16x5 FILLER_368_382 ();
 b15zdnd11an1n04x5 FILLER_368_398 ();
 b15zdnd00an1n02x5 FILLER_368_402 ();
 b15zdnd00an1n01x5 FILLER_368_404 ();
 b15zdnd11an1n32x5 FILLER_368_414 ();
 b15zdnd11an1n08x5 FILLER_368_446 ();
 b15zdnd11an1n04x5 FILLER_368_454 ();
 b15zdnd00an1n02x5 FILLER_368_458 ();
 b15zdnd11an1n64x5 FILLER_368_469 ();
 b15zdnd11an1n16x5 FILLER_368_533 ();
 b15zdnd11an1n04x5 FILLER_368_549 ();
 b15zdnd11an1n04x5 FILLER_368_567 ();
 b15zdnd11an1n64x5 FILLER_368_611 ();
 b15zdnd11an1n32x5 FILLER_368_675 ();
 b15zdnd11an1n08x5 FILLER_368_707 ();
 b15zdnd00an1n02x5 FILLER_368_715 ();
 b15zdnd00an1n01x5 FILLER_368_717 ();
 b15zdnd11an1n16x5 FILLER_368_726 ();
 b15zdnd11an1n04x5 FILLER_368_742 ();
 b15zdnd11an1n64x5 FILLER_368_749 ();
 b15zdnd11an1n32x5 FILLER_368_813 ();
 b15zdnd11an1n08x5 FILLER_368_845 ();
 b15zdnd00an1n02x5 FILLER_368_853 ();
 b15zdnd11an1n04x5 FILLER_368_858 ();
 b15zdnd11an1n04x5 FILLER_368_865 ();
 b15zdnd11an1n64x5 FILLER_368_921 ();
 b15zdnd11an1n64x5 FILLER_368_985 ();
 b15zdnd11an1n64x5 FILLER_368_1049 ();
 b15zdnd11an1n32x5 FILLER_368_1113 ();
 b15zdnd11an1n16x5 FILLER_368_1145 ();
 b15zdnd11an1n04x5 FILLER_368_1161 ();
 b15zdnd00an1n01x5 FILLER_368_1165 ();
 b15zdnd11an1n64x5 FILLER_368_1173 ();
 b15zdnd11an1n64x5 FILLER_368_1237 ();
 b15zdnd11an1n64x5 FILLER_368_1301 ();
 b15zdnd11an1n64x5 FILLER_368_1365 ();
 b15zdnd11an1n64x5 FILLER_368_1429 ();
 b15zdnd11an1n64x5 FILLER_368_1493 ();
 b15zdnd11an1n32x5 FILLER_368_1557 ();
 b15zdnd11an1n04x5 FILLER_368_1589 ();
 b15zdnd00an1n02x5 FILLER_368_1593 ();
 b15zdnd00an1n01x5 FILLER_368_1595 ();
 b15zdnd11an1n64x5 FILLER_368_1648 ();
 b15zdnd11an1n04x5 FILLER_368_1712 ();
 b15zdnd00an1n01x5 FILLER_368_1716 ();
 b15zdnd11an1n08x5 FILLER_368_1737 ();
 b15zdnd11an1n64x5 FILLER_368_1797 ();
 b15zdnd11an1n64x5 FILLER_368_1861 ();
 b15zdnd11an1n64x5 FILLER_368_1925 ();
 b15zdnd11an1n64x5 FILLER_368_1989 ();
 b15zdnd11an1n64x5 FILLER_368_2053 ();
 b15zdnd11an1n32x5 FILLER_368_2117 ();
 b15zdnd11an1n04x5 FILLER_368_2149 ();
 b15zdnd00an1n01x5 FILLER_368_2153 ();
 b15zdnd11an1n64x5 FILLER_368_2162 ();
 b15zdnd11an1n32x5 FILLER_368_2226 ();
 b15zdnd11an1n16x5 FILLER_368_2258 ();
 b15zdnd00an1n02x5 FILLER_368_2274 ();
 b15zdnd11an1n64x5 FILLER_369_0 ();
 b15zdnd11an1n64x5 FILLER_369_64 ();
 b15zdnd11an1n64x5 FILLER_369_128 ();
 b15zdnd11an1n32x5 FILLER_369_192 ();
 b15zdnd11an1n08x5 FILLER_369_224 ();
 b15zdnd00an1n02x5 FILLER_369_232 ();
 b15zdnd11an1n04x5 FILLER_369_237 ();
 b15zdnd11an1n08x5 FILLER_369_244 ();
 b15zdnd11an1n04x5 FILLER_369_252 ();
 b15zdnd00an1n01x5 FILLER_369_256 ();
 b15zdnd11an1n64x5 FILLER_369_299 ();
 b15zdnd11an1n32x5 FILLER_369_363 ();
 b15zdnd11an1n04x5 FILLER_369_395 ();
 b15zdnd11an1n64x5 FILLER_369_451 ();
 b15zdnd11an1n64x5 FILLER_369_515 ();
 b15zdnd11an1n08x5 FILLER_369_579 ();
 b15zdnd11an1n04x5 FILLER_369_587 ();
 b15zdnd00an1n02x5 FILLER_369_591 ();
 b15zdnd00an1n01x5 FILLER_369_593 ();
 b15zdnd11an1n04x5 FILLER_369_597 ();
 b15zdnd11an1n04x5 FILLER_369_604 ();
 b15zdnd11an1n64x5 FILLER_369_611 ();
 b15zdnd11an1n32x5 FILLER_369_675 ();
 b15zdnd11an1n08x5 FILLER_369_707 ();
 b15zdnd11an1n04x5 FILLER_369_715 ();
 b15zdnd11an1n64x5 FILLER_369_771 ();
 b15zdnd11an1n32x5 FILLER_369_835 ();
 b15zdnd11an1n16x5 FILLER_369_867 ();
 b15zdnd11an1n04x5 FILLER_369_883 ();
 b15zdnd00an1n01x5 FILLER_369_887 ();
 b15zdnd11an1n04x5 FILLER_369_891 ();
 b15zdnd11an1n64x5 FILLER_369_898 ();
 b15zdnd11an1n16x5 FILLER_369_962 ();
 b15zdnd11an1n08x5 FILLER_369_978 ();
 b15zdnd11an1n04x5 FILLER_369_986 ();
 b15zdnd11an1n04x5 FILLER_369_993 ();
 b15zdnd11an1n64x5 FILLER_369_1000 ();
 b15zdnd11an1n64x5 FILLER_369_1064 ();
 b15zdnd11an1n64x5 FILLER_369_1128 ();
 b15zdnd11an1n64x5 FILLER_369_1192 ();
 b15zdnd11an1n64x5 FILLER_369_1256 ();
 b15zdnd11an1n08x5 FILLER_369_1320 ();
 b15zdnd00an1n02x5 FILLER_369_1328 ();
 b15zdnd00an1n01x5 FILLER_369_1330 ();
 b15zdnd11an1n64x5 FILLER_369_1373 ();
 b15zdnd11an1n64x5 FILLER_369_1437 ();
 b15zdnd11an1n64x5 FILLER_369_1501 ();
 b15zdnd11an1n32x5 FILLER_369_1565 ();
 b15zdnd11an1n32x5 FILLER_369_1649 ();
 b15zdnd11an1n16x5 FILLER_369_1681 ();
 b15zdnd00an1n02x5 FILLER_369_1697 ();
 b15zdnd11an1n08x5 FILLER_369_1719 ();
 b15zdnd11an1n04x5 FILLER_369_1727 ();
 b15zdnd00an1n01x5 FILLER_369_1731 ();
 b15zdnd11an1n04x5 FILLER_369_1743 ();
 b15zdnd11an1n64x5 FILLER_369_1767 ();
 b15zdnd11an1n64x5 FILLER_369_1831 ();
 b15zdnd11an1n64x5 FILLER_369_1895 ();
 b15zdnd11an1n64x5 FILLER_369_1959 ();
 b15zdnd11an1n64x5 FILLER_369_2023 ();
 b15zdnd11an1n64x5 FILLER_369_2087 ();
 b15zdnd11an1n64x5 FILLER_369_2151 ();
 b15zdnd11an1n64x5 FILLER_369_2215 ();
 b15zdnd11an1n04x5 FILLER_369_2279 ();
 b15zdnd00an1n01x5 FILLER_369_2283 ();
 b15zdnd11an1n64x5 FILLER_370_8 ();
 b15zdnd11an1n64x5 FILLER_370_72 ();
 b15zdnd11an1n64x5 FILLER_370_136 ();
 b15zdnd11an1n08x5 FILLER_370_200 ();
 b15zdnd11an1n04x5 FILLER_370_208 ();
 b15zdnd00an1n02x5 FILLER_370_212 ();
 b15zdnd11an1n64x5 FILLER_370_266 ();
 b15zdnd11an1n64x5 FILLER_370_330 ();
 b15zdnd11an1n16x5 FILLER_370_394 ();
 b15zdnd11an1n08x5 FILLER_370_410 ();
 b15zdnd00an1n01x5 FILLER_370_418 ();
 b15zdnd11an1n16x5 FILLER_370_422 ();
 b15zdnd11an1n08x5 FILLER_370_438 ();
 b15zdnd00an1n01x5 FILLER_370_446 ();
 b15zdnd11an1n64x5 FILLER_370_474 ();
 b15zdnd11an1n64x5 FILLER_370_538 ();
 b15zdnd11an1n64x5 FILLER_370_602 ();
 b15zdnd11an1n32x5 FILLER_370_666 ();
 b15zdnd11an1n16x5 FILLER_370_698 ();
 b15zdnd11an1n04x5 FILLER_370_714 ();
 b15zdnd11an1n08x5 FILLER_370_726 ();
 b15zdnd00an1n02x5 FILLER_370_734 ();
 b15zdnd00an1n01x5 FILLER_370_736 ();
 b15zdnd11an1n04x5 FILLER_370_740 ();
 b15zdnd11an1n64x5 FILLER_370_747 ();
 b15zdnd11an1n64x5 FILLER_370_811 ();
 b15zdnd11an1n16x5 FILLER_370_875 ();
 b15zdnd11an1n04x5 FILLER_370_891 ();
 b15zdnd00an1n01x5 FILLER_370_895 ();
 b15zdnd11an1n16x5 FILLER_370_899 ();
 b15zdnd11an1n04x5 FILLER_370_915 ();
 b15zdnd00an1n02x5 FILLER_370_919 ();
 b15zdnd00an1n01x5 FILLER_370_921 ();
 b15zdnd11an1n16x5 FILLER_370_942 ();
 b15zdnd11an1n08x5 FILLER_370_958 ();
 b15zdnd00an1n01x5 FILLER_370_966 ();
 b15zdnd11an1n64x5 FILLER_370_1019 ();
 b15zdnd11an1n64x5 FILLER_370_1083 ();
 b15zdnd11an1n32x5 FILLER_370_1147 ();
 b15zdnd11an1n08x5 FILLER_370_1179 ();
 b15zdnd11an1n04x5 FILLER_370_1187 ();
 b15zdnd00an1n02x5 FILLER_370_1191 ();
 b15zdnd11an1n64x5 FILLER_370_1208 ();
 b15zdnd11an1n64x5 FILLER_370_1272 ();
 b15zdnd11an1n64x5 FILLER_370_1336 ();
 b15zdnd11an1n64x5 FILLER_370_1400 ();
 b15zdnd11an1n64x5 FILLER_370_1464 ();
 b15zdnd11an1n32x5 FILLER_370_1528 ();
 b15zdnd11an1n16x5 FILLER_370_1560 ();
 b15zdnd11an1n08x5 FILLER_370_1576 ();
 b15zdnd11an1n04x5 FILLER_370_1584 ();
 b15zdnd00an1n01x5 FILLER_370_1588 ();
 b15zdnd11an1n04x5 FILLER_370_1631 ();
 b15zdnd11an1n64x5 FILLER_370_1638 ();
 b15zdnd11an1n64x5 FILLER_370_1702 ();
 b15zdnd11an1n64x5 FILLER_370_1766 ();
 b15zdnd11an1n64x5 FILLER_370_1830 ();
 b15zdnd11an1n64x5 FILLER_370_1894 ();
 b15zdnd11an1n64x5 FILLER_370_1958 ();
 b15zdnd11an1n64x5 FILLER_370_2022 ();
 b15zdnd11an1n64x5 FILLER_370_2086 ();
 b15zdnd11an1n04x5 FILLER_370_2150 ();
 b15zdnd11an1n64x5 FILLER_370_2162 ();
 b15zdnd11an1n32x5 FILLER_370_2226 ();
 b15zdnd11an1n16x5 FILLER_370_2258 ();
 b15zdnd00an1n02x5 FILLER_370_2274 ();
 b15zdnd11an1n64x5 FILLER_371_0 ();
 b15zdnd11an1n64x5 FILLER_371_64 ();
 b15zdnd11an1n64x5 FILLER_371_128 ();
 b15zdnd11an1n32x5 FILLER_371_192 ();
 b15zdnd11an1n16x5 FILLER_371_224 ();
 b15zdnd11an1n04x5 FILLER_371_260 ();
 b15zdnd11an1n64x5 FILLER_371_284 ();
 b15zdnd11an1n64x5 FILLER_371_348 ();
 b15zdnd11an1n08x5 FILLER_371_412 ();
 b15zdnd11an1n04x5 FILLER_371_423 ();
 b15zdnd11an1n04x5 FILLER_371_479 ();
 b15zdnd11an1n64x5 FILLER_371_486 ();
 b15zdnd11an1n64x5 FILLER_371_550 ();
 b15zdnd11an1n64x5 FILLER_371_614 ();
 b15zdnd11an1n32x5 FILLER_371_678 ();
 b15zdnd11an1n04x5 FILLER_371_710 ();
 b15zdnd00an1n01x5 FILLER_371_714 ();
 b15zdnd11an1n32x5 FILLER_371_726 ();
 b15zdnd00an1n02x5 FILLER_371_758 ();
 b15zdnd00an1n01x5 FILLER_371_760 ();
 b15zdnd11an1n64x5 FILLER_371_764 ();
 b15zdnd11an1n64x5 FILLER_371_828 ();
 b15zdnd11an1n64x5 FILLER_371_892 ();
 b15zdnd11an1n32x5 FILLER_371_956 ();
 b15zdnd11an1n08x5 FILLER_371_988 ();
 b15zdnd00an1n02x5 FILLER_371_996 ();
 b15zdnd00an1n01x5 FILLER_371_998 ();
 b15zdnd11an1n32x5 FILLER_371_1002 ();
 b15zdnd11an1n16x5 FILLER_371_1034 ();
 b15zdnd00an1n01x5 FILLER_371_1050 ();
 b15zdnd11an1n64x5 FILLER_371_1093 ();
 b15zdnd11an1n32x5 FILLER_371_1157 ();
 b15zdnd11an1n16x5 FILLER_371_1189 ();
 b15zdnd11an1n08x5 FILLER_371_1205 ();
 b15zdnd11an1n04x5 FILLER_371_1213 ();
 b15zdnd00an1n01x5 FILLER_371_1217 ();
 b15zdnd11an1n64x5 FILLER_371_1232 ();
 b15zdnd11an1n64x5 FILLER_371_1296 ();
 b15zdnd11an1n64x5 FILLER_371_1360 ();
 b15zdnd11an1n64x5 FILLER_371_1424 ();
 b15zdnd11an1n64x5 FILLER_371_1488 ();
 b15zdnd11an1n32x5 FILLER_371_1552 ();
 b15zdnd11an1n16x5 FILLER_371_1584 ();
 b15zdnd11an1n08x5 FILLER_371_1600 ();
 b15zdnd11an1n04x5 FILLER_371_1608 ();
 b15zdnd00an1n02x5 FILLER_371_1612 ();
 b15zdnd00an1n01x5 FILLER_371_1614 ();
 b15zdnd11an1n04x5 FILLER_371_1618 ();
 b15zdnd11an1n64x5 FILLER_371_1664 ();
 b15zdnd11an1n64x5 FILLER_371_1728 ();
 b15zdnd11an1n64x5 FILLER_371_1792 ();
 b15zdnd11an1n64x5 FILLER_371_1856 ();
 b15zdnd11an1n64x5 FILLER_371_1920 ();
 b15zdnd11an1n64x5 FILLER_371_1984 ();
 b15zdnd11an1n64x5 FILLER_371_2048 ();
 b15zdnd11an1n64x5 FILLER_371_2112 ();
 b15zdnd11an1n64x5 FILLER_371_2176 ();
 b15zdnd11an1n32x5 FILLER_371_2240 ();
 b15zdnd11an1n08x5 FILLER_371_2272 ();
 b15zdnd11an1n04x5 FILLER_371_2280 ();
 b15zdnd11an1n64x5 FILLER_372_8 ();
 b15zdnd11an1n64x5 FILLER_372_72 ();
 b15zdnd11an1n64x5 FILLER_372_136 ();
 b15zdnd11an1n64x5 FILLER_372_200 ();
 b15zdnd00an1n02x5 FILLER_372_264 ();
 b15zdnd00an1n01x5 FILLER_372_266 ();
 b15zdnd11an1n64x5 FILLER_372_278 ();
 b15zdnd11an1n64x5 FILLER_372_342 ();
 b15zdnd11an1n16x5 FILLER_372_406 ();
 b15zdnd11an1n04x5 FILLER_372_422 ();
 b15zdnd00an1n02x5 FILLER_372_426 ();
 b15zdnd11an1n04x5 FILLER_372_480 ();
 b15zdnd11an1n64x5 FILLER_372_487 ();
 b15zdnd11an1n64x5 FILLER_372_551 ();
 b15zdnd11an1n64x5 FILLER_372_615 ();
 b15zdnd11an1n32x5 FILLER_372_679 ();
 b15zdnd11an1n04x5 FILLER_372_711 ();
 b15zdnd00an1n02x5 FILLER_372_715 ();
 b15zdnd00an1n01x5 FILLER_372_717 ();
 b15zdnd11an1n08x5 FILLER_372_726 ();
 b15zdnd11an1n64x5 FILLER_372_786 ();
 b15zdnd11an1n64x5 FILLER_372_850 ();
 b15zdnd11an1n64x5 FILLER_372_914 ();
 b15zdnd11an1n64x5 FILLER_372_978 ();
 b15zdnd11an1n64x5 FILLER_372_1042 ();
 b15zdnd11an1n64x5 FILLER_372_1106 ();
 b15zdnd11an1n32x5 FILLER_372_1170 ();
 b15zdnd00an1n02x5 FILLER_372_1202 ();
 b15zdnd00an1n01x5 FILLER_372_1204 ();
 b15zdnd11an1n32x5 FILLER_372_1247 ();
 b15zdnd11an1n16x5 FILLER_372_1279 ();
 b15zdnd11an1n04x5 FILLER_372_1295 ();
 b15zdnd00an1n02x5 FILLER_372_1299 ();
 b15zdnd00an1n01x5 FILLER_372_1301 ();
 b15zdnd11an1n16x5 FILLER_372_1344 ();
 b15zdnd11an1n04x5 FILLER_372_1360 ();
 b15zdnd00an1n02x5 FILLER_372_1364 ();
 b15zdnd00an1n01x5 FILLER_372_1366 ();
 b15zdnd11an1n64x5 FILLER_372_1377 ();
 b15zdnd11an1n64x5 FILLER_372_1441 ();
 b15zdnd11an1n64x5 FILLER_372_1505 ();
 b15zdnd11an1n04x5 FILLER_372_1569 ();
 b15zdnd11an1n16x5 FILLER_372_1604 ();
 b15zdnd00an1n02x5 FILLER_372_1620 ();
 b15zdnd00an1n01x5 FILLER_372_1622 ();
 b15zdnd11an1n64x5 FILLER_372_1626 ();
 b15zdnd11an1n64x5 FILLER_372_1690 ();
 b15zdnd11an1n64x5 FILLER_372_1754 ();
 b15zdnd11an1n64x5 FILLER_372_1818 ();
 b15zdnd11an1n64x5 FILLER_372_1882 ();
 b15zdnd11an1n64x5 FILLER_372_1946 ();
 b15zdnd11an1n64x5 FILLER_372_2010 ();
 b15zdnd11an1n64x5 FILLER_372_2074 ();
 b15zdnd11an1n16x5 FILLER_372_2138 ();
 b15zdnd11an1n64x5 FILLER_372_2162 ();
 b15zdnd11an1n32x5 FILLER_372_2226 ();
 b15zdnd11an1n16x5 FILLER_372_2258 ();
 b15zdnd00an1n02x5 FILLER_372_2274 ();
 b15zdnd11an1n64x5 FILLER_373_0 ();
 b15zdnd11an1n64x5 FILLER_373_64 ();
 b15zdnd11an1n64x5 FILLER_373_128 ();
 b15zdnd11an1n64x5 FILLER_373_192 ();
 b15zdnd11an1n64x5 FILLER_373_256 ();
 b15zdnd11an1n64x5 FILLER_373_320 ();
 b15zdnd11an1n16x5 FILLER_373_384 ();
 b15zdnd11an1n08x5 FILLER_373_400 ();
 b15zdnd11an1n04x5 FILLER_373_408 ();
 b15zdnd11an1n04x5 FILLER_373_464 ();
 b15zdnd11an1n64x5 FILLER_373_471 ();
 b15zdnd11an1n32x5 FILLER_373_535 ();
 b15zdnd11an1n08x5 FILLER_373_567 ();
 b15zdnd00an1n01x5 FILLER_373_575 ();
 b15zdnd11an1n64x5 FILLER_373_618 ();
 b15zdnd11an1n64x5 FILLER_373_682 ();
 b15zdnd11an1n04x5 FILLER_373_746 ();
 b15zdnd11an1n04x5 FILLER_373_753 ();
 b15zdnd00an1n02x5 FILLER_373_757 ();
 b15zdnd11an1n64x5 FILLER_373_762 ();
 b15zdnd11an1n32x5 FILLER_373_826 ();
 b15zdnd11an1n16x5 FILLER_373_858 ();
 b15zdnd11an1n08x5 FILLER_373_874 ();
 b15zdnd00an1n02x5 FILLER_373_882 ();
 b15zdnd11an1n64x5 FILLER_373_926 ();
 b15zdnd11an1n64x5 FILLER_373_990 ();
 b15zdnd11an1n64x5 FILLER_373_1054 ();
 b15zdnd11an1n32x5 FILLER_373_1118 ();
 b15zdnd11an1n16x5 FILLER_373_1150 ();
 b15zdnd00an1n01x5 FILLER_373_1166 ();
 b15zdnd11an1n64x5 FILLER_373_1209 ();
 b15zdnd11an1n32x5 FILLER_373_1273 ();
 b15zdnd11an1n16x5 FILLER_373_1305 ();
 b15zdnd11an1n08x5 FILLER_373_1321 ();
 b15zdnd11an1n08x5 FILLER_373_1371 ();
 b15zdnd00an1n02x5 FILLER_373_1379 ();
 b15zdnd11an1n64x5 FILLER_373_1396 ();
 b15zdnd11an1n64x5 FILLER_373_1460 ();
 b15zdnd11an1n16x5 FILLER_373_1524 ();
 b15zdnd11an1n08x5 FILLER_373_1540 ();
 b15zdnd11an1n32x5 FILLER_373_1563 ();
 b15zdnd11an1n16x5 FILLER_373_1595 ();
 b15zdnd11an1n04x5 FILLER_373_1611 ();
 b15zdnd11an1n64x5 FILLER_373_1657 ();
 b15zdnd11an1n64x5 FILLER_373_1721 ();
 b15zdnd11an1n64x5 FILLER_373_1785 ();
 b15zdnd11an1n64x5 FILLER_373_1849 ();
 b15zdnd11an1n64x5 FILLER_373_1913 ();
 b15zdnd11an1n64x5 FILLER_373_1977 ();
 b15zdnd11an1n64x5 FILLER_373_2041 ();
 b15zdnd11an1n64x5 FILLER_373_2105 ();
 b15zdnd11an1n64x5 FILLER_373_2169 ();
 b15zdnd11an1n32x5 FILLER_373_2233 ();
 b15zdnd11an1n16x5 FILLER_373_2265 ();
 b15zdnd00an1n02x5 FILLER_373_2281 ();
 b15zdnd00an1n01x5 FILLER_373_2283 ();
 b15zdnd11an1n64x5 FILLER_374_8 ();
 b15zdnd11an1n64x5 FILLER_374_72 ();
 b15zdnd11an1n64x5 FILLER_374_136 ();
 b15zdnd11an1n64x5 FILLER_374_200 ();
 b15zdnd11an1n64x5 FILLER_374_264 ();
 b15zdnd11an1n64x5 FILLER_374_328 ();
 b15zdnd11an1n16x5 FILLER_374_392 ();
 b15zdnd11an1n08x5 FILLER_374_408 ();
 b15zdnd00an1n02x5 FILLER_374_416 ();
 b15zdnd11an1n04x5 FILLER_374_421 ();
 b15zdnd11an1n04x5 FILLER_374_428 ();
 b15zdnd11an1n04x5 FILLER_374_435 ();
 b15zdnd11an1n04x5 FILLER_374_442 ();
 b15zdnd11an1n04x5 FILLER_374_455 ();
 b15zdnd11an1n04x5 FILLER_374_462 ();
 b15zdnd00an1n01x5 FILLER_374_466 ();
 b15zdnd11an1n04x5 FILLER_374_470 ();
 b15zdnd11an1n64x5 FILLER_374_477 ();
 b15zdnd11an1n32x5 FILLER_374_541 ();
 b15zdnd11an1n08x5 FILLER_374_573 ();
 b15zdnd11an1n64x5 FILLER_374_623 ();
 b15zdnd11an1n16x5 FILLER_374_687 ();
 b15zdnd11an1n08x5 FILLER_374_703 ();
 b15zdnd11an1n04x5 FILLER_374_711 ();
 b15zdnd00an1n02x5 FILLER_374_715 ();
 b15zdnd00an1n01x5 FILLER_374_717 ();
 b15zdnd11an1n64x5 FILLER_374_726 ();
 b15zdnd11an1n64x5 FILLER_374_790 ();
 b15zdnd11an1n64x5 FILLER_374_854 ();
 b15zdnd11an1n32x5 FILLER_374_918 ();
 b15zdnd11an1n16x5 FILLER_374_950 ();
 b15zdnd11an1n08x5 FILLER_374_966 ();
 b15zdnd00an1n02x5 FILLER_374_974 ();
 b15zdnd00an1n01x5 FILLER_374_976 ();
 b15zdnd11an1n64x5 FILLER_374_983 ();
 b15zdnd11an1n64x5 FILLER_374_1047 ();
 b15zdnd11an1n16x5 FILLER_374_1111 ();
 b15zdnd11an1n04x5 FILLER_374_1127 ();
 b15zdnd00an1n01x5 FILLER_374_1131 ();
 b15zdnd11an1n32x5 FILLER_374_1163 ();
 b15zdnd11an1n16x5 FILLER_374_1195 ();
 b15zdnd11an1n08x5 FILLER_374_1211 ();
 b15zdnd11an1n04x5 FILLER_374_1219 ();
 b15zdnd00an1n02x5 FILLER_374_1223 ();
 b15zdnd11an1n04x5 FILLER_374_1228 ();
 b15zdnd11an1n32x5 FILLER_374_1235 ();
 b15zdnd11an1n16x5 FILLER_374_1267 ();
 b15zdnd11an1n08x5 FILLER_374_1283 ();
 b15zdnd00an1n02x5 FILLER_374_1291 ();
 b15zdnd00an1n01x5 FILLER_374_1293 ();
 b15zdnd11an1n08x5 FILLER_374_1304 ();
 b15zdnd11an1n04x5 FILLER_374_1312 ();
 b15zdnd00an1n02x5 FILLER_374_1316 ();
 b15zdnd00an1n01x5 FILLER_374_1318 ();
 b15zdnd11an1n08x5 FILLER_374_1322 ();
 b15zdnd00an1n02x5 FILLER_374_1330 ();
 b15zdnd00an1n01x5 FILLER_374_1332 ();
 b15zdnd11an1n64x5 FILLER_374_1340 ();
 b15zdnd11an1n32x5 FILLER_374_1404 ();
 b15zdnd11an1n16x5 FILLER_374_1436 ();
 b15zdnd00an1n02x5 FILLER_374_1452 ();
 b15zdnd00an1n01x5 FILLER_374_1454 ();
 b15zdnd11an1n04x5 FILLER_374_1458 ();
 b15zdnd11an1n64x5 FILLER_374_1465 ();
 b15zdnd11an1n08x5 FILLER_374_1529 ();
 b15zdnd11an1n04x5 FILLER_374_1537 ();
 b15zdnd00an1n01x5 FILLER_374_1541 ();
 b15zdnd11an1n16x5 FILLER_374_1567 ();
 b15zdnd11an1n08x5 FILLER_374_1583 ();
 b15zdnd11an1n04x5 FILLER_374_1591 ();
 b15zdnd00an1n02x5 FILLER_374_1595 ();
 b15zdnd00an1n01x5 FILLER_374_1597 ();
 b15zdnd11an1n64x5 FILLER_374_1640 ();
 b15zdnd11an1n16x5 FILLER_374_1704 ();
 b15zdnd11an1n08x5 FILLER_374_1720 ();
 b15zdnd11an1n04x5 FILLER_374_1728 ();
 b15zdnd00an1n02x5 FILLER_374_1732 ();
 b15zdnd00an1n01x5 FILLER_374_1734 ();
 b15zdnd11an1n64x5 FILLER_374_1777 ();
 b15zdnd11an1n64x5 FILLER_374_1841 ();
 b15zdnd11an1n64x5 FILLER_374_1905 ();
 b15zdnd11an1n64x5 FILLER_374_1969 ();
 b15zdnd11an1n64x5 FILLER_374_2033 ();
 b15zdnd11an1n32x5 FILLER_374_2097 ();
 b15zdnd11an1n16x5 FILLER_374_2129 ();
 b15zdnd11an1n08x5 FILLER_374_2145 ();
 b15zdnd00an1n01x5 FILLER_374_2153 ();
 b15zdnd11an1n64x5 FILLER_374_2162 ();
 b15zdnd11an1n32x5 FILLER_374_2226 ();
 b15zdnd11an1n16x5 FILLER_374_2258 ();
 b15zdnd00an1n02x5 FILLER_374_2274 ();
 b15zdnd11an1n64x5 FILLER_375_0 ();
 b15zdnd11an1n64x5 FILLER_375_64 ();
 b15zdnd11an1n64x5 FILLER_375_128 ();
 b15zdnd11an1n64x5 FILLER_375_192 ();
 b15zdnd11an1n64x5 FILLER_375_256 ();
 b15zdnd11an1n64x5 FILLER_375_320 ();
 b15zdnd11an1n08x5 FILLER_375_384 ();
 b15zdnd00an1n02x5 FILLER_375_392 ();
 b15zdnd00an1n01x5 FILLER_375_394 ();
 b15zdnd11an1n04x5 FILLER_375_437 ();
 b15zdnd00an1n02x5 FILLER_375_441 ();
 b15zdnd11an1n64x5 FILLER_375_485 ();
 b15zdnd11an1n64x5 FILLER_375_549 ();
 b15zdnd11an1n64x5 FILLER_375_613 ();
 b15zdnd11an1n64x5 FILLER_375_677 ();
 b15zdnd11an1n64x5 FILLER_375_741 ();
 b15zdnd11an1n64x5 FILLER_375_805 ();
 b15zdnd11an1n64x5 FILLER_375_869 ();
 b15zdnd11an1n32x5 FILLER_375_933 ();
 b15zdnd11an1n08x5 FILLER_375_965 ();
 b15zdnd11an1n16x5 FILLER_375_1015 ();
 b15zdnd11an1n04x5 FILLER_375_1031 ();
 b15zdnd11an1n04x5 FILLER_375_1049 ();
 b15zdnd11an1n32x5 FILLER_375_1059 ();
 b15zdnd00an1n02x5 FILLER_375_1091 ();
 b15zdnd00an1n01x5 FILLER_375_1093 ();
 b15zdnd11an1n32x5 FILLER_375_1146 ();
 b15zdnd11an1n16x5 FILLER_375_1178 ();
 b15zdnd11an1n04x5 FILLER_375_1194 ();
 b15zdnd00an1n02x5 FILLER_375_1198 ();
 b15zdnd11an1n32x5 FILLER_375_1252 ();
 b15zdnd11an1n08x5 FILLER_375_1284 ();
 b15zdnd00an1n02x5 FILLER_375_1292 ();
 b15zdnd11an1n64x5 FILLER_375_1346 ();
 b15zdnd11an1n16x5 FILLER_375_1410 ();
 b15zdnd11an1n08x5 FILLER_375_1426 ();
 b15zdnd00an1n02x5 FILLER_375_1434 ();
 b15zdnd00an1n01x5 FILLER_375_1436 ();
 b15zdnd11an1n32x5 FILLER_375_1489 ();
 b15zdnd11an1n08x5 FILLER_375_1521 ();
 b15zdnd11an1n04x5 FILLER_375_1529 ();
 b15zdnd00an1n01x5 FILLER_375_1533 ();
 b15zdnd11an1n32x5 FILLER_375_1559 ();
 b15zdnd11an1n04x5 FILLER_375_1591 ();
 b15zdnd00an1n02x5 FILLER_375_1595 ();
 b15zdnd11an1n04x5 FILLER_375_1639 ();
 b15zdnd00an1n02x5 FILLER_375_1643 ();
 b15zdnd00an1n01x5 FILLER_375_1645 ();
 b15zdnd11an1n16x5 FILLER_375_1688 ();
 b15zdnd11an1n04x5 FILLER_375_1704 ();
 b15zdnd00an1n02x5 FILLER_375_1708 ();
 b15zdnd00an1n01x5 FILLER_375_1710 ();
 b15zdnd11an1n64x5 FILLER_375_1753 ();
 b15zdnd11an1n64x5 FILLER_375_1817 ();
 b15zdnd11an1n64x5 FILLER_375_1881 ();
 b15zdnd11an1n64x5 FILLER_375_1945 ();
 b15zdnd11an1n64x5 FILLER_375_2009 ();
 b15zdnd11an1n64x5 FILLER_375_2073 ();
 b15zdnd11an1n64x5 FILLER_375_2137 ();
 b15zdnd11an1n64x5 FILLER_375_2201 ();
 b15zdnd11an1n16x5 FILLER_375_2265 ();
 b15zdnd00an1n02x5 FILLER_375_2281 ();
 b15zdnd00an1n01x5 FILLER_375_2283 ();
 b15zdnd11an1n64x5 FILLER_376_8 ();
 b15zdnd11an1n64x5 FILLER_376_72 ();
 b15zdnd11an1n64x5 FILLER_376_136 ();
 b15zdnd11an1n64x5 FILLER_376_200 ();
 b15zdnd11an1n64x5 FILLER_376_264 ();
 b15zdnd11an1n64x5 FILLER_376_328 ();
 b15zdnd11an1n32x5 FILLER_376_392 ();
 b15zdnd11an1n08x5 FILLER_376_466 ();
 b15zdnd00an1n01x5 FILLER_376_474 ();
 b15zdnd11an1n64x5 FILLER_376_517 ();
 b15zdnd11an1n08x5 FILLER_376_581 ();
 b15zdnd11an1n04x5 FILLER_376_589 ();
 b15zdnd00an1n02x5 FILLER_376_593 ();
 b15zdnd00an1n01x5 FILLER_376_595 ();
 b15zdnd11an1n64x5 FILLER_376_638 ();
 b15zdnd11an1n16x5 FILLER_376_702 ();
 b15zdnd11an1n64x5 FILLER_376_726 ();
 b15zdnd11an1n64x5 FILLER_376_790 ();
 b15zdnd11an1n64x5 FILLER_376_854 ();
 b15zdnd11an1n64x5 FILLER_376_918 ();
 b15zdnd11an1n64x5 FILLER_376_982 ();
 b15zdnd11an1n32x5 FILLER_376_1046 ();
 b15zdnd11an1n16x5 FILLER_376_1078 ();
 b15zdnd11an1n04x5 FILLER_376_1094 ();
 b15zdnd00an1n02x5 FILLER_376_1098 ();
 b15zdnd11an1n64x5 FILLER_376_1142 ();
 b15zdnd11an1n08x5 FILLER_376_1206 ();
 b15zdnd11an1n04x5 FILLER_376_1214 ();
 b15zdnd00an1n01x5 FILLER_376_1218 ();
 b15zdnd11an1n04x5 FILLER_376_1222 ();
 b15zdnd11an1n04x5 FILLER_376_1246 ();
 b15zdnd00an1n01x5 FILLER_376_1250 ();
 b15zdnd11an1n16x5 FILLER_376_1277 ();
 b15zdnd11an1n08x5 FILLER_376_1293 ();
 b15zdnd00an1n02x5 FILLER_376_1301 ();
 b15zdnd11an1n04x5 FILLER_376_1306 ();
 b15zdnd11an1n64x5 FILLER_376_1352 ();
 b15zdnd11an1n32x5 FILLER_376_1416 ();
 b15zdnd11an1n08x5 FILLER_376_1448 ();
 b15zdnd11an1n04x5 FILLER_376_1456 ();
 b15zdnd00an1n02x5 FILLER_376_1460 ();
 b15zdnd11an1n64x5 FILLER_376_1465 ();
 b15zdnd11an1n64x5 FILLER_376_1529 ();
 b15zdnd11an1n64x5 FILLER_376_1593 ();
 b15zdnd11an1n64x5 FILLER_376_1657 ();
 b15zdnd11an1n64x5 FILLER_376_1721 ();
 b15zdnd11an1n64x5 FILLER_376_1785 ();
 b15zdnd11an1n64x5 FILLER_376_1849 ();
 b15zdnd11an1n64x5 FILLER_376_1913 ();
 b15zdnd11an1n64x5 FILLER_376_1977 ();
 b15zdnd11an1n64x5 FILLER_376_2041 ();
 b15zdnd11an1n32x5 FILLER_376_2105 ();
 b15zdnd11an1n16x5 FILLER_376_2137 ();
 b15zdnd00an1n01x5 FILLER_376_2153 ();
 b15zdnd11an1n64x5 FILLER_376_2162 ();
 b15zdnd11an1n32x5 FILLER_376_2226 ();
 b15zdnd11an1n16x5 FILLER_376_2258 ();
 b15zdnd00an1n02x5 FILLER_376_2274 ();
 b15zdnd11an1n64x5 FILLER_377_0 ();
 b15zdnd11an1n64x5 FILLER_377_64 ();
 b15zdnd11an1n64x5 FILLER_377_128 ();
 b15zdnd11an1n64x5 FILLER_377_192 ();
 b15zdnd11an1n64x5 FILLER_377_256 ();
 b15zdnd11an1n64x5 FILLER_377_320 ();
 b15zdnd11an1n32x5 FILLER_377_384 ();
 b15zdnd00an1n02x5 FILLER_377_416 ();
 b15zdnd00an1n01x5 FILLER_377_418 ();
 b15zdnd11an1n08x5 FILLER_377_461 ();
 b15zdnd11an1n64x5 FILLER_377_511 ();
 b15zdnd11an1n64x5 FILLER_377_575 ();
 b15zdnd11an1n64x5 FILLER_377_639 ();
 b15zdnd11an1n32x5 FILLER_377_703 ();
 b15zdnd11an1n16x5 FILLER_377_735 ();
 b15zdnd11an1n08x5 FILLER_377_751 ();
 b15zdnd00an1n02x5 FILLER_377_759 ();
 b15zdnd00an1n01x5 FILLER_377_761 ();
 b15zdnd11an1n64x5 FILLER_377_804 ();
 b15zdnd11an1n64x5 FILLER_377_868 ();
 b15zdnd11an1n64x5 FILLER_377_932 ();
 b15zdnd11an1n64x5 FILLER_377_996 ();
 b15zdnd11an1n32x5 FILLER_377_1060 ();
 b15zdnd11an1n08x5 FILLER_377_1092 ();
 b15zdnd00an1n02x5 FILLER_377_1100 ();
 b15zdnd00an1n01x5 FILLER_377_1102 ();
 b15zdnd11an1n04x5 FILLER_377_1110 ();
 b15zdnd11an1n04x5 FILLER_377_1117 ();
 b15zdnd11an1n04x5 FILLER_377_1124 ();
 b15zdnd11an1n16x5 FILLER_377_1131 ();
 b15zdnd00an1n02x5 FILLER_377_1147 ();
 b15zdnd00an1n01x5 FILLER_377_1149 ();
 b15zdnd11an1n64x5 FILLER_377_1175 ();
 b15zdnd11an1n32x5 FILLER_377_1239 ();
 b15zdnd11an1n16x5 FILLER_377_1271 ();
 b15zdnd11an1n08x5 FILLER_377_1287 ();
 b15zdnd11an1n04x5 FILLER_377_1295 ();
 b15zdnd00an1n02x5 FILLER_377_1299 ();
 b15zdnd11an1n64x5 FILLER_377_1343 ();
 b15zdnd11an1n64x5 FILLER_377_1407 ();
 b15zdnd11an1n08x5 FILLER_377_1471 ();
 b15zdnd00an1n02x5 FILLER_377_1479 ();
 b15zdnd00an1n01x5 FILLER_377_1481 ();
 b15zdnd11an1n64x5 FILLER_377_1513 ();
 b15zdnd11an1n64x5 FILLER_377_1577 ();
 b15zdnd11an1n64x5 FILLER_377_1641 ();
 b15zdnd11an1n64x5 FILLER_377_1705 ();
 b15zdnd11an1n64x5 FILLER_377_1769 ();
 b15zdnd11an1n64x5 FILLER_377_1833 ();
 b15zdnd11an1n64x5 FILLER_377_1897 ();
 b15zdnd11an1n64x5 FILLER_377_1961 ();
 b15zdnd11an1n64x5 FILLER_377_2025 ();
 b15zdnd11an1n64x5 FILLER_377_2089 ();
 b15zdnd11an1n64x5 FILLER_377_2153 ();
 b15zdnd11an1n64x5 FILLER_377_2217 ();
 b15zdnd00an1n02x5 FILLER_377_2281 ();
 b15zdnd00an1n01x5 FILLER_377_2283 ();
 b15zdnd11an1n64x5 FILLER_378_8 ();
 b15zdnd11an1n64x5 FILLER_378_72 ();
 b15zdnd11an1n64x5 FILLER_378_136 ();
 b15zdnd11an1n64x5 FILLER_378_200 ();
 b15zdnd11an1n64x5 FILLER_378_264 ();
 b15zdnd11an1n64x5 FILLER_378_328 ();
 b15zdnd11an1n16x5 FILLER_378_392 ();
 b15zdnd11an1n04x5 FILLER_378_408 ();
 b15zdnd00an1n02x5 FILLER_378_412 ();
 b15zdnd00an1n01x5 FILLER_378_414 ();
 b15zdnd11an1n04x5 FILLER_378_457 ();
 b15zdnd11an1n64x5 FILLER_378_503 ();
 b15zdnd11an1n16x5 FILLER_378_567 ();
 b15zdnd11an1n04x5 FILLER_378_583 ();
 b15zdnd00an1n01x5 FILLER_378_587 ();
 b15zdnd11an1n64x5 FILLER_378_630 ();
 b15zdnd00an1n02x5 FILLER_378_694 ();
 b15zdnd00an1n01x5 FILLER_378_696 ();
 b15zdnd11an1n08x5 FILLER_378_703 ();
 b15zdnd11an1n04x5 FILLER_378_711 ();
 b15zdnd00an1n02x5 FILLER_378_715 ();
 b15zdnd00an1n01x5 FILLER_378_717 ();
 b15zdnd11an1n32x5 FILLER_378_726 ();
 b15zdnd11an1n16x5 FILLER_378_758 ();
 b15zdnd11an1n08x5 FILLER_378_774 ();
 b15zdnd11an1n04x5 FILLER_378_782 ();
 b15zdnd00an1n02x5 FILLER_378_786 ();
 b15zdnd00an1n01x5 FILLER_378_788 ();
 b15zdnd11an1n32x5 FILLER_378_831 ();
 b15zdnd11an1n16x5 FILLER_378_863 ();
 b15zdnd11an1n08x5 FILLER_378_879 ();
 b15zdnd11an1n04x5 FILLER_378_887 ();
 b15zdnd00an1n02x5 FILLER_378_891 ();
 b15zdnd00an1n01x5 FILLER_378_893 ();
 b15zdnd11an1n64x5 FILLER_378_899 ();
 b15zdnd11an1n64x5 FILLER_378_963 ();
 b15zdnd11an1n64x5 FILLER_378_1027 ();
 b15zdnd11an1n32x5 FILLER_378_1091 ();
 b15zdnd11an1n04x5 FILLER_378_1123 ();
 b15zdnd00an1n02x5 FILLER_378_1127 ();
 b15zdnd11an1n04x5 FILLER_378_1134 ();
 b15zdnd11an1n08x5 FILLER_378_1141 ();
 b15zdnd11an1n04x5 FILLER_378_1149 ();
 b15zdnd00an1n02x5 FILLER_378_1153 ();
 b15zdnd11an1n64x5 FILLER_378_1197 ();
 b15zdnd11an1n32x5 FILLER_378_1261 ();
 b15zdnd11an1n16x5 FILLER_378_1293 ();
 b15zdnd11an1n08x5 FILLER_378_1309 ();
 b15zdnd00an1n02x5 FILLER_378_1317 ();
 b15zdnd11an1n64x5 FILLER_378_1322 ();
 b15zdnd11an1n32x5 FILLER_378_1386 ();
 b15zdnd11an1n16x5 FILLER_378_1418 ();
 b15zdnd11an1n08x5 FILLER_378_1434 ();
 b15zdnd11an1n04x5 FILLER_378_1442 ();
 b15zdnd11an1n32x5 FILLER_378_1466 ();
 b15zdnd11an1n16x5 FILLER_378_1498 ();
 b15zdnd00an1n01x5 FILLER_378_1514 ();
 b15zdnd11an1n08x5 FILLER_378_1557 ();
 b15zdnd00an1n01x5 FILLER_378_1565 ();
 b15zdnd11an1n04x5 FILLER_378_1578 ();
 b15zdnd11an1n08x5 FILLER_378_1587 ();
 b15zdnd11an1n04x5 FILLER_378_1595 ();
 b15zdnd00an1n02x5 FILLER_378_1599 ();
 b15zdnd00an1n01x5 FILLER_378_1601 ();
 b15zdnd11an1n64x5 FILLER_378_1644 ();
 b15zdnd11an1n64x5 FILLER_378_1708 ();
 b15zdnd11an1n64x5 FILLER_378_1772 ();
 b15zdnd11an1n64x5 FILLER_378_1836 ();
 b15zdnd11an1n64x5 FILLER_378_1900 ();
 b15zdnd11an1n64x5 FILLER_378_1964 ();
 b15zdnd11an1n64x5 FILLER_378_2028 ();
 b15zdnd11an1n32x5 FILLER_378_2092 ();
 b15zdnd11an1n16x5 FILLER_378_2124 ();
 b15zdnd11an1n08x5 FILLER_378_2140 ();
 b15zdnd11an1n04x5 FILLER_378_2148 ();
 b15zdnd00an1n02x5 FILLER_378_2152 ();
 b15zdnd11an1n64x5 FILLER_378_2162 ();
 b15zdnd11an1n32x5 FILLER_378_2226 ();
 b15zdnd11an1n16x5 FILLER_378_2258 ();
 b15zdnd00an1n02x5 FILLER_378_2274 ();
 b15zdnd11an1n64x5 FILLER_379_0 ();
 b15zdnd11an1n64x5 FILLER_379_64 ();
 b15zdnd11an1n64x5 FILLER_379_128 ();
 b15zdnd11an1n64x5 FILLER_379_192 ();
 b15zdnd11an1n64x5 FILLER_379_256 ();
 b15zdnd11an1n64x5 FILLER_379_320 ();
 b15zdnd00an1n02x5 FILLER_379_384 ();
 b15zdnd00an1n01x5 FILLER_379_386 ();
 b15zdnd11an1n04x5 FILLER_379_429 ();
 b15zdnd00an1n02x5 FILLER_379_433 ();
 b15zdnd11an1n64x5 FILLER_379_477 ();
 b15zdnd11an1n32x5 FILLER_379_541 ();
 b15zdnd11an1n08x5 FILLER_379_573 ();
 b15zdnd11an1n04x5 FILLER_379_596 ();
 b15zdnd00an1n01x5 FILLER_379_600 ();
 b15zdnd11an1n04x5 FILLER_379_611 ();
 b15zdnd11an1n64x5 FILLER_379_657 ();
 b15zdnd11an1n32x5 FILLER_379_721 ();
 b15zdnd11an1n08x5 FILLER_379_753 ();
 b15zdnd11an1n04x5 FILLER_379_761 ();
 b15zdnd00an1n02x5 FILLER_379_765 ();
 b15zdnd11an1n64x5 FILLER_379_772 ();
 b15zdnd11an1n32x5 FILLER_379_836 ();
 b15zdnd00an1n02x5 FILLER_379_868 ();
 b15zdnd11an1n08x5 FILLER_379_912 ();
 b15zdnd11an1n04x5 FILLER_379_920 ();
 b15zdnd00an1n02x5 FILLER_379_924 ();
 b15zdnd00an1n01x5 FILLER_379_926 ();
 b15zdnd11an1n16x5 FILLER_379_931 ();
 b15zdnd11an1n04x5 FILLER_379_959 ();
 b15zdnd00an1n02x5 FILLER_379_963 ();
 b15zdnd11an1n32x5 FILLER_379_980 ();
 b15zdnd11an1n16x5 FILLER_379_1012 ();
 b15zdnd11an1n08x5 FILLER_379_1028 ();
 b15zdnd11an1n04x5 FILLER_379_1036 ();
 b15zdnd00an1n01x5 FILLER_379_1040 ();
 b15zdnd11an1n04x5 FILLER_379_1051 ();
 b15zdnd00an1n02x5 FILLER_379_1055 ();
 b15zdnd00an1n01x5 FILLER_379_1057 ();
 b15zdnd11an1n32x5 FILLER_379_1061 ();
 b15zdnd11an1n16x5 FILLER_379_1093 ();
 b15zdnd11an1n08x5 FILLER_379_1109 ();
 b15zdnd11an1n04x5 FILLER_379_1117 ();
 b15zdnd00an1n01x5 FILLER_379_1121 ();
 b15zdnd11an1n08x5 FILLER_379_1153 ();
 b15zdnd11an1n04x5 FILLER_379_1161 ();
 b15zdnd00an1n01x5 FILLER_379_1165 ();
 b15zdnd11an1n08x5 FILLER_379_1172 ();
 b15zdnd00an1n02x5 FILLER_379_1180 ();
 b15zdnd11an1n32x5 FILLER_379_1224 ();
 b15zdnd00an1n02x5 FILLER_379_1256 ();
 b15zdnd00an1n01x5 FILLER_379_1258 ();
 b15zdnd11an1n08x5 FILLER_379_1301 ();
 b15zdnd11an1n04x5 FILLER_379_1309 ();
 b15zdnd00an1n02x5 FILLER_379_1313 ();
 b15zdnd00an1n01x5 FILLER_379_1315 ();
 b15zdnd11an1n04x5 FILLER_379_1358 ();
 b15zdnd11an1n32x5 FILLER_379_1404 ();
 b15zdnd11an1n04x5 FILLER_379_1436 ();
 b15zdnd00an1n01x5 FILLER_379_1440 ();
 b15zdnd11an1n08x5 FILLER_379_1483 ();
 b15zdnd11an1n32x5 FILLER_379_1533 ();
 b15zdnd11an1n04x5 FILLER_379_1607 ();
 b15zdnd11an1n64x5 FILLER_379_1653 ();
 b15zdnd11an1n64x5 FILLER_379_1717 ();
 b15zdnd11an1n64x5 FILLER_379_1781 ();
 b15zdnd11an1n64x5 FILLER_379_1845 ();
 b15zdnd11an1n64x5 FILLER_379_1909 ();
 b15zdnd11an1n64x5 FILLER_379_1973 ();
 b15zdnd11an1n64x5 FILLER_379_2037 ();
 b15zdnd11an1n64x5 FILLER_379_2101 ();
 b15zdnd11an1n64x5 FILLER_379_2165 ();
 b15zdnd11an1n32x5 FILLER_379_2229 ();
 b15zdnd11an1n16x5 FILLER_379_2261 ();
 b15zdnd11an1n04x5 FILLER_379_2277 ();
 b15zdnd00an1n02x5 FILLER_379_2281 ();
 b15zdnd00an1n01x5 FILLER_379_2283 ();
 b15zdnd11an1n64x5 FILLER_380_8 ();
 b15zdnd11an1n64x5 FILLER_380_72 ();
 b15zdnd11an1n64x5 FILLER_380_136 ();
 b15zdnd11an1n64x5 FILLER_380_200 ();
 b15zdnd11an1n64x5 FILLER_380_264 ();
 b15zdnd11an1n64x5 FILLER_380_328 ();
 b15zdnd11an1n16x5 FILLER_380_392 ();
 b15zdnd11an1n08x5 FILLER_380_408 ();
 b15zdnd11an1n08x5 FILLER_380_458 ();
 b15zdnd11an1n04x5 FILLER_380_466 ();
 b15zdnd00an1n02x5 FILLER_380_470 ();
 b15zdnd11an1n32x5 FILLER_380_514 ();
 b15zdnd11an1n16x5 FILLER_380_546 ();
 b15zdnd11an1n08x5 FILLER_380_577 ();
 b15zdnd00an1n01x5 FILLER_380_585 ();
 b15zdnd11an1n04x5 FILLER_380_628 ();
 b15zdnd11an1n04x5 FILLER_380_638 ();
 b15zdnd11an1n08x5 FILLER_380_645 ();
 b15zdnd11an1n04x5 FILLER_380_653 ();
 b15zdnd00an1n02x5 FILLER_380_657 ();
 b15zdnd11an1n32x5 FILLER_380_669 ();
 b15zdnd11an1n16x5 FILLER_380_701 ();
 b15zdnd00an1n01x5 FILLER_380_717 ();
 b15zdnd11an1n32x5 FILLER_380_726 ();
 b15zdnd11an1n04x5 FILLER_380_758 ();
 b15zdnd00an1n02x5 FILLER_380_762 ();
 b15zdnd11an1n64x5 FILLER_380_771 ();
 b15zdnd11an1n32x5 FILLER_380_835 ();
 b15zdnd11an1n08x5 FILLER_380_867 ();
 b15zdnd00an1n02x5 FILLER_380_875 ();
 b15zdnd11an1n04x5 FILLER_380_881 ();
 b15zdnd11an1n04x5 FILLER_380_890 ();
 b15zdnd11an1n16x5 FILLER_380_904 ();
 b15zdnd11an1n04x5 FILLER_380_920 ();
 b15zdnd11an1n04x5 FILLER_380_931 ();
 b15zdnd11an1n04x5 FILLER_380_944 ();
 b15zdnd11an1n16x5 FILLER_380_958 ();
 b15zdnd00an1n01x5 FILLER_380_974 ();
 b15zdnd11an1n16x5 FILLER_380_978 ();
 b15zdnd11an1n08x5 FILLER_380_994 ();
 b15zdnd11an1n04x5 FILLER_380_1002 ();
 b15zdnd00an1n01x5 FILLER_380_1006 ();
 b15zdnd11an1n64x5 FILLER_380_1015 ();
 b15zdnd00an1n02x5 FILLER_380_1079 ();
 b15zdnd11an1n16x5 FILLER_380_1096 ();
 b15zdnd11an1n04x5 FILLER_380_1112 ();
 b15zdnd00an1n02x5 FILLER_380_1116 ();
 b15zdnd00an1n01x5 FILLER_380_1118 ();
 b15zdnd11an1n04x5 FILLER_380_1136 ();
 b15zdnd00an1n02x5 FILLER_380_1140 ();
 b15zdnd00an1n01x5 FILLER_380_1142 ();
 b15zdnd11an1n04x5 FILLER_380_1160 ();
 b15zdnd11an1n04x5 FILLER_380_1195 ();
 b15zdnd11an1n16x5 FILLER_380_1230 ();
 b15zdnd00an1n02x5 FILLER_380_1246 ();
 b15zdnd11an1n04x5 FILLER_380_1272 ();
 b15zdnd11an1n16x5 FILLER_380_1288 ();
 b15zdnd00an1n01x5 FILLER_380_1304 ();
 b15zdnd11an1n08x5 FILLER_380_1320 ();
 b15zdnd11an1n04x5 FILLER_380_1328 ();
 b15zdnd00an1n01x5 FILLER_380_1332 ();
 b15zdnd11an1n32x5 FILLER_380_1337 ();
 b15zdnd11an1n04x5 FILLER_380_1389 ();
 b15zdnd11an1n08x5 FILLER_380_1398 ();
 b15zdnd11an1n04x5 FILLER_380_1406 ();
 b15zdnd00an1n02x5 FILLER_380_1410 ();
 b15zdnd00an1n01x5 FILLER_380_1412 ();
 b15zdnd11an1n04x5 FILLER_380_1430 ();
 b15zdnd11an1n04x5 FILLER_380_1438 ();
 b15zdnd00an1n02x5 FILLER_380_1442 ();
 b15zdnd00an1n01x5 FILLER_380_1444 ();
 b15zdnd11an1n04x5 FILLER_380_1487 ();
 b15zdnd11an1n04x5 FILLER_380_1522 ();
 b15zdnd11an1n32x5 FILLER_380_1532 ();
 b15zdnd11an1n16x5 FILLER_380_1564 ();
 b15zdnd11an1n04x5 FILLER_380_1580 ();
 b15zdnd11an1n08x5 FILLER_380_1629 ();
 b15zdnd11an1n04x5 FILLER_380_1637 ();
 b15zdnd00an1n02x5 FILLER_380_1641 ();
 b15zdnd11an1n64x5 FILLER_380_1685 ();
 b15zdnd11an1n64x5 FILLER_380_1749 ();
 b15zdnd11an1n64x5 FILLER_380_1813 ();
 b15zdnd11an1n64x5 FILLER_380_1877 ();
 b15zdnd11an1n64x5 FILLER_380_1941 ();
 b15zdnd11an1n64x5 FILLER_380_2005 ();
 b15zdnd11an1n64x5 FILLER_380_2069 ();
 b15zdnd11an1n16x5 FILLER_380_2133 ();
 b15zdnd11an1n04x5 FILLER_380_2149 ();
 b15zdnd00an1n01x5 FILLER_380_2153 ();
 b15zdnd11an1n64x5 FILLER_380_2162 ();
 b15zdnd11an1n32x5 FILLER_380_2226 ();
 b15zdnd11an1n16x5 FILLER_380_2258 ();
 b15zdnd00an1n02x5 FILLER_380_2274 ();
 b15zdnd11an1n64x5 FILLER_381_0 ();
 b15zdnd11an1n64x5 FILLER_381_64 ();
 b15zdnd11an1n64x5 FILLER_381_128 ();
 b15zdnd11an1n64x5 FILLER_381_192 ();
 b15zdnd11an1n64x5 FILLER_381_256 ();
 b15zdnd11an1n64x5 FILLER_381_320 ();
 b15zdnd11an1n16x5 FILLER_381_384 ();
 b15zdnd11an1n08x5 FILLER_381_400 ();
 b15zdnd11an1n04x5 FILLER_381_408 ();
 b15zdnd11an1n04x5 FILLER_381_454 ();
 b15zdnd11an1n32x5 FILLER_381_500 ();
 b15zdnd11an1n16x5 FILLER_381_532 ();
 b15zdnd11an1n16x5 FILLER_381_553 ();
 b15zdnd11an1n08x5 FILLER_381_569 ();
 b15zdnd00an1n02x5 FILLER_381_577 ();
 b15zdnd11an1n04x5 FILLER_381_589 ();
 b15zdnd11an1n04x5 FILLER_381_635 ();
 b15zdnd00an1n01x5 FILLER_381_639 ();
 b15zdnd11an1n04x5 FILLER_381_644 ();
 b15zdnd00an1n02x5 FILLER_381_648 ();
 b15zdnd00an1n01x5 FILLER_381_650 ();
 b15zdnd11an1n32x5 FILLER_381_654 ();
 b15zdnd11an1n04x5 FILLER_381_686 ();
 b15zdnd00an1n01x5 FILLER_381_690 ();
 b15zdnd11an1n04x5 FILLER_381_733 ();
 b15zdnd00an1n02x5 FILLER_381_737 ();
 b15zdnd11an1n64x5 FILLER_381_781 ();
 b15zdnd11an1n64x5 FILLER_381_845 ();
 b15zdnd11an1n32x5 FILLER_381_909 ();
 b15zdnd11an1n16x5 FILLER_381_941 ();
 b15zdnd11an1n04x5 FILLER_381_957 ();
 b15zdnd00an1n02x5 FILLER_381_961 ();
 b15zdnd00an1n01x5 FILLER_381_963 ();
 b15zdnd11an1n64x5 FILLER_381_970 ();
 b15zdnd11an1n64x5 FILLER_381_1034 ();
 b15zdnd11an1n16x5 FILLER_381_1098 ();
 b15zdnd11an1n08x5 FILLER_381_1114 ();
 b15zdnd11an1n04x5 FILLER_381_1122 ();
 b15zdnd00an1n01x5 FILLER_381_1126 ();
 b15zdnd11an1n04x5 FILLER_381_1169 ();
 b15zdnd11an1n08x5 FILLER_381_1180 ();
 b15zdnd11an1n04x5 FILLER_381_1188 ();
 b15zdnd00an1n02x5 FILLER_381_1192 ();
 b15zdnd00an1n01x5 FILLER_381_1194 ();
 b15zdnd11an1n64x5 FILLER_381_1201 ();
 b15zdnd11an1n32x5 FILLER_381_1265 ();
 b15zdnd11an1n04x5 FILLER_381_1297 ();
 b15zdnd00an1n01x5 FILLER_381_1301 ();
 b15zdnd11an1n64x5 FILLER_381_1307 ();
 b15zdnd11an1n08x5 FILLER_381_1371 ();
 b15zdnd00an1n02x5 FILLER_381_1379 ();
 b15zdnd00an1n01x5 FILLER_381_1381 ();
 b15zdnd11an1n16x5 FILLER_381_1402 ();
 b15zdnd11an1n04x5 FILLER_381_1418 ();
 b15zdnd00an1n02x5 FILLER_381_1422 ();
 b15zdnd00an1n01x5 FILLER_381_1424 ();
 b15zdnd11an1n04x5 FILLER_381_1429 ();
 b15zdnd00an1n02x5 FILLER_381_1433 ();
 b15zdnd11an1n04x5 FILLER_381_1459 ();
 b15zdnd11an1n04x5 FILLER_381_1483 ();
 b15zdnd11an1n04x5 FILLER_381_1491 ();
 b15zdnd11an1n16x5 FILLER_381_1499 ();
 b15zdnd11an1n08x5 FILLER_381_1515 ();
 b15zdnd00an1n02x5 FILLER_381_1523 ();
 b15zdnd11an1n04x5 FILLER_381_1532 ();
 b15zdnd11an1n08x5 FILLER_381_1553 ();
 b15zdnd11an1n04x5 FILLER_381_1561 ();
 b15zdnd11an1n08x5 FILLER_381_1569 ();
 b15zdnd11an1n04x5 FILLER_381_1582 ();
 b15zdnd00an1n01x5 FILLER_381_1586 ();
 b15zdnd11an1n04x5 FILLER_381_1629 ();
 b15zdnd11an1n64x5 FILLER_381_1639 ();
 b15zdnd11an1n64x5 FILLER_381_1703 ();
 b15zdnd11an1n64x5 FILLER_381_1767 ();
 b15zdnd11an1n64x5 FILLER_381_1831 ();
 b15zdnd11an1n64x5 FILLER_381_1895 ();
 b15zdnd11an1n64x5 FILLER_381_1959 ();
 b15zdnd11an1n64x5 FILLER_381_2023 ();
 b15zdnd11an1n64x5 FILLER_381_2087 ();
 b15zdnd11an1n64x5 FILLER_381_2151 ();
 b15zdnd11an1n64x5 FILLER_381_2215 ();
 b15zdnd11an1n04x5 FILLER_381_2279 ();
 b15zdnd00an1n01x5 FILLER_381_2283 ();
 b15zdnd11an1n64x5 FILLER_382_8 ();
 b15zdnd11an1n64x5 FILLER_382_72 ();
 b15zdnd11an1n64x5 FILLER_382_136 ();
 b15zdnd11an1n64x5 FILLER_382_200 ();
 b15zdnd11an1n64x5 FILLER_382_264 ();
 b15zdnd11an1n64x5 FILLER_382_328 ();
 b15zdnd11an1n08x5 FILLER_382_392 ();
 b15zdnd11an1n04x5 FILLER_382_400 ();
 b15zdnd00an1n01x5 FILLER_382_404 ();
 b15zdnd11an1n08x5 FILLER_382_447 ();
 b15zdnd11an1n04x5 FILLER_382_455 ();
 b15zdnd11an1n64x5 FILLER_382_501 ();
 b15zdnd11an1n16x5 FILLER_382_565 ();
 b15zdnd11an1n04x5 FILLER_382_581 ();
 b15zdnd11an1n64x5 FILLER_382_627 ();
 b15zdnd11an1n16x5 FILLER_382_691 ();
 b15zdnd11an1n08x5 FILLER_382_707 ();
 b15zdnd00an1n02x5 FILLER_382_715 ();
 b15zdnd00an1n01x5 FILLER_382_717 ();
 b15zdnd11an1n64x5 FILLER_382_726 ();
 b15zdnd11an1n64x5 FILLER_382_790 ();
 b15zdnd11an1n64x5 FILLER_382_854 ();
 b15zdnd11an1n64x5 FILLER_382_918 ();
 b15zdnd11an1n64x5 FILLER_382_982 ();
 b15zdnd11an1n16x5 FILLER_382_1046 ();
 b15zdnd11an1n08x5 FILLER_382_1062 ();
 b15zdnd00an1n01x5 FILLER_382_1070 ();
 b15zdnd11an1n32x5 FILLER_382_1091 ();
 b15zdnd11an1n08x5 FILLER_382_1123 ();
 b15zdnd00an1n01x5 FILLER_382_1131 ();
 b15zdnd11an1n04x5 FILLER_382_1156 ();
 b15zdnd11an1n64x5 FILLER_382_1202 ();
 b15zdnd11an1n16x5 FILLER_382_1308 ();
 b15zdnd11an1n08x5 FILLER_382_1324 ();
 b15zdnd00an1n02x5 FILLER_382_1332 ();
 b15zdnd11an1n04x5 FILLER_382_1376 ();
 b15zdnd11an1n16x5 FILLER_382_1422 ();
 b15zdnd11an1n04x5 FILLER_382_1438 ();
 b15zdnd11an1n08x5 FILLER_382_1484 ();
 b15zdnd00an1n01x5 FILLER_382_1492 ();
 b15zdnd11an1n64x5 FILLER_382_1535 ();
 b15zdnd11an1n64x5 FILLER_382_1599 ();
 b15zdnd11an1n64x5 FILLER_382_1663 ();
 b15zdnd11an1n64x5 FILLER_382_1727 ();
 b15zdnd11an1n64x5 FILLER_382_1791 ();
 b15zdnd11an1n64x5 FILLER_382_1855 ();
 b15zdnd11an1n64x5 FILLER_382_1919 ();
 b15zdnd11an1n64x5 FILLER_382_1983 ();
 b15zdnd11an1n64x5 FILLER_382_2047 ();
 b15zdnd11an1n32x5 FILLER_382_2111 ();
 b15zdnd11an1n08x5 FILLER_382_2143 ();
 b15zdnd00an1n02x5 FILLER_382_2151 ();
 b15zdnd00an1n01x5 FILLER_382_2153 ();
 b15zdnd11an1n64x5 FILLER_382_2162 ();
 b15zdnd11an1n32x5 FILLER_382_2226 ();
 b15zdnd11an1n16x5 FILLER_382_2258 ();
 b15zdnd00an1n02x5 FILLER_382_2274 ();
 b15zdnd11an1n64x5 FILLER_383_0 ();
 b15zdnd11an1n64x5 FILLER_383_64 ();
 b15zdnd11an1n64x5 FILLER_383_128 ();
 b15zdnd11an1n64x5 FILLER_383_192 ();
 b15zdnd11an1n64x5 FILLER_383_256 ();
 b15zdnd11an1n64x5 FILLER_383_320 ();
 b15zdnd11an1n64x5 FILLER_383_384 ();
 b15zdnd11an1n64x5 FILLER_383_448 ();
 b15zdnd11an1n64x5 FILLER_383_512 ();
 b15zdnd11an1n16x5 FILLER_383_576 ();
 b15zdnd00an1n02x5 FILLER_383_592 ();
 b15zdnd11an1n04x5 FILLER_383_600 ();
 b15zdnd00an1n01x5 FILLER_383_604 ();
 b15zdnd11an1n04x5 FILLER_383_620 ();
 b15zdnd11an1n64x5 FILLER_383_630 ();
 b15zdnd11an1n64x5 FILLER_383_694 ();
 b15zdnd11an1n64x5 FILLER_383_758 ();
 b15zdnd11an1n64x5 FILLER_383_822 ();
 b15zdnd11an1n64x5 FILLER_383_886 ();
 b15zdnd11an1n64x5 FILLER_383_950 ();
 b15zdnd11an1n64x5 FILLER_383_1014 ();
 b15zdnd11an1n64x5 FILLER_383_1078 ();
 b15zdnd11an1n64x5 FILLER_383_1142 ();
 b15zdnd11an1n64x5 FILLER_383_1206 ();
 b15zdnd11an1n64x5 FILLER_383_1270 ();
 b15zdnd11an1n64x5 FILLER_383_1334 ();
 b15zdnd11an1n64x5 FILLER_383_1398 ();
 b15zdnd11an1n04x5 FILLER_383_1462 ();
 b15zdnd00an1n02x5 FILLER_383_1466 ();
 b15zdnd00an1n01x5 FILLER_383_1468 ();
 b15zdnd11an1n64x5 FILLER_383_1489 ();
 b15zdnd11an1n64x5 FILLER_383_1553 ();
 b15zdnd11an1n64x5 FILLER_383_1617 ();
 b15zdnd11an1n64x5 FILLER_383_1681 ();
 b15zdnd11an1n64x5 FILLER_383_1745 ();
 b15zdnd11an1n64x5 FILLER_383_1809 ();
 b15zdnd11an1n64x5 FILLER_383_1873 ();
 b15zdnd11an1n64x5 FILLER_383_1937 ();
 b15zdnd11an1n64x5 FILLER_383_2001 ();
 b15zdnd11an1n64x5 FILLER_383_2065 ();
 b15zdnd11an1n64x5 FILLER_383_2129 ();
 b15zdnd11an1n64x5 FILLER_383_2193 ();
 b15zdnd11an1n16x5 FILLER_383_2257 ();
 b15zdnd11an1n08x5 FILLER_383_2273 ();
 b15zdnd00an1n02x5 FILLER_383_2281 ();
 b15zdnd00an1n01x5 FILLER_383_2283 ();
 b15zdnd11an1n64x5 FILLER_384_8 ();
 b15zdnd11an1n64x5 FILLER_384_72 ();
 b15zdnd11an1n64x5 FILLER_384_136 ();
 b15zdnd11an1n64x5 FILLER_384_200 ();
 b15zdnd11an1n64x5 FILLER_384_264 ();
 b15zdnd11an1n64x5 FILLER_384_328 ();
 b15zdnd11an1n64x5 FILLER_384_392 ();
 b15zdnd11an1n64x5 FILLER_384_456 ();
 b15zdnd11an1n64x5 FILLER_384_520 ();
 b15zdnd11an1n16x5 FILLER_384_584 ();
 b15zdnd11an1n04x5 FILLER_384_600 ();
 b15zdnd00an1n02x5 FILLER_384_604 ();
 b15zdnd00an1n01x5 FILLER_384_606 ();
 b15zdnd11an1n64x5 FILLER_384_649 ();
 b15zdnd11an1n04x5 FILLER_384_713 ();
 b15zdnd00an1n01x5 FILLER_384_717 ();
 b15zdnd11an1n64x5 FILLER_384_726 ();
 b15zdnd11an1n64x5 FILLER_384_790 ();
 b15zdnd11an1n64x5 FILLER_384_854 ();
 b15zdnd11an1n64x5 FILLER_384_918 ();
 b15zdnd11an1n32x5 FILLER_384_982 ();
 b15zdnd11an1n16x5 FILLER_384_1014 ();
 b15zdnd11an1n08x5 FILLER_384_1030 ();
 b15zdnd00an1n02x5 FILLER_384_1038 ();
 b15zdnd00an1n01x5 FILLER_384_1040 ();
 b15zdnd11an1n64x5 FILLER_384_1083 ();
 b15zdnd11an1n64x5 FILLER_384_1147 ();
 b15zdnd11an1n64x5 FILLER_384_1211 ();
 b15zdnd11an1n64x5 FILLER_384_1275 ();
 b15zdnd11an1n64x5 FILLER_384_1339 ();
 b15zdnd11an1n64x5 FILLER_384_1403 ();
 b15zdnd11an1n64x5 FILLER_384_1467 ();
 b15zdnd11an1n64x5 FILLER_384_1531 ();
 b15zdnd11an1n64x5 FILLER_384_1595 ();
 b15zdnd11an1n64x5 FILLER_384_1659 ();
 b15zdnd11an1n64x5 FILLER_384_1723 ();
 b15zdnd11an1n64x5 FILLER_384_1787 ();
 b15zdnd11an1n64x5 FILLER_384_1851 ();
 b15zdnd11an1n64x5 FILLER_384_1915 ();
 b15zdnd11an1n64x5 FILLER_384_1979 ();
 b15zdnd11an1n64x5 FILLER_384_2043 ();
 b15zdnd11an1n32x5 FILLER_384_2107 ();
 b15zdnd11an1n08x5 FILLER_384_2139 ();
 b15zdnd11an1n04x5 FILLER_384_2147 ();
 b15zdnd00an1n02x5 FILLER_384_2151 ();
 b15zdnd00an1n01x5 FILLER_384_2153 ();
 b15zdnd11an1n64x5 FILLER_384_2162 ();
 b15zdnd11an1n32x5 FILLER_384_2226 ();
 b15zdnd11an1n16x5 FILLER_384_2258 ();
 b15zdnd00an1n02x5 FILLER_384_2274 ();
 b15zdnd11an1n64x5 FILLER_385_0 ();
 b15zdnd11an1n64x5 FILLER_385_64 ();
 b15zdnd11an1n64x5 FILLER_385_128 ();
 b15zdnd11an1n64x5 FILLER_385_192 ();
 b15zdnd11an1n64x5 FILLER_385_256 ();
 b15zdnd11an1n64x5 FILLER_385_320 ();
 b15zdnd11an1n16x5 FILLER_385_384 ();
 b15zdnd00an1n02x5 FILLER_385_400 ();
 b15zdnd11an1n04x5 FILLER_385_406 ();
 b15zdnd11an1n04x5 FILLER_385_414 ();
 b15zdnd11an1n04x5 FILLER_385_422 ();
 b15zdnd11an1n04x5 FILLER_385_430 ();
 b15zdnd00an1n01x5 FILLER_385_434 ();
 b15zdnd11an1n04x5 FILLER_385_439 ();
 b15zdnd11an1n64x5 FILLER_385_447 ();
 b15zdnd11an1n64x5 FILLER_385_511 ();
 b15zdnd11an1n32x5 FILLER_385_575 ();
 b15zdnd11an1n08x5 FILLER_385_607 ();
 b15zdnd11an1n04x5 FILLER_385_615 ();
 b15zdnd00an1n02x5 FILLER_385_619 ();
 b15zdnd11an1n64x5 FILLER_385_663 ();
 b15zdnd11an1n64x5 FILLER_385_727 ();
 b15zdnd11an1n64x5 FILLER_385_791 ();
 b15zdnd11an1n64x5 FILLER_385_855 ();
 b15zdnd11an1n64x5 FILLER_385_919 ();
 b15zdnd11an1n64x5 FILLER_385_983 ();
 b15zdnd11an1n64x5 FILLER_385_1047 ();
 b15zdnd11an1n64x5 FILLER_385_1111 ();
 b15zdnd11an1n32x5 FILLER_385_1175 ();
 b15zdnd11an1n16x5 FILLER_385_1207 ();
 b15zdnd11an1n08x5 FILLER_385_1223 ();
 b15zdnd00an1n02x5 FILLER_385_1231 ();
 b15zdnd11an1n64x5 FILLER_385_1275 ();
 b15zdnd11an1n64x5 FILLER_385_1339 ();
 b15zdnd11an1n64x5 FILLER_385_1403 ();
 b15zdnd11an1n16x5 FILLER_385_1467 ();
 b15zdnd11an1n64x5 FILLER_385_1525 ();
 b15zdnd11an1n16x5 FILLER_385_1589 ();
 b15zdnd00an1n02x5 FILLER_385_1605 ();
 b15zdnd11an1n08x5 FILLER_385_1649 ();
 b15zdnd00an1n01x5 FILLER_385_1657 ();
 b15zdnd11an1n64x5 FILLER_385_1700 ();
 b15zdnd11an1n64x5 FILLER_385_1764 ();
 b15zdnd11an1n64x5 FILLER_385_1828 ();
 b15zdnd11an1n64x5 FILLER_385_1892 ();
 b15zdnd11an1n64x5 FILLER_385_1956 ();
 b15zdnd11an1n64x5 FILLER_385_2020 ();
 b15zdnd11an1n64x5 FILLER_385_2084 ();
 b15zdnd11an1n64x5 FILLER_385_2148 ();
 b15zdnd11an1n64x5 FILLER_385_2212 ();
 b15zdnd11an1n08x5 FILLER_385_2276 ();
 b15zdnd11an1n64x5 FILLER_386_8 ();
 b15zdnd11an1n64x5 FILLER_386_72 ();
 b15zdnd11an1n64x5 FILLER_386_136 ();
 b15zdnd11an1n64x5 FILLER_386_200 ();
 b15zdnd11an1n64x5 FILLER_386_264 ();
 b15zdnd11an1n32x5 FILLER_386_328 ();
 b15zdnd11an1n16x5 FILLER_386_360 ();
 b15zdnd00an1n02x5 FILLER_386_376 ();
 b15zdnd11an1n08x5 FILLER_386_382 ();
 b15zdnd11an1n04x5 FILLER_386_394 ();
 b15zdnd11an1n04x5 FILLER_386_440 ();
 b15zdnd00an1n01x5 FILLER_386_444 ();
 b15zdnd11an1n04x5 FILLER_386_449 ();
 b15zdnd11an1n04x5 FILLER_386_457 ();
 b15zdnd00an1n02x5 FILLER_386_461 ();
 b15zdnd00an1n01x5 FILLER_386_463 ();
 b15zdnd11an1n64x5 FILLER_386_468 ();
 b15zdnd11an1n64x5 FILLER_386_532 ();
 b15zdnd00an1n01x5 FILLER_386_596 ();
 b15zdnd11an1n04x5 FILLER_386_601 ();
 b15zdnd11an1n04x5 FILLER_386_609 ();
 b15zdnd00an1n01x5 FILLER_386_613 ();
 b15zdnd11an1n32x5 FILLER_386_656 ();
 b15zdnd11an1n16x5 FILLER_386_688 ();
 b15zdnd11an1n08x5 FILLER_386_704 ();
 b15zdnd11an1n04x5 FILLER_386_712 ();
 b15zdnd00an1n02x5 FILLER_386_716 ();
 b15zdnd11an1n64x5 FILLER_386_726 ();
 b15zdnd11an1n64x5 FILLER_386_790 ();
 b15zdnd11an1n64x5 FILLER_386_854 ();
 b15zdnd11an1n64x5 FILLER_386_918 ();
 b15zdnd11an1n64x5 FILLER_386_982 ();
 b15zdnd11an1n64x5 FILLER_386_1046 ();
 b15zdnd11an1n64x5 FILLER_386_1110 ();
 b15zdnd11an1n64x5 FILLER_386_1174 ();
 b15zdnd11an1n32x5 FILLER_386_1238 ();
 b15zdnd11an1n08x5 FILLER_386_1270 ();
 b15zdnd00an1n02x5 FILLER_386_1278 ();
 b15zdnd11an1n04x5 FILLER_386_1284 ();
 b15zdnd11an1n04x5 FILLER_386_1292 ();
 b15zdnd00an1n01x5 FILLER_386_1296 ();
 b15zdnd11an1n64x5 FILLER_386_1301 ();
 b15zdnd11an1n64x5 FILLER_386_1365 ();
 b15zdnd11an1n64x5 FILLER_386_1429 ();
 b15zdnd11an1n64x5 FILLER_386_1493 ();
 b15zdnd11an1n64x5 FILLER_386_1557 ();
 b15zdnd11an1n16x5 FILLER_386_1621 ();
 b15zdnd11an1n64x5 FILLER_386_1641 ();
 b15zdnd11an1n64x5 FILLER_386_1705 ();
 b15zdnd11an1n64x5 FILLER_386_1769 ();
 b15zdnd11an1n64x5 FILLER_386_1833 ();
 b15zdnd11an1n64x5 FILLER_386_1897 ();
 b15zdnd11an1n64x5 FILLER_386_1961 ();
 b15zdnd11an1n64x5 FILLER_386_2025 ();
 b15zdnd11an1n64x5 FILLER_386_2089 ();
 b15zdnd00an1n01x5 FILLER_386_2153 ();
 b15zdnd11an1n64x5 FILLER_386_2162 ();
 b15zdnd11an1n32x5 FILLER_386_2226 ();
 b15zdnd11an1n16x5 FILLER_386_2258 ();
 b15zdnd00an1n02x5 FILLER_386_2274 ();
 b15zdnd11an1n64x5 FILLER_387_0 ();
 b15zdnd11an1n64x5 FILLER_387_64 ();
 b15zdnd11an1n64x5 FILLER_387_128 ();
 b15zdnd11an1n64x5 FILLER_387_192 ();
 b15zdnd11an1n64x5 FILLER_387_256 ();
 b15zdnd11an1n32x5 FILLER_387_320 ();
 b15zdnd11an1n16x5 FILLER_387_352 ();
 b15zdnd11an1n08x5 FILLER_387_368 ();
 b15zdnd00an1n02x5 FILLER_387_376 ();
 b15zdnd00an1n01x5 FILLER_387_378 ();
 b15zdnd11an1n08x5 FILLER_387_421 ();
 b15zdnd00an1n02x5 FILLER_387_429 ();
 b15zdnd00an1n01x5 FILLER_387_431 ();
 b15zdnd11an1n64x5 FILLER_387_474 ();
 b15zdnd11an1n32x5 FILLER_387_538 ();
 b15zdnd11an1n16x5 FILLER_387_570 ();
 b15zdnd11an1n08x5 FILLER_387_586 ();
 b15zdnd11an1n04x5 FILLER_387_594 ();
 b15zdnd11an1n04x5 FILLER_387_602 ();
 b15zdnd11an1n04x5 FILLER_387_610 ();
 b15zdnd00an1n01x5 FILLER_387_614 ();
 b15zdnd11an1n16x5 FILLER_387_657 ();
 b15zdnd11an1n08x5 FILLER_387_673 ();
 b15zdnd00an1n01x5 FILLER_387_681 ();
 b15zdnd11an1n64x5 FILLER_387_724 ();
 b15zdnd11an1n64x5 FILLER_387_788 ();
 b15zdnd11an1n64x5 FILLER_387_852 ();
 b15zdnd11an1n64x5 FILLER_387_916 ();
 b15zdnd11an1n64x5 FILLER_387_980 ();
 b15zdnd11an1n64x5 FILLER_387_1044 ();
 b15zdnd11an1n08x5 FILLER_387_1108 ();
 b15zdnd11an1n04x5 FILLER_387_1120 ();
 b15zdnd11an1n08x5 FILLER_387_1135 ();
 b15zdnd00an1n01x5 FILLER_387_1143 ();
 b15zdnd11an1n16x5 FILLER_387_1148 ();
 b15zdnd11an1n04x5 FILLER_387_1164 ();
 b15zdnd00an1n01x5 FILLER_387_1168 ();
 b15zdnd11an1n64x5 FILLER_387_1173 ();
 b15zdnd11an1n16x5 FILLER_387_1237 ();
 b15zdnd00an1n02x5 FILLER_387_1253 ();
 b15zdnd11an1n04x5 FILLER_387_1259 ();
 b15zdnd11an1n04x5 FILLER_387_1267 ();
 b15zdnd00an1n01x5 FILLER_387_1271 ();
 b15zdnd11an1n04x5 FILLER_387_1276 ();
 b15zdnd00an1n02x5 FILLER_387_1280 ();
 b15zdnd00an1n01x5 FILLER_387_1282 ();
 b15zdnd11an1n04x5 FILLER_387_1287 ();
 b15zdnd11an1n04x5 FILLER_387_1295 ();
 b15zdnd11an1n04x5 FILLER_387_1303 ();
 b15zdnd11an1n04x5 FILLER_387_1311 ();
 b15zdnd11an1n64x5 FILLER_387_1319 ();
 b15zdnd11an1n32x5 FILLER_387_1383 ();
 b15zdnd11an1n08x5 FILLER_387_1415 ();
 b15zdnd11an1n04x5 FILLER_387_1423 ();
 b15zdnd00an1n02x5 FILLER_387_1427 ();
 b15zdnd00an1n01x5 FILLER_387_1429 ();
 b15zdnd11an1n04x5 FILLER_387_1434 ();
 b15zdnd11an1n04x5 FILLER_387_1442 ();
 b15zdnd11an1n16x5 FILLER_387_1450 ();
 b15zdnd11an1n08x5 FILLER_387_1466 ();
 b15zdnd00an1n02x5 FILLER_387_1474 ();
 b15zdnd11an1n04x5 FILLER_387_1480 ();
 b15zdnd11an1n08x5 FILLER_387_1488 ();
 b15zdnd00an1n01x5 FILLER_387_1496 ();
 b15zdnd11an1n64x5 FILLER_387_1501 ();
 b15zdnd11an1n32x5 FILLER_387_1565 ();
 b15zdnd11an1n04x5 FILLER_387_1597 ();
 b15zdnd00an1n01x5 FILLER_387_1601 ();
 b15zdnd11an1n08x5 FILLER_387_1606 ();
 b15zdnd11an1n04x5 FILLER_387_1614 ();
 b15zdnd00an1n02x5 FILLER_387_1618 ();
 b15zdnd11an1n08x5 FILLER_387_1624 ();
 b15zdnd11an1n04x5 FILLER_387_1632 ();
 b15zdnd00an1n01x5 FILLER_387_1636 ();
 b15zdnd11an1n64x5 FILLER_387_1679 ();
 b15zdnd11an1n64x5 FILLER_387_1743 ();
 b15zdnd11an1n64x5 FILLER_387_1807 ();
 b15zdnd11an1n64x5 FILLER_387_1871 ();
 b15zdnd11an1n64x5 FILLER_387_1935 ();
 b15zdnd11an1n64x5 FILLER_387_1999 ();
 b15zdnd11an1n64x5 FILLER_387_2063 ();
 b15zdnd11an1n64x5 FILLER_387_2127 ();
 b15zdnd11an1n64x5 FILLER_387_2191 ();
 b15zdnd11an1n16x5 FILLER_387_2255 ();
 b15zdnd11an1n08x5 FILLER_387_2271 ();
 b15zdnd11an1n04x5 FILLER_387_2279 ();
 b15zdnd00an1n01x5 FILLER_387_2283 ();
 b15zdnd11an1n64x5 FILLER_388_8 ();
 b15zdnd11an1n64x5 FILLER_388_72 ();
 b15zdnd11an1n64x5 FILLER_388_136 ();
 b15zdnd11an1n64x5 FILLER_388_200 ();
 b15zdnd11an1n64x5 FILLER_388_264 ();
 b15zdnd11an1n32x5 FILLER_388_328 ();
 b15zdnd11an1n04x5 FILLER_388_360 ();
 b15zdnd00an1n01x5 FILLER_388_364 ();
 b15zdnd11an1n04x5 FILLER_388_369 ();
 b15zdnd11an1n04x5 FILLER_388_377 ();
 b15zdnd11an1n04x5 FILLER_388_385 ();
 b15zdnd11an1n04x5 FILLER_388_393 ();
 b15zdnd11an1n04x5 FILLER_388_401 ();
 b15zdnd11an1n04x5 FILLER_388_447 ();
 b15zdnd11an1n64x5 FILLER_388_493 ();
 b15zdnd11an1n32x5 FILLER_388_557 ();
 b15zdnd11an1n04x5 FILLER_388_589 ();
 b15zdnd11an1n04x5 FILLER_388_597 ();
 b15zdnd11an1n04x5 FILLER_388_605 ();
 b15zdnd11an1n04x5 FILLER_388_613 ();
 b15zdnd11an1n04x5 FILLER_388_659 ();
 b15zdnd11an1n08x5 FILLER_388_667 ();
 b15zdnd11an1n04x5 FILLER_388_675 ();
 b15zdnd11an1n32x5 FILLER_388_683 ();
 b15zdnd00an1n02x5 FILLER_388_715 ();
 b15zdnd00an1n01x5 FILLER_388_717 ();
 b15zdnd11an1n32x5 FILLER_388_726 ();
 b15zdnd11an1n08x5 FILLER_388_758 ();
 b15zdnd11an1n04x5 FILLER_388_766 ();
 b15zdnd11an1n08x5 FILLER_388_774 ();
 b15zdnd11an1n04x5 FILLER_388_782 ();
 b15zdnd11an1n08x5 FILLER_388_790 ();
 b15zdnd11an1n04x5 FILLER_388_798 ();
 b15zdnd00an1n02x5 FILLER_388_802 ();
 b15zdnd11an1n16x5 FILLER_388_808 ();
 b15zdnd00an1n02x5 FILLER_388_824 ();
 b15zdnd11an1n08x5 FILLER_388_831 ();
 b15zdnd11an1n04x5 FILLER_388_839 ();
 b15zdnd00an1n01x5 FILLER_388_843 ();
 b15zdnd11an1n64x5 FILLER_388_848 ();
 b15zdnd11an1n64x5 FILLER_388_912 ();
 b15zdnd11an1n32x5 FILLER_388_976 ();
 b15zdnd11an1n16x5 FILLER_388_1008 ();
 b15zdnd11an1n08x5 FILLER_388_1024 ();
 b15zdnd00an1n02x5 FILLER_388_1032 ();
 b15zdnd11an1n04x5 FILLER_388_1038 ();
 b15zdnd11an1n08x5 FILLER_388_1046 ();
 b15zdnd11an1n04x5 FILLER_388_1054 ();
 b15zdnd00an1n01x5 FILLER_388_1058 ();
 b15zdnd11an1n32x5 FILLER_388_1067 ();
 b15zdnd00an1n02x5 FILLER_388_1099 ();
 b15zdnd00an1n01x5 FILLER_388_1101 ();
 b15zdnd11an1n08x5 FILLER_388_1106 ();
 b15zdnd00an1n02x5 FILLER_388_1114 ();
 b15zdnd00an1n01x5 FILLER_388_1116 ();
 b15zdnd11an1n04x5 FILLER_388_1159 ();
 b15zdnd11an1n08x5 FILLER_388_1167 ();
 b15zdnd00an1n02x5 FILLER_388_1175 ();
 b15zdnd11an1n04x5 FILLER_388_1185 ();
 b15zdnd11an1n04x5 FILLER_388_1193 ();
 b15zdnd00an1n02x5 FILLER_388_1197 ();
 b15zdnd11an1n04x5 FILLER_388_1203 ();
 b15zdnd11an1n08x5 FILLER_388_1218 ();
 b15zdnd11an1n08x5 FILLER_388_1230 ();
 b15zdnd11an1n04x5 FILLER_388_1238 ();
 b15zdnd11an1n04x5 FILLER_388_1246 ();
 b15zdnd00an1n02x5 FILLER_388_1250 ();
 b15zdnd00an1n01x5 FILLER_388_1252 ();
 b15zdnd11an1n08x5 FILLER_388_1259 ();
 b15zdnd00an1n02x5 FILLER_388_1267 ();
 b15zdnd11an1n04x5 FILLER_388_1274 ();
 b15zdnd00an1n02x5 FILLER_388_1278 ();
 b15zdnd00an1n01x5 FILLER_388_1280 ();
 b15zdnd11an1n08x5 FILLER_388_1323 ();
 b15zdnd00an1n02x5 FILLER_388_1331 ();
 b15zdnd00an1n01x5 FILLER_388_1333 ();
 b15zdnd11an1n08x5 FILLER_388_1376 ();
 b15zdnd00an1n02x5 FILLER_388_1384 ();
 b15zdnd11an1n04x5 FILLER_388_1390 ();
 b15zdnd11an1n08x5 FILLER_388_1398 ();
 b15zdnd11an1n04x5 FILLER_388_1406 ();
 b15zdnd11an1n04x5 FILLER_388_1414 ();
 b15zdnd11an1n08x5 FILLER_388_1422 ();
 b15zdnd00an1n02x5 FILLER_388_1430 ();
 b15zdnd00an1n01x5 FILLER_388_1432 ();
 b15zdnd11an1n04x5 FILLER_388_1475 ();
 b15zdnd00an1n02x5 FILLER_388_1479 ();
 b15zdnd00an1n01x5 FILLER_388_1481 ();
 b15zdnd11an1n32x5 FILLER_388_1524 ();
 b15zdnd11an1n16x5 FILLER_388_1556 ();
 b15zdnd11an1n08x5 FILLER_388_1572 ();
 b15zdnd11an1n04x5 FILLER_388_1580 ();
 b15zdnd00an1n01x5 FILLER_388_1584 ();
 b15zdnd11an1n08x5 FILLER_388_1589 ();
 b15zdnd11an1n04x5 FILLER_388_1597 ();
 b15zdnd00an1n02x5 FILLER_388_1601 ();
 b15zdnd00an1n01x5 FILLER_388_1603 ();
 b15zdnd11an1n04x5 FILLER_388_1611 ();
 b15zdnd00an1n01x5 FILLER_388_1615 ();
 b15zdnd11an1n32x5 FILLER_388_1658 ();
 b15zdnd00an1n01x5 FILLER_388_1690 ();
 b15zdnd11an1n04x5 FILLER_388_1695 ();
 b15zdnd11an1n08x5 FILLER_388_1703 ();
 b15zdnd11an1n64x5 FILLER_388_1753 ();
 b15zdnd11an1n64x5 FILLER_388_1817 ();
 b15zdnd11an1n64x5 FILLER_388_1881 ();
 b15zdnd11an1n64x5 FILLER_388_1945 ();
 b15zdnd11an1n64x5 FILLER_388_2009 ();
 b15zdnd11an1n64x5 FILLER_388_2073 ();
 b15zdnd11an1n16x5 FILLER_388_2137 ();
 b15zdnd00an1n01x5 FILLER_388_2153 ();
 b15zdnd11an1n64x5 FILLER_388_2162 ();
 b15zdnd11an1n32x5 FILLER_388_2226 ();
 b15zdnd11an1n16x5 FILLER_388_2258 ();
 b15zdnd00an1n02x5 FILLER_388_2274 ();
 b15zdnd11an1n64x5 FILLER_389_0 ();
 b15zdnd11an1n64x5 FILLER_389_64 ();
 b15zdnd11an1n64x5 FILLER_389_128 ();
 b15zdnd11an1n64x5 FILLER_389_192 ();
 b15zdnd11an1n64x5 FILLER_389_256 ();
 b15zdnd11an1n32x5 FILLER_389_320 ();
 b15zdnd11an1n08x5 FILLER_389_352 ();
 b15zdnd00an1n02x5 FILLER_389_360 ();
 b15zdnd11an1n04x5 FILLER_389_404 ();
 b15zdnd11an1n04x5 FILLER_389_450 ();
 b15zdnd11an1n04x5 FILLER_389_496 ();
 b15zdnd11an1n16x5 FILLER_389_507 ();
 b15zdnd11an1n08x5 FILLER_389_523 ();
 b15zdnd11an1n04x5 FILLER_389_531 ();
 b15zdnd00an1n02x5 FILLER_389_535 ();
 b15zdnd00an1n01x5 FILLER_389_537 ();
 b15zdnd11an1n16x5 FILLER_389_542 ();
 b15zdnd11an1n08x5 FILLER_389_565 ();
 b15zdnd00an1n02x5 FILLER_389_573 ();
 b15zdnd11an1n04x5 FILLER_389_617 ();
 b15zdnd11an1n04x5 FILLER_389_663 ();
 b15zdnd00an1n02x5 FILLER_389_667 ();
 b15zdnd11an1n08x5 FILLER_389_675 ();
 b15zdnd00an1n02x5 FILLER_389_683 ();
 b15zdnd00an1n01x5 FILLER_389_685 ();
 b15zdnd11an1n04x5 FILLER_389_690 ();
 b15zdnd11an1n16x5 FILLER_389_736 ();
 b15zdnd11an1n04x5 FILLER_389_752 ();
 b15zdnd00an1n02x5 FILLER_389_756 ();
 b15zdnd11an1n04x5 FILLER_389_800 ();
 b15zdnd11an1n08x5 FILLER_389_846 ();
 b15zdnd11an1n04x5 FILLER_389_858 ();
 b15zdnd00an1n02x5 FILLER_389_862 ();
 b15zdnd00an1n01x5 FILLER_389_864 ();
 b15zdnd11an1n64x5 FILLER_389_907 ();
 b15zdnd11an1n32x5 FILLER_389_971 ();
 b15zdnd11an1n16x5 FILLER_389_1003 ();
 b15zdnd11an1n04x5 FILLER_389_1023 ();
 b15zdnd11an1n32x5 FILLER_389_1069 ();
 b15zdnd11an1n04x5 FILLER_389_1105 ();
 b15zdnd11an1n04x5 FILLER_389_1115 ();
 b15zdnd11an1n08x5 FILLER_389_1123 ();
 b15zdnd11an1n04x5 FILLER_389_1131 ();
 b15zdnd00an1n02x5 FILLER_389_1135 ();
 b15zdnd00an1n01x5 FILLER_389_1137 ();
 b15zdnd11an1n04x5 FILLER_389_1142 ();
 b15zdnd00an1n01x5 FILLER_389_1146 ();
 b15zdnd11an1n04x5 FILLER_389_1151 ();
 b15zdnd11an1n08x5 FILLER_389_1197 ();
 b15zdnd00an1n02x5 FILLER_389_1205 ();
 b15zdnd11an1n04x5 FILLER_389_1249 ();
 b15zdnd11an1n04x5 FILLER_389_1295 ();
 b15zdnd11an1n04x5 FILLER_389_1341 ();
 b15zdnd11an1n04x5 FILLER_389_1349 ();
 b15zdnd11an1n04x5 FILLER_389_1357 ();
 b15zdnd00an1n02x5 FILLER_389_1361 ();
 b15zdnd11an1n04x5 FILLER_389_1367 ();
 b15zdnd11an1n04x5 FILLER_389_1413 ();
 b15zdnd11an1n04x5 FILLER_389_1459 ();
 b15zdnd11an1n04x5 FILLER_389_1505 ();
 b15zdnd11an1n08x5 FILLER_389_1551 ();
 b15zdnd11an1n04x5 FILLER_389_1559 ();
 b15zdnd00an1n01x5 FILLER_389_1563 ();
 b15zdnd11an1n16x5 FILLER_389_1569 ();
 b15zdnd00an1n02x5 FILLER_389_1585 ();
 b15zdnd11an1n04x5 FILLER_389_1629 ();
 b15zdnd11an1n04x5 FILLER_389_1675 ();
 b15zdnd11an1n04x5 FILLER_389_1721 ();
 b15zdnd11an1n64x5 FILLER_389_1729 ();
 b15zdnd11an1n64x5 FILLER_389_1793 ();
 b15zdnd11an1n64x5 FILLER_389_1857 ();
 b15zdnd11an1n64x5 FILLER_389_1921 ();
 b15zdnd11an1n64x5 FILLER_389_1985 ();
 b15zdnd11an1n64x5 FILLER_389_2049 ();
 b15zdnd11an1n64x5 FILLER_389_2113 ();
 b15zdnd11an1n64x5 FILLER_389_2177 ();
 b15zdnd11an1n32x5 FILLER_389_2241 ();
 b15zdnd11an1n08x5 FILLER_389_2273 ();
 b15zdnd00an1n02x5 FILLER_389_2281 ();
 b15zdnd00an1n01x5 FILLER_389_2283 ();
endmodule
