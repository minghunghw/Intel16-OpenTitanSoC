************************************************************************
* auCdl Netlist:
* 
* Library Name:  2305_tisar
* Top Cell Name: Noise_injection_block_modified_v13
* View Name:     schematic
* Netlisted on:  May 20 16:33:27 2023
************************************************************************

.INCLUDE  /afs/eecs.umich.edu/kits/Intel/P1222.4/2022.08/pdk224_r0.9HP3/libraries/custom/cdl/common/intel22custom.cdl
*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



*.EQUIV vss=vss!
*.EXPAND_ON_M_FACTOR

************************************************************************
* Library Name: intel22custom
* Cell Name:    mfc_s2s_ns_pcell_0
* View Name:    schematic
************************************************************************

.SUBCKT mfc_s2s_ns_pcell_0 a b
*.PININFO a:B b:B
XI0 a b  b88xp_mfcs2sns mtop=6 mbot=1 w=640.00n l=640.00n multx=1 multy=10 
+ fill=0 via=1 shield=0
.ENDS

************************************************************************
* Library Name: 2305_tisar
* Cell Name:    Noise_injection_block_v17
* View Name:    schematic
************************************************************************

.SUBCKT Noise_injection_block_v17 Iout Random S<0> S<1> S<2> S<3> VB vdd vss
*.PININFO Iout:B Random:B S<0>:B S<1>:B S<2>:B S<3>:B VB:B vdd:B vss:B
MMN43 net2 S<3> vss vss nulvt W=360n L=40n m=200
MMN42 net2 S<3> vss vss nulvt W=360n L=40n m=100
MMN41 net2 S<3> vss vss nulvt W=360n L=40n m=200
MMN38 net4 S<2> vss vss nulvt W=360n L=40n m=200
MMN37 net3 S<1> vss vss nulvt W=360n L=40n m=200
MMN36 net1 S<0> vss vss nulvt W=360n L=40n m=100
MMP23 Iout VB vdd vdd pulvt W=360n L=40n m=90
XI97 Random net2 / mfc_s2s_ns_pcell_0
XI96 net2 Random / mfc_s2s_ns_pcell_0
XI95 VB net2 / mfc_s2s_ns_pcell_0
XI94 net2 VB / mfc_s2s_ns_pcell_0
XI52 net3 VB / mfc_s2s_ns_pcell_0
XI51 net1 VB / mfc_s2s_ns_pcell_0
XI50 net3 VB / mfc_s2s_ns_pcell_0
XI49 net3 VB / mfc_s2s_ns_pcell_0
XI65 Random net1 / mfc_s2s_ns_pcell_0
XI47 Random net3 / mfc_s2s_ns_pcell_0
XI46 Random net3 / mfc_s2s_ns_pcell_0
XI45 Random net3 / mfc_s2s_ns_pcell_0
XI44 Random net4 / mfc_s2s_ns_pcell_0
XI43 Random net4 / mfc_s2s_ns_pcell_0
XI42 Random net4 / mfc_s2s_ns_pcell_0
XI41 net4 VB / mfc_s2s_ns_pcell_0
XI40 net4 VB / mfc_s2s_ns_pcell_0
XI39 net4 VB / mfc_s2s_ns_pcell_0
XI38 net4 VB / mfc_s2s_ns_pcell_0
XI37 Random net4 / mfc_s2s_ns_pcell_0
XI36 net4 Random / mfc_s2s_ns_pcell_0
XI35 VB net4 / mfc_s2s_ns_pcell_0
XI34 net4 Random / mfc_s2s_ns_pcell_0
XI33 VB net4 / mfc_s2s_ns_pcell_0
XI32 net4 Random / mfc_s2s_ns_pcell_0
XI31 VB net4 / mfc_s2s_ns_pcell_0
XI30 net4 Random / mfc_s2s_ns_pcell_0
XI29 VB net4 / mfc_s2s_ns_pcell_0
XI28 net3 Random / mfc_s2s_ns_pcell_0
XI27 VB net3 / mfc_s2s_ns_pcell_0
XI26 net3 Random / mfc_s2s_ns_pcell_0
XI25 VB net3 / mfc_s2s_ns_pcell_0
XI24 net3 Random / mfc_s2s_ns_pcell_0
XI23 VB net3 / mfc_s2s_ns_pcell_0
XI22 net1 Random / mfc_s2s_ns_pcell_0
XI21 VB net1 / mfc_s2s_ns_pcell_0
XI78 Random net2 / mfc_s2s_ns_pcell_0
XI93 net2 Random / mfc_s2s_ns_pcell_0
XI77 net2 Random / mfc_s2s_ns_pcell_0
XI76 net2 Random / mfc_s2s_ns_pcell_0
XI89 net2 VB / mfc_s2s_ns_pcell_0
XI67 net2 VB / mfc_s2s_ns_pcell_0
XI66 net2 VB / mfc_s2s_ns_pcell_0
XI68 net2 VB / mfc_s2s_ns_pcell_0
XI69 net2 VB / mfc_s2s_ns_pcell_0
XI70 VB net2 / mfc_s2s_ns_pcell_0
XI71 VB net2 / mfc_s2s_ns_pcell_0
XI72 VB net2 / mfc_s2s_ns_pcell_0
XI81 Random net2 / mfc_s2s_ns_pcell_0
XI80 Random net2 / mfc_s2s_ns_pcell_0
XI85 Random net2 / mfc_s2s_ns_pcell_0
XI73 VB net2 / mfc_s2s_ns_pcell_0
XI82 Random net2 / mfc_s2s_ns_pcell_0
XI74 net2 Random / mfc_s2s_ns_pcell_0
XI84 VB net2 / mfc_s2s_ns_pcell_0
XI92 net2 Random / mfc_s2s_ns_pcell_0
XI75 net2 Random / mfc_s2s_ns_pcell_0
XI88 VB net2 / mfc_s2s_ns_pcell_0
XI83 net2 Random / mfc_s2s_ns_pcell_0
XI91 net2 VB / mfc_s2s_ns_pcell_0
XI90 net2 VB / mfc_s2s_ns_pcell_0
XI87 VB net2 / mfc_s2s_ns_pcell_0
XI86 Random net2 / mfc_s2s_ns_pcell_0
XI79 Random net2 / mfc_s2s_ns_pcell_0
.ENDS

************************************************************************
* Library Name: 2305_tisar
* Cell Name:    Noise_injection_block_modified_v13
* View Name:    schematic
************************************************************************

.SUBCKT Noise_injection_block_modified_v13 Iout Random S<0> S<1> S<2> S<3> 
+ S<4> S<5> S<6> S<7> S<8> S<9> S<10> S<11> S<12> S<13> S<14> S<15> VB<0> 
+ VB<1> VB<2> VB<3> vdd vss
*.PININFO Iout:B Random:B S<0>:B S<1>:B S<2>:B S<3>:B S<4>:B S<5>:B S<6>:B 
*.PININFO S<7>:B S<8>:B S<9>:B S<10>:B S<11>:B S<12>:B S<13>:B S<14>:B S<15>:B 
*.PININFO VB<0>:B VB<1>:B VB<2>:B VB<3>:B vdd:B vss:B
XI101 Iout Random S<12> S<13> S<14> S<15> VB<3> vdd vss / 
+ Noise_injection_block_v17
XI98 Iout Random S<4> S<5> S<6> S<7> VB<1> vdd vss / Noise_injection_block_v17
XI99 Iout Random S<0> S<1> S<2> S<3> VB<0> vdd vss / Noise_injection_block_v17
XI100 Iout Random S<8> S<9> S<10> S<11> VB<2> vdd vss / 
+ Noise_injection_block_v17
.ENDS

