## ##############################################################################
## ## Intel Top Secret                                                         ##
## ##############################################################################
## ## Copyright © Intel Corporation.                                           ##
## ##                                                                          ##
## ## This is the property of Intel Corporation and may only be utilized       ##
## ## pursuant to a written Restricted Use Nondisclosure Agreement             ##
## ## with Intel Corporation.  It may not be used, reproduced, or              ##
## ## disclosed to others except in accordance with the terms and              ##
## ## conditions of such agreement.                                            ##
## ##                                                                          ##
## ## All products, processes, computer systems, dates, and figures            ##
## ## specified are preliminary based on current expectations, and are         ##
## ## subject to change without notice.                                        ##
## ##############################################################################
## ## Text_Tag % __Placeholder neutral1


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO b15cdiar2hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cdiar2hn1n04x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.158 3.166 0.472 ;
      LAYER v0 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.068 3.058 0.562 ;
      LAYER v0 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 2.99 0.138 3.058 0.182 ;
    END
  END clkout
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.2705 0.466 0.3145 ;
    END
  END d
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.95583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 3.716875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.202 ;
      LAYER v0 ;
        RECT 2.558 0.138 2.626 0.182 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.098 0.538 3.166 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.098 0.048 3.166 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.428 3.292 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.782 0.518 2.018 0.562 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 1.694 0.428 1.91 0.472 ;
      RECT 3.206 0.068 3.274 0.562 ;
    LAYER v1 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.186 0.428 0.246 0.472 ;
    LAYER v0 ;
      RECT 3.206 0.138 3.274 0.182 ;
      RECT 3.206 0.448 3.274 0.492 ;
      RECT 2.774 0.248 2.842 0.292 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.912 0.138 1.976 0.182 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.154 0.138 1.222 0.182 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.614 0.2705 0.682 0.3145 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.506 0.408 0.574 0.452 ;
      RECT 0.182 0.2705 0.25 0.3145 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.006 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.338 1.762 0.382 ;
      RECT 1.222 0.248 1.478 0.292 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 1.546 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.382 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 2.194 0.338 2.342 0.382 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 1.91 0.068 1.978 0.472 ;
      RECT 1.978 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.302 0.248 2.95 0.292 ;
  END
END b15cdiar2hn1n04x5

MACRO b15cdiar2hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cdiar2hn1n08x5 0 0 ;
  SIZE 3.996 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.068 3.706 0.382 ;
      LAYER v0 ;
        RECT 3.638 0.248 3.706 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.068 3.49 0.562 ;
      LAYER v0 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.422 0.138 3.49 0.182 ;
    END
  END clkout
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END d
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 3.256389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 2.170926 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.248 3.078 0.292 ;
        RECT 2.666 0.068 2.734 0.292 ;
        RECT 1.802 0.068 2.734 0.112 ;
        RECT 1.458 0.158 1.87 0.202 ;
        RECT 1.802 0.068 1.87 0.202 ;
      LAYER v0 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 2.99 0.248 3.058 0.292 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.03 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.45 0.248 2.518 0.472 ;
        RECT 2.234 0.248 2.518 0.292 ;
        RECT 2.234 0.248 2.302 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.45 0.408 2.518 0.452 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.53 0.448 3.598 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.03 0.022 ;
        RECT 3.53 -0.022 3.598 0.202 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 3.314 0.138 3.382 0.182 ;
        RECT 3.53 0.138 3.598 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.428 3.832 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 3.746 0.068 3.814 0.562 ;
    LAYER v1 ;
      RECT 3.75 0.428 3.81 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 0.726 0.428 0.786 0.472 ;
      RECT 0.186 0.428 0.246 0.472 ;
    LAYER v0 ;
      RECT 3.746 0.138 3.814 0.182 ;
      RECT 3.746 0.448 3.814 0.492 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 2.774 0.448 2.842 0.492 ;
      RECT 2.342 0.408 2.41 0.452 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.293 2.194 0.337 ;
      RECT 2.018 0.3965 2.086 0.4405 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.154 0.138 1.222 0.182 ;
      RECT 1.156 0.408 1.22 0.452 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.408 0.682 0.452 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.506 0.408 0.574 0.452 ;
      RECT 0.182 0.293 0.25 0.337 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.158 0.83 0.202 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.33 0.428 1.566 0.472 ;
      RECT 1.006 0.338 1.154 0.382 ;
      RECT 1.154 0.338 1.222 0.472 ;
      RECT 1.222 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.222 0.248 1.87 0.292 ;
      RECT 2.41 0.518 2.774 0.562 ;
      RECT 2.774 0.428 2.842 0.562 ;
      RECT 2.086 0.158 2.558 0.202 ;
      RECT 2.558 0.158 2.626 0.382 ;
      RECT 2.626 0.338 3.206 0.382 ;
      RECT 3.206 0.158 3.274 0.382 ;
  END
END b15cdiar2hn1n08x5

MACRO b15cdiyr2hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cdiyr2hn1n04x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.248 1.762 0.562 ;
      LAYER v0 ;
        RECT 1.694 0.338 1.762 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.342 0.178 2.41 0.222 ;
    END
  END clkout
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.2705 0.466 0.3145 ;
    END
  END d
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.046 0.338 1.114 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.046 0.408 1.114 0.452 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.234 -0.022 2.302 0.382 ;
        RECT 1.478 0.158 2.302 0.202 ;
        RECT 0.83 0.158 1.114 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.234 0.2585 2.302 0.3025 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.428 1.888 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 1.154 0.518 1.37 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.802 0.338 1.87 0.562 ;
    LAYER v1 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.186 0.428 0.246 0.472 ;
    LAYER v0 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.802 0.4445 1.87 0.4885 ;
      RECT 1.478 0.2705 1.546 0.3145 ;
      RECT 1.37 0.1535 1.438 0.1975 ;
      RECT 1.262 0.3155 1.33 0.3595 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.154 0.138 1.222 0.182 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.614 0.2705 0.682 0.3145 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.506 0.408 0.574 0.452 ;
      RECT 0.182 0.2705 0.25 0.3145 ;
    LAYER m1 ;
      RECT 0.938 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.472 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.438 0.068 1.998 0.112 ;
  END
END b15cdiyr2hn1n04x5

MACRO b15cdiyr2hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cdiyr2hn1n08x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.498 0.466 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.4645 2.518 0.5085 ;
        RECT 2.45 0.1205 2.518 0.1645 ;
    END
  END clkout
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.64666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.64666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.338 2.194 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.384 0.358 0.428 ;
        RECT 0.83 0.383 0.898 0.427 ;
        RECT 1.478 0.383 1.546 0.427 ;
        RECT 2.126 0.383 2.194 0.427 ;
        RECT 2.342 0.4645 2.41 0.5085 ;
        RECT 2.558 0.4645 2.626 0.5085 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.262 0.158 1.654 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
        RECT 0.83 0.198 0.898 0.242 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 2.126 0.203 2.194 0.247 ;
        RECT 2.342 0.1205 2.41 0.1645 ;
        RECT 2.558 0.1205 2.626 0.1645 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.244 0.338 1.688 0.382 ;
      RECT 0.164 0.158 1.78 0.202 ;
      RECT 1.768 0.338 2.428 0.382 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.154 0.158 1.222 0.382 ;
      RECT 1.262 0.248 1.33 0.382 ;
      RECT 1.586 0.428 1.802 0.472 ;
      RECT 1.586 0.248 1.654 0.382 ;
      RECT 1.694 0.158 1.762 0.382 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.018 0.068 2.086 0.382 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.342 0.248 2.41 0.382 ;
    LAYER v1 ;
      RECT 2.346 0.338 2.406 0.382 ;
      RECT 1.806 0.338 1.866 0.382 ;
      RECT 1.698 0.158 1.758 0.202 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 1.158 0.158 1.218 0.202 ;
      RECT 0.186 0.158 0.246 0.202 ;
    LAYER v0 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.234 0.1205 2.302 0.1645 ;
      RECT 2.234 0.4645 2.302 0.5085 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.088 1.978 0.132 ;
      RECT 1.91 0.498 1.978 0.542 ;
      RECT 1.802 0.203 1.87 0.247 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.198 1.114 0.242 ;
      RECT 0.938 0.198 1.006 0.242 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.182 0.203 0.25 0.247 ;
      RECT 0.182 0.384 0.25 0.428 ;
    LAYER m1 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 1.114 0.428 1.33 0.472 ;
      RECT 1.114 0.068 1.546 0.112 ;
      RECT 1.802 0.158 1.87 0.472 ;
  END
END b15cdiyr2hn1n08x5

MACRO b15cilao5hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilao5hn1n02x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.338 2.086 0.382 ;
        RECT 1.478 0.518 1.762 0.562 ;
        RECT 1.694 0.338 1.762 0.562 ;
        RECT 1.478 0.248 1.546 0.562 ;
        RECT 0.702 0.248 1.546 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.91 0.338 1.978 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.342 0.138 2.41 0.182 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.594 0.382 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.486 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.586 0.248 1.87 0.292 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.586 0.158 1.654 0.292 ;
        RECT 1.242 0.158 1.654 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 2.234 0.138 2.302 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.562 ;
      RECT 0.398 0.158 1.134 0.202 ;
      RECT 0.81 0.068 1.694 0.112 ;
      RECT 1.91 0.158 2.126 0.202 ;
    LAYER v0 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.696 0.138 1.76 0.182 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.724 0.408 0.788 0.452 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.338 1.026 0.382 ;
      RECT 0.142 0.248 0.182 0.292 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.142 0.518 0.29 0.562 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.518 1.154 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.338 1.35 0.382 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 2.126 0.158 2.194 0.562 ;
  END
END b15cilao5hn1n02x5

MACRO b15cilao5hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilao5hn1n04x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.338 2.086 0.382 ;
        RECT 1.478 0.518 1.762 0.562 ;
        RECT 1.694 0.338 1.762 0.562 ;
        RECT 1.478 0.248 1.546 0.562 ;
        RECT 0.702 0.248 1.546 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.91 0.338 1.978 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.342 0.138 2.41 0.182 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.594 0.382 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.486 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.586 0.248 1.87 0.292 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.586 0.158 1.654 0.292 ;
        RECT 1.242 0.158 1.654 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 2.234 0.138 2.302 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.562 ;
      RECT 0.398 0.158 1.134 0.202 ;
      RECT 0.81 0.068 1.694 0.112 ;
      RECT 1.91 0.158 2.126 0.202 ;
    LAYER v0 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.696 0.138 1.76 0.182 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.724 0.408 0.788 0.452 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.338 1.026 0.382 ;
      RECT 0.142 0.248 0.182 0.292 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.142 0.518 0.29 0.562 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.518 1.154 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.338 1.35 0.382 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 2.126 0.158 2.194 0.562 ;
  END
END b15cilao5hn1n04x5

MACRO b15cilao5hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilao5hn1n06x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.64666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.338 2.086 0.382 ;
        RECT 1.478 0.518 1.762 0.562 ;
        RECT 1.694 0.338 1.762 0.562 ;
        RECT 1.478 0.248 1.546 0.562 ;
        RECT 0.702 0.248 1.546 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.91 0.338 1.978 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
        RECT 2.342 0.338 2.626 0.382 ;
        RECT 2.342 0.068 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.558 0.138 2.626 0.182 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.594 0.382 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.486 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.586 0.248 1.87 0.292 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.586 0.158 1.654 0.292 ;
        RECT 1.242 0.158 1.654 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.562 ;
      RECT 0.398 0.158 1.134 0.202 ;
      RECT 0.81 0.068 1.694 0.112 ;
      RECT 1.91 0.158 2.126 0.202 ;
    LAYER v0 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.694 0.138 1.762 0.182 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.724 0.408 0.788 0.452 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.338 1.026 0.382 ;
      RECT 0.142 0.248 0.182 0.292 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.142 0.518 0.29 0.562 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.518 1.154 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.338 1.35 0.382 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 2.126 0.158 2.194 0.562 ;
  END
END b15cilao5hn1n06x5

MACRO b15cilao5hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilao5hn1n08x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.338 2.086 0.382 ;
        RECT 1.478 0.518 1.762 0.562 ;
        RECT 1.694 0.338 1.762 0.562 ;
        RECT 1.478 0.248 1.546 0.562 ;
        RECT 0.702 0.248 1.546 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.91 0.338 1.978 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
        RECT 2.342 0.338 2.626 0.382 ;
        RECT 2.342 0.068 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.558 0.138 2.626 0.182 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.594 0.382 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.486 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.586 0.248 1.87 0.292 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.586 0.158 1.654 0.292 ;
        RECT 1.242 0.158 1.654 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.562 ;
      RECT 0.398 0.158 1.134 0.202 ;
      RECT 0.81 0.068 1.694 0.112 ;
      RECT 1.91 0.158 2.126 0.202 ;
    LAYER v0 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.694 0.138 1.762 0.182 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.724 0.408 0.788 0.452 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.338 1.026 0.382 ;
      RECT 0.142 0.248 0.182 0.292 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.142 0.518 0.29 0.562 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.518 1.154 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.338 1.35 0.382 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 2.126 0.158 2.194 0.562 ;
  END
END b15cilao5hn1n08x5

MACRO b15cilao5hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilao5hn1n12x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 5.09833325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.54916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.518 1.87 0.562 ;
        RECT 1.802 0.338 1.87 0.562 ;
        RECT 1.478 0.248 1.546 0.562 ;
        RECT 0.702 0.248 1.546 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.802 0.358 1.87 0.402 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.562 ;
        RECT 2.666 0.338 2.95 0.382 ;
        RECT 2.666 0.068 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.666 0.138 2.734 0.182 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 2.882 0.138 2.95 0.182 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.594 0.382 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.486 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.774 0.448 2.842 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.586 0.248 1.87 0.292 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.586 0.158 1.654 0.292 ;
        RECT 1.242 0.158 1.654 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.562 ;
      RECT 0.398 0.158 1.134 0.202 ;
      RECT 0.81 0.068 1.694 0.112 ;
      RECT 1.91 0.068 1.978 0.202 ;
      RECT 2.018 0.158 2.086 0.472 ;
    LAYER v0 ;
      RECT 2.558 0.338 2.626 0.382 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.128 0.138 2.192 0.182 ;
      RECT 2.018 0.228 2.086 0.272 ;
      RECT 1.912 0.138 1.976 0.182 ;
      RECT 1.696 0.138 1.76 0.182 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.724 0.408 0.788 0.452 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.338 1.026 0.382 ;
      RECT 0.142 0.248 0.182 0.292 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.142 0.518 0.29 0.562 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.518 1.154 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.338 1.35 0.382 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.978 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.194 0.248 2.45 0.292 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.086 0.428 2.558 0.472 ;
      RECT 2.558 0.248 2.626 0.472 ;
  END
END b15cilao5hn1n12x5

MACRO b15cilao5hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilao5hn1n16x5 0 0 ;
  SIZE 3.132 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.805 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.338 1.978 0.382 ;
        RECT 1.478 0.518 1.762 0.562 ;
        RECT 1.694 0.338 1.762 0.562 ;
        RECT 1.478 0.248 1.546 0.562 ;
        RECT 0.702 0.248 1.546 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.562 ;
        RECT 2.666 0.338 2.95 0.382 ;
        RECT 2.666 0.068 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.666 0.138 2.734 0.182 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 2.882 0.138 2.95 0.182 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.594 0.382 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.486 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.166 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.166 0.022 ;
        RECT 2.99 -0.022 3.058 0.382 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.586 0.248 1.87 0.292 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.586 0.158 1.654 0.292 ;
        RECT 1.242 0.158 1.654 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 2.99 0.138 3.058 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.562 ;
      RECT 0.398 0.158 1.134 0.202 ;
      RECT 0.81 0.068 1.694 0.112 ;
      RECT 1.91 0.068 1.978 0.202 ;
      RECT 2.018 0.158 2.086 0.562 ;
    LAYER v0 ;
      RECT 2.558 0.293 2.626 0.337 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.128 0.138 2.192 0.182 ;
      RECT 2.018 0.223 2.086 0.267 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.912 0.138 1.976 0.182 ;
      RECT 1.696 0.138 1.76 0.182 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.724 0.408 0.788 0.452 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.338 1.026 0.382 ;
      RECT 0.142 0.248 0.182 0.292 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.142 0.518 0.29 0.562 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.518 1.154 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.338 1.35 0.382 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.978 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.194 0.248 2.45 0.292 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.086 0.338 2.234 0.382 ;
      RECT 2.234 0.338 2.302 0.472 ;
      RECT 2.302 0.428 2.558 0.472 ;
      RECT 2.558 0.248 2.626 0.472 ;
  END
END b15cilao5hn1n16x5

MACRO b15cilb01hn1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n02x3 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.248 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.498 1.978 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.158 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.203 2.734 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.478 0.4705 1.546 0.5145 ;
        RECT 2.018 0.403 2.086 0.447 ;
        RECT 2.342 0.403 2.41 0.447 ;
        RECT 2.774 0.428 2.842 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.018 -0.022 2.086 0.292 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 2.018 0.203 2.086 0.247 ;
        RECT 2.774 0.203 2.842 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 2.126 0.158 2.194 0.472 ;
    LAYER v0 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.403 2.194 0.447 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.2035 1.87 0.2475 ;
      RECT 1.802 0.403 1.87 0.447 ;
      RECT 1.586 0.171 1.654 0.215 ;
      RECT 1.586 0.4705 1.654 0.5145 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.508 0.408 0.572 0.452 ;
      RECT 0.398 0.293 0.466 0.337 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.068 1.438 0.112 ;
      RECT 0.574 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.654 0.068 1.89 0.112 ;
      RECT 2.194 0.158 2.45 0.202 ;
      RECT 2.45 0.068 2.518 0.202 ;
      RECT 2.518 0.068 2.734 0.112 ;
  END
END b15cilb01hn1n02x3

MACRO b15cilb01hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n02x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37071425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.248 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.498 1.978 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.158 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.203 2.734 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.478 0.4705 1.546 0.5145 ;
        RECT 2.018 0.403 2.086 0.447 ;
        RECT 2.342 0.403 2.41 0.447 ;
        RECT 2.774 0.428 2.842 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.018 -0.022 2.086 0.292 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 2.018 0.203 2.086 0.247 ;
        RECT 2.774 0.203 2.842 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.158 1.87 0.472 ;
    LAYER v0 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.403 2.194 0.447 ;
      RECT 1.802 0.2035 1.87 0.2475 ;
      RECT 1.802 0.403 1.87 0.447 ;
      RECT 1.586 0.171 1.654 0.215 ;
      RECT 1.586 0.4705 1.654 0.5145 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.508 0.408 0.572 0.452 ;
      RECT 0.398 0.293 0.466 0.337 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.068 1.438 0.112 ;
      RECT 0.574 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 2.194 0.158 2.45 0.202 ;
      RECT 2.45 0.068 2.518 0.202 ;
      RECT 2.518 0.068 2.734 0.112 ;
  END
END b15cilb01hn1n02x5

MACRO b15cilb01hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n03x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37071425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.498 2.302 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.158 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.4675 2.734 0.5115 ;
        RECT 2.666 0.203 2.734 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.478 0.4705 1.546 0.5145 ;
        RECT 2.018 0.473 2.086 0.517 ;
        RECT 2.342 0.403 2.41 0.447 ;
        RECT 2.774 0.4675 2.842 0.5115 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.882 -0.022 2.95 0.292 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.882 0.203 2.95 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 2.126 0.158 2.194 0.472 ;
    LAYER v0 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.383 2.194 0.427 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.802 0.2035 1.87 0.2475 ;
      RECT 1.802 0.403 1.87 0.447 ;
      RECT 1.586 0.171 1.654 0.215 ;
      RECT 1.586 0.4705 1.654 0.5145 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.068 1.438 0.112 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.654 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.202 ;
      RECT 1.978 0.158 2.018 0.202 ;
      RECT 2.018 0.158 2.086 0.382 ;
      RECT 2.194 0.158 2.45 0.202 ;
      RECT 2.45 0.068 2.518 0.202 ;
      RECT 2.518 0.068 2.842 0.112 ;
  END
END b15cilb01hn1n03x5

MACRO b15cilb01hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n04x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37071425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.498 2.302 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.158 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.4725 2.95 0.5165 ;
        RECT 2.882 0.203 2.95 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.478 0.4705 1.546 0.5145 ;
        RECT 2.018 0.473 2.086 0.517 ;
        RECT 2.342 0.403 2.41 0.447 ;
        RECT 2.558 0.428 2.626 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.666 0.048 2.734 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 2.126 0.158 2.194 0.472 ;
    LAYER v0 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.383 2.194 0.427 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.802 0.2035 1.87 0.2475 ;
      RECT 1.802 0.403 1.87 0.447 ;
      RECT 1.586 0.171 1.654 0.215 ;
      RECT 1.586 0.4705 1.654 0.5145 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.068 1.438 0.112 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.654 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.202 ;
      RECT 1.978 0.158 2.018 0.202 ;
      RECT 2.018 0.158 2.086 0.382 ;
      RECT 2.194 0.158 2.666 0.202 ;
      RECT 2.666 0.158 2.734 0.382 ;
  END
END b15cilb01hn1n04x5

MACRO b15cilb01hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n06x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37071425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.498 2.302 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06732 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.158 2.95 0.562 ;
        RECT 2.558 0.338 2.95 0.382 ;
        RECT 2.558 0.158 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.4715 2.626 0.5155 ;
        RECT 2.558 0.203 2.626 0.247 ;
        RECT 2.882 0.4725 2.95 0.5165 ;
        RECT 2.882 0.203 2.95 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.478 0.4705 1.546 0.5145 ;
        RECT 2.018 0.473 2.086 0.517 ;
        RECT 2.342 0.403 2.41 0.447 ;
        RECT 2.666 0.4715 2.734 0.5155 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.666 0.203 2.734 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 2.126 0.158 2.194 0.472 ;
    LAYER v0 ;
      RECT 2.45 0.293 2.518 0.337 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.383 2.194 0.427 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.802 0.2035 1.87 0.2475 ;
      RECT 1.802 0.403 1.87 0.447 ;
      RECT 1.586 0.171 1.654 0.215 ;
      RECT 1.586 0.4705 1.654 0.5145 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.068 1.438 0.112 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.654 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.202 ;
      RECT 1.978 0.158 2.018 0.202 ;
      RECT 2.018 0.158 2.086 0.382 ;
      RECT 2.194 0.158 2.45 0.202 ;
      RECT 2.45 0.158 2.518 0.382 ;
  END
END b15cilb01hn1n06x5

MACRO b15cilb01hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n08x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37071425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.498 2.302 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.158 2.95 0.562 ;
        RECT 2.558 0.338 2.95 0.382 ;
        RECT 2.558 0.158 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.4715 2.626 0.5155 ;
        RECT 2.558 0.203 2.626 0.247 ;
        RECT 2.882 0.4725 2.95 0.5165 ;
        RECT 2.882 0.203 2.95 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.478 0.4705 1.546 0.5145 ;
        RECT 2.018 0.473 2.086 0.517 ;
        RECT 2.342 0.403 2.41 0.447 ;
        RECT 2.666 0.4715 2.734 0.5155 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.666 0.203 2.734 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 2.126 0.158 2.194 0.472 ;
    LAYER v0 ;
      RECT 2.45 0.293 2.518 0.337 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.383 2.194 0.427 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.802 0.2035 1.87 0.2475 ;
      RECT 1.802 0.403 1.87 0.447 ;
      RECT 1.586 0.171 1.654 0.215 ;
      RECT 1.586 0.4705 1.654 0.5145 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.068 1.438 0.112 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.654 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.202 ;
      RECT 1.978 0.158 2.018 0.202 ;
      RECT 2.018 0.158 2.086 0.382 ;
      RECT 2.194 0.158 2.45 0.202 ;
      RECT 2.45 0.158 2.518 0.382 ;
  END
END b15cilb01hn1n08x5

MACRO b15cilb01hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n12x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.248 2.646 0.292 ;
        RECT 1.91 0.338 2.518 0.382 ;
        RECT 2.45 0.248 2.518 0.382 ;
        RECT 1.91 0.338 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.498 1.978 0.542 ;
        RECT 2.558 0.248 2.626 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.068 3.382 0.562 ;
        RECT 2.99 0.338 3.382 0.382 ;
        RECT 2.99 0.068 3.058 0.562 ;
      LAYER v0 ;
        RECT 2.99 0.4715 3.058 0.5155 ;
        RECT 2.99 0.113 3.058 0.157 ;
        RECT 3.314 0.4725 3.382 0.5165 ;
        RECT 3.314 0.113 3.382 0.157 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.45 0.538 2.518 0.582 ;
        RECT 2.666 0.538 2.734 0.582 ;
        RECT 2.882 0.4715 2.95 0.5155 ;
        RECT 3.098 0.4715 3.166 0.5155 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.234 0.048 2.302 0.092 ;
        RECT 2.882 0.113 2.95 0.157 ;
        RECT 3.098 0.113 3.166 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 2.322 0.428 2.774 0.472 ;
      RECT 2.018 0.158 2.646 0.202 ;
    LAYER v0 ;
      RECT 2.774 0.248 2.842 0.292 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.586 0.203 1.654 0.247 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.068 1.438 0.112 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.654 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.292 ;
      RECT 1.978 0.248 2.322 0.292 ;
      RECT 2.43 0.068 2.774 0.112 ;
      RECT 2.774 0.068 2.842 0.472 ;
  END
END b15cilb01hn1n12x5

MACRO b15cilb01hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n16x5 0 0 ;
  SIZE 3.564 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.248 2.646 0.292 ;
        RECT 1.91 0.338 2.518 0.382 ;
        RECT 2.45 0.248 2.518 0.382 ;
        RECT 1.91 0.338 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.498 1.978 0.542 ;
        RECT 2.558 0.248 2.626 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.068 3.274 0.562 ;
        RECT 2.99 0.338 3.274 0.382 ;
        RECT 2.99 0.068 3.058 0.562 ;
      LAYER v0 ;
        RECT 2.99 0.4715 3.058 0.5155 ;
        RECT 2.99 0.113 3.058 0.157 ;
        RECT 3.206 0.4715 3.274 0.5155 ;
        RECT 3.206 0.113 3.274 0.157 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.45 0.538 2.518 0.582 ;
        RECT 2.666 0.538 2.734 0.582 ;
        RECT 2.882 0.4715 2.95 0.5155 ;
        RECT 3.098 0.4715 3.166 0.5155 ;
        RECT 3.314 0.4715 3.382 0.5155 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.598 0.022 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.234 0.048 2.302 0.092 ;
        RECT 2.882 0.113 2.95 0.157 ;
        RECT 3.098 0.113 3.166 0.157 ;
        RECT 3.314 0.113 3.382 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 2.322 0.428 2.774 0.472 ;
      RECT 2.018 0.158 2.646 0.202 ;
    LAYER v0 ;
      RECT 2.774 0.248 2.842 0.292 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.586 0.203 1.654 0.247 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.068 1.438 0.112 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.654 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.292 ;
      RECT 1.978 0.248 2.322 0.292 ;
      RECT 2.43 0.068 2.774 0.112 ;
      RECT 2.774 0.068 2.842 0.472 ;
  END
END b15cilb01hn1n16x5

MACRO b15cilb01hn1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n24x5 0 0 ;
  SIZE 3.888 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.980625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0189 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6684615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.248 2.95 0.562 ;
        RECT 2.666 0.248 2.95 0.292 ;
      LAYER v0 ;
        RECT 2.774 0.248 2.842 0.292 ;
        RECT 2.882 0.383 2.95 0.427 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.428 3.834 0.472 ;
        RECT 3.638 0.248 3.706 0.472 ;
        RECT 3.098 0.248 3.706 0.292 ;
        RECT 3.53 0.068 3.598 0.292 ;
        RECT 3.314 0.068 3.382 0.292 ;
        RECT 3.098 0.068 3.166 0.292 ;
      LAYER v0 ;
        RECT 3.098 0.428 3.166 0.472 ;
        RECT 3.098 0.138 3.166 0.182 ;
        RECT 3.314 0.428 3.382 0.472 ;
        RECT 3.314 0.138 3.382 0.182 ;
        RECT 3.53 0.428 3.598 0.472 ;
        RECT 3.53 0.138 3.598 0.182 ;
        RECT 3.746 0.428 3.814 0.472 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.922 0.652 ;
        RECT 3.638 0.518 3.706 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 3.206 0.518 3.274 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.478 0.4705 1.546 0.5145 ;
        RECT 1.694 0.4705 1.762 0.5145 ;
        RECT 2.126 0.473 2.194 0.517 ;
        RECT 2.45 0.473 2.518 0.517 ;
        RECT 2.774 0.383 2.842 0.427 ;
        RECT 2.992 0.538 3.056 0.582 ;
        RECT 3.208 0.538 3.272 0.582 ;
        RECT 3.424 0.538 3.488 0.582 ;
        RECT 3.64 0.538 3.704 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.922 0.022 ;
        RECT 3.638 -0.022 3.706 0.112 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 3.206 -0.022 3.274 0.112 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 2.126 0.048 2.194 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
        RECT 3.208 0.048 3.272 0.092 ;
        RECT 3.424 0.048 3.488 0.092 ;
        RECT 3.64 0.048 3.704 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.91 0.248 1.978 0.562 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 3.746 0.248 3.814 0.382 ;
    LAYER v0 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 3.098 0.338 3.166 0.382 ;
      RECT 2.774 0.068 2.842 0.112 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.558 0.473 2.626 0.517 ;
      RECT 2.452 0.1445 2.516 0.1885 ;
      RECT 2.234 0.1445 2.302 0.1885 ;
      RECT 2.234 0.473 2.302 0.517 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 1.91 0.29 1.978 0.334 ;
      RECT 1.91 0.4705 1.978 0.5145 ;
      RECT 1.586 0.1365 1.654 0.1805 ;
      RECT 1.586 0.4705 1.654 0.5145 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.068 1.438 0.112 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.654 0.248 1.802 0.292 ;
      RECT 1.802 0.158 1.87 0.292 ;
      RECT 1.87 0.158 2.126 0.202 ;
      RECT 2.126 0.158 2.194 0.382 ;
      RECT 2.302 0.248 2.45 0.292 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.518 0.068 2.95 0.112 ;
      RECT 2.302 0.338 2.558 0.382 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 2.626 0.158 2.99 0.202 ;
      RECT 2.99 0.158 3.058 0.382 ;
      RECT 3.058 0.338 3.402 0.382 ;
  END
END b15cilb01hn1n24x5

MACRO b15cilb01hn1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n32x5 0 0 ;
  SIZE 4.428 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0189 LAYER m1 ;
      ANTENNAMAXAREACAR 2.18047625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.027 LAYER m1 ;
      ANTENNAMAXAREACAR 7.63166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.248 3.166 0.292 ;
        RECT 2.882 0.248 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.473 2.95 0.517 ;
        RECT 2.99 0.248 3.058 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.294 0.428 4.374 0.472 ;
        RECT 3.314 0.158 4.374 0.202 ;
        RECT 4.178 0.158 4.246 0.472 ;
        RECT 3.962 0.158 4.03 0.472 ;
      LAYER v0 ;
        RECT 3.422 0.428 3.49 0.472 ;
        RECT 3.422 0.158 3.49 0.202 ;
        RECT 3.638 0.428 3.706 0.472 ;
        RECT 3.638 0.158 3.706 0.202 ;
        RECT 3.854 0.428 3.922 0.472 ;
        RECT 3.854 0.158 3.922 0.202 ;
        RECT 4.07 0.428 4.138 0.472 ;
        RECT 4.07 0.158 4.138 0.202 ;
        RECT 4.286 0.428 4.354 0.472 ;
        RECT 4.286 0.158 4.354 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.462 0.652 ;
        RECT 4.178 0.518 4.246 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.478 0.4705 1.546 0.5145 ;
        RECT 1.694 0.4705 1.762 0.5145 ;
        RECT 2.126 0.473 2.194 0.517 ;
        RECT 2.45 0.473 2.518 0.517 ;
        RECT 2.774 0.473 2.842 0.517 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 4.18 0.538 4.244 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.462 0.022 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.748 0.048 3.812 0.092 ;
        RECT 3.964 0.048 4.028 0.092 ;
        RECT 4.18 0.048 4.244 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.91 0.248 1.978 0.562 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 4.286 0.248 4.354 0.382 ;
    LAYER v0 ;
      RECT 3.638 0.338 3.706 0.382 ;
      RECT 3.422 0.338 3.49 0.382 ;
      RECT 3.098 0.158 3.166 0.202 ;
      RECT 2.99 0.068 3.058 0.112 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.668 0.1445 2.732 0.1885 ;
      RECT 2.558 0.473 2.626 0.517 ;
      RECT 2.45 0.1445 2.518 0.1885 ;
      RECT 2.234 0.1445 2.302 0.1885 ;
      RECT 2.234 0.473 2.302 0.517 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 1.91 0.29 1.978 0.334 ;
      RECT 1.91 0.4705 1.978 0.5145 ;
      RECT 1.586 0.1365 1.654 0.1805 ;
      RECT 1.586 0.4705 1.654 0.5145 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.068 1.438 0.112 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.654 0.248 1.802 0.292 ;
      RECT 1.802 0.158 1.87 0.292 ;
      RECT 1.87 0.158 2.126 0.202 ;
      RECT 2.126 0.158 2.194 0.382 ;
      RECT 2.302 0.248 2.45 0.292 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.518 0.248 2.666 0.292 ;
      RECT 2.666 0.068 2.734 0.292 ;
      RECT 2.734 0.068 3.166 0.112 ;
      RECT 2.302 0.338 2.558 0.382 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 2.626 0.338 2.774 0.382 ;
      RECT 2.774 0.158 2.842 0.382 ;
      RECT 2.842 0.158 3.206 0.202 ;
      RECT 3.206 0.158 3.274 0.382 ;
      RECT 3.274 0.338 3.814 0.382 ;
  END
END b15cilb01hn1n32x5

MACRO b15cilb01hn1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n48x5 0 0 ;
  SIZE 5.292 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0261 LAYER m1 ;
      ANTENNAMAXAREACAR 1.0268445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0342 LAYER m1 ;
      ANTENNAMAXAREACAR 0.80222225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.338 3.598 0.382 ;
        RECT 2.342 0.338 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.338 2.626 0.382 ;
        RECT 2.99 0.338 3.058 0.382 ;
        RECT 3.206 0.338 3.274 0.382 ;
        RECT 3.422 0.338 3.49 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16524 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.428 5.238 0.472 ;
        RECT 3.746 0.158 5.238 0.202 ;
        RECT 5.042 0.158 5.11 0.472 ;
        RECT 4.826 0.158 4.894 0.472 ;
        RECT 4.61 0.158 4.678 0.472 ;
      LAYER v0 ;
        RECT 3.854 0.428 3.922 0.472 ;
        RECT 3.854 0.158 3.922 0.202 ;
        RECT 4.07 0.428 4.138 0.472 ;
        RECT 4.07 0.158 4.138 0.202 ;
        RECT 4.286 0.428 4.354 0.472 ;
        RECT 4.286 0.158 4.354 0.202 ;
        RECT 4.502 0.428 4.57 0.472 ;
        RECT 4.502 0.158 4.57 0.202 ;
        RECT 4.718 0.428 4.786 0.472 ;
        RECT 4.718 0.158 4.786 0.202 ;
        RECT 4.934 0.428 5.002 0.472 ;
        RECT 4.934 0.158 5.002 0.202 ;
        RECT 5.15 0.428 5.218 0.472 ;
        RECT 5.15 0.158 5.218 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68158725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.19277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.268 0.574 0.312 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.326 0.652 ;
        RECT 5.042 0.518 5.11 0.652 ;
        RECT 4.826 0.518 4.894 0.652 ;
        RECT 4.61 0.518 4.678 0.652 ;
        RECT 4.394 0.518 4.462 0.652 ;
        RECT 4.178 0.518 4.246 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 3.206 0.518 3.274 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 1.262 0.4705 1.33 0.5145 ;
        RECT 1.802 0.4705 1.87 0.5145 ;
        RECT 2.018 0.4705 2.086 0.5145 ;
        RECT 2.558 0.538 2.626 0.582 ;
        RECT 2.774 0.538 2.842 0.582 ;
        RECT 2.99 0.538 3.058 0.582 ;
        RECT 3.206 0.538 3.274 0.582 ;
        RECT 3.422 0.538 3.49 0.582 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 4.18 0.538 4.244 0.582 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 4.612 0.538 4.676 0.582 ;
        RECT 4.828 0.538 4.892 0.582 ;
        RECT 5.044 0.538 5.108 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.326 0.022 ;
        RECT 5.042 -0.022 5.11 0.112 ;
        RECT 4.826 -0.022 4.894 0.112 ;
        RECT 4.61 -0.022 4.678 0.112 ;
        RECT 4.394 -0.022 4.462 0.112 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
        RECT 3.748 0.048 3.812 0.092 ;
        RECT 3.964 0.048 4.028 0.092 ;
        RECT 4.18 0.048 4.244 0.092 ;
        RECT 4.396 0.048 4.46 0.092 ;
        RECT 4.612 0.048 4.676 0.092 ;
        RECT 4.828 0.048 4.892 0.092 ;
        RECT 5.044 0.048 5.108 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.398 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 0.722 0.428 0.938 0.472 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.558 0.158 3.206 0.202 ;
      RECT 3.098 0.248 3.314 0.292 ;
      RECT 5.15 0.248 5.218 0.382 ;
    LAYER v0 ;
      RECT 4.394 0.338 4.462 0.382 ;
      RECT 4.178 0.338 4.246 0.382 ;
      RECT 3.854 0.338 3.922 0.382 ;
      RECT 3.53 0.068 3.598 0.112 ;
      RECT 3.53 0.428 3.598 0.472 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.314 0.068 3.382 0.112 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 3.098 0.158 3.166 0.202 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.882 0.248 2.95 0.292 ;
      RECT 2.882 0.428 2.95 0.472 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.4705 2.194 0.5145 ;
      RECT 1.91 0.1365 1.978 0.1805 ;
      RECT 1.91 0.4705 1.978 0.5145 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.203 1.006 0.247 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.616 0.088 0.68 0.132 ;
      RECT 0.616 0.3855 0.68 0.4295 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.4 0.3855 0.464 0.4295 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.518 0.682 0.562 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 0.79 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.248 1.37 0.292 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.438 0.068 1.762 0.112 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.006 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.518 1.586 0.562 ;
      RECT 1.586 0.158 1.654 0.562 ;
      RECT 1.654 0.158 1.802 0.202 ;
      RECT 1.802 0.158 1.87 0.382 ;
      RECT 1.978 0.248 2.126 0.292 ;
      RECT 2.126 0.068 2.194 0.562 ;
      RECT 2.194 0.248 2.97 0.292 ;
      RECT 3.206 0.068 3.274 0.202 ;
      RECT 3.274 0.068 3.706 0.112 ;
      RECT 3.314 0.158 3.382 0.292 ;
      RECT 2.558 0.428 3.638 0.472 ;
      RECT 3.382 0.158 3.638 0.202 ;
      RECT 3.638 0.158 3.706 0.472 ;
      RECT 3.706 0.338 4.57 0.382 ;
  END
END b15cilb01hn1n48x5

MACRO b15cilb01hn1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n64x5 0 0 ;
  SIZE 6.156 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0324 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0414 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.248 4.03 0.292 ;
        RECT 2.558 0.338 3.382 0.382 ;
        RECT 3.314 0.248 3.382 0.382 ;
        RECT 2.558 0.338 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 3.53 0.248 3.598 0.292 ;
        RECT 3.854 0.248 3.922 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.428 6.102 0.472 ;
        RECT 4.178 0.158 6.102 0.202 ;
        RECT 5.906 0.158 5.974 0.472 ;
        RECT 5.258 0.158 5.326 0.472 ;
        RECT 5.042 0.158 5.11 0.472 ;
        RECT 4.826 0.158 4.894 0.472 ;
        RECT 4.178 0.158 4.246 0.472 ;
      LAYER v0 ;
        RECT 4.286 0.428 4.354 0.472 ;
        RECT 4.286 0.158 4.354 0.202 ;
        RECT 4.502 0.428 4.57 0.472 ;
        RECT 4.502 0.158 4.57 0.202 ;
        RECT 4.718 0.428 4.786 0.472 ;
        RECT 4.718 0.158 4.786 0.202 ;
        RECT 4.934 0.428 5.002 0.472 ;
        RECT 4.934 0.158 5.002 0.202 ;
        RECT 5.15 0.428 5.218 0.472 ;
        RECT 5.15 0.158 5.218 0.202 ;
        RECT 5.366 0.428 5.434 0.472 ;
        RECT 5.366 0.158 5.434 0.202 ;
        RECT 5.582 0.428 5.65 0.472 ;
        RECT 5.582 0.158 5.65 0.202 ;
        RECT 5.798 0.428 5.866 0.472 ;
        RECT 5.798 0.158 5.866 0.202 ;
        RECT 6.014 0.428 6.082 0.472 ;
        RECT 6.014 0.158 6.082 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 0.477111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.268 0.574 0.312 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.19 0.652 ;
        RECT 5.906 0.518 5.974 0.652 ;
        RECT 5.69 0.518 5.758 0.652 ;
        RECT 5.474 0.518 5.542 0.652 ;
        RECT 5.258 0.518 5.326 0.652 ;
        RECT 5.042 0.518 5.11 0.652 ;
        RECT 4.826 0.518 4.894 0.652 ;
        RECT 4.61 0.518 4.678 0.652 ;
        RECT 4.394 0.518 4.462 0.652 ;
        RECT 4.178 0.518 4.246 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 1.262 0.4705 1.33 0.5145 ;
        RECT 1.802 0.4705 1.87 0.5145 ;
        RECT 2.018 0.4705 2.086 0.5145 ;
        RECT 2.234 0.4705 2.302 0.5145 ;
        RECT 2.666 0.538 2.734 0.582 ;
        RECT 2.882 0.538 2.95 0.582 ;
        RECT 3.098 0.538 3.166 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 4.18 0.538 4.244 0.582 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 4.612 0.538 4.676 0.582 ;
        RECT 4.828 0.538 4.892 0.582 ;
        RECT 5.044 0.538 5.108 0.582 ;
        RECT 5.26 0.538 5.324 0.582 ;
        RECT 5.476 0.538 5.54 0.582 ;
        RECT 5.692 0.538 5.756 0.582 ;
        RECT 5.908 0.538 5.972 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.19 0.022 ;
        RECT 5.906 -0.022 5.974 0.112 ;
        RECT 5.69 -0.022 5.758 0.112 ;
        RECT 5.474 -0.022 5.542 0.112 ;
        RECT 5.258 -0.022 5.326 0.112 ;
        RECT 5.042 -0.022 5.11 0.112 ;
        RECT 4.826 -0.022 4.894 0.112 ;
        RECT 4.61 -0.022 4.678 0.112 ;
        RECT 4.394 -0.022 4.462 0.112 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.018 0.1365 2.086 0.1805 ;
        RECT 2.234 0.1365 2.302 0.1805 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.316 0.048 3.38 0.092 ;
        RECT 4.18 0.048 4.244 0.092 ;
        RECT 4.396 0.048 4.46 0.092 ;
        RECT 4.612 0.048 4.676 0.092 ;
        RECT 4.828 0.048 4.892 0.092 ;
        RECT 5.044 0.048 5.108 0.092 ;
        RECT 5.26 0.048 5.324 0.092 ;
        RECT 5.476 0.048 5.54 0.092 ;
        RECT 5.692 0.048 5.756 0.092 ;
        RECT 5.908 0.048 5.972 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.398 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 0.722 0.428 0.938 0.472 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.666 0.428 3.422 0.472 ;
      RECT 2.666 0.158 4.03 0.202 ;
      RECT 4.286 0.248 4.786 0.292 ;
      RECT 5.366 0.248 5.866 0.292 ;
      RECT 6.014 0.248 6.082 0.382 ;
    LAYER v0 ;
      RECT 5.69 0.248 5.758 0.292 ;
      RECT 5.474 0.248 5.542 0.292 ;
      RECT 4.61 0.248 4.678 0.292 ;
      RECT 4.394 0.248 4.462 0.292 ;
      RECT 4.07 0.246 4.138 0.29 ;
      RECT 3.962 0.068 4.03 0.112 ;
      RECT 3.854 0.158 3.922 0.202 ;
      RECT 3.854 0.424 3.922 0.468 ;
      RECT 3.746 0.068 3.814 0.112 ;
      RECT 3.638 0.158 3.706 0.202 ;
      RECT 3.638 0.424 3.706 0.468 ;
      RECT 3.53 0.068 3.598 0.112 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.99 0.248 3.058 0.292 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.248 2.842 0.292 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.126 0.1365 2.194 0.1805 ;
      RECT 2.126 0.4705 2.194 0.5145 ;
      RECT 1.91 0.1365 1.978 0.1805 ;
      RECT 1.91 0.4705 1.978 0.5145 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.203 1.006 0.247 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.616 0.088 0.68 0.132 ;
      RECT 0.616 0.3855 0.68 0.4295 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.4 0.3855 0.464 0.4295 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.518 0.682 0.562 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 0.79 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.248 1.37 0.292 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.438 0.068 1.762 0.112 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.006 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.518 1.586 0.562 ;
      RECT 1.586 0.158 1.654 0.562 ;
      RECT 1.654 0.158 1.802 0.202 ;
      RECT 1.802 0.158 1.87 0.382 ;
      RECT 1.978 0.248 2.126 0.292 ;
      RECT 2.126 0.068 2.194 0.562 ;
      RECT 2.194 0.248 3.078 0.292 ;
      RECT 3.422 0.338 3.49 0.472 ;
      RECT 3.49 0.338 3.638 0.382 ;
      RECT 3.638 0.338 3.706 0.562 ;
      RECT 3.706 0.338 3.854 0.382 ;
      RECT 3.854 0.338 3.922 0.562 ;
      RECT 3.922 0.518 4.07 0.562 ;
      RECT 3.422 0.068 4.07 0.112 ;
      RECT 4.07 0.068 4.138 0.562 ;
  END
END b15cilb01hn1n64x5

MACRO b15cilb01hn1n80x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb01hn1n80x5 0 0 ;
  SIZE 7.128 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0405 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0558 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.248 5.002 0.292 ;
        RECT 3.098 0.338 4.462 0.382 ;
        RECT 4.394 0.248 4.462 0.382 ;
        RECT 3.098 0.338 3.166 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.338 3.274 0.382 ;
        RECT 3.854 0.338 3.922 0.382 ;
        RECT 4.07 0.338 4.138 0.382 ;
        RECT 4.502 0.248 4.57 0.292 ;
        RECT 4.718 0.248 4.786 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.26622 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.428 7.054 0.472 ;
        RECT 6.986 0.158 7.054 0.472 ;
        RECT 5.69 0.158 7.054 0.202 ;
        RECT 6.338 0.158 6.406 0.472 ;
        RECT 6.122 0.158 6.19 0.472 ;
        RECT 5.906 0.158 5.974 0.472 ;
        RECT 5.69 0.158 5.758 0.472 ;
        RECT 5.15 0.248 5.758 0.292 ;
        RECT 5.474 0.248 5.542 0.472 ;
        RECT 5.258 0.248 5.326 0.472 ;
        RECT 5.15 0.068 5.218 0.292 ;
      LAYER v0 ;
        RECT 4.718 0.428 4.786 0.472 ;
        RECT 4.934 0.428 5.002 0.472 ;
        RECT 5.15 0.428 5.218 0.472 ;
        RECT 5.15 0.138 5.218 0.182 ;
        RECT 5.366 0.428 5.434 0.472 ;
        RECT 5.366 0.248 5.434 0.292 ;
        RECT 5.582 0.428 5.65 0.472 ;
        RECT 5.582 0.248 5.65 0.292 ;
        RECT 5.798 0.428 5.866 0.472 ;
        RECT 5.798 0.158 5.866 0.202 ;
        RECT 6.014 0.428 6.082 0.472 ;
        RECT 6.014 0.158 6.082 0.202 ;
        RECT 6.23 0.428 6.298 0.472 ;
        RECT 6.23 0.158 6.298 0.202 ;
        RECT 6.446 0.428 6.514 0.472 ;
        RECT 6.446 0.158 6.514 0.202 ;
        RECT 6.662 0.428 6.73 0.472 ;
        RECT 6.662 0.158 6.73 0.202 ;
        RECT 6.878 0.428 6.946 0.472 ;
        RECT 6.878 0.158 6.946 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5301235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.378 0.292 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0252 LAYER m1 ;
      ANTENNAMAXAREACAR 0.666508 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 1.09777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.268 0.898 0.312 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 7.162 0.652 ;
        RECT 6.986 0.518 7.054 0.652 ;
        RECT 6.77 0.518 6.838 0.652 ;
        RECT 6.554 0.518 6.622 0.652 ;
        RECT 6.338 0.518 6.406 0.652 ;
        RECT 6.122 0.518 6.19 0.652 ;
        RECT 5.906 0.518 5.974 0.652 ;
        RECT 5.69 0.518 5.758 0.652 ;
        RECT 5.474 0.518 5.542 0.652 ;
        RECT 5.258 0.518 5.326 0.652 ;
        RECT 5.042 0.518 5.11 0.652 ;
        RECT 4.826 0.518 4.894 0.652 ;
        RECT 4.502 0.518 4.57 0.652 ;
        RECT 4.286 0.518 4.354 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.854 0.518 3.922 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.586 0.4705 1.654 0.5145 ;
        RECT 2.126 0.4705 2.194 0.5145 ;
        RECT 2.342 0.4705 2.41 0.5145 ;
        RECT 2.558 0.4705 2.626 0.5145 ;
        RECT 2.774 0.4705 2.842 0.5145 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
        RECT 3.856 0.538 3.92 0.582 ;
        RECT 4.07 0.538 4.138 0.582 ;
        RECT 4.288 0.538 4.352 0.582 ;
        RECT 4.504 0.538 4.568 0.582 ;
        RECT 4.828 0.538 4.892 0.582 ;
        RECT 5.044 0.538 5.108 0.582 ;
        RECT 5.26 0.538 5.324 0.582 ;
        RECT 5.476 0.538 5.54 0.582 ;
        RECT 5.692 0.538 5.756 0.582 ;
        RECT 5.908 0.538 5.972 0.582 ;
        RECT 6.124 0.538 6.188 0.582 ;
        RECT 6.34 0.538 6.404 0.582 ;
        RECT 6.556 0.538 6.62 0.582 ;
        RECT 6.772 0.538 6.836 0.582 ;
        RECT 6.988 0.538 7.052 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 7.162 0.022 ;
        RECT 6.986 -0.022 7.054 0.112 ;
        RECT 6.77 -0.022 6.838 0.112 ;
        RECT 6.554 -0.022 6.622 0.112 ;
        RECT 6.338 -0.022 6.406 0.112 ;
        RECT 6.122 -0.022 6.19 0.112 ;
        RECT 5.906 -0.022 5.974 0.112 ;
        RECT 5.69 -0.022 5.758 0.112 ;
        RECT 5.474 -0.022 5.542 0.112 ;
        RECT 5.258 -0.022 5.326 0.112 ;
        RECT 4.07 -0.022 4.138 0.112 ;
        RECT 3.854 -0.022 3.922 0.112 ;
        RECT 3.638 -0.022 3.706 0.112 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 3.206 -0.022 3.274 0.112 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.342 0.1365 2.41 0.1805 ;
        RECT 2.558 0.1365 2.626 0.1805 ;
        RECT 2.774 0.1365 2.842 0.1805 ;
        RECT 3.208 0.048 3.272 0.092 ;
        RECT 3.424 0.048 3.488 0.092 ;
        RECT 3.64 0.048 3.704 0.092 ;
        RECT 3.856 0.048 3.92 0.092 ;
        RECT 4.072 0.048 4.136 0.092 ;
        RECT 5.26 0.048 5.324 0.092 ;
        RECT 5.476 0.048 5.54 0.092 ;
        RECT 5.692 0.048 5.756 0.092 ;
        RECT 5.908 0.048 5.972 0.092 ;
        RECT 6.124 0.048 6.188 0.092 ;
        RECT 6.34 0.048 6.404 0.092 ;
        RECT 6.556 0.048 6.62 0.092 ;
        RECT 6.772 0.048 6.836 0.092 ;
        RECT 6.988 0.048 7.052 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 4.916 0.338 6.964 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.506 0.202 ;
      RECT 1.046 0.068 1.114 0.382 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 1.046 0.428 1.262 0.472 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 3.314 0.428 4.502 0.472 ;
      RECT 3.206 0.158 5.002 0.202 ;
      RECT 6.446 0.338 6.946 0.382 ;
    LAYER v1 ;
      RECT 6.774 0.338 6.834 0.382 ;
      RECT 5.046 0.338 5.106 0.382 ;
    LAYER v0 ;
      RECT 6.77 0.338 6.838 0.382 ;
      RECT 6.554 0.338 6.622 0.382 ;
      RECT 4.934 0.068 5.002 0.112 ;
      RECT 4.934 0.338 5.002 0.382 ;
      RECT 4.826 0.158 4.894 0.202 ;
      RECT 4.718 0.068 4.786 0.112 ;
      RECT 4.718 0.338 4.786 0.382 ;
      RECT 4.61 0.158 4.678 0.202 ;
      RECT 4.502 0.068 4.57 0.112 ;
      RECT 4.394 0.158 4.462 0.202 ;
      RECT 4.394 0.428 4.462 0.472 ;
      RECT 4.286 0.068 4.354 0.112 ;
      RECT 4.178 0.158 4.246 0.202 ;
      RECT 4.178 0.428 4.246 0.472 ;
      RECT 3.962 0.158 4.03 0.202 ;
      RECT 3.962 0.248 4.03 0.292 ;
      RECT 3.962 0.428 4.03 0.472 ;
      RECT 3.746 0.158 3.814 0.202 ;
      RECT 3.746 0.248 3.814 0.292 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.53 0.158 3.598 0.202 ;
      RECT 3.53 0.248 3.598 0.292 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.314 0.248 3.382 0.292 ;
      RECT 2.666 0.1365 2.734 0.1805 ;
      RECT 2.666 0.4705 2.734 0.5145 ;
      RECT 2.45 0.1365 2.518 0.1805 ;
      RECT 2.45 0.4705 2.518 0.5145 ;
      RECT 2.234 0.1365 2.302 0.1805 ;
      RECT 2.234 0.4705 2.302 0.5145 ;
      RECT 2.126 0.293 2.194 0.337 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.383 1.87 0.427 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.203 1.33 0.247 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.94 0.088 1.004 0.132 ;
      RECT 0.94 0.3855 1.004 0.4295 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.3855 0.79 0.4295 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.508 0.3855 0.572 0.4295 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.398 0.472 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.518 1.006 0.562 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.79 0.158 0.938 0.202 ;
      RECT 0.938 0.068 1.006 0.472 ;
      RECT 1.114 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.438 0.248 1.694 0.292 ;
      RECT 1.694 0.068 1.762 0.292 ;
      RECT 1.762 0.068 2.086 0.112 ;
      RECT 1.262 0.158 1.33 0.472 ;
      RECT 1.33 0.338 1.694 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.762 0.518 1.91 0.562 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 1.978 0.158 2.126 0.202 ;
      RECT 2.126 0.158 2.194 0.382 ;
      RECT 2.302 0.248 2.45 0.292 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 2.518 0.248 2.666 0.292 ;
      RECT 2.666 0.068 2.734 0.562 ;
      RECT 2.734 0.248 4.05 0.292 ;
      RECT 4.502 0.338 4.57 0.472 ;
      RECT 4.57 0.338 5.042 0.382 ;
      RECT 4.178 0.068 5.042 0.112 ;
      RECT 5.042 0.068 5.11 0.382 ;
  END
END b15cilb01hn1n80x5

MACRO b15cilb05hn1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n02x3 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.562 ;
        RECT 1.478 0.068 1.87 0.112 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.478 0.068 1.546 0.202 ;
        RECT 1.262 0.068 1.33 0.202 ;
        RECT 1.046 0.068 1.33 0.112 ;
        RECT 0.722 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.398 0.068 0.79 0.112 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.802 0.498 1.87 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.158 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.428 2.626 0.472 ;
        RECT 2.558 0.203 2.626 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.37 0.4255 1.438 0.4695 ;
        RECT 1.91 0.403 1.978 0.447 ;
        RECT 2.234 0.403 2.302 0.447 ;
        RECT 2.666 0.428 2.734 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.91 0.203 1.978 0.247 ;
        RECT 2.666 0.203 2.734 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
    LAYER v0 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.403 2.086 0.447 ;
      RECT 1.694 0.178 1.762 0.222 ;
      RECT 1.694 0.403 1.762 0.447 ;
      RECT 1.586 0.178 1.654 0.222 ;
      RECT 1.478 0.4255 1.546 0.4695 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.508 0.408 0.572 0.452 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.574 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.546 0.338 1.586 0.382 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 2.086 0.158 2.342 0.202 ;
      RECT 2.342 0.068 2.41 0.202 ;
      RECT 2.41 0.068 2.626 0.112 ;
  END
END b15cilb05hn1n02x3

MACRO b15cilb05hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n02x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37071425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.562 ;
        RECT 1.478 0.068 1.87 0.112 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.478 0.068 1.546 0.202 ;
        RECT 1.262 0.068 1.33 0.202 ;
        RECT 1.046 0.068 1.33 0.112 ;
        RECT 0.722 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.398 0.068 0.79 0.112 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.802 0.498 1.87 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.158 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.428 2.626 0.472 ;
        RECT 2.558 0.203 2.626 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.91 0.403 1.978 0.447 ;
        RECT 2.234 0.403 2.302 0.447 ;
        RECT 2.666 0.428 2.734 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.91 0.203 1.978 0.247 ;
        RECT 2.666 0.203 2.734 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
    LAYER v0 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.403 2.086 0.447 ;
      RECT 1.694 0.178 1.762 0.222 ;
      RECT 1.694 0.403 1.762 0.447 ;
      RECT 1.586 0.178 1.654 0.222 ;
      RECT 1.478 0.408 1.546 0.452 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.508 0.408 0.572 0.452 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.574 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.546 0.338 1.586 0.382 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 2.086 0.158 2.342 0.202 ;
      RECT 2.342 0.068 2.41 0.202 ;
      RECT 2.41 0.068 2.626 0.112 ;
  END
END b15cilb05hn1n02x5

MACRO b15cilb05hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n03x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37071425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.562 ;
        RECT 1.478 0.068 1.87 0.112 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.478 0.068 1.546 0.202 ;
        RECT 1.262 0.068 1.33 0.202 ;
        RECT 1.046 0.068 1.33 0.112 ;
        RECT 0.722 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.802 0.498 1.87 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.158 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.451 2.518 0.495 ;
        RECT 2.45 0.209 2.518 0.253 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.91 0.403 1.978 0.447 ;
        RECT 2.234 0.403 2.302 0.447 ;
        RECT 2.666 0.451 2.734 0.495 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.91 0.203 1.978 0.247 ;
        RECT 2.666 0.1795 2.734 0.2235 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
    LAYER v0 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.403 2.086 0.447 ;
      RECT 1.694 0.2035 1.762 0.2475 ;
      RECT 1.694 0.403 1.762 0.447 ;
      RECT 1.586 0.2035 1.654 0.2475 ;
      RECT 1.478 0.408 1.546 0.452 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.546 0.338 1.586 0.382 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 2.086 0.158 2.234 0.202 ;
      RECT 2.234 0.068 2.302 0.202 ;
      RECT 2.302 0.068 2.626 0.112 ;
  END
END b15cilb05hn1n03x5

MACRO b15cilb05hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n04x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37071425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.562 ;
        RECT 1.478 0.068 1.87 0.112 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.478 0.068 1.546 0.202 ;
        RECT 1.262 0.068 1.33 0.202 ;
        RECT 1.046 0.068 1.33 0.112 ;
        RECT 0.722 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.802 0.498 1.87 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.158 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.4725 2.842 0.5165 ;
        RECT 2.774 0.203 2.842 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 2.234 0.403 2.302 0.447 ;
        RECT 2.558 0.448 2.626 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.558 0.048 2.626 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
    LAYER v0 ;
      RECT 2.558 0.293 2.626 0.337 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.383 2.086 0.427 ;
      RECT 1.694 0.2035 1.762 0.2475 ;
      RECT 1.694 0.403 1.762 0.447 ;
      RECT 1.586 0.2035 1.654 0.2475 ;
      RECT 1.478 0.408 1.546 0.452 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.546 0.338 1.586 0.382 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 2.086 0.158 2.558 0.202 ;
      RECT 2.558 0.158 2.626 0.382 ;
  END
END b15cilb05hn1n04x5

MACRO b15cilb05hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n06x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37071425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.562 ;
        RECT 1.478 0.068 1.87 0.112 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.478 0.068 1.546 0.202 ;
        RECT 1.262 0.068 1.33 0.202 ;
        RECT 1.046 0.068 1.33 0.112 ;
        RECT 0.722 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.802 0.498 1.87 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 4.62333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 4.62333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.158 2.842 0.562 ;
        RECT 2.45 0.338 2.842 0.382 ;
        RECT 2.45 0.158 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.4715 2.518 0.5155 ;
        RECT 2.45 0.203 2.518 0.247 ;
        RECT 2.774 0.4725 2.842 0.5165 ;
        RECT 2.774 0.203 2.842 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 2.234 0.403 2.302 0.447 ;
        RECT 2.558 0.4715 2.626 0.5155 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.558 -0.022 2.626 0.292 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.558 0.203 2.626 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
    LAYER v0 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.383 2.086 0.427 ;
      RECT 1.694 0.2035 1.762 0.2475 ;
      RECT 1.694 0.403 1.762 0.447 ;
      RECT 1.586 0.2035 1.654 0.2475 ;
      RECT 1.478 0.408 1.546 0.452 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.546 0.338 1.586 0.382 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 2.086 0.158 2.342 0.202 ;
      RECT 2.342 0.158 2.41 0.382 ;
  END
END b15cilb05hn1n06x5

MACRO b15cilb05hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n08x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.39875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37071425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.562 ;
        RECT 1.478 0.068 1.87 0.112 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.478 0.068 1.546 0.202 ;
        RECT 1.262 0.068 1.33 0.202 ;
        RECT 1.046 0.068 1.33 0.112 ;
        RECT 0.722 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.802 0.498 1.87 0.542 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.158 2.842 0.562 ;
        RECT 2.45 0.338 2.842 0.382 ;
        RECT 2.45 0.158 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.4715 2.518 0.5155 ;
        RECT 2.45 0.203 2.518 0.247 ;
        RECT 2.774 0.4725 2.842 0.5165 ;
        RECT 2.774 0.203 2.842 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 2.234 0.403 2.302 0.447 ;
        RECT 2.558 0.4715 2.626 0.5155 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.558 -0.022 2.626 0.292 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.558 0.203 2.626 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
    LAYER v0 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.383 2.086 0.427 ;
      RECT 1.694 0.2035 1.762 0.2475 ;
      RECT 1.694 0.403 1.762 0.447 ;
      RECT 1.586 0.2035 1.654 0.2475 ;
      RECT 1.478 0.408 1.546 0.452 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.546 0.338 1.586 0.382 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 2.086 0.158 2.342 0.202 ;
      RECT 2.342 0.158 2.41 0.382 ;
  END
END b15cilb05hn1n08x5

MACRO b15cilb05hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n12x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.248 2.538 0.292 ;
        RECT 1.478 0.338 2.41 0.382 ;
        RECT 2.342 0.248 2.41 0.382 ;
        RECT 1.802 0.338 1.87 0.562 ;
        RECT 1.478 0.158 1.546 0.382 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.262 0.068 1.33 0.202 ;
        RECT 1.046 0.068 1.33 0.112 ;
        RECT 0.722 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.802 0.498 1.87 0.542 ;
        RECT 2.45 0.248 2.518 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.068 3.274 0.562 ;
        RECT 2.882 0.338 3.274 0.382 ;
        RECT 2.882 0.068 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.4715 2.95 0.5155 ;
        RECT 2.882 0.113 2.95 0.157 ;
        RECT 3.206 0.4725 3.274 0.5165 ;
        RECT 3.206 0.113 3.274 0.157 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.342 0.538 2.41 0.582 ;
        RECT 2.558 0.538 2.626 0.582 ;
        RECT 2.774 0.4715 2.842 0.5155 ;
        RECT 2.99 0.4715 3.058 0.5155 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.126 0.048 2.194 0.092 ;
        RECT 2.774 0.113 2.842 0.157 ;
        RECT 2.99 0.113 3.058 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.586 0.158 1.654 0.292 ;
      RECT 2.214 0.428 2.666 0.472 ;
      RECT 1.91 0.158 2.538 0.202 ;
    LAYER v0 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.342 0.068 2.41 0.112 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.588 0.178 1.652 0.222 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.654 0.248 2.214 0.292 ;
      RECT 2.322 0.068 2.666 0.112 ;
      RECT 2.666 0.068 2.734 0.472 ;
  END
END b15cilb05hn1n12x5

MACRO b15cilb05hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n16x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.248 2.538 0.292 ;
        RECT 1.478 0.338 2.41 0.382 ;
        RECT 2.342 0.248 2.41 0.382 ;
        RECT 1.802 0.338 1.87 0.562 ;
        RECT 1.478 0.158 1.546 0.382 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.262 0.068 1.33 0.202 ;
        RECT 1.046 0.068 1.33 0.112 ;
        RECT 0.722 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.802 0.498 1.87 0.542 ;
        RECT 2.45 0.248 2.518 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.068 3.166 0.562 ;
        RECT 2.882 0.338 3.166 0.382 ;
        RECT 2.882 0.068 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.4715 2.95 0.5155 ;
        RECT 2.882 0.113 2.95 0.157 ;
        RECT 3.098 0.4715 3.166 0.5155 ;
        RECT 3.098 0.113 3.166 0.157 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.342 0.538 2.41 0.582 ;
        RECT 2.558 0.538 2.626 0.582 ;
        RECT 2.774 0.4715 2.842 0.5155 ;
        RECT 2.99 0.4715 3.058 0.5155 ;
        RECT 3.206 0.4715 3.274 0.5155 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.126 0.048 2.194 0.092 ;
        RECT 2.774 0.113 2.842 0.157 ;
        RECT 2.99 0.113 3.058 0.157 ;
        RECT 3.206 0.113 3.274 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.586 0.158 1.654 0.292 ;
      RECT 2.214 0.428 2.666 0.472 ;
      RECT 1.91 0.158 2.538 0.202 ;
    LAYER v0 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.342 0.068 2.41 0.112 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.588 0.178 1.652 0.222 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.654 0.248 2.214 0.292 ;
      RECT 2.322 0.068 2.666 0.112 ;
      RECT 2.666 0.068 2.734 0.472 ;
  END
END b15cilb05hn1n16x5

MACRO b15cilb05hn1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n24x5 0 0 ;
  SIZE 3.78 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 1.64666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.248 2.842 0.292 ;
        RECT 1.802 0.338 2.626 0.382 ;
        RECT 2.558 0.248 2.626 0.382 ;
        RECT 1.802 0.248 1.87 0.382 ;
        RECT 1.262 0.248 1.87 0.292 ;
        RECT 1.262 0.068 1.33 0.292 ;
        RECT 1.046 0.068 1.33 0.112 ;
        RECT 0.722 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.342 0.338 2.41 0.382 ;
        RECT 2.666 0.248 2.734 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.428 3.726 0.472 ;
        RECT 3.53 0.248 3.598 0.472 ;
        RECT 2.99 0.248 3.598 0.292 ;
        RECT 3.422 0.068 3.49 0.292 ;
        RECT 3.206 0.068 3.274 0.292 ;
        RECT 2.99 0.068 3.058 0.292 ;
      LAYER v0 ;
        RECT 2.99 0.428 3.058 0.472 ;
        RECT 2.99 0.138 3.058 0.182 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.206 0.138 3.274 0.182 ;
        RECT 3.422 0.428 3.49 0.472 ;
        RECT 3.422 0.138 3.49 0.182 ;
        RECT 3.638 0.428 3.706 0.472 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.814 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.37 0.383 1.438 0.427 ;
        RECT 1.586 0.4705 1.654 0.5145 ;
        RECT 2.018 0.538 2.086 0.582 ;
        RECT 2.234 0.538 2.302 0.582 ;
        RECT 2.558 0.538 2.626 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.814 0.022 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.316 0.048 3.38 0.092 ;
        RECT 3.532 0.048 3.596 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.37 0.158 1.91 0.202 ;
      RECT 2.018 0.158 2.342 0.202 ;
      RECT 2.018 0.428 2.666 0.472 ;
      RECT 3.638 0.248 3.706 0.382 ;
    LAYER v0 ;
      RECT 3.206 0.338 3.274 0.382 ;
      RECT 2.99 0.338 3.058 0.382 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.4705 1.762 0.5145 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.4705 1.546 0.5145 ;
      RECT 1.262 0.383 1.33 0.427 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.546 0.338 1.694 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.91 0.158 1.978 0.292 ;
      RECT 1.978 0.248 2.41 0.292 ;
      RECT 2.342 0.068 2.41 0.202 ;
      RECT 2.41 0.068 2.842 0.112 ;
      RECT 2.666 0.338 2.734 0.472 ;
      RECT 2.734 0.338 2.882 0.382 ;
      RECT 2.45 0.158 2.882 0.202 ;
      RECT 2.882 0.158 2.95 0.382 ;
      RECT 2.95 0.338 3.294 0.382 ;
  END
END b15cilb05hn1n24x5

MACRO b15cilb05hn1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n32x5 0 0 ;
  SIZE 4.32 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.248 3.058 0.292 ;
        RECT 1.802 0.338 2.734 0.382 ;
        RECT 2.666 0.248 2.734 0.382 ;
        RECT 1.802 0.248 1.87 0.382 ;
        RECT 1.262 0.248 1.87 0.292 ;
        RECT 1.262 0.068 1.33 0.292 ;
        RECT 1.046 0.068 1.33 0.112 ;
        RECT 0.722 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.45 0.338 2.518 0.382 ;
        RECT 2.882 0.248 2.95 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.186 0.428 4.266 0.472 ;
        RECT 3.206 0.158 4.266 0.202 ;
        RECT 4.07 0.158 4.138 0.472 ;
        RECT 3.854 0.158 3.922 0.472 ;
      LAYER v0 ;
        RECT 3.314 0.428 3.382 0.472 ;
        RECT 3.314 0.158 3.382 0.202 ;
        RECT 3.53 0.428 3.598 0.472 ;
        RECT 3.53 0.158 3.598 0.202 ;
        RECT 3.746 0.428 3.814 0.472 ;
        RECT 3.746 0.158 3.814 0.202 ;
        RECT 3.962 0.428 4.03 0.472 ;
        RECT 3.962 0.158 4.03 0.202 ;
        RECT 4.178 0.428 4.246 0.472 ;
        RECT 4.178 0.158 4.246 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.354 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.854 0.518 3.922 0.652 ;
        RECT 3.638 0.518 3.706 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 3.206 0.518 3.274 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.938 0.4705 1.006 0.5145 ;
        RECT 1.37 0.383 1.438 0.427 ;
        RECT 1.586 0.4705 1.654 0.5145 ;
        RECT 2.018 0.538 2.086 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 3.208 0.538 3.272 0.582 ;
        RECT 3.424 0.538 3.488 0.582 ;
        RECT 3.64 0.538 3.704 0.582 ;
        RECT 3.856 0.538 3.92 0.582 ;
        RECT 4.072 0.538 4.136 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.354 0.022 ;
        RECT 4.07 -0.022 4.138 0.112 ;
        RECT 3.854 -0.022 3.922 0.112 ;
        RECT 3.638 -0.022 3.706 0.112 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 3.424 0.048 3.488 0.092 ;
        RECT 3.64 0.048 3.704 0.092 ;
        RECT 3.856 0.048 3.92 0.092 ;
        RECT 4.072 0.048 4.136 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.37 0.158 1.91 0.202 ;
      RECT 2.018 0.428 2.882 0.472 ;
      RECT 2.018 0.158 3.058 0.202 ;
      RECT 4.178 0.248 4.246 0.382 ;
    LAYER v0 ;
      RECT 3.53 0.338 3.598 0.382 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 2.99 0.068 3.058 0.112 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.774 0.068 2.842 0.112 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.342 0.248 2.41 0.292 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.4705 1.762 0.5145 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.4705 1.546 0.5145 ;
      RECT 1.262 0.383 1.33 0.427 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.466 0.562 ;
      RECT 0.25 0.158 0.466 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.546 0.338 1.694 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.91 0.158 1.978 0.292 ;
      RECT 1.978 0.248 2.518 0.292 ;
      RECT 2.882 0.338 2.95 0.472 ;
      RECT 2.95 0.338 3.098 0.382 ;
      RECT 2.666 0.068 3.098 0.112 ;
      RECT 3.098 0.068 3.166 0.382 ;
      RECT 3.166 0.338 3.706 0.382 ;
  END
END b15cilb05hn1n32x5

MACRO b15cilb05hn1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n48x5 0 0 ;
  SIZE 5.184 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0315 LAYER m1 ;
      ANTENNAMAXAREACAR 1.0268445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0387 LAYER m1 ;
      ANTENNAMAXAREACAR 0.80222225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.338 3.49 0.382 ;
        RECT 2.234 0.248 2.302 0.382 ;
        RECT 1.586 0.248 2.302 0.292 ;
        RECT 1.586 0.068 1.654 0.292 ;
        RECT 1.37 0.068 1.654 0.112 ;
        RECT 1.046 0.248 1.438 0.292 ;
        RECT 1.37 0.068 1.438 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 1.114 0.112 ;
        RECT 0.722 0.068 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 2.45 0.338 2.518 0.382 ;
        RECT 2.882 0.338 2.95 0.382 ;
        RECT 3.098 0.338 3.166 0.382 ;
        RECT 3.314 0.338 3.382 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16524 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.428 5.13 0.472 ;
        RECT 3.638 0.158 5.13 0.202 ;
        RECT 4.934 0.158 5.002 0.472 ;
        RECT 4.718 0.158 4.786 0.472 ;
        RECT 4.502 0.158 4.57 0.472 ;
        RECT 4.286 0.158 4.354 0.472 ;
      LAYER v0 ;
        RECT 3.746 0.428 3.814 0.472 ;
        RECT 3.746 0.158 3.814 0.202 ;
        RECT 3.962 0.428 4.03 0.472 ;
        RECT 3.962 0.158 4.03 0.202 ;
        RECT 4.178 0.428 4.246 0.472 ;
        RECT 4.178 0.158 4.246 0.202 ;
        RECT 4.394 0.428 4.462 0.472 ;
        RECT 4.394 0.158 4.462 0.202 ;
        RECT 4.61 0.428 4.678 0.472 ;
        RECT 4.61 0.158 4.678 0.202 ;
        RECT 4.826 0.428 4.894 0.472 ;
        RECT 4.826 0.158 4.894 0.202 ;
        RECT 5.042 0.428 5.11 0.472 ;
        RECT 5.042 0.158 5.11 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68158725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.19277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.268 0.574 0.312 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.218 0.652 ;
        RECT 4.934 0.518 5.002 0.652 ;
        RECT 4.718 0.518 4.786 0.652 ;
        RECT 4.502 0.518 4.57 0.652 ;
        RECT 4.286 0.518 4.354 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.854 0.518 3.922 0.652 ;
        RECT 3.638 0.518 3.706 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 1.262 0.4705 1.33 0.5145 ;
        RECT 1.694 0.383 1.762 0.427 ;
        RECT 1.91 0.4705 1.978 0.5145 ;
        RECT 2.45 0.538 2.518 0.582 ;
        RECT 2.666 0.538 2.734 0.582 ;
        RECT 2.882 0.538 2.95 0.582 ;
        RECT 3.098 0.538 3.166 0.582 ;
        RECT 3.314 0.538 3.382 0.582 ;
        RECT 3.64 0.538 3.704 0.582 ;
        RECT 3.856 0.538 3.92 0.582 ;
        RECT 4.072 0.538 4.136 0.582 ;
        RECT 4.288 0.538 4.352 0.582 ;
        RECT 4.504 0.538 4.568 0.582 ;
        RECT 4.72 0.538 4.784 0.582 ;
        RECT 4.936 0.538 5 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.218 0.022 ;
        RECT 4.934 -0.022 5.002 0.112 ;
        RECT 4.718 -0.022 4.786 0.112 ;
        RECT 4.502 -0.022 4.57 0.112 ;
        RECT 4.286 -0.022 4.354 0.112 ;
        RECT 4.07 -0.022 4.138 0.112 ;
        RECT 3.854 -0.022 3.922 0.112 ;
        RECT 3.638 -0.022 3.706 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 1.91 0.048 1.978 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.638 0.048 3.706 0.092 ;
        RECT 3.854 0.048 3.922 0.092 ;
        RECT 4.07 0.048 4.138 0.092 ;
        RECT 4.286 0.048 4.354 0.092 ;
        RECT 4.502 0.048 4.57 0.092 ;
        RECT 4.718 0.048 4.786 0.092 ;
        RECT 4.934 0.048 5.002 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.398 0.202 ;
      RECT 0.722 0.428 0.938 0.472 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.694 0.158 2.342 0.202 ;
      RECT 2.45 0.158 3.098 0.202 ;
      RECT 2.99 0.248 3.206 0.292 ;
      RECT 5.042 0.248 5.11 0.382 ;
    LAYER v0 ;
      RECT 4.07 0.338 4.138 0.382 ;
      RECT 3.854 0.338 3.922 0.382 ;
      RECT 3.638 0.338 3.706 0.382 ;
      RECT 3.422 0.068 3.49 0.112 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.206 0.068 3.274 0.112 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.248 3.166 0.292 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.248 2.842 0.292 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.4705 2.194 0.5145 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.4705 1.87 0.5145 ;
      RECT 1.586 0.383 1.654 0.427 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 0.938 0.203 1.006 0.247 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.616 0.088 0.68 0.132 ;
      RECT 0.616 0.3855 0.68 0.4295 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.4 0.3855 0.464 0.4295 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.518 0.682 0.562 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.006 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.518 1.586 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.87 0.338 2.126 0.382 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.342 0.158 2.41 0.292 ;
      RECT 2.41 0.248 2.862 0.292 ;
      RECT 3.098 0.068 3.166 0.202 ;
      RECT 3.166 0.068 3.598 0.112 ;
      RECT 3.206 0.158 3.274 0.292 ;
      RECT 2.45 0.428 3.53 0.472 ;
      RECT 3.274 0.158 3.53 0.202 ;
      RECT 3.53 0.158 3.598 0.472 ;
      RECT 3.598 0.338 4.246 0.382 ;
  END
END b15cilb05hn1n48x5

MACRO b15cilb05hn1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n64x5 0 0 ;
  SIZE 6.048 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0396 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0468 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.248 3.922 0.292 ;
        RECT 2.342 0.338 3.274 0.382 ;
        RECT 3.206 0.248 3.274 0.382 ;
        RECT 2.342 0.248 2.41 0.382 ;
        RECT 1.586 0.248 2.41 0.292 ;
        RECT 1.586 0.068 1.654 0.292 ;
        RECT 1.37 0.068 1.654 0.112 ;
        RECT 1.046 0.248 1.438 0.292 ;
        RECT 1.37 0.068 1.438 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.722 0.068 1.114 0.112 ;
        RECT 0.722 0.068 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 2.558 0.338 2.626 0.382 ;
        RECT 3.422 0.248 3.49 0.292 ;
        RECT 3.746 0.248 3.814 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.428 5.994 0.472 ;
        RECT 4.07 0.158 5.994 0.202 ;
        RECT 5.798 0.158 5.866 0.472 ;
        RECT 5.582 0.158 5.65 0.472 ;
        RECT 5.366 0.158 5.434 0.472 ;
        RECT 5.15 0.158 5.218 0.472 ;
        RECT 4.934 0.158 5.002 0.472 ;
        RECT 4.718 0.158 4.786 0.472 ;
        RECT 4.07 0.158 4.138 0.472 ;
      LAYER v0 ;
        RECT 4.178 0.428 4.246 0.472 ;
        RECT 4.178 0.158 4.246 0.202 ;
        RECT 4.394 0.428 4.462 0.472 ;
        RECT 4.394 0.158 4.462 0.202 ;
        RECT 4.61 0.428 4.678 0.472 ;
        RECT 4.61 0.158 4.678 0.202 ;
        RECT 4.826 0.428 4.894 0.472 ;
        RECT 4.826 0.158 4.894 0.202 ;
        RECT 5.042 0.428 5.11 0.472 ;
        RECT 5.042 0.158 5.11 0.202 ;
        RECT 5.258 0.428 5.326 0.472 ;
        RECT 5.258 0.158 5.326 0.202 ;
        RECT 5.474 0.428 5.542 0.472 ;
        RECT 5.474 0.158 5.542 0.202 ;
        RECT 5.69 0.428 5.758 0.472 ;
        RECT 5.69 0.158 5.758 0.202 ;
        RECT 5.906 0.428 5.974 0.472 ;
        RECT 5.906 0.158 5.974 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 0.477111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.268 0.574 0.312 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.082 0.652 ;
        RECT 5.798 0.518 5.866 0.652 ;
        RECT 5.582 0.518 5.65 0.652 ;
        RECT 5.366 0.518 5.434 0.652 ;
        RECT 5.15 0.518 5.218 0.652 ;
        RECT 4.934 0.518 5.002 0.652 ;
        RECT 4.718 0.518 4.786 0.652 ;
        RECT 4.502 0.518 4.57 0.652 ;
        RECT 4.286 0.518 4.354 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.638 0.518 3.706 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 1.262 0.4705 1.33 0.5145 ;
        RECT 1.694 0.383 1.762 0.427 ;
        RECT 1.91 0.4705 1.978 0.5145 ;
        RECT 2.126 0.4705 2.194 0.5145 ;
        RECT 2.558 0.538 2.626 0.582 ;
        RECT 2.774 0.538 2.842 0.582 ;
        RECT 2.99 0.538 3.058 0.582 ;
        RECT 3.424 0.538 3.488 0.582 ;
        RECT 3.64 0.538 3.704 0.582 ;
        RECT 4.072 0.538 4.136 0.582 ;
        RECT 4.288 0.538 4.352 0.582 ;
        RECT 4.504 0.538 4.568 0.582 ;
        RECT 4.72 0.538 4.784 0.582 ;
        RECT 4.936 0.538 5 0.582 ;
        RECT 5.152 0.538 5.216 0.582 ;
        RECT 5.368 0.538 5.432 0.582 ;
        RECT 5.584 0.538 5.648 0.582 ;
        RECT 5.8 0.538 5.864 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.082 0.022 ;
        RECT 5.798 -0.022 5.866 0.112 ;
        RECT 5.582 -0.022 5.65 0.112 ;
        RECT 5.366 -0.022 5.434 0.112 ;
        RECT 5.15 -0.022 5.218 0.112 ;
        RECT 4.934 -0.022 5.002 0.112 ;
        RECT 4.718 -0.022 4.786 0.112 ;
        RECT 4.502 -0.022 4.57 0.112 ;
        RECT 4.286 -0.022 4.354 0.112 ;
        RECT 4.07 -0.022 4.138 0.112 ;
        RECT 3.206 -0.022 3.274 0.112 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 1.91 0.048 1.978 0.092 ;
        RECT 2.126 0.048 2.194 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
        RECT 3.208 0.048 3.272 0.092 ;
        RECT 4.072 0.048 4.136 0.092 ;
        RECT 4.288 0.048 4.352 0.092 ;
        RECT 4.504 0.048 4.568 0.092 ;
        RECT 4.72 0.048 4.784 0.092 ;
        RECT 4.936 0.048 5 0.092 ;
        RECT 5.152 0.048 5.216 0.092 ;
        RECT 5.368 0.048 5.432 0.092 ;
        RECT 5.584 0.048 5.648 0.092 ;
        RECT 5.8 0.048 5.864 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.398 0.202 ;
      RECT 0.722 0.428 0.938 0.472 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.694 0.158 2.45 0.202 ;
      RECT 2.558 0.428 3.314 0.472 ;
      RECT 2.558 0.158 3.922 0.202 ;
      RECT 4.178 0.248 4.678 0.292 ;
      RECT 5.906 0.248 5.974 0.382 ;
    LAYER v0 ;
      RECT 4.502 0.248 4.57 0.292 ;
      RECT 4.286 0.248 4.354 0.292 ;
      RECT 3.962 0.246 4.03 0.29 ;
      RECT 3.854 0.068 3.922 0.112 ;
      RECT 3.746 0.158 3.814 0.202 ;
      RECT 3.746 0.424 3.814 0.468 ;
      RECT 3.638 0.068 3.706 0.112 ;
      RECT 3.53 0.158 3.598 0.202 ;
      RECT 3.53 0.424 3.598 0.468 ;
      RECT 3.422 0.068 3.49 0.112 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.098 0.158 3.166 0.202 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.882 0.248 2.95 0.292 ;
      RECT 2.882 0.428 2.95 0.472 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.4705 2.302 0.5145 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 2.018 0.4705 2.086 0.5145 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.4705 1.87 0.5145 ;
      RECT 1.586 0.383 1.654 0.427 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 0.938 0.203 1.006 0.247 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.616 0.088 0.68 0.132 ;
      RECT 0.616 0.3855 0.68 0.4295 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.4 0.3855 0.464 0.4295 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.518 0.682 0.562 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.006 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.518 1.586 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.87 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.086 0.338 2.234 0.382 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 2.45 0.158 2.518 0.292 ;
      RECT 2.518 0.248 2.97 0.292 ;
      RECT 3.314 0.338 3.382 0.472 ;
      RECT 3.382 0.338 3.53 0.382 ;
      RECT 3.53 0.338 3.598 0.562 ;
      RECT 3.598 0.338 3.746 0.382 ;
      RECT 3.746 0.338 3.814 0.562 ;
      RECT 3.814 0.518 3.962 0.562 ;
      RECT 3.314 0.068 3.962 0.112 ;
      RECT 3.962 0.068 4.03 0.562 ;
  END
END b15cilb05hn1n64x5

MACRO b15cilb05hn1n80x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb05hn1n80x5 0 0 ;
  SIZE 7.02 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0477 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0612 LAYER m1 ;
      ANTENNAMAXAREACAR 1.17166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.248 4.894 0.292 ;
        RECT 2.882 0.338 4.354 0.382 ;
        RECT 4.286 0.248 4.354 0.382 ;
        RECT 2.882 0.248 2.95 0.382 ;
        RECT 1.91 0.248 2.95 0.292 ;
        RECT 1.91 0.068 1.978 0.292 ;
        RECT 1.694 0.068 1.978 0.112 ;
        RECT 1.37 0.248 1.762 0.292 ;
        RECT 1.694 0.068 1.762 0.292 ;
        RECT 1.37 0.068 1.438 0.292 ;
        RECT 1.046 0.068 1.438 0.112 ;
        RECT 1.046 0.068 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.262 0.068 1.33 0.112 ;
        RECT 3.098 0.338 3.166 0.382 ;
        RECT 3.746 0.338 3.814 0.382 ;
        RECT 3.962 0.338 4.03 0.382 ;
        RECT 4.61 0.248 4.678 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.26622 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.502 0.428 6.946 0.472 ;
        RECT 6.878 0.158 6.946 0.472 ;
        RECT 5.582 0.158 6.946 0.202 ;
        RECT 6.23 0.158 6.298 0.472 ;
        RECT 6.014 0.158 6.082 0.472 ;
        RECT 5.798 0.158 5.866 0.472 ;
        RECT 5.582 0.158 5.65 0.472 ;
        RECT 5.042 0.248 5.65 0.292 ;
        RECT 5.366 0.248 5.434 0.472 ;
        RECT 5.15 0.248 5.218 0.472 ;
        RECT 5.042 0.068 5.11 0.292 ;
      LAYER v0 ;
        RECT 4.61 0.428 4.678 0.472 ;
        RECT 4.826 0.428 4.894 0.472 ;
        RECT 5.042 0.428 5.11 0.472 ;
        RECT 5.042 0.138 5.11 0.182 ;
        RECT 5.258 0.428 5.326 0.472 ;
        RECT 5.258 0.248 5.326 0.292 ;
        RECT 5.474 0.428 5.542 0.472 ;
        RECT 5.474 0.248 5.542 0.292 ;
        RECT 5.69 0.428 5.758 0.472 ;
        RECT 5.69 0.158 5.758 0.202 ;
        RECT 5.906 0.428 5.974 0.472 ;
        RECT 5.906 0.158 5.974 0.202 ;
        RECT 6.122 0.428 6.19 0.472 ;
        RECT 6.122 0.158 6.19 0.202 ;
        RECT 6.338 0.428 6.406 0.472 ;
        RECT 6.338 0.158 6.406 0.202 ;
        RECT 6.554 0.428 6.622 0.472 ;
        RECT 6.554 0.158 6.622 0.202 ;
        RECT 6.77 0.428 6.838 0.472 ;
        RECT 6.77 0.158 6.838 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5301235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.378 0.292 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0252 LAYER m1 ;
      ANTENNAMAXAREACAR 0.666508 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 1.09777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.268 0.898 0.312 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 7.054 0.652 ;
        RECT 6.878 0.518 6.946 0.652 ;
        RECT 6.662 0.518 6.73 0.652 ;
        RECT 6.446 0.518 6.514 0.652 ;
        RECT 6.23 0.518 6.298 0.652 ;
        RECT 6.014 0.518 6.082 0.652 ;
        RECT 5.798 0.518 5.866 0.652 ;
        RECT 5.582 0.518 5.65 0.652 ;
        RECT 5.366 0.518 5.434 0.652 ;
        RECT 5.15 0.518 5.218 0.652 ;
        RECT 4.934 0.518 5.002 0.652 ;
        RECT 4.718 0.518 4.786 0.652 ;
        RECT 4.394 0.518 4.462 0.652 ;
        RECT 4.178 0.518 4.246 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 3.206 0.518 3.274 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 2.018 0.383 2.086 0.427 ;
        RECT 2.234 0.4705 2.302 0.5145 ;
        RECT 2.45 0.4705 2.518 0.5145 ;
        RECT 2.666 0.4705 2.734 0.5145 ;
        RECT 3.208 0.538 3.272 0.582 ;
        RECT 3.424 0.538 3.488 0.582 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 3.962 0.538 4.03 0.582 ;
        RECT 4.18 0.538 4.244 0.582 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 4.72 0.538 4.784 0.582 ;
        RECT 4.936 0.538 5 0.582 ;
        RECT 5.152 0.538 5.216 0.582 ;
        RECT 5.368 0.538 5.432 0.582 ;
        RECT 5.584 0.538 5.648 0.582 ;
        RECT 5.8 0.538 5.864 0.582 ;
        RECT 6.016 0.538 6.08 0.582 ;
        RECT 6.232 0.538 6.296 0.582 ;
        RECT 6.448 0.538 6.512 0.582 ;
        RECT 6.664 0.538 6.728 0.582 ;
        RECT 6.88 0.538 6.944 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 7.054 0.022 ;
        RECT 6.878 -0.022 6.946 0.112 ;
        RECT 6.662 -0.022 6.73 0.112 ;
        RECT 6.446 -0.022 6.514 0.112 ;
        RECT 6.23 -0.022 6.298 0.112 ;
        RECT 6.014 -0.022 6.082 0.112 ;
        RECT 5.798 -0.022 5.866 0.112 ;
        RECT 5.582 -0.022 5.65 0.112 ;
        RECT 5.366 -0.022 5.434 0.112 ;
        RECT 5.15 -0.022 5.218 0.112 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.234 0.048 2.302 0.092 ;
        RECT 2.45 0.048 2.518 0.092 ;
        RECT 2.666 0.048 2.734 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.316 0.048 3.38 0.092 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.748 0.048 3.812 0.092 ;
        RECT 3.964 0.048 4.028 0.092 ;
        RECT 5.152 0.048 5.216 0.092 ;
        RECT 5.368 0.048 5.432 0.092 ;
        RECT 5.584 0.048 5.648 0.092 ;
        RECT 5.8 0.048 5.864 0.092 ;
        RECT 6.016 0.048 6.08 0.092 ;
        RECT 6.232 0.048 6.296 0.092 ;
        RECT 6.448 0.048 6.512 0.092 ;
        RECT 6.664 0.048 6.728 0.092 ;
        RECT 6.88 0.048 6.944 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 4.808 0.338 6.856 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.506 0.202 ;
      RECT 1.046 0.428 1.262 0.472 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.018 0.158 2.99 0.202 ;
      RECT 3.206 0.428 4.394 0.472 ;
      RECT 3.098 0.158 4.894 0.202 ;
      RECT 6.338 0.338 6.838 0.382 ;
    LAYER v1 ;
      RECT 6.666 0.338 6.726 0.382 ;
      RECT 4.938 0.338 4.998 0.382 ;
    LAYER v0 ;
      RECT 6.662 0.338 6.73 0.382 ;
      RECT 6.446 0.338 6.514 0.382 ;
      RECT 4.826 0.068 4.894 0.112 ;
      RECT 4.826 0.338 4.894 0.382 ;
      RECT 4.718 0.158 4.786 0.202 ;
      RECT 4.61 0.068 4.678 0.112 ;
      RECT 4.61 0.338 4.678 0.382 ;
      RECT 4.502 0.158 4.57 0.202 ;
      RECT 4.394 0.068 4.462 0.112 ;
      RECT 4.286 0.158 4.354 0.202 ;
      RECT 4.286 0.428 4.354 0.472 ;
      RECT 4.178 0.068 4.246 0.112 ;
      RECT 4.07 0.158 4.138 0.202 ;
      RECT 4.07 0.428 4.138 0.472 ;
      RECT 3.854 0.158 3.922 0.202 ;
      RECT 3.854 0.248 3.922 0.292 ;
      RECT 3.854 0.428 3.922 0.472 ;
      RECT 3.638 0.158 3.706 0.202 ;
      RECT 3.638 0.248 3.706 0.292 ;
      RECT 3.53 0.428 3.598 0.472 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.422 0.248 3.49 0.292 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.4705 2.842 0.5145 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.558 0.338 2.626 0.382 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.4705 2.194 0.5145 ;
      RECT 1.91 0.383 1.978 0.427 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.383 1.87 0.427 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.262 0.203 1.33 0.247 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.94 0.088 1.004 0.132 ;
      RECT 0.94 0.3855 1.004 0.4295 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.3855 0.79 0.4295 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.508 0.3855 0.572 0.4295 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.398 0.472 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.518 1.006 0.562 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.79 0.158 0.938 0.202 ;
      RECT 0.938 0.068 1.006 0.472 ;
      RECT 1.262 0.158 1.33 0.472 ;
      RECT 1.33 0.338 1.694 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.762 0.518 1.91 0.562 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 2.194 0.338 2.774 0.382 ;
      RECT 2.774 0.338 2.842 0.562 ;
      RECT 2.99 0.158 3.058 0.292 ;
      RECT 3.058 0.248 3.942 0.292 ;
      RECT 4.394 0.338 4.462 0.472 ;
      RECT 4.462 0.338 4.934 0.382 ;
      RECT 4.07 0.068 4.934 0.112 ;
      RECT 4.934 0.068 5.002 0.382 ;
  END
END b15cilb05hn1n80x5

MACRO b15cilb81hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb81hn1n02x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.248 2.302 0.292 ;
        RECT 2.018 0.068 2.086 0.292 ;
      LAYER v0 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.126 0.248 2.194 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.666 0.158 2.734 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.428 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.262 0.338 1.33 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.45 0.4725 2.518 0.5165 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.37 0.093 1.438 0.137 ;
        RECT 1.694 0.093 1.762 0.137 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.158 1.888 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.398 0.068 0.614 0.112 ;
      RECT 0.378 0.428 0.722 0.472 ;
      RECT 0.594 0.248 0.938 0.292 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 2.126 0.338 2.342 0.382 ;
    LAYER v1 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 0.402 0.158 0.462 0.202 ;
    LAYER v0 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.018 0.466 2.086 0.51 ;
      RECT 1.802 0.093 1.87 0.137 ;
      RECT 1.586 0.093 1.654 0.137 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.154 0.2685 1.222 0.3125 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.046 0.2685 1.114 0.3125 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.134 0.112 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.518 1.154 0.562 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.33 0.248 1.546 0.292 ;
      RECT 1.654 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.342 0.068 2.41 0.382 ;
      RECT 2.41 0.338 2.538 0.382 ;
  END
END b15cilb81hn1n02x5

MACRO b15cilb81hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb81hn1n03x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.48622225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.248 2.302 0.292 ;
        RECT 2.018 0.068 2.086 0.292 ;
      LAYER v0 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.126 0.248 2.194 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.666 0.158 2.734 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.428 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.262 0.338 1.33 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.45 0.4725 2.518 0.5165 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.37 0.093 1.438 0.137 ;
        RECT 1.694 0.093 1.762 0.137 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.158 1.888 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.398 0.068 0.614 0.112 ;
      RECT 0.378 0.428 0.722 0.472 ;
      RECT 0.594 0.248 0.938 0.292 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 2.126 0.338 2.342 0.382 ;
    LAYER v1 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 0.402 0.158 0.462 0.202 ;
    LAYER v0 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.018 0.466 2.086 0.51 ;
      RECT 1.802 0.093 1.87 0.137 ;
      RECT 1.586 0.093 1.654 0.137 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.154 0.2685 1.222 0.3125 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.046 0.2685 1.114 0.3125 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.134 0.112 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.518 1.154 0.562 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.33 0.248 1.546 0.292 ;
      RECT 1.654 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.342 0.068 2.41 0.382 ;
      RECT 2.41 0.338 2.538 0.382 ;
  END
END b15cilb81hn1n03x5

MACRO b15cilb81hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb81hn1n04x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.48622225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.248 2.302 0.292 ;
        RECT 2.018 0.068 2.086 0.292 ;
      LAYER v0 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.126 0.248 2.194 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.666 0.158 2.734 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.428 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.262 0.338 1.33 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.45 0.4725 2.518 0.5165 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.37 0.093 1.438 0.137 ;
        RECT 1.694 0.093 1.762 0.137 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.158 1.888 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.398 0.068 0.614 0.112 ;
      RECT 0.378 0.428 0.722 0.472 ;
      RECT 0.594 0.248 0.938 0.292 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 2.126 0.338 2.342 0.382 ;
    LAYER v1 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 0.402 0.158 0.462 0.202 ;
    LAYER v0 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.018 0.466 2.086 0.51 ;
      RECT 1.802 0.093 1.87 0.137 ;
      RECT 1.586 0.093 1.654 0.137 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.154 0.2685 1.222 0.3125 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.046 0.2685 1.114 0.3125 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.134 0.112 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.518 1.154 0.562 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.33 0.248 1.546 0.292 ;
      RECT 1.654 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.342 0.068 2.41 0.382 ;
      RECT 2.41 0.338 2.558 0.382 ;
      RECT 2.558 0.158 2.626 0.382 ;
  END
END b15cilb81hn1n04x5

MACRO b15cilb81hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb81hn1n08x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.248 2.302 0.292 ;
        RECT 2.018 0.068 2.086 0.292 ;
      LAYER v0 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.126 0.248 2.194 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 2.842 0.382 ;
        RECT 2.774 0.158 2.842 0.382 ;
        RECT 2.45 0.158 2.842 0.202 ;
        RECT 2.558 0.338 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.4725 2.626 0.5165 ;
        RECT 2.558 0.158 2.626 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.428 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.262 0.338 1.33 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.45 0.4725 2.518 0.5165 ;
        RECT 2.666 0.4725 2.734 0.5165 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.37 0.093 1.438 0.137 ;
        RECT 1.694 0.093 1.762 0.137 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.158 1.888 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.398 0.068 0.614 0.112 ;
      RECT 0.378 0.428 0.722 0.472 ;
      RECT 0.594 0.248 0.938 0.292 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 2.126 0.338 2.342 0.382 ;
    LAYER v1 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 0.402 0.158 0.462 0.202 ;
    LAYER v0 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.018 0.466 2.086 0.51 ;
      RECT 1.802 0.093 1.87 0.137 ;
      RECT 1.586 0.093 1.654 0.137 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.154 0.2685 1.222 0.3125 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.046 0.2685 1.114 0.3125 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.134 0.112 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.518 1.154 0.562 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.33 0.248 1.546 0.292 ;
      RECT 1.654 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.342 0.068 2.41 0.382 ;
      RECT 2.41 0.248 2.646 0.292 ;
  END
END b15cilb81hn1n08x5

MACRO b15cilb81hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb81hn1n12x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.00918 LAYER m1 ;
    ANTENNADIFFAREA 0.03672 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.068 2.842 0.562 ;
        RECT 2.45 0.338 2.842 0.382 ;
        RECT 2.45 0.158 2.734 0.202 ;
      LAYER m2 ;
        RECT 2.416 0.158 2.984 0.202 ;
      LAYER v1 ;
        RECT 2.562 0.158 2.622 0.202 ;
        RECT 2.778 0.158 2.838 0.202 ;
      LAYER v0 ;
        RECT 2.558 0.338 2.626 0.382 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 2.774 0.45 2.842 0.494 ;
        RECT 2.774 0.138 2.842 0.182 ;
    END
  END clkout
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.82076925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.667 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.068 2.086 0.382 ;
      LAYER v0 ;
        RECT 2.018 0.133 2.086 0.177 ;
    END
  END clk
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.428 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.262 0.338 1.33 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.45 0.45 2.518 0.494 ;
        RECT 2.666 0.45 2.734 0.494 ;
        RECT 2.882 0.45 2.95 0.494 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.37 0.093 1.438 0.137 ;
        RECT 1.694 0.133 1.762 0.177 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.45 0.048 2.518 0.092 ;
        RECT 2.666 0.048 2.734 0.092 ;
        RECT 2.882 0.048 2.95 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.158 1.996 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.398 0.068 0.614 0.112 ;
      RECT 0.378 0.428 0.722 0.472 ;
      RECT 0.594 0.248 0.938 0.292 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.91 0.068 1.978 0.202 ;
      RECT 2.126 0.428 2.342 0.472 ;
      RECT 2.45 0.338 2.774 0.382 ;
      RECT 2.45 0.158 2.734 0.202 ;
    LAYER v1 ;
      RECT 1.914 0.158 1.974 0.202 ;
      RECT 0.402 0.158 0.462 0.202 ;
    LAYER v0 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.91 0.133 1.978 0.177 ;
      RECT 1.586 0.133 1.654 0.177 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.154 0.2685 1.222 0.3125 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.046 0.2685 1.114 0.3125 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.134 0.112 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.518 1.154 0.562 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.33 0.248 1.546 0.292 ;
      RECT 1.654 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.978 0.518 2.194 0.562 ;
      RECT 2.342 0.068 2.41 0.472 ;
      RECT 2.41 0.248 2.734 0.292 ;
      RECT 2.774 0.068 2.842 0.562 ;
  END
END b15cilb81hn1n12x5

MACRO b15cilb81hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb81hn1n16x5 0 0 ;
  SIZE 3.132 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 1.42617275 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 1.97470075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 2.194 0.292 ;
        RECT 2.126 0.068 2.194 0.292 ;
      LAYER v0 ;
        RECT 1.91 0.248 1.978 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.338 3.058 0.382 ;
        RECT 2.99 0.158 3.058 0.382 ;
        RECT 2.558 0.158 3.058 0.202 ;
        RECT 2.882 0.338 2.95 0.562 ;
        RECT 2.666 0.338 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 2.882 0.158 2.95 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.428 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.166 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.166 0.022 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 2.018 0.133 2.086 0.177 ;
        RECT 2.342 0.133 2.41 0.177 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.158 1.888 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.398 0.068 0.614 0.112 ;
      RECT 0.378 0.428 0.722 0.472 ;
      RECT 0.594 0.248 0.938 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 2.234 0.068 2.302 0.472 ;
    LAYER v1 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 0.402 0.158 0.462 0.202 ;
    LAYER v0 ;
      RECT 2.774 0.248 2.842 0.292 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.45 0.133 2.518 0.177 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.133 2.302 0.177 ;
      RECT 1.91 0.498 1.978 0.542 ;
      RECT 1.802 0.133 1.87 0.177 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.262 0.2705 1.33 0.3145 ;
      RECT 1.154 0.2705 1.222 0.3145 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.046 0.2705 1.114 0.3145 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.134 0.112 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.518 1.154 0.562 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.382 ;
      RECT 1.546 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 2.302 0.428 2.45 0.472 ;
      RECT 2.45 0.068 2.518 0.472 ;
      RECT 2.518 0.248 2.862 0.292 ;
  END
END b15cilb81hn1n16x5

MACRO b15cilb81hn1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb81hn1n24x5 0 0 ;
  SIZE 3.564 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 1.56222225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 2.163077 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.248 2.41 0.292 ;
        RECT 2.342 0.068 2.41 0.292 ;
      LAYER v0 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.234 0.248 2.302 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07956 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.338 3.49 0.382 ;
        RECT 3.422 0.158 3.49 0.382 ;
        RECT 2.774 0.158 3.49 0.202 ;
        RECT 3.314 0.338 3.382 0.562 ;
        RECT 3.098 0.338 3.166 0.562 ;
        RECT 2.882 0.338 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 2.882 0.158 2.95 0.202 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.098 0.158 3.166 0.202 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.314 0.158 3.382 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.428 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.598 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.802 0.428 2.518 0.472 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.774 0.364 2.842 0.408 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.422 0.448 3.49 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.598 0.022 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 3.206 -0.022 3.274 0.112 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.37 0.093 1.438 0.137 ;
        RECT 1.91 0.093 1.978 0.137 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
        RECT 3.208 0.048 3.272 0.092 ;
        RECT 3.424 0.048 3.488 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.158 1.888 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.398 0.068 0.614 0.112 ;
      RECT 0.378 0.428 0.722 0.472 ;
      RECT 0.594 0.248 0.938 0.292 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 2.018 0.338 2.45 0.382 ;
    LAYER v1 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 0.402 0.158 0.462 0.202 ;
    LAYER v0 ;
      RECT 3.098 0.248 3.166 0.292 ;
      RECT 2.882 0.248 2.95 0.292 ;
      RECT 2.666 0.138 2.734 0.182 ;
      RECT 2.558 0.338 2.626 0.382 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.802 0.093 1.87 0.137 ;
      RECT 1.586 0.113 1.654 0.157 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.154 0.2685 1.222 0.3125 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.046 0.2685 1.114 0.3125 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.134 0.112 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.518 1.154 0.562 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.33 0.248 1.546 0.292 ;
      RECT 1.546 0.338 1.586 0.382 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.654 0.338 1.694 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.762 0.518 2.106 0.562 ;
      RECT 2.45 0.068 2.518 0.382 ;
      RECT 2.518 0.338 2.666 0.382 ;
      RECT 2.666 0.068 2.734 0.382 ;
      RECT 2.734 0.248 3.274 0.292 ;
  END
END b15cilb81hn1n24x5

MACRO b15cilb81hn1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb81hn1n32x5 0 0 ;
  SIZE 3.888 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.027 LAYER m1 ;
      ANTENNAMAXAREACAR 1.98233325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0189 LAYER m1 ;
      ANTENNAMAXAREACAR 2.83190475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.292 ;
      LAYER v0 ;
        RECT 1.91 0.138 1.978 0.182 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.10404 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.338 3.814 0.382 ;
        RECT 3.746 0.158 3.814 0.382 ;
        RECT 2.882 0.158 3.814 0.202 ;
        RECT 3.638 0.338 3.706 0.562 ;
        RECT 3.206 0.338 3.274 0.562 ;
        RECT 2.99 0.338 3.058 0.562 ;
      LAYER v0 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.206 0.158 3.274 0.202 ;
        RECT 3.422 0.338 3.49 0.382 ;
        RECT 3.422 0.158 3.49 0.202 ;
        RECT 3.638 0.448 3.706 0.492 ;
        RECT 3.638 0.158 3.706 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.428 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.922 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 3.746 0.448 3.814 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.922 0.022 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.316 0.048 3.38 0.092 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.748 0.048 3.812 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.158 1.78 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.398 0.068 0.614 0.112 ;
      RECT 0.378 0.428 0.722 0.472 ;
      RECT 0.594 0.248 0.938 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.018 0.068 2.086 0.292 ;
    LAYER v1 ;
      RECT 1.698 0.158 1.758 0.202 ;
      RECT 0.402 0.158 0.462 0.202 ;
    LAYER v0 ;
      RECT 3.53 0.248 3.598 0.292 ;
      RECT 3.314 0.248 3.382 0.292 ;
      RECT 3.098 0.248 3.166 0.292 ;
      RECT 2.882 0.248 2.95 0.292 ;
      RECT 2.774 0.448 2.842 0.492 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.558 0.448 2.626 0.492 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.138 2.086 0.182 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.694 0.138 1.762 0.182 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.262 0.2705 1.33 0.3145 ;
      RECT 1.154 0.2705 1.222 0.3145 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.046 0.2705 1.114 0.3145 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.2255 0.466 0.2695 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.134 0.112 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.518 1.154 0.562 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.382 ;
      RECT 1.546 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 2.194 0.338 2.342 0.382 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.41 0.338 2.558 0.382 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 2.626 0.338 2.774 0.382 ;
      RECT 2.774 0.338 2.842 0.562 ;
      RECT 2.086 0.248 3.618 0.292 ;
  END
END b15cilb81hn1n32x5

MACRO b15cilb81hn1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cilb81hn1n64x5 0 0 ;
  SIZE 5.508 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0396 LAYER m1 ;
      ANTENNAMAXAREACAR 0.893 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0324 LAYER m1 ;
      ANTENNAMAXAREACAR 1.11625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.518 2.41 0.562 ;
        RECT 2.126 0.338 2.194 0.562 ;
        RECT 1.91 0.338 2.194 0.382 ;
      LAYER v0 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.234 0.518 2.302 0.562 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.20196 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.338 5.434 0.382 ;
        RECT 5.366 0.158 5.434 0.382 ;
        RECT 3.638 0.158 5.434 0.202 ;
        RECT 5.258 0.338 5.326 0.562 ;
        RECT 4.826 0.338 4.894 0.562 ;
        RECT 4.394 0.338 4.462 0.562 ;
        RECT 3.962 0.338 4.03 0.562 ;
        RECT 3.746 0.338 3.814 0.562 ;
      LAYER v0 ;
        RECT 3.746 0.448 3.814 0.492 ;
        RECT 3.746 0.158 3.814 0.202 ;
        RECT 3.962 0.448 4.03 0.492 ;
        RECT 3.962 0.158 4.03 0.202 ;
        RECT 4.178 0.338 4.246 0.382 ;
        RECT 4.178 0.158 4.246 0.202 ;
        RECT 4.394 0.448 4.462 0.492 ;
        RECT 4.394 0.158 4.462 0.202 ;
        RECT 4.61 0.338 4.678 0.382 ;
        RECT 4.61 0.158 4.678 0.202 ;
        RECT 4.826 0.448 4.894 0.492 ;
        RECT 4.826 0.158 4.894 0.202 ;
        RECT 5.042 0.338 5.11 0.382 ;
        RECT 5.042 0.158 5.11 0.202 ;
        RECT 5.258 0.448 5.326 0.492 ;
        RECT 5.258 0.158 5.326 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END en
  PIN te
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.2255 0.358 0.2695 ;
    END
  END te
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.542 0.652 ;
        RECT 5.366 0.428 5.434 0.652 ;
        RECT 5.15 0.428 5.218 0.652 ;
        RECT 4.934 0.428 5.002 0.652 ;
        RECT 4.718 0.428 4.786 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 4.286 0.428 4.354 0.652 ;
        RECT 4.07 0.428 4.138 0.652 ;
        RECT 3.854 0.428 3.922 0.652 ;
        RECT 3.638 0.338 3.706 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.638 0.448 3.706 0.492 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 4.07 0.448 4.138 0.492 ;
        RECT 4.286 0.448 4.354 0.492 ;
        RECT 4.502 0.448 4.57 0.492 ;
        RECT 4.718 0.448 4.786 0.492 ;
        RECT 4.934 0.448 5.002 0.492 ;
        RECT 5.15 0.448 5.218 0.492 ;
        RECT 5.366 0.448 5.434 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.542 0.022 ;
        RECT 5.366 -0.022 5.434 0.112 ;
        RECT 5.15 -0.022 5.218 0.112 ;
        RECT 4.934 -0.022 5.002 0.112 ;
        RECT 4.718 -0.022 4.786 0.112 ;
        RECT 4.502 -0.022 4.57 0.112 ;
        RECT 4.286 -0.022 4.354 0.112 ;
        RECT 4.07 -0.022 4.138 0.112 ;
        RECT 3.854 -0.022 3.922 0.112 ;
        RECT 3.638 -0.022 3.706 0.112 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.133 0.142 0.177 ;
        RECT 0.398 0.116 0.466 0.16 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.91 0.048 1.978 0.092 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 3.424 0.048 3.488 0.092 ;
        RECT 3.64 0.048 3.704 0.092 ;
        RECT 3.856 0.048 3.92 0.092 ;
        RECT 4.072 0.048 4.136 0.092 ;
        RECT 4.288 0.048 4.352 0.092 ;
        RECT 4.504 0.048 4.568 0.092 ;
        RECT 4.72 0.048 4.784 0.092 ;
        RECT 4.936 0.048 5 0.092 ;
        RECT 5.152 0.048 5.216 0.092 ;
        RECT 5.368 0.048 5.432 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.158 2.104 0.202 ;
      RECT 2.432 0.158 3.616 0.202 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.292 ;
      RECT 0.506 0.068 0.722 0.112 ;
      RECT 0.486 0.428 0.83 0.472 ;
      RECT 0.702 0.248 1.046 0.292 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 2.018 0.068 2.086 0.202 ;
      RECT 2.45 0.068 2.518 0.202 ;
      RECT 2.666 0.068 2.734 0.202 ;
      RECT 2.234 0.428 2.95 0.472 ;
      RECT 2.882 0.068 2.95 0.202 ;
      RECT 3.314 0.068 3.382 0.202 ;
      RECT 2.43 0.338 3.098 0.382 ;
      RECT 3.53 0.068 3.598 0.292 ;
    LAYER v1 ;
      RECT 3.534 0.158 3.594 0.202 ;
      RECT 3.318 0.158 3.378 0.202 ;
      RECT 2.886 0.158 2.946 0.202 ;
      RECT 2.67 0.158 2.73 0.202 ;
      RECT 2.454 0.158 2.514 0.202 ;
      RECT 2.022 0.158 2.082 0.202 ;
      RECT 0.51 0.158 0.57 0.202 ;
    LAYER v0 ;
      RECT 5.042 0.248 5.11 0.292 ;
      RECT 4.826 0.248 4.894 0.292 ;
      RECT 4.61 0.248 4.678 0.292 ;
      RECT 4.394 0.248 4.462 0.292 ;
      RECT 4.178 0.248 4.246 0.292 ;
      RECT 3.962 0.248 4.03 0.292 ;
      RECT 3.746 0.248 3.814 0.292 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.532 0.138 3.596 0.182 ;
      RECT 3.314 0.138 3.382 0.182 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 3.098 0.448 3.166 0.492 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.138 2.734 0.182 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.018 0.138 2.086 0.182 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.262 0.268 1.33 0.312 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.268 1.222 0.312 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.506 0.2255 0.574 0.2695 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.473 0.358 0.517 ;
      RECT 0.182 0.133 0.25 0.177 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.29 0.382 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.358 0.338 0.938 0.382 ;
      RECT 0.938 0.338 1.006 0.472 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.79 0.158 0.938 0.202 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.006 0.068 1.242 0.112 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.898 0.518 1.262 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 1.114 0.158 1.37 0.202 ;
      RECT 1.37 0.158 1.438 0.292 ;
      RECT 1.438 0.248 1.654 0.292 ;
      RECT 1.546 0.338 1.694 0.382 ;
      RECT 1.478 0.158 1.694 0.202 ;
      RECT 1.694 0.158 1.762 0.562 ;
      RECT 1.762 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.292 ;
      RECT 1.978 0.248 3.402 0.292 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 3.166 0.338 3.53 0.382 ;
      RECT 3.53 0.338 3.598 0.562 ;
      RECT 3.598 0.248 5.238 0.292 ;
  END
END b15cilb81hn1n64x5

MACRO b15fdw003hn1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fdw003hn1n05x5 0 0 ;
  SIZE 4.536 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.5669135 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.17518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.158 1.438 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.293 1.438 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.158 3.49 0.472 ;
      LAYER v0 ;
        RECT 3.422 0.2705 3.49 0.3145 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 6.09583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 5.225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
    END
  END rb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.248 4.354 0.382 ;
      LAYER v0 ;
        RECT 4.286 0.293 4.354 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2731625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.13777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.518 3.618 0.562 ;
        RECT 3.314 0.158 3.382 0.562 ;
      LAYER v0 ;
        RECT 3.314 0.2705 3.382 0.3145 ;
        RECT 3.53 0.518 3.598 0.562 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.57 0.652 ;
        RECT 3.746 0.338 3.814 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.45 0.473 2.518 0.517 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.746 0.3855 3.814 0.4295 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.57 0.022 ;
        RECT 4.286 -0.022 4.354 0.202 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.746 0.113 3.814 0.157 ;
        RECT 4.286 0.1185 4.354 0.1625 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.028 0.248 1.688 0.292 ;
      RECT 1.768 0.248 2.86 0.292 ;
      RECT 3.188 0.248 4.048 0.292 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 1.586 0.248 1.694 0.292 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.802 0.248 1.87 0.382 ;
      RECT 2.234 0.248 2.666 0.292 ;
      RECT 2.558 0.158 2.774 0.202 ;
      RECT 2.99 0.158 3.058 0.382 ;
      RECT 2.882 0.068 2.95 0.562 ;
      RECT 3.206 0.248 3.274 0.562 ;
      RECT 3.638 0.248 3.854 0.292 ;
      RECT 3.962 0.248 4.03 0.472 ;
      RECT 3.854 0.338 3.922 0.562 ;
      RECT 4.394 0.068 4.462 0.472 ;
    LAYER v1 ;
      RECT 3.966 0.248 4.026 0.292 ;
      RECT 3.21 0.248 3.27 0.292 ;
      RECT 2.778 0.248 2.838 0.292 ;
      RECT 1.806 0.248 1.866 0.292 ;
      RECT 1.59 0.248 1.65 0.292 ;
      RECT 1.266 0.248 1.326 0.292 ;
      RECT 1.05 0.248 1.11 0.292 ;
    LAYER v0 ;
      RECT 4.394 0.1185 4.462 0.1625 ;
      RECT 4.394 0.408 4.462 0.452 ;
      RECT 4.286 0.518 4.354 0.562 ;
      RECT 4.178 0.428 4.246 0.472 ;
      RECT 4.07 0.172 4.138 0.216 ;
      RECT 3.962 0.3855 4.03 0.4295 ;
      RECT 3.854 0.3855 3.922 0.4295 ;
      RECT 3.746 0.248 3.814 0.292 ;
      RECT 3.53 0.363 3.598 0.407 ;
      RECT 3.532 0.138 3.596 0.182 ;
      RECT 3.206 0.498 3.274 0.542 ;
      RECT 2.99 0.293 3.058 0.337 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.882 0.448 2.95 0.492 ;
      RECT 2.774 0.448 2.842 0.492 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.342 0.248 2.41 0.292 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.2705 0.574 0.3145 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.79 0.158 0.938 0.202 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.006 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.472 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 0.898 0.518 1.262 0.562 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.694 0.158 1.762 0.562 ;
      RECT 1.762 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 1.978 0.338 2.626 0.382 ;
      RECT 2.666 0.248 2.734 0.472 ;
      RECT 2.774 0.158 2.842 0.562 ;
      RECT 3.058 0.158 3.206 0.202 ;
      RECT 3.206 0.068 3.274 0.202 ;
      RECT 3.274 0.068 3.53 0.112 ;
      RECT 3.53 0.068 3.598 0.472 ;
      RECT 3.854 0.068 3.922 0.292 ;
      RECT 3.922 0.068 4.07 0.112 ;
      RECT 4.07 0.068 4.138 0.472 ;
      RECT 4.138 0.428 4.354 0.472 ;
      RECT 3.922 0.518 4.462 0.562 ;
  END
END b15fdw003hn1n05x5

MACRO b15fdw003hn1n10x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fdw003hn1n10x5 0 0 ;
  SIZE 4.86 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0117 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 3.29925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0117 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 3.29925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.158 3.814 0.382 ;
        RECT 3.314 0.158 3.382 0.382 ;
      LAYER m2 ;
        RECT 3.296 0.158 3.832 0.202 ;
      LAYER v1 ;
        RECT 3.318 0.158 3.378 0.202 ;
        RECT 3.75 0.158 3.81 0.202 ;
      LAYER v0 ;
        RECT 3.314 0.248 3.382 0.292 ;
        RECT 3.746 0.248 3.814 0.292 ;
    END
  END d
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.211 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.006875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.37 0.178 1.438 0.222 ;
    END
  END clk
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 3.04 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.518 1.546 0.562 ;
        RECT 0.938 0.248 1.006 0.562 ;
        RECT 0.614 0.338 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.37 0.518 1.438 0.562 ;
    END
  END rb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.248 4.678 0.382 ;
      LAYER v0 ;
        RECT 4.61 0.293 4.678 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2731625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 4.13777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.518 3.942 0.562 ;
        RECT 3.638 0.248 3.706 0.562 ;
        RECT 3.422 0.248 3.706 0.292 ;
      LAYER v0 ;
        RECT 3.53 0.248 3.598 0.292 ;
        RECT 3.854 0.518 3.922 0.562 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.894 0.652 ;
        RECT 4.07 0.338 4.138 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.558 0.473 2.626 0.517 ;
        RECT 3.098 0.473 3.166 0.517 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 4.07 0.3855 4.138 0.4295 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.894 0.022 ;
        RECT 4.61 -0.022 4.678 0.202 ;
        RECT 4.07 -0.022 4.138 0.202 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 1.694 0.1215 1.762 0.1655 ;
        RECT 2.126 0.1915 2.194 0.2355 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 3.098 0.138 3.166 0.182 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 4.07 0.113 4.138 0.157 ;
        RECT 4.61 0.1185 4.678 0.1625 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.158 1.364 0.202 ;
      RECT 1.444 0.158 2.32 0.202 ;
      RECT 1.028 0.428 2.336 0.472 ;
      RECT 2.416 0.428 2.86 0.472 ;
      RECT 3.188 0.428 4.372 0.472 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 2.234 0.428 2.342 0.472 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 2.234 0.068 2.302 0.202 ;
      RECT 2.45 0.428 2.518 0.562 ;
      RECT 1.802 0.068 2.018 0.112 ;
      RECT 2.774 0.248 2.842 0.472 ;
      RECT 3.206 0.068 3.274 0.382 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.206 0.428 3.274 0.562 ;
      RECT 3.314 0.158 3.382 0.382 ;
      RECT 3.746 0.158 3.814 0.382 ;
      RECT 3.962 0.248 4.394 0.292 ;
      RECT 4.286 0.338 4.354 0.472 ;
      RECT 4.178 0.338 4.246 0.562 ;
      RECT 4.718 0.068 4.786 0.472 ;
    LAYER v1 ;
      RECT 4.29 0.428 4.35 0.472 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.454 0.428 2.514 0.472 ;
      RECT 2.238 0.158 2.298 0.202 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.482 0.158 1.542 0.202 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 1.158 0.158 1.218 0.202 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.402 0.158 0.462 0.202 ;
    LAYER v0 ;
      RECT 4.718 0.1185 4.786 0.1625 ;
      RECT 4.718 0.408 4.786 0.452 ;
      RECT 4.61 0.518 4.678 0.562 ;
      RECT 4.502 0.428 4.57 0.472 ;
      RECT 4.396 0.172 4.46 0.216 ;
      RECT 4.286 0.3855 4.354 0.4295 ;
      RECT 4.178 0.3855 4.246 0.4295 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 3.854 0.363 3.922 0.407 ;
      RECT 3.856 0.138 3.92 0.182 ;
      RECT 3.314 0.068 3.382 0.112 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 3.206 0.473 3.274 0.517 ;
      RECT 2.99 0.138 3.058 0.182 ;
      RECT 2.99 0.473 3.058 0.517 ;
      RECT 2.882 0.473 2.95 0.517 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.338 2.842 0.382 ;
      RECT 2.558 0.338 2.626 0.382 ;
      RECT 2.45 0.473 2.518 0.517 ;
      RECT 2.234 0.088 2.302 0.132 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.91 0.268 1.978 0.312 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.398 0.338 0.466 0.382 ;
    LAYER m1 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 0.898 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.292 ;
      RECT 1.87 0.338 1.91 0.382 ;
      RECT 1.91 0.158 1.978 0.382 ;
      RECT 2.342 0.338 2.41 0.472 ;
      RECT 2.41 0.338 2.734 0.382 ;
      RECT 2.018 0.068 2.086 0.382 ;
      RECT 2.086 0.338 2.234 0.382 ;
      RECT 2.234 0.248 2.302 0.382 ;
      RECT 2.302 0.248 2.666 0.292 ;
      RECT 2.666 0.158 2.734 0.292 ;
      RECT 2.734 0.158 2.882 0.202 ;
      RECT 2.882 0.158 2.95 0.562 ;
      RECT 3.274 0.068 3.422 0.112 ;
      RECT 3.422 0.068 3.49 0.202 ;
      RECT 3.49 0.158 3.638 0.202 ;
      RECT 3.638 0.068 3.706 0.202 ;
      RECT 3.706 0.068 3.854 0.112 ;
      RECT 3.854 0.068 3.922 0.472 ;
      RECT 4.394 0.068 4.462 0.472 ;
      RECT 4.462 0.428 4.678 0.472 ;
      RECT 4.246 0.518 4.786 0.562 ;
  END
END b15fdw003hn1n10x5

MACRO b15fdw003hn1n20x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fdw003hn1n20x5 0 0 ;
  SIZE 5.724 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    ANTENNADIFFAREA 0.0612 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER m2 ;
        RECT 0.164 0.428 0.7 0.472 ;
      LAYER v1 ;
        RECT 0.294 0.428 0.354 0.472 ;
        RECT 0.51 0.428 0.57 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.29 0.178 0.358 0.222 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.506 0.178 0.574 0.222 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 3.861111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 3.861111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.474 0.248 5.542 0.382 ;
      LAYER m2 ;
        RECT 5.132 0.248 5.56 0.292 ;
      LAYER v1 ;
        RECT 5.478 0.248 5.538 0.292 ;
      LAYER v0 ;
        RECT 5.474 0.293 5.542 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 2.222963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.5214815 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0252 LAYER m2 ;
      ANTENNAMAXAREACAR 6.668889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.826 0.428 4.894 0.562 ;
        RECT 4.394 0.248 4.462 0.472 ;
        RECT 3.962 0.248 4.462 0.292 ;
      LAYER m2 ;
        RECT 4.376 0.428 4.912 0.472 ;
      LAYER v1 ;
        RECT 4.398 0.428 4.458 0.472 ;
        RECT 4.83 0.428 4.89 0.472 ;
      LAYER v0 ;
        RECT 4.07 0.248 4.138 0.292 ;
        RECT 4.826 0.498 4.894 0.542 ;
    END
  END ssb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 3.33363625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0252 LAYER m1 ;
      ANTENNAMAXAREACAR 1.30964275 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.292 ;
      LAYER v0 ;
        RECT 1.046 0.178 1.114 0.222 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.068 4.678 0.382 ;
      LAYER v0 ;
        RECT 4.61 0.293 4.678 0.337 ;
    END
  END d
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 2.6125 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 2.0096155 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.363 1.978 0.407 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.758 0.652 ;
        RECT 4.934 0.338 5.002 0.652 ;
        RECT 3.854 0.428 4.354 0.472 ;
        RECT 3.854 0.428 3.922 0.652 ;
        RECT 3.638 0.428 3.706 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 3.098 0.473 3.166 0.517 ;
        RECT 3.638 0.448 3.706 0.492 ;
        RECT 3.962 0.428 4.03 0.472 ;
        RECT 4.178 0.428 4.246 0.472 ;
        RECT 4.934 0.3855 5.002 0.4295 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.758 0.022 ;
        RECT 5.474 -0.022 5.542 0.202 ;
        RECT 4.934 -0.022 5.002 0.202 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 3.638 -0.022 3.706 0.112 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.126 0.158 2.41 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 0.938 -0.022 1.006 0.292 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.178 0.25 0.222 ;
        RECT 0.398 0.178 0.466 0.222 ;
        RECT 0.614 0.178 0.682 0.222 ;
        RECT 0.938 0.178 1.006 0.222 ;
        RECT 1.802 0.203 1.87 0.247 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.666 0.136 2.734 0.18 ;
        RECT 3.098 0.138 3.166 0.182 ;
        RECT 3.64 0.048 3.704 0.092 ;
        RECT 3.964 0.048 4.028 0.092 ;
        RECT 4.18 0.048 4.244 0.092 ;
        RECT 4.934 0.113 5.002 0.157 ;
        RECT 5.474 0.1185 5.542 0.1625 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.248 1.78 0.292 ;
      RECT 0.812 0.338 2.984 0.382 ;
      RECT 1.028 0.428 3.416 0.472 ;
      RECT 3.064 0.338 3.416 0.382 ;
      RECT 2.54 0.248 3.524 0.292 ;
      RECT 3.496 0.428 3.832 0.472 ;
      RECT 3.604 0.248 4.804 0.292 ;
      RECT 4.052 0.338 5.236 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.83 0.068 0.898 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.586 0.158 1.654 0.562 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.694 0.068 1.762 0.292 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 2.45 0.158 2.518 0.382 ;
      RECT 2.342 0.338 2.41 0.472 ;
      RECT 2.234 0.068 2.558 0.112 ;
      RECT 2.99 0.338 3.058 0.562 ;
      RECT 2.774 0.068 2.842 0.562 ;
      RECT 2.882 0.248 2.95 0.382 ;
      RECT 3.206 0.158 3.422 0.202 ;
      RECT 3.206 0.248 3.274 0.472 ;
      RECT 3.314 0.248 3.382 0.382 ;
      RECT 3.962 0.248 4.394 0.292 ;
      RECT 3.53 0.068 3.598 0.562 ;
      RECT 3.638 0.158 3.706 0.382 ;
      RECT 3.746 0.068 3.814 0.562 ;
      RECT 3.962 0.338 4.246 0.382 ;
      RECT 4.826 0.248 5.042 0.292 ;
      RECT 3.962 0.158 4.462 0.202 ;
      RECT 4.502 0.068 4.57 0.472 ;
      RECT 3.962 0.518 4.786 0.562 ;
      RECT 4.718 0.068 4.786 0.472 ;
      RECT 4.826 0.428 4.894 0.562 ;
      RECT 5.15 0.338 5.218 0.472 ;
      RECT 5.042 0.338 5.11 0.562 ;
      RECT 5.474 0.248 5.542 0.382 ;
      RECT 5.582 0.068 5.65 0.472 ;
    LAYER v1 ;
      RECT 5.154 0.338 5.214 0.382 ;
      RECT 4.722 0.248 4.782 0.292 ;
      RECT 4.506 0.248 4.566 0.292 ;
      RECT 4.074 0.338 4.134 0.382 ;
      RECT 3.75 0.428 3.81 0.472 ;
      RECT 3.642 0.248 3.702 0.292 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 3.426 0.248 3.486 0.292 ;
      RECT 3.318 0.338 3.378 0.382 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 3.102 0.338 3.162 0.382 ;
      RECT 2.886 0.338 2.946 0.382 ;
      RECT 2.562 0.248 2.622 0.292 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.698 0.248 1.758 0.292 ;
      RECT 1.482 0.338 1.542 0.382 ;
      RECT 1.158 0.428 1.218 0.472 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.078 0.248 0.138 0.292 ;
    LAYER v0 ;
      RECT 5.582 0.1185 5.65 0.1625 ;
      RECT 5.582 0.408 5.65 0.452 ;
      RECT 5.474 0.518 5.542 0.562 ;
      RECT 5.366 0.428 5.434 0.472 ;
      RECT 5.258 0.172 5.326 0.216 ;
      RECT 5.15 0.3855 5.218 0.4295 ;
      RECT 5.042 0.3855 5.11 0.4295 ;
      RECT 4.934 0.248 5.002 0.292 ;
      RECT 4.718 0.138 4.786 0.182 ;
      RECT 4.718 0.403 4.786 0.447 ;
      RECT 4.61 0.518 4.678 0.562 ;
      RECT 4.502 0.402 4.57 0.446 ;
      RECT 4.504 0.138 4.568 0.182 ;
      RECT 4.286 0.158 4.354 0.202 ;
      RECT 4.286 0.518 4.354 0.562 ;
      RECT 4.07 0.158 4.138 0.202 ;
      RECT 4.07 0.338 4.138 0.382 ;
      RECT 4.07 0.518 4.138 0.562 ;
      RECT 3.746 0.138 3.814 0.182 ;
      RECT 3.746 0.448 3.814 0.492 ;
      RECT 3.638 0.2705 3.706 0.3145 ;
      RECT 3.53 0.138 3.598 0.182 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.422 0.448 3.49 0.492 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.314 0.293 3.382 0.337 ;
      RECT 3.206 0.293 3.274 0.337 ;
      RECT 2.99 0.473 3.058 0.517 ;
      RECT 2.882 0.3155 2.95 0.3595 ;
      RECT 2.774 0.136 2.842 0.18 ;
      RECT 2.774 0.448 2.842 0.492 ;
      RECT 2.558 0.448 2.626 0.492 ;
      RECT 2.45 0.184 2.518 0.228 ;
      RECT 2.342 0.068 2.41 0.112 ;
      RECT 2.342 0.363 2.41 0.407 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.694 0.088 1.762 0.132 ;
      RECT 1.586 0.203 1.654 0.247 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.178 1.438 0.222 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.074 0.178 0.142 0.222 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 1.046 0.428 1.262 0.472 ;
      RECT 1.262 0.158 1.33 0.472 ;
      RECT 1.006 0.338 1.154 0.382 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.222 0.068 1.37 0.112 ;
      RECT 1.006 0.518 1.438 0.562 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 2.086 0.248 2.126 0.292 ;
      RECT 2.126 0.248 2.194 0.562 ;
      RECT 2.518 0.338 2.558 0.382 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 2.558 0.068 2.626 0.292 ;
      RECT 3.058 0.338 3.166 0.382 ;
      RECT 3.422 0.158 3.49 0.562 ;
      RECT 4.394 0.248 4.462 0.472 ;
      RECT 5.042 0.068 5.11 0.292 ;
      RECT 5.11 0.068 5.258 0.112 ;
      RECT 5.258 0.068 5.326 0.472 ;
      RECT 5.326 0.428 5.542 0.472 ;
      RECT 5.11 0.518 5.65 0.562 ;
  END
END b15fdw003hn1n20x5

MACRO b15fdw003hn1n30x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fdw003hn1n30x5 0 0 ;
  SIZE 6.804 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    ANTENNADIFFAREA 0.08874 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.562 ;
        RECT 0.506 0.068 0.574 0.562 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER m2 ;
        RECT 0.164 0.428 0.808 0.472 ;
      LAYER v1 ;
        RECT 0.294 0.428 0.354 0.472 ;
        RECT 0.51 0.428 0.57 0.472 ;
        RECT 0.726 0.428 0.786 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.29 0.178 0.358 0.222 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.506 0.178 0.574 0.222 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.722 0.178 0.79 0.222 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 3.861111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 3.861111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 6.554 0.248 6.622 0.382 ;
      LAYER m2 ;
        RECT 6.212 0.248 6.64 0.292 ;
      LAYER v1 ;
        RECT 6.558 0.248 6.618 0.292 ;
      LAYER v0 ;
        RECT 6.554 0.293 6.622 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 2.222963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.5214815 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0342 LAYER m2 ;
      ANTENNAMAXAREACAR 6.668889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.906 0.428 5.974 0.562 ;
        RECT 5.258 0.248 5.326 0.472 ;
        RECT 4.61 0.248 5.326 0.292 ;
      LAYER m2 ;
        RECT 5.24 0.428 5.992 0.472 ;
      LAYER v1 ;
        RECT 5.262 0.428 5.322 0.472 ;
        RECT 5.91 0.428 5.97 0.472 ;
      LAYER v0 ;
        RECT 4.718 0.248 4.786 0.292 ;
        RECT 4.934 0.248 5.002 0.292 ;
        RECT 5.906 0.498 5.974 0.542 ;
    END
  END ssb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 3.1715385 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.03075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.292 ;
      LAYER v0 ;
        RECT 1.262 0.178 1.33 0.222 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.746489 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.69 0.068 5.758 0.382 ;
      LAYER v0 ;
        RECT 5.69 0.293 5.758 0.337 ;
    END
  END d
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0279 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9796775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0342 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.068 2.302 0.472 ;
      LAYER v0 ;
        RECT 2.234 0.363 2.302 0.407 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.838 0.652 ;
        RECT 6.014 0.338 6.082 0.652 ;
        RECT 5.042 0.518 5.11 0.652 ;
        RECT 4.826 0.518 4.894 0.652 ;
        RECT 4.61 0.518 4.678 0.652 ;
        RECT 4.394 0.428 4.462 0.652 ;
        RECT 3.638 0.428 3.706 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.638 0.473 3.706 0.517 ;
        RECT 4.394 0.448 4.462 0.492 ;
        RECT 4.612 0.538 4.676 0.582 ;
        RECT 4.826 0.538 4.894 0.582 ;
        RECT 5.044 0.538 5.108 0.582 ;
        RECT 6.014 0.3855 6.082 0.4295 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.838 0.022 ;
        RECT 6.554 -0.022 6.622 0.202 ;
        RECT 6.014 -0.022 6.082 0.202 ;
        RECT 5.042 -0.022 5.11 0.112 ;
        RECT 4.826 -0.022 4.894 0.112 ;
        RECT 4.61 -0.022 4.678 0.112 ;
        RECT 4.394 -0.022 4.462 0.112 ;
        RECT 3.638 -0.022 3.706 0.202 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.666 0.158 2.95 0.202 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.342 -0.022 2.41 0.292 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.178 0.25 0.222 ;
        RECT 0.398 0.178 0.466 0.222 ;
        RECT 0.614 0.178 0.682 0.222 ;
        RECT 0.83 0.178 0.898 0.222 ;
        RECT 1.154 0.178 1.222 0.222 ;
        RECT 2.126 0.203 2.194 0.247 ;
        RECT 2.342 0.203 2.41 0.247 ;
        RECT 2.774 0.158 2.842 0.202 ;
        RECT 3.206 0.136 3.274 0.18 ;
        RECT 3.638 0.138 3.706 0.182 ;
        RECT 4.396 0.048 4.46 0.092 ;
        RECT 4.612 0.048 4.676 0.092 ;
        RECT 4.828 0.048 4.892 0.092 ;
        RECT 5.044 0.048 5.108 0.092 ;
        RECT 6.014 0.113 6.082 0.157 ;
        RECT 6.554 0.1185 6.622 0.1625 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.248 2.104 0.292 ;
      RECT 1.136 0.338 3.524 0.382 ;
      RECT 1.244 0.428 3.956 0.472 ;
      RECT 3.604 0.338 4.172 0.382 ;
      RECT 3.08 0.248 4.28 0.292 ;
      RECT 4.036 0.428 4.588 0.472 ;
      RECT 4.36 0.248 5.884 0.292 ;
      RECT 4.916 0.338 6.316 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 1.154 0.428 1.37 0.472 ;
      RECT 0.938 0.248 1.006 0.562 ;
      RECT 1.802 0.068 2.018 0.112 ;
      RECT 1.802 0.248 1.87 0.382 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 2.558 0.068 2.626 0.292 ;
      RECT 2.45 0.428 2.518 0.562 ;
      RECT 2.99 0.158 3.058 0.382 ;
      RECT 2.882 0.338 2.95 0.472 ;
      RECT 2.774 0.068 3.098 0.112 ;
      RECT 3.53 0.338 3.598 0.562 ;
      RECT 3.314 0.068 3.382 0.562 ;
      RECT 3.422 0.248 3.49 0.382 ;
      RECT 3.746 0.158 3.962 0.202 ;
      RECT 3.746 0.248 3.814 0.472 ;
      RECT 3.854 0.248 3.922 0.382 ;
      RECT 4.07 0.428 4.138 0.562 ;
      RECT 4.07 0.248 4.138 0.382 ;
      RECT 4.61 0.248 5.258 0.292 ;
      RECT 4.286 0.068 4.354 0.562 ;
      RECT 4.394 0.158 4.462 0.382 ;
      RECT 4.502 0.068 4.57 0.562 ;
      RECT 4.61 0.338 5.11 0.382 ;
      RECT 4.61 0.158 5.258 0.202 ;
      RECT 5.366 0.158 5.434 0.472 ;
      RECT 5.582 0.158 5.65 0.472 ;
      RECT 4.61 0.428 5.15 0.472 ;
      RECT 5.906 0.248 6.122 0.292 ;
      RECT 5.798 0.158 5.866 0.472 ;
      RECT 5.906 0.428 5.974 0.562 ;
      RECT 6.23 0.338 6.298 0.472 ;
      RECT 6.122 0.338 6.19 0.562 ;
      RECT 6.554 0.248 6.622 0.382 ;
      RECT 6.662 0.068 6.73 0.472 ;
    LAYER v1 ;
      RECT 6.234 0.338 6.294 0.382 ;
      RECT 5.802 0.248 5.862 0.292 ;
      RECT 5.586 0.248 5.646 0.292 ;
      RECT 5.37 0.248 5.43 0.292 ;
      RECT 4.938 0.338 4.998 0.382 ;
      RECT 4.506 0.428 4.566 0.472 ;
      RECT 4.398 0.248 4.458 0.292 ;
      RECT 4.29 0.428 4.35 0.472 ;
      RECT 4.182 0.248 4.242 0.292 ;
      RECT 4.074 0.338 4.134 0.382 ;
      RECT 4.074 0.428 4.134 0.472 ;
      RECT 3.966 0.248 4.026 0.292 ;
      RECT 3.858 0.338 3.918 0.382 ;
      RECT 3.75 0.428 3.81 0.472 ;
      RECT 3.642 0.338 3.702 0.382 ;
      RECT 3.426 0.338 3.486 0.382 ;
      RECT 3.102 0.248 3.162 0.292 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 2.67 0.428 2.73 0.472 ;
      RECT 2.454 0.428 2.514 0.472 ;
      RECT 2.022 0.248 2.082 0.292 ;
      RECT 1.806 0.338 1.866 0.382 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.078 0.248 0.138 0.292 ;
    LAYER v0 ;
      RECT 6.662 0.1185 6.73 0.1625 ;
      RECT 6.662 0.408 6.73 0.452 ;
      RECT 6.554 0.518 6.622 0.562 ;
      RECT 6.446 0.428 6.514 0.472 ;
      RECT 6.338 0.172 6.406 0.216 ;
      RECT 6.23 0.3855 6.298 0.4295 ;
      RECT 6.122 0.3855 6.19 0.4295 ;
      RECT 6.014 0.248 6.082 0.292 ;
      RECT 5.798 0.403 5.866 0.447 ;
      RECT 5.8 0.184 5.864 0.228 ;
      RECT 5.69 0.518 5.758 0.562 ;
      RECT 5.582 0.184 5.65 0.228 ;
      RECT 5.582 0.402 5.65 0.446 ;
      RECT 5.474 0.068 5.542 0.112 ;
      RECT 5.474 0.518 5.542 0.562 ;
      RECT 5.366 0.402 5.434 0.446 ;
      RECT 5.368 0.184 5.432 0.228 ;
      RECT 5.258 0.518 5.326 0.562 ;
      RECT 5.15 0.158 5.218 0.202 ;
      RECT 4.934 0.158 5.002 0.202 ;
      RECT 4.934 0.338 5.002 0.382 ;
      RECT 4.934 0.428 5.002 0.472 ;
      RECT 4.718 0.158 4.786 0.202 ;
      RECT 4.718 0.338 4.786 0.382 ;
      RECT 4.718 0.428 4.786 0.472 ;
      RECT 4.502 0.138 4.57 0.182 ;
      RECT 4.502 0.448 4.57 0.492 ;
      RECT 4.394 0.248 4.462 0.292 ;
      RECT 4.286 0.138 4.354 0.182 ;
      RECT 4.286 0.448 4.354 0.492 ;
      RECT 4.178 0.448 4.246 0.492 ;
      RECT 4.07 0.158 4.138 0.202 ;
      RECT 4.07 0.293 4.138 0.337 ;
      RECT 4.07 0.448 4.138 0.492 ;
      RECT 3.962 0.448 4.03 0.492 ;
      RECT 3.854 0.158 3.922 0.202 ;
      RECT 3.854 0.293 3.922 0.337 ;
      RECT 3.746 0.293 3.814 0.337 ;
      RECT 3.53 0.473 3.598 0.517 ;
      RECT 3.422 0.3155 3.49 0.3595 ;
      RECT 3.314 0.136 3.382 0.18 ;
      RECT 3.314 0.448 3.382 0.492 ;
      RECT 3.098 0.448 3.166 0.492 ;
      RECT 2.99 0.184 3.058 0.228 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.882 0.363 2.95 0.407 ;
      RECT 2.666 0.448 2.734 0.492 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.91 0.203 1.978 0.247 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.802 0.3155 1.87 0.3595 ;
      RECT 1.694 0.178 1.762 0.222 ;
      RECT 1.586 0.178 1.654 0.222 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.178 1.438 0.222 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.074 0.178 0.142 0.222 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 1.046 0.068 1.114 0.382 ;
      RECT 1.114 0.338 1.33 0.382 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.478 0.068 1.546 0.382 ;
      RECT 1.006 0.518 1.694 0.562 ;
      RECT 1.546 0.068 1.694 0.112 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 1.978 0.338 2.126 0.382 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.626 0.248 2.666 0.292 ;
      RECT 2.666 0.248 2.734 0.562 ;
      RECT 3.058 0.338 3.098 0.382 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 3.098 0.068 3.166 0.292 ;
      RECT 3.598 0.338 3.706 0.382 ;
      RECT 3.962 0.158 4.03 0.562 ;
      RECT 4.03 0.158 4.178 0.202 ;
      RECT 4.178 0.158 4.246 0.562 ;
      RECT 5.258 0.248 5.326 0.472 ;
      RECT 5.258 0.068 5.326 0.202 ;
      RECT 5.326 0.068 5.65 0.112 ;
      RECT 5.15 0.428 5.218 0.562 ;
      RECT 5.218 0.518 5.866 0.562 ;
      RECT 6.122 0.068 6.19 0.292 ;
      RECT 6.19 0.068 6.338 0.112 ;
      RECT 6.338 0.068 6.406 0.472 ;
      RECT 6.406 0.428 6.622 0.472 ;
      RECT 6.19 0.518 6.73 0.562 ;
  END
END b15fdw003hn1n30x5

MACRO b15fhw000hn1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fhw000hn1n05x5 0 0 ;
  SIZE 4.104 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 3.959111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 3.29925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
        RECT 0.29 0.248 0.358 0.382 ;
      LAYER m2 ;
        RECT 0.272 0.248 1.024 0.292 ;
      LAYER v1 ;
        RECT 0.294 0.248 0.354 0.292 ;
        RECT 0.942 0.248 1.002 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.158 3.058 0.472 ;
      LAYER v0 ;
        RECT 2.99 0.2705 3.058 0.3145 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.248 3.922 0.382 ;
      LAYER v0 ;
        RECT 3.854 0.293 3.922 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2731625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.13777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.518 3.186 0.562 ;
        RECT 2.882 0.158 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.2705 2.95 0.3145 ;
        RECT 3.098 0.518 3.166 0.562 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.138 0.652 ;
        RECT 3.314 0.338 3.382 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 2.018 0.473 2.086 0.517 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 3.314 0.3855 3.382 0.4295 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.138 0.022 ;
        RECT 3.854 -0.022 3.922 0.202 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.722 0.113 0.79 0.157 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 3.314 0.113 3.382 0.157 ;
        RECT 3.854 0.1185 3.922 0.1625 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.352 0.248 2.428 0.292 ;
      RECT 2.756 0.248 3.616 0.292 ;
    LAYER m1 ;
      RECT 0.29 0.248 0.358 0.382 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.83 0.158 1.046 0.202 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.154 0.068 1.222 0.472 ;
      RECT 1.37 0.248 1.438 0.382 ;
      RECT 1.802 0.248 2.234 0.292 ;
      RECT 2.126 0.158 2.342 0.202 ;
      RECT 2.558 0.158 2.626 0.382 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 2.774 0.248 2.842 0.562 ;
      RECT 3.206 0.248 3.422 0.292 ;
      RECT 3.53 0.248 3.598 0.472 ;
      RECT 3.422 0.338 3.49 0.562 ;
      RECT 3.962 0.068 4.03 0.472 ;
    LAYER v1 ;
      RECT 3.534 0.248 3.594 0.292 ;
      RECT 2.778 0.248 2.838 0.292 ;
      RECT 2.346 0.248 2.406 0.292 ;
      RECT 1.374 0.248 1.434 0.292 ;
    LAYER v0 ;
      RECT 3.962 0.1185 4.03 0.1625 ;
      RECT 3.962 0.408 4.03 0.452 ;
      RECT 3.854 0.518 3.922 0.562 ;
      RECT 3.746 0.428 3.814 0.472 ;
      RECT 3.638 0.172 3.706 0.216 ;
      RECT 3.53 0.3855 3.598 0.4295 ;
      RECT 3.422 0.3855 3.49 0.4295 ;
      RECT 3.314 0.248 3.382 0.292 ;
      RECT 3.098 0.363 3.166 0.407 ;
      RECT 3.1 0.138 3.164 0.182 ;
      RECT 2.774 0.498 2.842 0.542 ;
      RECT 2.558 0.293 2.626 0.337 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.408 0.682 0.452 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
    LAYER m1 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.682 0.248 0.898 0.292 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.546 0.338 2.194 0.382 ;
      RECT 2.234 0.248 2.302 0.472 ;
      RECT 2.342 0.158 2.41 0.562 ;
      RECT 2.626 0.158 2.774 0.202 ;
      RECT 2.774 0.068 2.842 0.202 ;
      RECT 2.842 0.068 3.098 0.112 ;
      RECT 3.098 0.068 3.166 0.472 ;
      RECT 3.422 0.068 3.49 0.292 ;
      RECT 3.49 0.068 3.638 0.112 ;
      RECT 3.638 0.068 3.706 0.472 ;
      RECT 3.706 0.428 3.922 0.472 ;
      RECT 3.49 0.518 4.03 0.562 ;
  END
END b15fhw000hn1n05x5

MACRO b15fhw000hn1n10x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fhw000hn1n10x5 0 0 ;
  SIZE 4.428 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
      ANTENNAMAXAREACAR 3.3244445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER m2 ;
        RECT 0.38 0.428 1.132 0.472 ;
      LAYER v1 ;
        RECT 0.402 0.428 0.462 0.472 ;
        RECT 1.05 0.428 1.11 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.3155 0.466 0.3595 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0117 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 3.29925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0117 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 3.29925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.158 3.382 0.382 ;
        RECT 2.882 0.158 2.95 0.382 ;
      LAYER m2 ;
        RECT 2.864 0.158 3.4 0.202 ;
      LAYER v1 ;
        RECT 2.886 0.158 2.946 0.202 ;
        RECT 3.318 0.158 3.378 0.202 ;
      LAYER v0 ;
        RECT 2.882 0.248 2.95 0.292 ;
        RECT 3.314 0.248 3.382 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.248 4.246 0.382 ;
      LAYER v0 ;
        RECT 4.178 0.293 4.246 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2731625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 4.13777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.518 3.51 0.562 ;
        RECT 3.206 0.248 3.274 0.562 ;
        RECT 2.99 0.248 3.274 0.292 ;
      LAYER v0 ;
        RECT 3.098 0.248 3.166 0.292 ;
        RECT 3.422 0.518 3.49 0.562 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.462 0.652 ;
        RECT 3.638 0.338 3.706 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.83 0.408 0.898 0.452 ;
        RECT 1.694 0.473 1.762 0.517 ;
        RECT 2.126 0.473 2.194 0.517 ;
        RECT 2.666 0.473 2.734 0.517 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.638 0.3855 3.706 0.4295 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.462 0.022 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.638 -0.022 3.706 0.202 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.113 0.898 0.157 ;
        RECT 1.478 0.113 1.546 0.157 ;
        RECT 1.694 0.113 1.762 0.157 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.666 0.138 2.734 0.182 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.638 0.113 3.706 0.157 ;
        RECT 4.178 0.1185 4.246 0.1625 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.46 0.428 2.552 0.472 ;
      RECT 2.632 0.428 3.94 0.472 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.938 0.158 1.154 0.202 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.262 0.068 1.33 0.562 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.91 0.248 2.342 0.292 ;
      RECT 2.234 0.158 2.45 0.202 ;
      RECT 2.774 0.068 2.842 0.382 ;
      RECT 2.558 0.068 2.626 0.562 ;
      RECT 2.774 0.428 2.842 0.562 ;
      RECT 2.882 0.158 2.95 0.382 ;
      RECT 3.314 0.158 3.382 0.382 ;
      RECT 3.53 0.248 3.962 0.292 ;
      RECT 3.854 0.338 3.922 0.472 ;
      RECT 3.746 0.338 3.814 0.562 ;
      RECT 4.286 0.068 4.354 0.472 ;
    LAYER v1 ;
      RECT 3.858 0.428 3.918 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.454 0.428 2.514 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
    LAYER v0 ;
      RECT 4.286 0.1185 4.354 0.1625 ;
      RECT 4.286 0.408 4.354 0.452 ;
      RECT 4.178 0.518 4.246 0.562 ;
      RECT 4.07 0.428 4.138 0.472 ;
      RECT 3.964 0.172 4.028 0.216 ;
      RECT 3.854 0.3855 3.922 0.4295 ;
      RECT 3.746 0.3855 3.814 0.4295 ;
      RECT 3.638 0.248 3.706 0.292 ;
      RECT 3.422 0.363 3.49 0.407 ;
      RECT 3.424 0.138 3.488 0.182 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.774 0.248 2.842 0.292 ;
      RECT 2.774 0.473 2.842 0.517 ;
      RECT 2.558 0.138 2.626 0.182 ;
      RECT 2.558 0.473 2.626 0.517 ;
      RECT 2.45 0.473 2.518 0.517 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.586 0.113 1.654 0.157 ;
      RECT 1.478 0.2705 1.546 0.3145 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.262 0.138 1.33 0.182 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.722 0.408 0.79 0.452 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.448 0.574 0.492 ;
    LAYER m1 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 0.79 0.248 1.006 0.292 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 1.33 0.518 1.586 0.562 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.654 0.338 2.302 0.382 ;
      RECT 2.342 0.248 2.41 0.472 ;
      RECT 2.45 0.158 2.518 0.562 ;
      RECT 2.842 0.068 2.99 0.112 ;
      RECT 2.99 0.068 3.058 0.202 ;
      RECT 3.058 0.158 3.206 0.202 ;
      RECT 3.206 0.068 3.274 0.202 ;
      RECT 3.274 0.068 3.422 0.112 ;
      RECT 3.422 0.068 3.49 0.472 ;
      RECT 3.962 0.068 4.03 0.472 ;
      RECT 4.03 0.428 4.246 0.472 ;
      RECT 3.814 0.518 4.354 0.562 ;
  END
END b15fhw000hn1n10x5

MACRO b15fhw000hn1n20x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fhw000hn1n20x5 0 0 ;
  SIZE 5.184 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 1.3004445 LAYER m1 ;
      ANTENNAMAXAREACAR 4.68533325 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.2515555 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.0243 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 2.2244445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.248 1.654 0.292 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER m2 ;
        RECT 0.704 0.248 1.564 0.292 ;
      LAYER v1 ;
        RECT 0.726 0.248 0.786 0.292 ;
        RECT 1.482 0.248 1.542 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.3155 0.79 0.3595 ;
        RECT 1.478 0.248 1.546 0.292 ;
    END
  END clk
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 3.861111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 3.861111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.934 0.248 5.002 0.382 ;
      LAYER m2 ;
        RECT 4.592 0.248 5.02 0.292 ;
      LAYER v1 ;
        RECT 4.938 0.248 4.998 0.292 ;
      LAYER v0 ;
        RECT 4.934 0.293 5.002 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 2.222963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.5214815 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0252 LAYER m2 ;
      ANTENNAMAXAREACAR 6.668889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.428 4.354 0.562 ;
        RECT 3.854 0.248 3.922 0.472 ;
        RECT 3.422 0.248 3.922 0.292 ;
      LAYER m2 ;
        RECT 3.836 0.428 4.372 0.472 ;
      LAYER v1 ;
        RECT 3.858 0.428 3.918 0.472 ;
        RECT 4.29 0.428 4.35 0.472 ;
      LAYER v0 ;
        RECT 3.53 0.248 3.598 0.292 ;
        RECT 4.286 0.498 4.354 0.542 ;
    END
  END ssb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.068 4.138 0.382 ;
      LAYER v0 ;
        RECT 4.07 0.293 4.138 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06732 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
        RECT 0.074 0.248 0.574 0.292 ;
        RECT 0.29 0.068 0.358 0.562 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.218 0.652 ;
        RECT 4.394 0.338 4.462 0.652 ;
        RECT 3.314 0.428 3.814 0.472 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 1.154 0.473 1.222 0.517 ;
        RECT 1.91 0.538 1.978 0.582 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.558 0.473 2.626 0.517 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.422 0.428 3.49 0.472 ;
        RECT 3.638 0.428 3.706 0.472 ;
        RECT 4.394 0.3855 4.462 0.4295 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.218 0.022 ;
        RECT 4.934 -0.022 5.002 0.202 ;
        RECT 4.394 -0.022 4.462 0.202 ;
        RECT 3.638 -0.022 3.706 0.112 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 1.154 0.113 1.222 0.157 ;
        RECT 1.91 0.136 1.978 0.18 ;
        RECT 2.126 0.136 2.194 0.18 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.424 0.048 3.488 0.092 ;
        RECT 3.64 0.048 3.704 0.092 ;
        RECT 4.394 0.113 4.462 0.157 ;
        RECT 4.934 0.1185 5.002 0.1625 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.812 0.338 2.444 0.382 ;
      RECT 1.568 0.428 2.768 0.472 ;
      RECT 2.524 0.338 2.876 0.382 ;
      RECT 1.892 0.248 2.984 0.292 ;
      RECT 2.848 0.428 3.292 0.472 ;
      RECT 3.064 0.248 4.264 0.292 ;
      RECT 3.512 0.338 4.696 0.382 ;
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 0.83 0.068 0.898 0.562 ;
      RECT 0.938 0.248 1.006 0.562 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.37 0.338 1.654 0.382 ;
      RECT 1.37 0.248 1.654 0.292 ;
      RECT 1.37 0.068 1.802 0.112 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 2.018 0.068 2.086 0.562 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.342 0.248 2.41 0.472 ;
      RECT 2.666 0.158 2.882 0.202 ;
      RECT 2.666 0.248 2.734 0.472 ;
      RECT 2.774 0.248 2.842 0.382 ;
      RECT 3.422 0.248 3.854 0.292 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.098 0.158 3.166 0.382 ;
      RECT 3.206 0.068 3.274 0.562 ;
      RECT 3.422 0.338 3.706 0.382 ;
      RECT 4.286 0.248 4.502 0.292 ;
      RECT 3.422 0.158 3.922 0.202 ;
      RECT 3.962 0.068 4.03 0.472 ;
      RECT 3.422 0.518 4.246 0.562 ;
      RECT 4.178 0.068 4.246 0.472 ;
      RECT 4.286 0.428 4.354 0.562 ;
      RECT 4.61 0.338 4.678 0.472 ;
      RECT 4.502 0.338 4.57 0.562 ;
      RECT 4.934 0.248 5.002 0.382 ;
      RECT 5.042 0.068 5.11 0.472 ;
    LAYER v1 ;
      RECT 4.614 0.338 4.674 0.382 ;
      RECT 4.182 0.248 4.242 0.292 ;
      RECT 3.966 0.248 4.026 0.292 ;
      RECT 3.534 0.338 3.594 0.382 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 3.102 0.248 3.162 0.292 ;
      RECT 2.994 0.428 3.054 0.472 ;
      RECT 2.886 0.248 2.946 0.292 ;
      RECT 2.778 0.338 2.838 0.382 ;
      RECT 2.67 0.428 2.73 0.472 ;
      RECT 2.562 0.338 2.622 0.382 ;
      RECT 2.346 0.338 2.406 0.382 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.914 0.248 1.974 0.292 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.482 0.338 1.542 0.382 ;
      RECT 0.834 0.338 0.894 0.382 ;
    LAYER v0 ;
      RECT 5.042 0.1185 5.11 0.1625 ;
      RECT 5.042 0.408 5.11 0.452 ;
      RECT 4.934 0.518 5.002 0.562 ;
      RECT 4.826 0.428 4.894 0.472 ;
      RECT 4.718 0.172 4.786 0.216 ;
      RECT 4.61 0.3855 4.678 0.4295 ;
      RECT 4.502 0.3855 4.57 0.4295 ;
      RECT 4.394 0.248 4.462 0.292 ;
      RECT 4.178 0.138 4.246 0.182 ;
      RECT 4.178 0.403 4.246 0.447 ;
      RECT 4.07 0.518 4.138 0.562 ;
      RECT 3.962 0.402 4.03 0.446 ;
      RECT 3.964 0.138 4.028 0.182 ;
      RECT 3.746 0.158 3.814 0.202 ;
      RECT 3.746 0.518 3.814 0.562 ;
      RECT 3.53 0.158 3.598 0.202 ;
      RECT 3.53 0.338 3.598 0.382 ;
      RECT 3.53 0.518 3.598 0.562 ;
      RECT 3.206 0.138 3.274 0.182 ;
      RECT 3.206 0.448 3.274 0.492 ;
      RECT 3.098 0.2705 3.166 0.3145 ;
      RECT 2.99 0.138 3.058 0.182 ;
      RECT 2.99 0.448 3.058 0.492 ;
      RECT 2.882 0.448 2.95 0.492 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.45 0.473 2.518 0.517 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.234 0.136 2.302 0.18 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.136 2.086 0.18 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 1.046 0.473 1.114 0.517 ;
      RECT 0.938 0.473 1.006 0.517 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.83 0.473 0.898 0.517 ;
    LAYER m1 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.338 1.33 0.382 ;
      RECT 1.006 0.248 1.262 0.292 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.33 0.158 1.694 0.202 ;
      RECT 1.694 0.158 1.762 0.562 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 2.518 0.338 2.626 0.382 ;
      RECT 2.882 0.158 2.95 0.562 ;
      RECT 3.854 0.248 3.922 0.472 ;
      RECT 4.502 0.068 4.57 0.292 ;
      RECT 4.57 0.068 4.718 0.112 ;
      RECT 4.718 0.068 4.786 0.472 ;
      RECT 4.786 0.428 5.002 0.472 ;
      RECT 4.57 0.518 5.11 0.562 ;
  END
END b15fhw000hn1n20x5

MACRO b15fhw000hn1n30x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fhw000hn1n30x5 0 0 ;
  SIZE 6.156 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 3.83166675 LAYER m1 ;
      ANTENNAMAXAREACAR 6.6524075 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAGATEAREA 0.036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.436875 LAYER m1 ;
      ANTENNAMAXAREACAR 2.49465275 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.391111 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.782 0.248 1.978 0.292 ;
        RECT 1.154 0.068 1.222 0.292 ;
      LAYER m2 ;
        RECT 1.136 0.248 1.888 0.292 ;
      LAYER v1 ;
        RECT 1.158 0.248 1.218 0.292 ;
        RECT 1.806 0.248 1.866 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.802 0.248 1.87 0.292 ;
    END
  END clk
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 3.861111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 3.861111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.906 0.248 5.974 0.382 ;
      LAYER m2 ;
        RECT 5.564 0.248 5.992 0.292 ;
      LAYER v1 ;
        RECT 5.91 0.248 5.97 0.292 ;
      LAYER v0 ;
        RECT 5.906 0.293 5.974 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 2.222963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.5214815 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0342 LAYER m2 ;
      ANTENNAMAXAREACAR 6.668889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.258 0.428 5.326 0.562 ;
        RECT 4.61 0.248 4.678 0.472 ;
        RECT 3.962 0.248 4.678 0.292 ;
      LAYER m2 ;
        RECT 4.592 0.428 5.344 0.472 ;
      LAYER v1 ;
        RECT 4.614 0.428 4.674 0.472 ;
        RECT 5.262 0.428 5.322 0.472 ;
      LAYER v0 ;
        RECT 4.07 0.248 4.138 0.292 ;
        RECT 4.286 0.248 4.354 0.292 ;
        RECT 5.258 0.498 5.326 0.542 ;
    END
  END ssb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.746489 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.042 0.068 5.11 0.382 ;
      LAYER v0 ;
        RECT 5.042 0.293 5.11 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.182 0.248 0.682 0.292 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.19 0.652 ;
        RECT 5.366 0.338 5.434 0.652 ;
        RECT 4.394 0.518 4.462 0.652 ;
        RECT 4.178 0.518 4.246 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.99 0.473 3.058 0.517 ;
        RECT 3.746 0.448 3.814 0.492 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 4.178 0.538 4.246 0.582 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 5.366 0.3855 5.434 0.4295 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.19 0.022 ;
        RECT 5.906 -0.022 5.974 0.202 ;
        RECT 5.366 -0.022 5.434 0.202 ;
        RECT 4.394 -0.022 4.462 0.112 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.37 0.1215 1.438 0.1655 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.45 0.136 2.518 0.18 ;
        RECT 2.99 0.138 3.058 0.182 ;
        RECT 3.748 0.048 3.812 0.092 ;
        RECT 3.964 0.048 4.028 0.092 ;
        RECT 4.18 0.048 4.244 0.092 ;
        RECT 4.396 0.048 4.46 0.092 ;
        RECT 5.366 0.113 5.434 0.157 ;
        RECT 5.906 0.1185 5.974 0.1625 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.428 1.796 0.472 ;
      RECT 1.028 0.338 2.644 0.382 ;
      RECT 1.876 0.428 3.308 0.472 ;
      RECT 2.972 0.338 3.508 0.382 ;
      RECT 2.216 0.248 3.632 0.292 ;
      RECT 3.388 0.428 3.94 0.472 ;
      RECT 3.712 0.248 5.236 0.292 ;
      RECT 4.268 0.338 5.668 0.382 ;
    LAYER m1 ;
      RECT 0.722 0.338 0.938 0.382 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.91 0.428 1.978 0.562 ;
      RECT 1.782 0.338 1.978 0.382 ;
      RECT 1.782 0.248 1.978 0.292 ;
      RECT 1.694 0.068 2.126 0.112 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 2.234 0.248 2.302 0.472 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.558 0.248 2.626 0.472 ;
      RECT 2.666 0.068 2.734 0.562 ;
      RECT 3.098 0.158 3.314 0.202 ;
      RECT 3.098 0.248 3.166 0.472 ;
      RECT 3.206 0.248 3.274 0.382 ;
      RECT 3.422 0.428 3.49 0.562 ;
      RECT 3.422 0.248 3.49 0.382 ;
      RECT 3.962 0.248 4.61 0.292 ;
      RECT 3.638 0.068 3.706 0.562 ;
      RECT 3.746 0.158 3.814 0.382 ;
      RECT 3.854 0.068 3.922 0.562 ;
      RECT 3.962 0.338 4.462 0.382 ;
      RECT 3.962 0.158 4.61 0.202 ;
      RECT 4.718 0.158 4.786 0.472 ;
      RECT 4.934 0.158 5.002 0.472 ;
      RECT 3.962 0.428 4.502 0.472 ;
      RECT 5.258 0.248 5.474 0.292 ;
      RECT 5.15 0.158 5.218 0.472 ;
      RECT 5.258 0.428 5.326 0.562 ;
      RECT 5.582 0.338 5.65 0.472 ;
      RECT 5.474 0.338 5.542 0.562 ;
      RECT 5.906 0.248 5.974 0.382 ;
      RECT 6.014 0.068 6.082 0.472 ;
    LAYER v1 ;
      RECT 5.586 0.338 5.646 0.382 ;
      RECT 5.154 0.248 5.214 0.292 ;
      RECT 4.938 0.248 4.998 0.292 ;
      RECT 4.722 0.248 4.782 0.292 ;
      RECT 4.29 0.338 4.35 0.382 ;
      RECT 3.858 0.428 3.918 0.472 ;
      RECT 3.75 0.248 3.81 0.292 ;
      RECT 3.642 0.428 3.702 0.472 ;
      RECT 3.534 0.248 3.594 0.292 ;
      RECT 3.426 0.338 3.486 0.382 ;
      RECT 3.426 0.428 3.486 0.472 ;
      RECT 3.318 0.248 3.378 0.292 ;
      RECT 3.21 0.338 3.27 0.382 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.994 0.338 3.054 0.382 ;
      RECT 2.562 0.338 2.622 0.382 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.238 0.248 2.298 0.292 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.806 0.338 1.866 0.382 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.482 0.338 1.542 0.382 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.942 0.428 1.002 0.472 ;
    LAYER v0 ;
      RECT 6.014 0.1185 6.082 0.1625 ;
      RECT 6.014 0.408 6.082 0.452 ;
      RECT 5.906 0.518 5.974 0.562 ;
      RECT 5.798 0.428 5.866 0.472 ;
      RECT 5.69 0.172 5.758 0.216 ;
      RECT 5.582 0.3855 5.65 0.4295 ;
      RECT 5.474 0.3855 5.542 0.4295 ;
      RECT 5.366 0.248 5.434 0.292 ;
      RECT 5.15 0.403 5.218 0.447 ;
      RECT 5.152 0.184 5.216 0.228 ;
      RECT 5.042 0.518 5.11 0.562 ;
      RECT 4.934 0.184 5.002 0.228 ;
      RECT 4.934 0.402 5.002 0.446 ;
      RECT 4.826 0.068 4.894 0.112 ;
      RECT 4.826 0.518 4.894 0.562 ;
      RECT 4.718 0.402 4.786 0.446 ;
      RECT 4.72 0.184 4.784 0.228 ;
      RECT 4.61 0.518 4.678 0.562 ;
      RECT 4.502 0.158 4.57 0.202 ;
      RECT 4.286 0.158 4.354 0.202 ;
      RECT 4.286 0.338 4.354 0.382 ;
      RECT 4.286 0.428 4.354 0.472 ;
      RECT 4.07 0.158 4.138 0.202 ;
      RECT 4.07 0.338 4.138 0.382 ;
      RECT 4.07 0.428 4.138 0.472 ;
      RECT 3.854 0.138 3.922 0.182 ;
      RECT 3.854 0.448 3.922 0.492 ;
      RECT 3.746 0.248 3.814 0.292 ;
      RECT 3.638 0.138 3.706 0.182 ;
      RECT 3.638 0.448 3.706 0.492 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.422 0.293 3.49 0.337 ;
      RECT 3.422 0.448 3.49 0.492 ;
      RECT 3.314 0.448 3.382 0.492 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.206 0.293 3.274 0.337 ;
      RECT 3.098 0.293 3.166 0.337 ;
      RECT 2.882 0.473 2.95 0.517 ;
      RECT 2.666 0.136 2.734 0.18 ;
      RECT 2.666 0.448 2.734 0.492 ;
      RECT 2.558 0.338 2.626 0.382 ;
      RECT 2.342 0.136 2.41 0.18 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.588 0.088 1.652 0.132 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.338 0.898 0.382 ;
    LAYER m1 ;
      RECT 0.722 0.248 1.046 0.292 ;
      RECT 1.046 0.248 1.114 0.382 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.006 0.518 1.242 0.562 ;
      RECT 1.654 0.158 2.018 0.202 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 2.126 0.068 2.194 0.562 ;
      RECT 2.95 0.338 3.058 0.382 ;
      RECT 3.314 0.158 3.382 0.562 ;
      RECT 3.382 0.158 3.53 0.202 ;
      RECT 3.53 0.158 3.598 0.562 ;
      RECT 4.61 0.248 4.678 0.472 ;
      RECT 4.61 0.068 4.678 0.202 ;
      RECT 4.678 0.068 5.002 0.112 ;
      RECT 4.502 0.428 4.57 0.562 ;
      RECT 4.57 0.518 5.218 0.562 ;
      RECT 5.474 0.068 5.542 0.292 ;
      RECT 5.542 0.068 5.69 0.112 ;
      RECT 5.69 0.068 5.758 0.472 ;
      RECT 5.758 0.428 5.974 0.472 ;
      RECT 5.542 0.518 6.082 0.562 ;
  END
END b15fhw000hn1n30x5

MACRO b15fmm200hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fmm200hn1n04x5 0 0 ;
  SIZE 7.128 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.70571425 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 6.986 0.068 7.054 0.562 ;
      LAYER v0 ;
        RECT 6.986 0.428 7.054 0.472 ;
        RECT 6.986 0.178 7.054 0.222 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 8.93 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.97666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 7.162 0.652 ;
        RECT 6.878 0.338 6.946 0.652 ;
        RECT 6.554 0.428 6.622 0.652 ;
        RECT 5.906 0.428 5.974 0.652 ;
        RECT 5.69 0.428 5.758 0.652 ;
        RECT 5.15 0.428 5.218 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 4.286 0.428 4.354 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.854 0.428 3.922 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4725 0.25 0.5165 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 4.07 0.538 4.138 0.582 ;
        RECT 4.286 0.448 4.354 0.492 ;
        RECT 4.502 0.448 4.57 0.492 ;
        RECT 5.15 0.448 5.218 0.492 ;
        RECT 5.69 0.448 5.758 0.492 ;
        RECT 5.906 0.448 5.974 0.492 ;
        RECT 6.554 0.493 6.622 0.537 ;
        RECT 6.878 0.428 6.946 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 7.162 0.022 ;
        RECT 6.878 -0.022 6.946 0.292 ;
        RECT 6.554 -0.022 6.622 0.292 ;
        RECT 5.906 -0.022 5.974 0.292 ;
        RECT 5.69 -0.022 5.758 0.292 ;
        RECT 5.15 -0.022 5.218 0.202 ;
        RECT 4.502 -0.022 4.57 0.202 ;
        RECT 4.286 -0.022 4.354 0.202 ;
        RECT 4.07 -0.022 4.138 0.202 ;
        RECT 3.854 -0.022 3.922 0.202 ;
        RECT 3.314 -0.022 3.382 0.292 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.074 0.158 0.27 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.45 0.1805 2.518 0.2245 ;
        RECT 2.666 0.1805 2.734 0.2245 ;
        RECT 3.314 0.1805 3.382 0.2245 ;
        RECT 3.854 0.138 3.922 0.182 ;
        RECT 4.07 0.138 4.138 0.182 ;
        RECT 4.286 0.138 4.354 0.182 ;
        RECT 4.502 0.138 4.57 0.182 ;
        RECT 5.15 0.138 5.218 0.182 ;
        RECT 5.69 0.203 5.758 0.247 ;
        RECT 5.906 0.203 5.974 0.247 ;
        RECT 6.554 0.158 6.622 0.202 ;
        RECT 6.878 0.178 6.946 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.892 0.518 2.644 0.562 ;
      RECT 2.108 0.428 4.696 0.472 ;
      RECT 1.244 0.068 6.424 0.112 ;
    LAYER m1 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.262 0.068 1.33 0.562 ;
      RECT 2.99 0.338 3.058 0.562 ;
      RECT 2.018 0.248 2.086 0.562 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 2.774 0.158 2.842 0.562 ;
      RECT 2.882 0.068 2.95 0.562 ;
      RECT 3.746 0.338 3.814 0.562 ;
      RECT 3.638 0.068 3.706 0.562 ;
      RECT 4.178 0.158 4.246 0.562 ;
      RECT 4.394 0.068 4.462 0.202 ;
      RECT 4.61 0.428 4.678 0.562 ;
      RECT 4.718 0.068 4.786 0.202 ;
      RECT 4.826 0.338 4.894 0.562 ;
      RECT 5.474 0.068 5.542 0.202 ;
      RECT 5.474 0.338 5.542 0.562 ;
      RECT 6.122 0.158 6.19 0.472 ;
      RECT 6.014 0.158 6.082 0.562 ;
      RECT 6.338 0.068 6.406 0.382 ;
      RECT 6.662 0.068 6.73 0.292 ;
    LAYER v1 ;
      RECT 6.342 0.068 6.402 0.112 ;
      RECT 5.478 0.068 5.538 0.112 ;
      RECT 4.722 0.068 4.782 0.112 ;
      RECT 4.614 0.428 4.674 0.472 ;
      RECT 4.398 0.068 4.458 0.112 ;
      RECT 3.642 0.068 3.702 0.112 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 2.562 0.518 2.622 0.562 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 2.022 0.518 2.082 0.562 ;
      RECT 1.266 0.068 1.326 0.112 ;
    LAYER v0 ;
      RECT 6.77 0.428 6.838 0.472 ;
      RECT 6.662 0.158 6.73 0.202 ;
      RECT 6.554 0.338 6.622 0.382 ;
      RECT 6.338 0.088 6.406 0.132 ;
      RECT 6.338 0.3155 6.406 0.3595 ;
      RECT 6.23 0.428 6.298 0.472 ;
      RECT 6.122 0.203 6.19 0.247 ;
      RECT 6.014 0.203 6.082 0.247 ;
      RECT 6.014 0.448 6.082 0.492 ;
      RECT 5.798 0.203 5.866 0.247 ;
      RECT 5.798 0.448 5.866 0.492 ;
      RECT 5.582 0.113 5.65 0.157 ;
      RECT 5.474 0.113 5.542 0.157 ;
      RECT 5.474 0.448 5.542 0.492 ;
      RECT 5.366 0.113 5.434 0.157 ;
      RECT 5.366 0.448 5.434 0.492 ;
      RECT 4.934 0.138 5.002 0.182 ;
      RECT 4.826 0.138 4.894 0.182 ;
      RECT 4.826 0.448 4.894 0.492 ;
      RECT 4.718 0.138 4.786 0.182 ;
      RECT 4.718 0.448 4.786 0.492 ;
      RECT 4.61 0.448 4.678 0.492 ;
      RECT 4.394 0.138 4.462 0.182 ;
      RECT 4.178 0.223 4.246 0.267 ;
      RECT 4.178 0.448 4.246 0.492 ;
      RECT 3.962 0.138 4.03 0.182 ;
      RECT 3.962 0.448 4.03 0.492 ;
      RECT 3.746 0.448 3.814 0.492 ;
      RECT 3.638 0.448 3.706 0.492 ;
      RECT 3.53 0.138 3.598 0.182 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.098 0.191 3.166 0.235 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.882 0.088 2.95 0.132 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.774 0.1805 2.842 0.2245 ;
      RECT 2.774 0.448 2.842 0.492 ;
      RECT 2.558 0.1805 2.626 0.2245 ;
      RECT 2.558 0.448 2.626 0.492 ;
      RECT 2.234 0.138 2.302 0.182 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.478 0.191 1.546 0.235 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.133 1.33 0.177 ;
      RECT 1.262 0.3155 1.33 0.3595 ;
      RECT 1.154 0.133 1.222 0.177 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 0.938 0.138 1.006 0.182 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.898 0.338 1.114 0.382 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.438 0.338 1.478 0.382 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.546 0.338 1.91 0.382 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 3.058 0.338 3.098 0.382 ;
      RECT 3.098 0.158 3.166 0.382 ;
      RECT 3.166 0.338 3.53 0.382 ;
      RECT 3.53 0.068 3.598 0.562 ;
      RECT 3.814 0.338 3.962 0.382 ;
      RECT 3.962 0.068 4.03 0.562 ;
      RECT 4.246 0.338 4.718 0.382 ;
      RECT 4.718 0.248 4.786 0.562 ;
      RECT 4.786 0.248 4.826 0.292 ;
      RECT 4.826 0.068 4.894 0.292 ;
      RECT 4.894 0.338 4.934 0.382 ;
      RECT 4.934 0.068 5.002 0.382 ;
      RECT 5.002 0.338 5.366 0.382 ;
      RECT 5.366 0.068 5.434 0.562 ;
      RECT 5.434 0.248 5.582 0.292 ;
      RECT 5.582 0.068 5.65 0.292 ;
      RECT 5.542 0.338 5.798 0.382 ;
      RECT 5.798 0.158 5.866 0.562 ;
      RECT 6.19 0.428 6.446 0.472 ;
      RECT 6.446 0.338 6.514 0.472 ;
      RECT 6.514 0.338 6.73 0.382 ;
      RECT 6.73 0.248 6.77 0.292 ;
      RECT 6.77 0.248 6.838 0.562 ;
  END
END b15fmm200hn1n04x5

MACRO b15fmm203hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fmm203hn1n04x5 0 0 ;
  SIZE 8.64 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAGATEAREA 0.0504 LAYER m2 ;
      ANTENNAMAXAREACAR 1.946923 LAYER m1 ;
      ANTENNAMAXAREACAR 3.2488035 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4813675 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAGATEAREA 0.0612 LAYER m2 ;
      ANTENNAMAXAREACAR 1.82 LAYER m1 ;
      ANTENNAMAXAREACAR 2.8155555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.3681045 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 6.338 0.428 6.406 0.562 ;
        RECT 3.962 0.428 4.03 0.562 ;
        RECT 3.206 0.338 3.274 0.562 ;
      LAYER m2 ;
        RECT 3.188 0.518 6.424 0.562 ;
      LAYER v1 ;
        RECT 3.21 0.518 3.27 0.562 ;
        RECT 3.966 0.518 4.026 0.562 ;
        RECT 6.342 0.518 6.402 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.364 3.274 0.408 ;
        RECT 3.962 0.448 4.03 0.492 ;
        RECT 6.338 0.448 6.406 0.492 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53079375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.31901225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 8.498 0.068 8.566 0.562 ;
      LAYER v0 ;
        RECT 8.498 0.428 8.566 0.472 ;
        RECT 8.498 0.152 8.566 0.196 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 8.93 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.97666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
        RECT 0.182 0.068 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 8.674 0.652 ;
        RECT 8.39 0.338 8.458 0.652 ;
        RECT 7.634 0.428 7.702 0.652 ;
        RECT 7.094 0.428 7.162 0.652 ;
        RECT 6.878 0.338 6.946 0.652 ;
        RECT 6.662 0.428 6.73 0.652 ;
        RECT 6.446 0.428 6.514 0.652 ;
        RECT 5.906 0.428 5.974 0.652 ;
        RECT 5.258 0.428 5.326 0.652 ;
        RECT 5.042 0.428 5.11 0.652 ;
        RECT 4.826 0.518 4.894 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 4.286 0.338 4.354 0.652 ;
        RECT 4.07 0.428 4.138 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4725 0.25 0.5165 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 4.07 0.448 4.138 0.492 ;
        RECT 4.286 0.448 4.354 0.492 ;
        RECT 4.502 0.448 4.57 0.492 ;
        RECT 4.826 0.538 4.894 0.582 ;
        RECT 5.042 0.448 5.11 0.492 ;
        RECT 5.258 0.448 5.326 0.492 ;
        RECT 5.906 0.448 5.974 0.492 ;
        RECT 6.446 0.448 6.514 0.492 ;
        RECT 6.662 0.448 6.73 0.492 ;
        RECT 6.878 0.448 6.946 0.492 ;
        RECT 7.094 0.448 7.162 0.492 ;
        RECT 7.634 0.448 7.702 0.492 ;
        RECT 8.39 0.428 8.458 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 8.674 0.022 ;
        RECT 8.39 -0.022 8.458 0.202 ;
        RECT 7.526 -0.022 7.594 0.202 ;
        RECT 6.878 -0.022 6.946 0.202 ;
        RECT 6.446 -0.022 6.514 0.202 ;
        RECT 5.906 -0.022 5.974 0.202 ;
        RECT 5.258 -0.022 5.326 0.202 ;
        RECT 5.042 -0.022 5.11 0.112 ;
        RECT 4.826 -0.022 4.894 0.202 ;
        RECT 4.61 -0.022 4.678 0.202 ;
        RECT 4.07 -0.022 4.138 0.112 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 4.072 0.048 4.136 0.092 ;
        RECT 4.61 0.138 4.678 0.182 ;
        RECT 4.826 0.138 4.894 0.182 ;
        RECT 5.042 0.048 5.11 0.092 ;
        RECT 5.258 0.138 5.326 0.182 ;
        RECT 5.906 0.138 5.974 0.182 ;
        RECT 6.446 0.138 6.514 0.182 ;
        RECT 6.878 0.138 6.946 0.182 ;
        RECT 7.526 0.138 7.594 0.182 ;
        RECT 8.39 0.068 8.458 0.112 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.784 0.518 2.86 0.562 ;
      RECT 2.216 0.428 8.152 0.472 ;
      RECT 1.244 0.068 8.26 0.112 ;
      RECT 7.184 0.518 8.6 0.562 ;
    LAYER m1 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 1.262 0.428 1.586 0.472 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.99 0.338 3.058 0.562 ;
      RECT 3.206 0.338 3.274 0.562 ;
      RECT 3.314 0.338 3.382 0.562 ;
      RECT 3.638 0.158 3.706 0.562 ;
      RECT 3.962 0.428 4.03 0.562 ;
      RECT 3.962 0.068 4.03 0.202 ;
      RECT 3.314 0.158 3.53 0.202 ;
      RECT 4.934 0.068 5.002 0.562 ;
      RECT 4.718 0.068 4.786 0.562 ;
      RECT 5.15 0.068 5.218 0.202 ;
      RECT 5.366 0.428 5.434 0.562 ;
      RECT 5.474 0.068 5.542 0.202 ;
      RECT 5.582 0.338 5.65 0.562 ;
      RECT 6.23 0.068 6.298 0.202 ;
      RECT 6.338 0.428 6.406 0.562 ;
      RECT 6.23 0.338 6.298 0.562 ;
      RECT 7.526 0.338 7.594 0.562 ;
      RECT 7.31 0.158 7.378 0.562 ;
      RECT 7.418 0.338 7.486 0.562 ;
      RECT 7.85 0.248 7.918 0.562 ;
      RECT 8.066 0.428 8.134 0.562 ;
      RECT 6.986 0.338 7.054 0.562 ;
      RECT 8.282 0.158 8.35 0.562 ;
      RECT 7.958 0.068 8.35 0.112 ;
    LAYER v1 ;
      RECT 8.286 0.518 8.346 0.562 ;
      RECT 8.178 0.068 8.238 0.112 ;
      RECT 8.07 0.428 8.13 0.472 ;
      RECT 7.854 0.518 7.914 0.562 ;
      RECT 7.422 0.518 7.482 0.562 ;
      RECT 6.234 0.068 6.294 0.112 ;
      RECT 5.478 0.068 5.538 0.112 ;
      RECT 5.37 0.428 5.43 0.472 ;
      RECT 5.154 0.068 5.214 0.112 ;
      RECT 3.966 0.068 4.026 0.112 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 2.778 0.518 2.838 0.562 ;
      RECT 2.562 0.518 2.622 0.562 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.266 0.068 1.326 0.112 ;
    LAYER v0 ;
      RECT 8.282 0.248 8.35 0.292 ;
      RECT 8.174 0.068 8.242 0.112 ;
      RECT 8.066 0.158 8.134 0.202 ;
      RECT 8.066 0.448 8.134 0.492 ;
      RECT 7.958 0.248 8.026 0.292 ;
      RECT 7.958 0.448 8.026 0.492 ;
      RECT 7.85 0.448 7.918 0.492 ;
      RECT 7.742 0.448 7.81 0.492 ;
      RECT 7.526 0.448 7.594 0.492 ;
      RECT 7.418 0.448 7.486 0.492 ;
      RECT 7.31 0.178 7.378 0.222 ;
      RECT 7.31 0.448 7.378 0.492 ;
      RECT 7.094 0.248 7.162 0.292 ;
      RECT 6.986 0.448 7.054 0.492 ;
      RECT 6.77 0.448 6.838 0.492 ;
      RECT 6.662 0.158 6.73 0.202 ;
      RECT 6.554 0.448 6.622 0.492 ;
      RECT 6.338 0.138 6.406 0.182 ;
      RECT 6.23 0.138 6.298 0.182 ;
      RECT 6.23 0.448 6.298 0.492 ;
      RECT 6.122 0.138 6.19 0.182 ;
      RECT 6.122 0.448 6.19 0.492 ;
      RECT 5.69 0.138 5.758 0.182 ;
      RECT 5.582 0.138 5.65 0.182 ;
      RECT 5.582 0.448 5.65 0.492 ;
      RECT 5.474 0.138 5.542 0.182 ;
      RECT 5.474 0.448 5.542 0.492 ;
      RECT 5.366 0.448 5.434 0.492 ;
      RECT 5.15 0.138 5.218 0.182 ;
      RECT 4.934 0.138 5.002 0.182 ;
      RECT 4.934 0.448 5.002 0.492 ;
      RECT 4.718 0.138 4.786 0.182 ;
      RECT 4.718 0.428 4.786 0.472 ;
      RECT 4.502 0.293 4.57 0.337 ;
      RECT 4.394 0.448 4.462 0.492 ;
      RECT 4.286 0.248 4.354 0.292 ;
      RECT 4.178 0.448 4.246 0.492 ;
      RECT 3.962 0.138 4.03 0.182 ;
      RECT 3.746 0.178 3.814 0.222 ;
      RECT 3.746 0.408 3.814 0.452 ;
      RECT 3.638 0.178 3.706 0.222 ;
      RECT 3.638 0.408 3.706 0.452 ;
      RECT 3.53 0.408 3.598 0.452 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.422 0.493 3.49 0.537 ;
      RECT 3.314 0.493 3.382 0.537 ;
      RECT 3.098 0.178 3.166 0.222 ;
      RECT 2.99 0.448 3.058 0.492 ;
      RECT 2.774 0.448 2.842 0.492 ;
      RECT 2.666 0.178 2.734 0.222 ;
      RECT 2.558 0.448 2.626 0.492 ;
      RECT 2.234 0.138 2.302 0.182 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.088 1.33 0.132 ;
      RECT 1.262 0.3155 1.33 0.3595 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.94 0.178 1.004 0.222 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.4725 0.574 0.5165 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.898 0.338 1.114 0.382 ;
      RECT 0.83 0.428 1.154 0.472 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 1.222 0.518 1.438 0.562 ;
      RECT 1.87 0.428 1.91 0.472 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 1.37 0.158 1.586 0.202 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.158 1.87 0.382 ;
      RECT 1.87 0.158 2.086 0.202 ;
      RECT 2.626 0.338 2.666 0.382 ;
      RECT 2.666 0.158 2.734 0.382 ;
      RECT 2.734 0.338 2.774 0.382 ;
      RECT 2.774 0.338 2.842 0.562 ;
      RECT 3.058 0.338 3.098 0.382 ;
      RECT 3.098 0.158 3.166 0.382 ;
      RECT 3.166 0.248 3.422 0.292 ;
      RECT 3.422 0.248 3.49 0.562 ;
      RECT 3.706 0.518 3.854 0.562 ;
      RECT 3.854 0.338 3.922 0.562 ;
      RECT 3.922 0.338 4.178 0.382 ;
      RECT 4.178 0.248 4.246 0.562 ;
      RECT 4.246 0.248 4.394 0.292 ;
      RECT 4.394 0.248 4.462 0.562 ;
      RECT 3.53 0.068 3.598 0.562 ;
      RECT 3.598 0.068 3.746 0.112 ;
      RECT 3.746 0.068 3.814 0.472 ;
      RECT 3.814 0.248 4.07 0.292 ;
      RECT 4.07 0.158 4.138 0.292 ;
      RECT 4.138 0.158 4.502 0.202 ;
      RECT 4.502 0.158 4.57 0.382 ;
      RECT 5.002 0.248 5.474 0.292 ;
      RECT 5.474 0.248 5.542 0.562 ;
      RECT 5.542 0.248 5.582 0.292 ;
      RECT 5.582 0.068 5.65 0.292 ;
      RECT 5.65 0.338 5.69 0.382 ;
      RECT 5.69 0.068 5.758 0.382 ;
      RECT 5.758 0.338 6.122 0.382 ;
      RECT 6.122 0.068 6.19 0.562 ;
      RECT 6.19 0.248 6.338 0.292 ;
      RECT 6.338 0.068 6.406 0.292 ;
      RECT 6.298 0.338 6.554 0.382 ;
      RECT 6.554 0.158 6.622 0.562 ;
      RECT 6.622 0.158 6.77 0.202 ;
      RECT 6.77 0.158 6.838 0.562 ;
      RECT 7.594 0.338 7.742 0.382 ;
      RECT 7.742 0.338 7.81 0.562 ;
      RECT 7.918 0.248 8.134 0.292 ;
      RECT 7.054 0.338 7.094 0.382 ;
      RECT 7.094 0.068 7.162 0.382 ;
      RECT 7.162 0.068 7.418 0.112 ;
      RECT 7.418 0.068 7.486 0.292 ;
      RECT 7.486 0.248 7.742 0.292 ;
      RECT 7.742 0.158 7.81 0.292 ;
      RECT 7.958 0.338 8.026 0.562 ;
      RECT 8.026 0.338 8.174 0.382 ;
      RECT 7.81 0.158 8.174 0.202 ;
      RECT 8.174 0.158 8.242 0.382 ;
  END
END b15fmm203hn1n04x5

MACRO b15fmm20chn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fmm20chn1n04x5 0 0 ;
  SIZE 8.532 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAGATEAREA 0.0504 LAYER m2 ;
      ANTENNAMAXAREACAR 1.946923 LAYER m1 ;
      ANTENNAMAXAREACAR 3.2488035 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4813675 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAGATEAREA 0.0612 LAYER m2 ;
      ANTENNAMAXAREACAR 1.82 LAYER m1 ;
      ANTENNAMAXAREACAR 2.8155555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.3681045 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 6.23 0.428 6.298 0.562 ;
        RECT 3.854 0.428 3.922 0.562 ;
        RECT 3.098 0.338 3.166 0.562 ;
      LAYER m2 ;
        RECT 3.08 0.518 6.316 0.562 ;
      LAYER v1 ;
        RECT 3.102 0.518 3.162 0.562 ;
        RECT 3.858 0.518 3.918 0.562 ;
        RECT 6.234 0.518 6.294 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.364 3.166 0.408 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 6.23 0.448 6.298 0.492 ;
    END
  END psb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53079375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.158 2.302 0.472 ;
      LAYER v0 ;
        RECT 2.234 0.293 2.302 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.92239325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.856508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 8.39 0.068 8.458 0.562 ;
      LAYER v0 ;
        RECT 8.39 0.403 8.458 0.447 ;
        RECT 8.39 0.178 8.458 0.222 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 12.35 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 2.7444445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
        RECT 0.182 0.068 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 8.566 0.652 ;
        RECT 8.282 0.338 8.35 0.652 ;
        RECT 7.526 0.428 7.594 0.652 ;
        RECT 6.986 0.428 7.054 0.652 ;
        RECT 6.77 0.338 6.838 0.652 ;
        RECT 6.554 0.428 6.622 0.652 ;
        RECT 6.338 0.428 6.406 0.652 ;
        RECT 5.798 0.428 5.866 0.652 ;
        RECT 5.15 0.428 5.218 0.652 ;
        RECT 4.934 0.428 5.002 0.652 ;
        RECT 4.718 0.518 4.786 0.652 ;
        RECT 4.394 0.428 4.462 0.652 ;
        RECT 4.178 0.338 4.246 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4725 0.25 0.5165 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.962 0.448 4.03 0.492 ;
        RECT 4.178 0.448 4.246 0.492 ;
        RECT 4.394 0.448 4.462 0.492 ;
        RECT 4.718 0.538 4.786 0.582 ;
        RECT 4.934 0.448 5.002 0.492 ;
        RECT 5.15 0.448 5.218 0.492 ;
        RECT 5.798 0.448 5.866 0.492 ;
        RECT 6.338 0.448 6.406 0.492 ;
        RECT 6.554 0.448 6.622 0.492 ;
        RECT 6.77 0.448 6.838 0.492 ;
        RECT 6.986 0.448 7.054 0.492 ;
        RECT 7.526 0.448 7.594 0.492 ;
        RECT 8.282 0.403 8.35 0.447 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 8.566 0.022 ;
        RECT 8.282 -0.022 8.35 0.292 ;
        RECT 7.418 -0.022 7.486 0.202 ;
        RECT 6.77 -0.022 6.838 0.202 ;
        RECT 6.338 -0.022 6.406 0.202 ;
        RECT 5.798 -0.022 5.866 0.202 ;
        RECT 5.15 -0.022 5.218 0.202 ;
        RECT 4.934 -0.022 5.002 0.112 ;
        RECT 4.718 -0.022 4.786 0.112 ;
        RECT 4.502 -0.022 4.57 0.202 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.074 0.158 0.27 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 3.964 0.048 4.028 0.092 ;
        RECT 4.502 0.138 4.57 0.182 ;
        RECT 4.72 0.048 4.784 0.092 ;
        RECT 4.934 0.048 5.002 0.092 ;
        RECT 5.15 0.138 5.218 0.182 ;
        RECT 5.798 0.138 5.866 0.182 ;
        RECT 6.338 0.138 6.406 0.182 ;
        RECT 6.77 0.138 6.838 0.182 ;
        RECT 7.418 0.138 7.486 0.182 ;
        RECT 8.282 0.178 8.35 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.676 0.518 2.752 0.562 ;
      RECT 2.108 0.428 8.044 0.472 ;
      RECT 7.076 0.518 8.152 0.562 ;
      RECT 1.136 0.068 8.152 0.112 ;
    LAYER m1 ;
      RECT 1.694 0.428 1.762 0.562 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.154 0.428 1.37 0.472 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.126 0.068 2.194 0.562 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 3.206 0.338 3.274 0.562 ;
      RECT 3.53 0.158 3.598 0.562 ;
      RECT 3.854 0.428 3.922 0.562 ;
      RECT 3.854 0.068 3.922 0.202 ;
      RECT 3.206 0.158 3.422 0.202 ;
      RECT 4.826 0.068 4.894 0.562 ;
      RECT 4.61 0.068 4.678 0.562 ;
      RECT 5.042 0.068 5.11 0.202 ;
      RECT 5.258 0.428 5.326 0.562 ;
      RECT 5.366 0.068 5.434 0.202 ;
      RECT 5.474 0.338 5.542 0.562 ;
      RECT 6.122 0.068 6.19 0.202 ;
      RECT 6.23 0.428 6.298 0.562 ;
      RECT 6.122 0.338 6.19 0.562 ;
      RECT 7.418 0.338 7.486 0.562 ;
      RECT 7.202 0.158 7.27 0.562 ;
      RECT 7.31 0.338 7.378 0.562 ;
      RECT 7.742 0.248 7.81 0.562 ;
      RECT 7.958 0.428 8.026 0.562 ;
      RECT 6.878 0.338 6.946 0.562 ;
      RECT 8.066 0.428 8.134 0.562 ;
      RECT 7.85 0.068 8.242 0.112 ;
    LAYER v1 ;
      RECT 8.07 0.068 8.13 0.112 ;
      RECT 8.07 0.518 8.13 0.562 ;
      RECT 7.962 0.428 8.022 0.472 ;
      RECT 7.746 0.518 7.806 0.562 ;
      RECT 7.314 0.518 7.374 0.562 ;
      RECT 6.126 0.068 6.186 0.112 ;
      RECT 5.37 0.068 5.43 0.112 ;
      RECT 5.262 0.428 5.322 0.472 ;
      RECT 5.046 0.068 5.106 0.112 ;
      RECT 3.858 0.068 3.918 0.112 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 2.67 0.518 2.73 0.562 ;
      RECT 2.454 0.518 2.514 0.562 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.698 0.518 1.758 0.562 ;
      RECT 1.158 0.068 1.218 0.112 ;
    LAYER v0 ;
      RECT 8.066 0.068 8.134 0.112 ;
      RECT 8.066 0.448 8.134 0.492 ;
      RECT 7.958 0.158 8.026 0.202 ;
      RECT 7.958 0.448 8.026 0.492 ;
      RECT 7.85 0.248 7.918 0.292 ;
      RECT 7.85 0.448 7.918 0.492 ;
      RECT 7.742 0.448 7.81 0.492 ;
      RECT 7.634 0.448 7.702 0.492 ;
      RECT 7.418 0.448 7.486 0.492 ;
      RECT 7.31 0.448 7.378 0.492 ;
      RECT 7.202 0.178 7.27 0.222 ;
      RECT 7.202 0.448 7.27 0.492 ;
      RECT 6.986 0.248 7.054 0.292 ;
      RECT 6.878 0.448 6.946 0.492 ;
      RECT 6.662 0.448 6.73 0.492 ;
      RECT 6.554 0.158 6.622 0.202 ;
      RECT 6.446 0.448 6.514 0.492 ;
      RECT 6.23 0.138 6.298 0.182 ;
      RECT 6.122 0.138 6.19 0.182 ;
      RECT 6.122 0.448 6.19 0.492 ;
      RECT 6.014 0.138 6.082 0.182 ;
      RECT 6.014 0.448 6.082 0.492 ;
      RECT 5.582 0.138 5.65 0.182 ;
      RECT 5.474 0.138 5.542 0.182 ;
      RECT 5.474 0.448 5.542 0.492 ;
      RECT 5.366 0.138 5.434 0.182 ;
      RECT 5.366 0.448 5.434 0.492 ;
      RECT 5.258 0.448 5.326 0.492 ;
      RECT 5.042 0.138 5.11 0.182 ;
      RECT 4.826 0.448 4.894 0.492 ;
      RECT 4.828 0.168 4.892 0.212 ;
      RECT 4.61 0.138 4.678 0.182 ;
      RECT 4.61 0.428 4.678 0.472 ;
      RECT 4.394 0.293 4.462 0.337 ;
      RECT 4.286 0.448 4.354 0.492 ;
      RECT 4.178 0.248 4.246 0.292 ;
      RECT 4.07 0.448 4.138 0.492 ;
      RECT 3.854 0.138 3.922 0.182 ;
      RECT 3.638 0.178 3.706 0.222 ;
      RECT 3.638 0.408 3.706 0.452 ;
      RECT 3.53 0.178 3.598 0.222 ;
      RECT 3.53 0.408 3.598 0.452 ;
      RECT 3.422 0.408 3.49 0.452 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.314 0.493 3.382 0.537 ;
      RECT 3.206 0.493 3.274 0.537 ;
      RECT 2.99 0.178 3.058 0.222 ;
      RECT 2.882 0.448 2.95 0.492 ;
      RECT 2.666 0.448 2.734 0.492 ;
      RECT 2.558 0.178 2.626 0.222 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.37 0.191 1.438 0.235 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.3155 1.222 0.3595 ;
      RECT 1.046 0.4355 1.114 0.4795 ;
      RECT 1.048 0.178 1.112 0.222 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.456 0.574 0.5 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.762 0.428 1.802 0.472 ;
      RECT 1.802 0.248 1.87 0.472 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 1.438 0.338 1.694 0.382 ;
      RECT 1.694 0.158 1.762 0.382 ;
      RECT 1.762 0.158 1.978 0.202 ;
      RECT 2.518 0.338 2.558 0.382 ;
      RECT 2.558 0.158 2.626 0.382 ;
      RECT 2.626 0.338 2.666 0.382 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.95 0.338 2.99 0.382 ;
      RECT 2.99 0.158 3.058 0.382 ;
      RECT 3.058 0.248 3.314 0.292 ;
      RECT 3.314 0.248 3.382 0.562 ;
      RECT 3.598 0.518 3.746 0.562 ;
      RECT 3.746 0.338 3.814 0.562 ;
      RECT 3.814 0.338 4.07 0.382 ;
      RECT 4.07 0.248 4.138 0.562 ;
      RECT 4.138 0.248 4.286 0.292 ;
      RECT 4.286 0.248 4.354 0.562 ;
      RECT 3.422 0.068 3.49 0.562 ;
      RECT 3.49 0.068 3.638 0.112 ;
      RECT 3.638 0.068 3.706 0.472 ;
      RECT 3.706 0.248 3.962 0.292 ;
      RECT 3.962 0.158 4.03 0.292 ;
      RECT 4.03 0.158 4.394 0.202 ;
      RECT 4.394 0.158 4.462 0.382 ;
      RECT 4.894 0.248 5.366 0.292 ;
      RECT 5.366 0.248 5.434 0.562 ;
      RECT 5.434 0.248 5.474 0.292 ;
      RECT 5.474 0.068 5.542 0.292 ;
      RECT 5.542 0.338 5.582 0.382 ;
      RECT 5.582 0.068 5.65 0.382 ;
      RECT 5.65 0.338 6.014 0.382 ;
      RECT 6.014 0.068 6.082 0.562 ;
      RECT 6.082 0.248 6.23 0.292 ;
      RECT 6.23 0.068 6.298 0.292 ;
      RECT 6.19 0.338 6.446 0.382 ;
      RECT 6.446 0.158 6.514 0.562 ;
      RECT 6.514 0.158 6.662 0.202 ;
      RECT 6.662 0.158 6.73 0.562 ;
      RECT 7.486 0.338 7.634 0.382 ;
      RECT 7.634 0.338 7.702 0.562 ;
      RECT 7.81 0.248 8.026 0.292 ;
      RECT 6.946 0.338 6.986 0.382 ;
      RECT 6.986 0.068 7.054 0.382 ;
      RECT 7.054 0.068 7.31 0.112 ;
      RECT 7.31 0.068 7.378 0.292 ;
      RECT 7.378 0.248 7.634 0.292 ;
      RECT 7.634 0.158 7.702 0.292 ;
      RECT 7.85 0.338 7.918 0.562 ;
      RECT 7.918 0.338 8.066 0.382 ;
      RECT 7.702 0.158 8.066 0.202 ;
      RECT 8.066 0.158 8.134 0.382 ;
  END
END b15fmm20chn1n04x5

MACRO b15fmm300hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fmm300hn1n04x5 0 0 ;
  SIZE 10.26 BY 0.63 ;
  SYMMETRY Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.84941175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.84941175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.158 2.518 0.472 ;
      LAYER v0 ;
        RECT 2.45 0.293 2.518 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 10.118 0.068 10.186 0.562 ;
      LAYER v0 ;
        RECT 10.118 0.428 10.186 0.472 ;
        RECT 10.118 0.138 10.186 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 8.93 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.97666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 10.294 0.652 ;
        RECT 10.01 0.338 10.078 0.652 ;
        RECT 9.686 0.428 9.754 0.652 ;
        RECT 9.038 0.428 9.106 0.652 ;
        RECT 8.822 0.428 8.89 0.652 ;
        RECT 8.39 0.428 8.458 0.652 ;
        RECT 7.742 0.428 7.81 0.652 ;
        RECT 7.526 0.428 7.594 0.652 ;
        RECT 7.31 0.428 7.378 0.652 ;
        RECT 6.878 0.428 6.946 0.652 ;
        RECT 6.23 0.428 6.298 0.652 ;
        RECT 6.014 0.428 6.082 0.652 ;
        RECT 5.474 0.428 5.542 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 4.394 0.428 4.462 0.652 ;
        RECT 4.178 0.518 4.246 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4725 0.25 0.5165 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.962 0.448 4.03 0.492 ;
        RECT 4.178 0.538 4.246 0.582 ;
        RECT 4.394 0.448 4.462 0.492 ;
        RECT 4.61 0.448 4.678 0.492 ;
        RECT 5.474 0.448 5.542 0.492 ;
        RECT 6.014 0.448 6.082 0.492 ;
        RECT 6.23 0.448 6.298 0.492 ;
        RECT 6.878 0.448 6.946 0.492 ;
        RECT 7.31 0.448 7.378 0.492 ;
        RECT 7.526 0.448 7.594 0.492 ;
        RECT 7.742 0.448 7.81 0.492 ;
        RECT 8.39 0.448 8.458 0.492 ;
        RECT 8.822 0.448 8.89 0.492 ;
        RECT 9.038 0.448 9.106 0.492 ;
        RECT 9.686 0.493 9.754 0.537 ;
        RECT 10.01 0.428 10.078 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 10.294 0.022 ;
        RECT 10.01 -0.022 10.078 0.202 ;
        RECT 9.686 -0.022 9.754 0.202 ;
        RECT 9.038 -0.022 9.106 0.202 ;
        RECT 8.822 -0.022 8.89 0.202 ;
        RECT 8.39 -0.022 8.458 0.202 ;
        RECT 7.742 -0.022 7.81 0.202 ;
        RECT 7.526 -0.022 7.594 0.202 ;
        RECT 7.31 -0.022 7.378 0.202 ;
        RECT 6.878 -0.022 6.946 0.202 ;
        RECT 6.23 -0.022 6.298 0.292 ;
        RECT 6.014 -0.022 6.082 0.292 ;
        RECT 5.474 -0.022 5.542 0.202 ;
        RECT 4.826 -0.022 4.894 0.202 ;
        RECT 4.61 -0.022 4.678 0.202 ;
        RECT 4.394 -0.022 4.462 0.202 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.422 -0.022 3.49 0.292 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.558 -0.022 2.626 0.292 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.074 0.158 0.27 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.558 0.1805 2.626 0.2245 ;
        RECT 2.774 0.1805 2.842 0.2245 ;
        RECT 3.422 0.1805 3.49 0.2245 ;
        RECT 3.962 0.138 4.03 0.182 ;
        RECT 4.178 0.138 4.246 0.182 ;
        RECT 4.394 0.138 4.462 0.182 ;
        RECT 4.61 0.138 4.678 0.182 ;
        RECT 4.826 0.138 4.894 0.182 ;
        RECT 5.474 0.138 5.542 0.182 ;
        RECT 6.014 0.203 6.082 0.247 ;
        RECT 6.23 0.203 6.298 0.247 ;
        RECT 6.878 0.138 6.946 0.182 ;
        RECT 7.31 0.138 7.378 0.182 ;
        RECT 7.526 0.138 7.594 0.182 ;
        RECT 7.742 0.138 7.81 0.182 ;
        RECT 8.39 0.138 8.458 0.182 ;
        RECT 8.822 0.113 8.89 0.157 ;
        RECT 9.038 0.113 9.106 0.157 ;
        RECT 9.686 0.138 9.754 0.182 ;
        RECT 10.01 0.138 10.078 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 2 0.518 2.752 0.562 ;
      RECT 2.108 0.428 9.34 0.472 ;
      RECT 1.244 0.068 9.556 0.112 ;
    LAYER m1 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.262 0.068 1.33 0.562 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 2.018 0.248 2.086 0.562 ;
      RECT 2.126 0.068 2.194 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.666 0.158 2.734 0.562 ;
      RECT 2.882 0.158 2.95 0.562 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.854 0.338 3.922 0.562 ;
      RECT 3.746 0.068 3.814 0.562 ;
      RECT 4.286 0.158 4.354 0.562 ;
      RECT 4.502 0.068 4.57 0.202 ;
      RECT 4.934 0.428 5.002 0.562 ;
      RECT 5.042 0.068 5.11 0.202 ;
      RECT 5.15 0.338 5.218 0.562 ;
      RECT 5.798 0.068 5.866 0.202 ;
      RECT 5.798 0.338 5.866 0.562 ;
      RECT 6.446 0.068 6.514 0.562 ;
      RECT 6.338 0.158 6.406 0.562 ;
      RECT 6.554 0.158 6.622 0.562 ;
      RECT 7.202 0.338 7.27 0.562 ;
      RECT 7.634 0.068 7.702 0.562 ;
      RECT 7.85 0.068 7.918 0.202 ;
      RECT 8.066 0.338 8.134 0.562 ;
      RECT 8.714 0.338 8.782 0.562 ;
      RECT 9.254 0.068 9.322 0.292 ;
      RECT 9.146 0.068 9.214 0.562 ;
      RECT 9.254 0.338 9.322 0.562 ;
      RECT 9.47 0.068 9.538 0.382 ;
      RECT 9.794 0.068 9.862 0.292 ;
    LAYER v1 ;
      RECT 9.474 0.068 9.534 0.112 ;
      RECT 9.258 0.428 9.318 0.472 ;
      RECT 7.854 0.068 7.914 0.112 ;
      RECT 6.45 0.428 6.51 0.472 ;
      RECT 5.802 0.068 5.862 0.112 ;
      RECT 5.046 0.068 5.106 0.112 ;
      RECT 4.938 0.428 4.998 0.472 ;
      RECT 4.506 0.068 4.566 0.112 ;
      RECT 3.75 0.068 3.81 0.112 ;
      RECT 2.994 0.428 3.054 0.472 ;
      RECT 2.67 0.518 2.73 0.562 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 2.022 0.518 2.082 0.562 ;
      RECT 1.266 0.068 1.326 0.112 ;
    LAYER v0 ;
      RECT 9.902 0.428 9.97 0.472 ;
      RECT 9.794 0.138 9.862 0.182 ;
      RECT 9.686 0.338 9.754 0.382 ;
      RECT 9.47 0.088 9.538 0.132 ;
      RECT 9.47 0.293 9.538 0.337 ;
      RECT 9.362 0.403 9.43 0.447 ;
      RECT 9.254 0.113 9.322 0.157 ;
      RECT 9.254 0.498 9.322 0.542 ;
      RECT 9.146 0.113 9.214 0.157 ;
      RECT 9.146 0.363 9.214 0.407 ;
      RECT 8.93 0.113 8.998 0.157 ;
      RECT 8.93 0.448 8.998 0.492 ;
      RECT 8.714 0.448 8.782 0.492 ;
      RECT 8.606 0.158 8.674 0.202 ;
      RECT 8.606 0.448 8.674 0.492 ;
      RECT 8.174 0.138 8.242 0.182 ;
      RECT 8.066 0.138 8.134 0.182 ;
      RECT 8.066 0.448 8.134 0.492 ;
      RECT 7.958 0.448 8.026 0.492 ;
      RECT 7.85 0.138 7.918 0.182 ;
      RECT 7.634 0.138 7.702 0.182 ;
      RECT 7.634 0.448 7.702 0.492 ;
      RECT 7.418 0.138 7.486 0.182 ;
      RECT 7.418 0.448 7.486 0.492 ;
      RECT 7.202 0.448 7.27 0.492 ;
      RECT 7.094 0.158 7.162 0.202 ;
      RECT 7.094 0.448 7.162 0.492 ;
      RECT 6.662 0.158 6.73 0.202 ;
      RECT 6.554 0.068 6.622 0.112 ;
      RECT 6.554 0.448 6.622 0.492 ;
      RECT 6.446 0.293 6.514 0.337 ;
      RECT 6.338 0.203 6.406 0.247 ;
      RECT 6.338 0.448 6.406 0.492 ;
      RECT 6.122 0.203 6.19 0.247 ;
      RECT 6.122 0.448 6.19 0.492 ;
      RECT 5.906 0.113 5.974 0.157 ;
      RECT 5.798 0.113 5.866 0.157 ;
      RECT 5.798 0.448 5.866 0.492 ;
      RECT 5.69 0.113 5.758 0.157 ;
      RECT 5.69 0.448 5.758 0.492 ;
      RECT 5.258 0.138 5.326 0.182 ;
      RECT 5.15 0.138 5.218 0.182 ;
      RECT 5.15 0.448 5.218 0.492 ;
      RECT 5.042 0.138 5.11 0.182 ;
      RECT 5.042 0.448 5.11 0.492 ;
      RECT 4.934 0.448 5.002 0.492 ;
      RECT 4.502 0.138 4.57 0.182 ;
      RECT 4.286 0.223 4.354 0.267 ;
      RECT 4.286 0.448 4.354 0.492 ;
      RECT 4.07 0.138 4.138 0.182 ;
      RECT 4.07 0.448 4.138 0.492 ;
      RECT 3.854 0.448 3.922 0.492 ;
      RECT 3.746 0.448 3.814 0.492 ;
      RECT 3.638 0.138 3.706 0.182 ;
      RECT 3.638 0.448 3.706 0.492 ;
      RECT 3.206 0.191 3.274 0.235 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.99 0.088 3.058 0.132 ;
      RECT 2.99 0.338 3.058 0.382 ;
      RECT 2.882 0.1805 2.95 0.2245 ;
      RECT 2.882 0.448 2.95 0.492 ;
      RECT 2.666 0.1805 2.734 0.2245 ;
      RECT 2.666 0.448 2.734 0.492 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.478 0.191 1.546 0.235 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.133 1.33 0.177 ;
      RECT 1.262 0.3155 1.33 0.3595 ;
      RECT 1.154 0.133 1.222 0.177 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 0.938 0.138 1.006 0.182 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.898 0.338 1.114 0.382 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.438 0.338 1.478 0.382 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.546 0.338 1.91 0.382 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 3.166 0.338 3.206 0.382 ;
      RECT 3.206 0.158 3.274 0.382 ;
      RECT 3.274 0.338 3.638 0.382 ;
      RECT 3.638 0.068 3.706 0.562 ;
      RECT 3.922 0.338 4.07 0.382 ;
      RECT 4.07 0.068 4.138 0.562 ;
      RECT 4.354 0.338 5.042 0.382 ;
      RECT 5.042 0.248 5.11 0.562 ;
      RECT 5.11 0.248 5.15 0.292 ;
      RECT 5.15 0.068 5.218 0.292 ;
      RECT 5.218 0.338 5.258 0.382 ;
      RECT 5.258 0.068 5.326 0.382 ;
      RECT 5.326 0.338 5.69 0.382 ;
      RECT 5.69 0.068 5.758 0.562 ;
      RECT 5.758 0.248 5.906 0.292 ;
      RECT 5.906 0.068 5.974 0.292 ;
      RECT 5.866 0.338 6.122 0.382 ;
      RECT 6.122 0.158 6.19 0.562 ;
      RECT 6.514 0.068 6.73 0.112 ;
      RECT 6.622 0.158 6.77 0.202 ;
      RECT 6.77 0.158 6.838 0.382 ;
      RECT 6.838 0.338 7.094 0.382 ;
      RECT 7.094 0.068 7.162 0.562 ;
      RECT 7.27 0.338 7.418 0.382 ;
      RECT 7.418 0.068 7.486 0.562 ;
      RECT 7.702 0.338 7.958 0.382 ;
      RECT 7.958 0.248 8.026 0.562 ;
      RECT 8.026 0.248 8.066 0.292 ;
      RECT 8.066 0.068 8.134 0.292 ;
      RECT 8.134 0.338 8.174 0.382 ;
      RECT 8.174 0.068 8.242 0.382 ;
      RECT 8.242 0.338 8.606 0.382 ;
      RECT 8.606 0.068 8.674 0.562 ;
      RECT 8.782 0.338 8.93 0.382 ;
      RECT 8.93 0.068 8.998 0.562 ;
      RECT 9.322 0.248 9.362 0.292 ;
      RECT 9.362 0.248 9.43 0.562 ;
      RECT 9.43 0.518 9.578 0.562 ;
      RECT 9.578 0.338 9.646 0.562 ;
      RECT 9.646 0.338 9.862 0.382 ;
      RECT 9.862 0.248 9.902 0.292 ;
      RECT 9.902 0.248 9.97 0.562 ;
  END
END b15fmm300hn1n04x5

MACRO b15fmm303hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fmm303hn1n04x5 0 0 ;
  SIZE 12.312 BY 0.63 ;
  SYMMETRY Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAGATEAREA 0.0765 LAYER m2 ;
      ANTENNAMAXAREACAR 1.946923 LAYER m1 ;
      ANTENNAMAXAREACAR 3.2488035 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4813675 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAGATEAREA 0.0963 LAYER m2 ;
      ANTENNAMAXAREACAR 1.67462975 LAYER m1 ;
      ANTENNAMAXAREACAR 2.67018525 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.3681045 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 10.766 0.428 10.834 0.562 ;
        RECT 6.662 0.428 6.73 0.562 ;
        RECT 4.07 0.428 4.138 0.562 ;
        RECT 3.314 0.338 3.382 0.562 ;
      LAYER m2 ;
        RECT 3.296 0.518 10.868 0.562 ;
      LAYER v1 ;
        RECT 3.318 0.518 3.378 0.562 ;
        RECT 4.074 0.518 4.134 0.562 ;
        RECT 6.666 0.518 6.726 0.562 ;
        RECT 10.77 0.518 10.83 0.562 ;
      LAYER v0 ;
        RECT 3.314 0.364 3.382 0.408 ;
        RECT 4.07 0.448 4.138 0.492 ;
        RECT 6.662 0.448 6.73 0.492 ;
        RECT 10.766 0.448 10.834 0.492 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.158 2.518 0.472 ;
      LAYER v0 ;
        RECT 2.45 0.293 2.518 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.31901225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 12.17 0.068 12.238 0.562 ;
      LAYER v0 ;
        RECT 12.17 0.428 12.238 0.472 ;
        RECT 12.17 0.152 12.238 0.196 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 8.93 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.97666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
        RECT 0.182 0.068 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 12.346 0.652 ;
        RECT 12.062 0.518 12.13 0.652 ;
        RECT 11.306 0.428 11.374 0.652 ;
        RECT 11.09 0.428 11.158 0.652 ;
        RECT 10.874 0.428 10.942 0.652 ;
        RECT 10.658 0.338 10.726 0.652 ;
        RECT 10.442 0.428 10.51 0.652 ;
        RECT 10.226 0.428 10.294 0.652 ;
        RECT 9.794 0.428 9.862 0.652 ;
        RECT 9.254 0.518 9.322 0.652 ;
        RECT 8.174 0.428 8.242 0.652 ;
        RECT 7.85 0.428 7.918 0.652 ;
        RECT 7.634 0.428 7.702 0.652 ;
        RECT 7.418 0.428 7.486 0.652 ;
        RECT 7.202 0.338 7.27 0.652 ;
        RECT 6.986 0.428 7.054 0.652 ;
        RECT 6.77 0.428 6.838 0.652 ;
        RECT 6.23 0.428 6.298 0.652 ;
        RECT 5.366 0.428 5.434 0.652 ;
        RECT 5.15 0.428 5.218 0.652 ;
        RECT 4.934 0.518 5.002 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 4.394 0.338 4.462 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.338 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4725 0.25 0.5165 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 4.178 0.448 4.246 0.492 ;
        RECT 4.394 0.448 4.462 0.492 ;
        RECT 4.61 0.448 4.678 0.492 ;
        RECT 4.934 0.538 5.002 0.582 ;
        RECT 5.15 0.448 5.218 0.492 ;
        RECT 5.366 0.448 5.434 0.492 ;
        RECT 6.23 0.448 6.298 0.492 ;
        RECT 6.77 0.448 6.838 0.492 ;
        RECT 6.986 0.448 7.054 0.492 ;
        RECT 7.202 0.448 7.27 0.492 ;
        RECT 7.418 0.448 7.486 0.492 ;
        RECT 7.634 0.448 7.702 0.492 ;
        RECT 7.85 0.448 7.918 0.492 ;
        RECT 8.174 0.448 8.242 0.492 ;
        RECT 9.254 0.538 9.322 0.582 ;
        RECT 9.794 0.448 9.862 0.492 ;
        RECT 10.226 0.448 10.294 0.492 ;
        RECT 10.442 0.448 10.51 0.492 ;
        RECT 10.658 0.448 10.726 0.492 ;
        RECT 10.874 0.448 10.942 0.492 ;
        RECT 11.09 0.448 11.158 0.492 ;
        RECT 11.306 0.448 11.374 0.492 ;
        RECT 12.064 0.538 12.128 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 12.346 0.022 ;
        RECT 12.062 -0.022 12.13 0.112 ;
        RECT 11.09 -0.022 11.158 0.112 ;
        RECT 10.658 -0.022 10.726 0.112 ;
        RECT 10.226 -0.022 10.294 0.112 ;
        RECT 9.794 -0.022 9.862 0.202 ;
        RECT 9.254 -0.022 9.322 0.202 ;
        RECT 8.066 -0.022 8.134 0.202 ;
        RECT 7.85 -0.022 7.918 0.202 ;
        RECT 7.634 -0.022 7.702 0.202 ;
        RECT 7.202 -0.022 7.27 0.202 ;
        RECT 6.77 -0.022 6.838 0.202 ;
        RECT 6.23 -0.022 6.298 0.202 ;
        RECT 5.69 -0.022 5.758 0.202 ;
        RECT 5.366 -0.022 5.434 0.202 ;
        RECT 5.15 -0.022 5.218 0.112 ;
        RECT 4.934 -0.022 5.002 0.112 ;
        RECT 4.718 -0.022 4.786 0.202 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.99 0.138 3.058 0.182 ;
        RECT 4.18 0.048 4.244 0.092 ;
        RECT 4.718 0.138 4.786 0.182 ;
        RECT 4.936 0.048 5 0.092 ;
        RECT 5.15 0.048 5.218 0.092 ;
        RECT 5.366 0.138 5.434 0.182 ;
        RECT 5.69 0.138 5.758 0.182 ;
        RECT 6.23 0.138 6.298 0.182 ;
        RECT 6.77 0.138 6.838 0.182 ;
        RECT 7.202 0.138 7.27 0.182 ;
        RECT 7.634 0.138 7.702 0.182 ;
        RECT 7.85 0.138 7.918 0.182 ;
        RECT 8.066 0.138 8.134 0.182 ;
        RECT 9.254 0.138 9.322 0.182 ;
        RECT 9.794 0.138 9.862 0.182 ;
        RECT 10.228 0.048 10.292 0.092 ;
        RECT 10.66 0.048 10.724 0.092 ;
        RECT 11.09 0.048 11.158 0.092 ;
        RECT 12.064 0.048 12.128 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.784 0.518 2.968 0.562 ;
      RECT 6.644 0.248 8.044 0.292 ;
      RECT 7.4 0.158 8.924 0.202 ;
      RECT 7.94 0.338 9.448 0.382 ;
      RECT 9.004 0.158 10.96 0.202 ;
      RECT 2.108 0.428 11.5 0.472 ;
      RECT 1.244 0.068 11.824 0.112 ;
      RECT 10.948 0.518 11.932 0.562 ;
      RECT 11.288 0.338 12.04 0.382 ;
      RECT 11.396 0.158 12.148 0.202 ;
    LAYER m1 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 1.262 0.428 1.586 0.472 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.126 0.068 2.194 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 3.314 0.338 3.382 0.562 ;
      RECT 3.422 0.338 3.49 0.562 ;
      RECT 3.746 0.158 3.814 0.562 ;
      RECT 4.07 0.428 4.138 0.562 ;
      RECT 4.07 0.068 4.138 0.202 ;
      RECT 3.422 0.158 3.638 0.202 ;
      RECT 5.042 0.068 5.11 0.562 ;
      RECT 4.826 0.068 4.894 0.562 ;
      RECT 5.258 0.068 5.326 0.202 ;
      RECT 5.69 0.428 5.758 0.562 ;
      RECT 5.798 0.068 5.866 0.202 ;
      RECT 5.906 0.338 5.974 0.562 ;
      RECT 6.554 0.068 6.622 0.202 ;
      RECT 6.662 0.428 6.73 0.562 ;
      RECT 6.554 0.338 6.622 0.562 ;
      RECT 7.31 0.248 7.378 0.562 ;
      RECT 8.066 0.338 8.134 0.562 ;
      RECT 7.742 0.068 7.81 0.562 ;
      RECT 7.958 0.338 8.026 0.472 ;
      RECT 7.958 0.068 8.026 0.292 ;
      RECT 8.282 0.068 8.498 0.112 ;
      RECT 8.39 0.248 8.458 0.472 ;
      RECT 8.606 0.248 8.674 0.562 ;
      RECT 8.714 0.338 8.782 0.562 ;
      RECT 8.822 0.428 8.89 0.562 ;
      RECT 9.038 0.428 9.47 0.472 ;
      RECT 8.93 0.068 8.998 0.562 ;
      RECT 9.038 0.068 9.106 0.202 ;
      RECT 9.038 0.338 9.43 0.382 ;
      RECT 9.362 0.518 9.686 0.562 ;
      RECT 9.47 0.068 9.538 0.202 ;
      RECT 9.578 0.158 9.646 0.472 ;
      RECT 9.902 0.248 9.97 0.472 ;
      RECT 10.01 0.068 10.078 0.202 ;
      RECT 10.422 0.248 10.55 0.292 ;
      RECT 10.854 0.068 10.982 0.112 ;
      RECT 10.766 0.428 10.834 0.562 ;
      RECT 10.874 0.158 10.942 0.382 ;
      RECT 11.198 0.158 11.266 0.562 ;
      RECT 11.306 0.248 11.374 0.382 ;
      RECT 11.414 0.338 11.482 0.562 ;
      RECT 11.522 0.428 11.59 0.562 ;
      RECT 11.306 0.068 11.59 0.112 ;
      RECT 11.63 0.068 11.698 0.202 ;
      RECT 11.738 0.068 11.806 0.292 ;
      RECT 11.954 0.068 12.022 0.562 ;
      RECT 12.062 0.158 12.13 0.472 ;
    LAYER v1 ;
      RECT 12.066 0.158 12.126 0.202 ;
      RECT 11.958 0.338 12.018 0.382 ;
      RECT 11.85 0.518 11.91 0.562 ;
      RECT 11.634 0.158 11.694 0.202 ;
      RECT 11.526 0.518 11.586 0.562 ;
      RECT 11.418 0.068 11.478 0.112 ;
      RECT 11.418 0.428 11.478 0.472 ;
      RECT 11.31 0.338 11.37 0.382 ;
      RECT 10.986 0.518 11.046 0.562 ;
      RECT 10.878 0.158 10.938 0.202 ;
      RECT 10.554 0.158 10.614 0.202 ;
      RECT 10.014 0.158 10.074 0.202 ;
      RECT 9.69 0.428 9.75 0.472 ;
      RECT 9.582 0.158 9.642 0.202 ;
      RECT 9.474 0.068 9.534 0.112 ;
      RECT 9.258 0.338 9.318 0.382 ;
      RECT 9.042 0.158 9.102 0.202 ;
      RECT 8.934 0.068 8.994 0.112 ;
      RECT 8.826 0.428 8.886 0.472 ;
      RECT 8.718 0.158 8.778 0.202 ;
      RECT 8.718 0.338 8.778 0.382 ;
      RECT 8.502 0.338 8.562 0.382 ;
      RECT 8.394 0.428 8.454 0.472 ;
      RECT 7.962 0.248 8.022 0.292 ;
      RECT 7.962 0.338 8.022 0.382 ;
      RECT 7.422 0.158 7.482 0.202 ;
      RECT 6.666 0.248 6.726 0.292 ;
      RECT 6.558 0.068 6.618 0.112 ;
      RECT 5.802 0.068 5.862 0.112 ;
      RECT 5.694 0.428 5.754 0.472 ;
      RECT 5.262 0.068 5.322 0.112 ;
      RECT 4.074 0.068 4.134 0.112 ;
      RECT 3.426 0.428 3.486 0.472 ;
      RECT 2.886 0.518 2.946 0.562 ;
      RECT 2.67 0.518 2.73 0.562 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.266 0.068 1.326 0.112 ;
    LAYER v0 ;
      RECT 12.062 0.338 12.13 0.382 ;
      RECT 11.954 0.158 12.022 0.202 ;
      RECT 11.954 0.454 12.022 0.498 ;
      RECT 11.738 0.114 11.806 0.158 ;
      RECT 11.74 0.408 11.804 0.452 ;
      RECT 11.63 0.114 11.698 0.158 ;
      RECT 11.522 0.248 11.59 0.292 ;
      RECT 11.522 0.448 11.59 0.492 ;
      RECT 11.414 0.068 11.482 0.112 ;
      RECT 11.414 0.448 11.482 0.492 ;
      RECT 11.306 0.158 11.374 0.202 ;
      RECT 11.306 0.293 11.374 0.337 ;
      RECT 11.198 0.448 11.266 0.492 ;
      RECT 10.982 0.448 11.05 0.492 ;
      RECT 10.874 0.068 10.942 0.112 ;
      RECT 10.874 0.2705 10.942 0.3145 ;
      RECT 10.55 0.448 10.618 0.492 ;
      RECT 10.442 0.248 10.51 0.292 ;
      RECT 10.444 0.088 10.508 0.132 ;
      RECT 10.334 0.338 10.402 0.382 ;
      RECT 10.01 0.138 10.078 0.182 ;
      RECT 9.902 0.293 9.97 0.337 ;
      RECT 9.578 0.248 9.646 0.292 ;
      RECT 9.47 0.113 9.538 0.157 ;
      RECT 9.47 0.518 9.538 0.562 ;
      RECT 9.362 0.248 9.43 0.292 ;
      RECT 9.362 0.428 9.43 0.472 ;
      RECT 9.254 0.338 9.322 0.382 ;
      RECT 9.146 0.248 9.214 0.292 ;
      RECT 9.146 0.428 9.214 0.472 ;
      RECT 9.038 0.138 9.106 0.182 ;
      RECT 8.93 0.448 8.998 0.492 ;
      RECT 8.822 0.09 8.89 0.134 ;
      RECT 8.822 0.448 8.89 0.492 ;
      RECT 8.714 0.09 8.782 0.134 ;
      RECT 8.714 0.448 8.782 0.492 ;
      RECT 8.606 0.448 8.674 0.492 ;
      RECT 8.498 0.448 8.566 0.492 ;
      RECT 8.39 0.068 8.458 0.112 ;
      RECT 8.39 0.293 8.458 0.337 ;
      RECT 8.282 0.1805 8.35 0.2245 ;
      RECT 8.282 0.448 8.35 0.492 ;
      RECT 8.066 0.448 8.134 0.492 ;
      RECT 7.958 0.138 8.026 0.182 ;
      RECT 7.958 0.358 8.026 0.402 ;
      RECT 7.742 0.138 7.81 0.182 ;
      RECT 7.742 0.448 7.81 0.492 ;
      RECT 7.526 0.448 7.594 0.492 ;
      RECT 7.418 0.138 7.486 0.182 ;
      RECT 7.31 0.448 7.378 0.492 ;
      RECT 7.094 0.448 7.162 0.492 ;
      RECT 6.986 0.158 7.054 0.202 ;
      RECT 6.878 0.448 6.946 0.492 ;
      RECT 6.662 0.138 6.73 0.182 ;
      RECT 6.554 0.138 6.622 0.182 ;
      RECT 6.554 0.448 6.622 0.492 ;
      RECT 6.446 0.138 6.514 0.182 ;
      RECT 6.446 0.448 6.514 0.492 ;
      RECT 6.014 0.138 6.082 0.182 ;
      RECT 5.906 0.138 5.974 0.182 ;
      RECT 5.906 0.448 5.974 0.492 ;
      RECT 5.798 0.138 5.866 0.182 ;
      RECT 5.798 0.448 5.866 0.492 ;
      RECT 5.69 0.448 5.758 0.492 ;
      RECT 5.258 0.138 5.326 0.182 ;
      RECT 5.042 0.448 5.11 0.492 ;
      RECT 5.044 0.168 5.108 0.212 ;
      RECT 4.826 0.138 4.894 0.182 ;
      RECT 4.826 0.428 4.894 0.472 ;
      RECT 4.61 0.293 4.678 0.337 ;
      RECT 4.502 0.448 4.57 0.492 ;
      RECT 4.394 0.248 4.462 0.292 ;
      RECT 4.286 0.448 4.354 0.492 ;
      RECT 4.07 0.138 4.138 0.182 ;
      RECT 3.854 0.178 3.922 0.222 ;
      RECT 3.854 0.408 3.922 0.452 ;
      RECT 3.746 0.178 3.814 0.222 ;
      RECT 3.746 0.408 3.814 0.452 ;
      RECT 3.638 0.408 3.706 0.452 ;
      RECT 3.53 0.158 3.598 0.202 ;
      RECT 3.53 0.493 3.598 0.537 ;
      RECT 3.422 0.493 3.49 0.537 ;
      RECT 3.206 0.178 3.274 0.222 ;
      RECT 3.098 0.448 3.166 0.492 ;
      RECT 2.882 0.448 2.95 0.492 ;
      RECT 2.774 0.178 2.842 0.222 ;
      RECT 2.666 0.448 2.734 0.492 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.088 1.33 0.132 ;
      RECT 1.262 0.3155 1.33 0.3595 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.94 0.178 1.004 0.222 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.4725 0.574 0.5165 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.898 0.338 1.114 0.382 ;
      RECT 0.83 0.428 1.154 0.472 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 1.222 0.518 1.438 0.562 ;
      RECT 1.87 0.428 1.91 0.472 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 1.37 0.158 1.586 0.202 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.158 1.87 0.382 ;
      RECT 1.87 0.158 2.086 0.202 ;
      RECT 2.734 0.338 2.774 0.382 ;
      RECT 2.774 0.158 2.842 0.382 ;
      RECT 2.842 0.338 2.882 0.382 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 3.166 0.338 3.206 0.382 ;
      RECT 3.206 0.158 3.274 0.382 ;
      RECT 3.274 0.248 3.53 0.292 ;
      RECT 3.53 0.248 3.598 0.562 ;
      RECT 3.814 0.518 3.962 0.562 ;
      RECT 3.962 0.338 4.03 0.562 ;
      RECT 4.03 0.338 4.286 0.382 ;
      RECT 4.286 0.248 4.354 0.562 ;
      RECT 4.354 0.248 4.502 0.292 ;
      RECT 4.502 0.248 4.57 0.562 ;
      RECT 3.638 0.068 3.706 0.562 ;
      RECT 3.706 0.068 3.854 0.112 ;
      RECT 3.854 0.068 3.922 0.472 ;
      RECT 3.922 0.248 4.178 0.292 ;
      RECT 4.178 0.158 4.246 0.292 ;
      RECT 4.246 0.158 4.61 0.202 ;
      RECT 4.61 0.158 4.678 0.382 ;
      RECT 5.11 0.248 5.798 0.292 ;
      RECT 5.798 0.248 5.866 0.562 ;
      RECT 5.866 0.248 5.906 0.292 ;
      RECT 5.906 0.068 5.974 0.292 ;
      RECT 5.974 0.338 6.014 0.382 ;
      RECT 6.014 0.068 6.082 0.382 ;
      RECT 6.082 0.338 6.446 0.382 ;
      RECT 6.446 0.068 6.514 0.562 ;
      RECT 6.514 0.248 6.662 0.292 ;
      RECT 6.662 0.068 6.73 0.292 ;
      RECT 6.622 0.338 6.878 0.382 ;
      RECT 6.878 0.158 6.946 0.562 ;
      RECT 6.946 0.158 7.094 0.202 ;
      RECT 7.094 0.158 7.162 0.562 ;
      RECT 7.378 0.248 7.418 0.292 ;
      RECT 7.418 0.068 7.486 0.292 ;
      RECT 7.486 0.248 7.526 0.292 ;
      RECT 7.526 0.248 7.594 0.562 ;
      RECT 8.134 0.338 8.282 0.382 ;
      RECT 8.282 0.158 8.35 0.562 ;
      RECT 8.498 0.068 8.566 0.562 ;
      RECT 8.674 0.248 8.714 0.292 ;
      RECT 8.714 0.068 8.782 0.292 ;
      RECT 8.782 0.338 8.822 0.382 ;
      RECT 8.822 0.068 8.89 0.382 ;
      RECT 9.038 0.248 9.47 0.292 ;
      RECT 9.47 0.248 9.538 0.472 ;
      RECT 9.686 0.428 9.754 0.562 ;
      RECT 9.97 0.428 10.118 0.472 ;
      RECT 10.118 0.158 10.186 0.472 ;
      RECT 10.186 0.158 10.442 0.202 ;
      RECT 10.442 0.068 10.51 0.202 ;
      RECT 10.186 0.338 10.55 0.382 ;
      RECT 10.55 0.338 10.618 0.562 ;
      RECT 10.55 0.158 10.618 0.292 ;
      RECT 10.982 0.068 11.05 0.562 ;
      RECT 11.266 0.158 11.414 0.202 ;
      RECT 11.414 0.158 11.482 0.292 ;
      RECT 11.482 0.248 11.63 0.292 ;
      RECT 11.63 0.248 11.698 0.382 ;
      RECT 11.698 0.338 11.738 0.382 ;
      RECT 11.738 0.338 11.806 0.472 ;
      RECT 11.806 0.248 11.846 0.292 ;
      RECT 11.846 0.248 11.914 0.562 ;
  END
END b15fmm303hn1n04x5

MACRO b15fmm30chn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fmm30chn1n04x5 0 0 ;
  SIZE 12.636 BY 0.63 ;
  SYMMETRY Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0819 LAYER m2 ;
      ANTENNAMAXAREACAR 2.185 LAYER m1 ;
      ANTENNAMAXAREACAR 4.3005555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0882 LAYER m2 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
      ANTENNAMAXAREACAR 5.734074 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 10.766 0.428 10.834 0.562 ;
        RECT 7.958 0.338 8.026 0.562 ;
        RECT 6.662 0.428 6.73 0.562 ;
        RECT 4.61 0.338 4.678 0.562 ;
        RECT 3.962 0.428 4.03 0.562 ;
        RECT 3.206 0.338 3.274 0.562 ;
      LAYER m2 ;
        RECT 3.188 0.518 10.868 0.562 ;
      LAYER v1 ;
        RECT 3.21 0.518 3.27 0.562 ;
        RECT 3.966 0.518 4.026 0.562 ;
        RECT 4.614 0.518 4.674 0.562 ;
        RECT 6.666 0.518 6.726 0.562 ;
        RECT 7.962 0.518 8.022 0.562 ;
        RECT 10.77 0.518 10.83 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.364 3.274 0.408 ;
        RECT 3.962 0.448 4.03 0.492 ;
        RECT 4.61 0.448 4.678 0.492 ;
        RECT 6.662 0.448 6.73 0.492 ;
        RECT 7.958 0.448 8.026 0.492 ;
        RECT 10.766 0.448 10.834 0.492 ;
    END
  END psb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.856508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 12.494 0.068 12.562 0.562 ;
      LAYER v0 ;
        RECT 12.494 0.493 12.562 0.537 ;
        RECT 12.494 0.093 12.562 0.137 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 12.35 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 2.7444445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
        RECT 0.182 0.068 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 12.67 0.652 ;
        RECT 12.386 0.428 12.454 0.652 ;
        RECT 12.062 0.518 12.13 0.652 ;
        RECT 11.306 0.428 11.374 0.652 ;
        RECT 11.09 0.428 11.158 0.652 ;
        RECT 10.874 0.428 10.942 0.652 ;
        RECT 10.658 0.338 10.726 0.652 ;
        RECT 10.442 0.428 10.51 0.652 ;
        RECT 10.226 0.428 10.294 0.652 ;
        RECT 9.794 0.428 9.862 0.652 ;
        RECT 9.254 0.518 9.322 0.652 ;
        RECT 8.174 0.428 8.242 0.652 ;
        RECT 7.85 0.428 7.918 0.652 ;
        RECT 7.634 0.428 7.702 0.652 ;
        RECT 7.418 0.428 7.486 0.652 ;
        RECT 7.202 0.338 7.27 0.652 ;
        RECT 6.986 0.428 7.054 0.652 ;
        RECT 6.77 0.428 6.838 0.652 ;
        RECT 6.23 0.428 6.298 0.652 ;
        RECT 5.366 0.428 5.434 0.652 ;
        RECT 5.15 0.428 5.218 0.652 ;
        RECT 4.934 0.518 5.002 0.652 ;
        RECT 4.718 0.338 4.786 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 4.286 0.338 4.354 0.652 ;
        RECT 4.07 0.428 4.138 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4725 0.25 0.5165 ;
        RECT 0.83 0.4055 0.898 0.4495 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 4.07 0.448 4.138 0.492 ;
        RECT 4.286 0.448 4.354 0.492 ;
        RECT 4.502 0.448 4.57 0.492 ;
        RECT 4.718 0.448 4.786 0.492 ;
        RECT 4.934 0.538 5.002 0.582 ;
        RECT 5.15 0.448 5.218 0.492 ;
        RECT 5.366 0.448 5.434 0.492 ;
        RECT 6.23 0.448 6.298 0.492 ;
        RECT 6.77 0.448 6.838 0.492 ;
        RECT 6.986 0.448 7.054 0.492 ;
        RECT 7.202 0.448 7.27 0.492 ;
        RECT 7.418 0.448 7.486 0.492 ;
        RECT 7.634 0.448 7.702 0.492 ;
        RECT 7.85 0.448 7.918 0.492 ;
        RECT 8.174 0.448 8.242 0.492 ;
        RECT 9.254 0.538 9.322 0.582 ;
        RECT 9.794 0.448 9.862 0.492 ;
        RECT 10.226 0.448 10.294 0.492 ;
        RECT 10.442 0.448 10.51 0.492 ;
        RECT 10.658 0.448 10.726 0.492 ;
        RECT 10.874 0.448 10.942 0.492 ;
        RECT 11.09 0.448 11.158 0.492 ;
        RECT 11.306 0.448 11.374 0.492 ;
        RECT 12.062 0.538 12.13 0.582 ;
        RECT 12.386 0.493 12.454 0.537 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 12.67 0.022 ;
        RECT 12.386 -0.022 12.454 0.202 ;
        RECT 12.062 -0.022 12.13 0.112 ;
        RECT 11.09 -0.022 11.158 0.112 ;
        RECT 10.658 -0.022 10.726 0.112 ;
        RECT 10.226 -0.022 10.294 0.112 ;
        RECT 9.794 -0.022 9.862 0.202 ;
        RECT 9.254 -0.022 9.322 0.202 ;
        RECT 8.066 -0.022 8.134 0.202 ;
        RECT 7.85 -0.022 7.918 0.202 ;
        RECT 7.634 -0.022 7.702 0.202 ;
        RECT 7.202 -0.022 7.27 0.202 ;
        RECT 6.77 -0.022 6.838 0.202 ;
        RECT 6.23 -0.022 6.298 0.202 ;
        RECT 5.69 -0.022 5.758 0.202 ;
        RECT 5.366 -0.022 5.434 0.202 ;
        RECT 5.15 -0.022 5.218 0.112 ;
        RECT 4.934 -0.022 5.002 0.112 ;
        RECT 4.718 -0.022 4.786 0.202 ;
        RECT 4.07 -0.022 4.138 0.112 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.074 0.158 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.832 0.138 0.896 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 4.072 0.048 4.136 0.092 ;
        RECT 4.718 0.138 4.786 0.182 ;
        RECT 4.936 0.048 5 0.092 ;
        RECT 5.15 0.048 5.218 0.092 ;
        RECT 5.366 0.138 5.434 0.182 ;
        RECT 5.69 0.138 5.758 0.182 ;
        RECT 6.23 0.138 6.298 0.182 ;
        RECT 6.77 0.138 6.838 0.182 ;
        RECT 7.202 0.138 7.27 0.182 ;
        RECT 7.634 0.138 7.702 0.182 ;
        RECT 7.85 0.138 7.918 0.182 ;
        RECT 8.066 0.138 8.134 0.182 ;
        RECT 9.254 0.138 9.322 0.182 ;
        RECT 9.794 0.138 9.862 0.182 ;
        RECT 10.228 0.048 10.292 0.092 ;
        RECT 10.66 0.048 10.724 0.092 ;
        RECT 11.09 0.048 11.158 0.092 ;
        RECT 12.062 0.048 12.13 0.092 ;
        RECT 12.386 0.093 12.454 0.137 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.676 0.518 2.86 0.562 ;
      RECT 6.644 0.248 8.044 0.292 ;
      RECT 7.4 0.158 8.924 0.202 ;
      RECT 7.832 0.338 9.448 0.382 ;
      RECT 9.004 0.158 10.96 0.202 ;
      RECT 2 0.428 11.5 0.472 ;
      RECT 1.136 0.068 11.5 0.112 ;
      RECT 10.948 0.518 11.932 0.562 ;
      RECT 11.288 0.338 12.04 0.382 ;
      RECT 11.396 0.158 12.148 0.202 ;
    LAYER m1 ;
      RECT 1.694 0.428 1.762 0.562 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.154 0.428 1.478 0.472 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 2.018 0.068 2.086 0.562 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.99 0.338 3.058 0.562 ;
      RECT 3.206 0.338 3.274 0.562 ;
      RECT 3.314 0.338 3.382 0.562 ;
      RECT 3.638 0.158 3.706 0.562 ;
      RECT 3.962 0.428 4.03 0.562 ;
      RECT 3.962 0.068 4.03 0.202 ;
      RECT 3.314 0.158 3.53 0.202 ;
      RECT 5.042 0.068 5.11 0.562 ;
      RECT 4.61 0.338 4.678 0.562 ;
      RECT 4.826 0.068 4.894 0.562 ;
      RECT 5.258 0.068 5.326 0.202 ;
      RECT 5.69 0.428 5.758 0.562 ;
      RECT 5.798 0.068 5.866 0.202 ;
      RECT 5.906 0.338 5.974 0.562 ;
      RECT 6.554 0.068 6.622 0.202 ;
      RECT 6.662 0.428 6.73 0.562 ;
      RECT 6.554 0.338 6.622 0.562 ;
      RECT 7.31 0.248 7.378 0.562 ;
      RECT 8.066 0.338 8.134 0.562 ;
      RECT 7.742 0.068 7.81 0.562 ;
      RECT 7.85 0.248 7.918 0.382 ;
      RECT 7.958 0.338 8.026 0.562 ;
      RECT 7.958 0.068 8.026 0.292 ;
      RECT 8.282 0.068 8.498 0.112 ;
      RECT 8.39 0.248 8.458 0.472 ;
      RECT 8.606 0.248 8.674 0.562 ;
      RECT 8.714 0.338 8.782 0.562 ;
      RECT 8.822 0.428 8.89 0.562 ;
      RECT 9.038 0.428 9.47 0.472 ;
      RECT 8.93 0.068 8.998 0.562 ;
      RECT 9.038 0.068 9.106 0.202 ;
      RECT 9.038 0.338 9.43 0.382 ;
      RECT 9.362 0.518 9.686 0.562 ;
      RECT 9.47 0.068 9.538 0.202 ;
      RECT 9.578 0.158 9.646 0.472 ;
      RECT 9.902 0.248 9.97 0.472 ;
      RECT 10.01 0.068 10.078 0.202 ;
      RECT 10.422 0.248 10.55 0.292 ;
      RECT 10.854 0.068 10.982 0.112 ;
      RECT 10.766 0.428 10.834 0.562 ;
      RECT 10.874 0.158 10.942 0.382 ;
      RECT 11.198 0.158 11.266 0.562 ;
      RECT 11.306 0.248 11.374 0.382 ;
      RECT 11.414 0.338 11.482 0.562 ;
      RECT 11.522 0.428 11.59 0.562 ;
      RECT 11.306 0.068 11.59 0.112 ;
      RECT 11.63 0.068 11.698 0.202 ;
      RECT 11.738 0.068 11.806 0.292 ;
      RECT 11.954 0.068 12.022 0.562 ;
      RECT 12.062 0.158 12.13 0.472 ;
      RECT 12.17 0.068 12.238 0.562 ;
    LAYER v1 ;
      RECT 12.066 0.158 12.126 0.202 ;
      RECT 11.958 0.338 12.018 0.382 ;
      RECT 11.85 0.518 11.91 0.562 ;
      RECT 11.634 0.158 11.694 0.202 ;
      RECT 11.526 0.518 11.586 0.562 ;
      RECT 11.418 0.068 11.478 0.112 ;
      RECT 11.418 0.428 11.478 0.472 ;
      RECT 11.31 0.338 11.37 0.382 ;
      RECT 10.986 0.518 11.046 0.562 ;
      RECT 10.878 0.158 10.938 0.202 ;
      RECT 10.554 0.158 10.614 0.202 ;
      RECT 10.014 0.158 10.074 0.202 ;
      RECT 9.69 0.428 9.75 0.472 ;
      RECT 9.582 0.158 9.642 0.202 ;
      RECT 9.474 0.068 9.534 0.112 ;
      RECT 9.258 0.338 9.318 0.382 ;
      RECT 9.042 0.158 9.102 0.202 ;
      RECT 8.934 0.068 8.994 0.112 ;
      RECT 8.826 0.338 8.886 0.382 ;
      RECT 8.826 0.428 8.886 0.472 ;
      RECT 8.718 0.158 8.778 0.202 ;
      RECT 8.502 0.338 8.562 0.382 ;
      RECT 8.394 0.428 8.454 0.472 ;
      RECT 7.962 0.248 8.022 0.292 ;
      RECT 7.854 0.338 7.914 0.382 ;
      RECT 7.422 0.158 7.482 0.202 ;
      RECT 6.666 0.248 6.726 0.292 ;
      RECT 6.558 0.068 6.618 0.112 ;
      RECT 5.802 0.068 5.862 0.112 ;
      RECT 5.694 0.428 5.754 0.472 ;
      RECT 5.262 0.068 5.322 0.112 ;
      RECT 3.966 0.068 4.026 0.112 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 2.778 0.518 2.838 0.562 ;
      RECT 2.562 0.518 2.622 0.562 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.698 0.518 1.758 0.562 ;
      RECT 1.158 0.068 1.218 0.112 ;
    LAYER v0 ;
      RECT 12.17 0.158 12.238 0.202 ;
      RECT 12.17 0.454 12.238 0.498 ;
      RECT 12.062 0.338 12.13 0.382 ;
      RECT 11.954 0.158 12.022 0.202 ;
      RECT 11.954 0.454 12.022 0.498 ;
      RECT 11.738 0.114 11.806 0.158 ;
      RECT 11.74 0.408 11.804 0.452 ;
      RECT 11.63 0.114 11.698 0.158 ;
      RECT 11.522 0.248 11.59 0.292 ;
      RECT 11.522 0.448 11.59 0.492 ;
      RECT 11.414 0.068 11.482 0.112 ;
      RECT 11.414 0.448 11.482 0.492 ;
      RECT 11.306 0.158 11.374 0.202 ;
      RECT 11.306 0.293 11.374 0.337 ;
      RECT 11.198 0.448 11.266 0.492 ;
      RECT 10.982 0.448 11.05 0.492 ;
      RECT 10.874 0.068 10.942 0.112 ;
      RECT 10.874 0.2705 10.942 0.3145 ;
      RECT 10.55 0.448 10.618 0.492 ;
      RECT 10.442 0.248 10.51 0.292 ;
      RECT 10.444 0.088 10.508 0.132 ;
      RECT 10.334 0.338 10.402 0.382 ;
      RECT 10.01 0.138 10.078 0.182 ;
      RECT 9.902 0.293 9.97 0.337 ;
      RECT 9.578 0.248 9.646 0.292 ;
      RECT 9.47 0.113 9.538 0.157 ;
      RECT 9.47 0.518 9.538 0.562 ;
      RECT 9.362 0.248 9.43 0.292 ;
      RECT 9.362 0.428 9.43 0.472 ;
      RECT 9.254 0.338 9.322 0.382 ;
      RECT 9.146 0.248 9.214 0.292 ;
      RECT 9.146 0.428 9.214 0.472 ;
      RECT 9.038 0.138 9.106 0.182 ;
      RECT 8.93 0.448 8.998 0.492 ;
      RECT 8.822 0.09 8.89 0.134 ;
      RECT 8.822 0.448 8.89 0.492 ;
      RECT 8.714 0.09 8.782 0.134 ;
      RECT 8.714 0.448 8.782 0.492 ;
      RECT 8.606 0.448 8.674 0.492 ;
      RECT 8.498 0.448 8.566 0.492 ;
      RECT 8.39 0.068 8.458 0.112 ;
      RECT 8.39 0.293 8.458 0.337 ;
      RECT 8.282 0.1805 8.35 0.2245 ;
      RECT 8.282 0.448 8.35 0.492 ;
      RECT 8.066 0.448 8.134 0.492 ;
      RECT 7.958 0.138 8.026 0.182 ;
      RECT 7.85 0.293 7.918 0.337 ;
      RECT 7.742 0.138 7.81 0.182 ;
      RECT 7.742 0.448 7.81 0.492 ;
      RECT 7.526 0.448 7.594 0.492 ;
      RECT 7.418 0.138 7.486 0.182 ;
      RECT 7.31 0.448 7.378 0.492 ;
      RECT 7.094 0.448 7.162 0.492 ;
      RECT 6.986 0.158 7.054 0.202 ;
      RECT 6.878 0.448 6.946 0.492 ;
      RECT 6.662 0.138 6.73 0.182 ;
      RECT 6.554 0.138 6.622 0.182 ;
      RECT 6.554 0.448 6.622 0.492 ;
      RECT 6.446 0.138 6.514 0.182 ;
      RECT 6.446 0.448 6.514 0.492 ;
      RECT 6.014 0.138 6.082 0.182 ;
      RECT 5.906 0.138 5.974 0.182 ;
      RECT 5.906 0.448 5.974 0.492 ;
      RECT 5.798 0.138 5.866 0.182 ;
      RECT 5.798 0.448 5.866 0.492 ;
      RECT 5.69 0.448 5.758 0.492 ;
      RECT 5.258 0.138 5.326 0.182 ;
      RECT 5.042 0.448 5.11 0.492 ;
      RECT 5.044 0.168 5.108 0.212 ;
      RECT 4.826 0.138 4.894 0.182 ;
      RECT 4.826 0.448 4.894 0.492 ;
      RECT 4.502 0.293 4.57 0.337 ;
      RECT 4.394 0.448 4.462 0.492 ;
      RECT 4.286 0.248 4.354 0.292 ;
      RECT 4.178 0.448 4.246 0.492 ;
      RECT 3.962 0.138 4.03 0.182 ;
      RECT 3.746 0.178 3.814 0.222 ;
      RECT 3.746 0.408 3.814 0.452 ;
      RECT 3.638 0.178 3.706 0.222 ;
      RECT 3.638 0.408 3.706 0.452 ;
      RECT 3.53 0.408 3.598 0.452 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.422 0.493 3.49 0.537 ;
      RECT 3.314 0.493 3.382 0.537 ;
      RECT 3.098 0.178 3.166 0.222 ;
      RECT 2.99 0.448 3.058 0.492 ;
      RECT 2.774 0.448 2.842 0.492 ;
      RECT 2.666 0.178 2.734 0.222 ;
      RECT 2.558 0.448 2.626 0.492 ;
      RECT 2.234 0.138 2.302 0.182 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.138 2.086 0.182 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.154 0.3155 1.222 0.3595 ;
      RECT 1.046 0.4505 1.114 0.4945 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.4505 0.574 0.4945 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.292 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.762 0.428 1.802 0.472 ;
      RECT 1.802 0.248 1.87 0.472 ;
      RECT 1.262 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.546 0.338 1.694 0.382 ;
      RECT 1.694 0.158 1.762 0.382 ;
      RECT 1.762 0.158 1.978 0.202 ;
      RECT 2.626 0.338 2.666 0.382 ;
      RECT 2.666 0.158 2.734 0.382 ;
      RECT 2.734 0.338 2.774 0.382 ;
      RECT 2.774 0.338 2.842 0.562 ;
      RECT 3.058 0.338 3.098 0.382 ;
      RECT 3.098 0.158 3.166 0.382 ;
      RECT 3.166 0.248 3.422 0.292 ;
      RECT 3.422 0.248 3.49 0.562 ;
      RECT 3.706 0.518 3.854 0.562 ;
      RECT 3.854 0.338 3.922 0.562 ;
      RECT 3.922 0.338 4.178 0.382 ;
      RECT 4.178 0.248 4.246 0.562 ;
      RECT 4.246 0.248 4.394 0.292 ;
      RECT 4.394 0.248 4.462 0.562 ;
      RECT 3.53 0.068 3.598 0.562 ;
      RECT 3.598 0.068 3.746 0.112 ;
      RECT 3.746 0.068 3.814 0.472 ;
      RECT 3.814 0.248 4.07 0.292 ;
      RECT 4.07 0.158 4.138 0.292 ;
      RECT 4.138 0.158 4.502 0.202 ;
      RECT 4.502 0.158 4.57 0.382 ;
      RECT 5.11 0.248 5.798 0.292 ;
      RECT 5.798 0.248 5.866 0.562 ;
      RECT 5.866 0.248 5.906 0.292 ;
      RECT 5.906 0.068 5.974 0.292 ;
      RECT 5.974 0.338 6.014 0.382 ;
      RECT 6.014 0.068 6.082 0.382 ;
      RECT 6.082 0.338 6.446 0.382 ;
      RECT 6.446 0.068 6.514 0.562 ;
      RECT 6.514 0.248 6.662 0.292 ;
      RECT 6.662 0.068 6.73 0.292 ;
      RECT 6.622 0.338 6.878 0.382 ;
      RECT 6.878 0.158 6.946 0.562 ;
      RECT 6.946 0.158 7.094 0.202 ;
      RECT 7.094 0.158 7.162 0.562 ;
      RECT 7.378 0.248 7.418 0.292 ;
      RECT 7.418 0.068 7.486 0.292 ;
      RECT 7.486 0.248 7.526 0.292 ;
      RECT 7.526 0.248 7.594 0.562 ;
      RECT 8.134 0.338 8.282 0.382 ;
      RECT 8.282 0.158 8.35 0.562 ;
      RECT 8.498 0.068 8.566 0.562 ;
      RECT 8.674 0.248 8.714 0.292 ;
      RECT 8.714 0.068 8.782 0.292 ;
      RECT 8.782 0.338 8.822 0.382 ;
      RECT 8.822 0.068 8.89 0.382 ;
      RECT 9.038 0.248 9.47 0.292 ;
      RECT 9.47 0.248 9.538 0.472 ;
      RECT 9.686 0.428 9.754 0.562 ;
      RECT 9.97 0.428 10.118 0.472 ;
      RECT 10.118 0.158 10.186 0.472 ;
      RECT 10.186 0.158 10.442 0.202 ;
      RECT 10.442 0.068 10.51 0.202 ;
      RECT 10.186 0.338 10.55 0.382 ;
      RECT 10.55 0.338 10.618 0.562 ;
      RECT 10.55 0.158 10.618 0.292 ;
      RECT 10.982 0.068 11.05 0.562 ;
      RECT 11.266 0.158 11.414 0.202 ;
      RECT 11.414 0.158 11.482 0.292 ;
      RECT 11.482 0.248 11.63 0.292 ;
      RECT 11.63 0.248 11.698 0.382 ;
      RECT 11.698 0.338 11.738 0.382 ;
      RECT 11.738 0.338 11.806 0.472 ;
      RECT 11.806 0.248 11.846 0.292 ;
      RECT 11.846 0.248 11.914 0.562 ;
  END
END b15fmm30chn1n04x5

MACRO b15fpn000hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn000hn1n02x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.158 1.762 0.472 ;
      LAYER v0 ;
        RECT 1.694 0.338 1.762 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.018 0.178 2.086 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.91 0.178 1.978 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.338 1.672 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.182 0.158 0.25 0.382 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.722 0.248 0.79 0.382 ;
      RECT 1.046 0.518 1.262 0.562 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.37 0.248 1.438 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.158 1.87 0.562 ;
    LAYER v1 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.2705 1.438 0.3145 ;
      RECT 1.262 0.1535 1.33 0.1975 ;
      RECT 1.154 0.3155 1.222 0.3595 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.83 0.3155 0.898 0.3595 ;
      RECT 0.722 0.3155 0.79 0.3595 ;
      RECT 0.614 0.1575 0.682 0.2015 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.248 0.25 0.292 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 1.262 0.068 1.33 0.562 ;
  END
END b15fpn000hn1n02x5

MACRO b15fpn000hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn000hn1n03x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.158 1.762 0.472 ;
      LAYER v0 ;
        RECT 1.694 0.338 1.762 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.018 0.178 2.086 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.91 0.178 1.978 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.338 1.672 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.182 0.158 0.25 0.382 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.722 0.248 0.79 0.382 ;
      RECT 1.046 0.518 1.262 0.562 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.37 0.248 1.438 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.158 1.87 0.562 ;
    LAYER v1 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.2705 1.438 0.3145 ;
      RECT 1.262 0.1535 1.33 0.1975 ;
      RECT 1.154 0.3155 1.222 0.3595 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.83 0.3155 0.898 0.3595 ;
      RECT 0.722 0.3155 0.79 0.3595 ;
      RECT 0.614 0.1575 0.682 0.2015 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.248 0.25 0.292 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 1.262 0.068 1.33 0.562 ;
  END
END b15fpn000hn1n03x5

MACRO b15fpn000hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn000hn1n04x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.158 1.762 0.472 ;
      LAYER v0 ;
        RECT 1.694 0.338 1.762 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.018 0.178 2.086 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.91 0.178 1.978 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.338 1.672 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.182 0.158 0.25 0.382 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.722 0.248 0.79 0.382 ;
      RECT 1.046 0.518 1.262 0.562 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.37 0.248 1.438 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.158 1.87 0.562 ;
    LAYER v1 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.2705 1.438 0.3145 ;
      RECT 1.262 0.1535 1.33 0.1975 ;
      RECT 1.154 0.3155 1.222 0.3595 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.83 0.3155 0.898 0.3595 ;
      RECT 0.722 0.3155 0.79 0.3595 ;
      RECT 0.614 0.1575 0.682 0.2015 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.248 0.25 0.292 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 1.262 0.068 1.33 0.562 ;
  END
END b15fpn000hn1n04x5

MACRO b15fpn000hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn000hn1n06x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.068 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.4055 2.086 0.4495 ;
        RECT 2.018 0.203 2.086 0.247 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.126 0.338 2.194 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.586 0.338 1.654 0.652 ;
        RECT 1.046 0.338 1.114 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.384 0.25 0.428 ;
        RECT 0.506 0.383 0.574 0.427 ;
        RECT 1.046 0.383 1.114 0.427 ;
        RECT 1.586 0.383 1.654 0.427 ;
        RECT 1.91 0.4055 1.978 0.4495 ;
        RECT 2.126 0.4055 2.194 0.4495 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.198 0.574 0.242 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.586 0.203 1.654 0.247 ;
        RECT 1.91 0.203 1.978 0.247 ;
        RECT 2.126 0.203 2.194 0.247 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.338 1.256 0.382 ;
      RECT 0.04 0.158 1.348 0.202 ;
      RECT 1.336 0.338 1.78 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.154 0.428 1.37 0.472 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.262 0.158 1.33 0.382 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.802 0.068 1.87 0.562 ;
    LAYER v1 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.158 0.894 0.202 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 1.802 0.203 1.87 0.247 ;
      RECT 1.802 0.4055 1.87 0.4495 ;
      RECT 1.694 0.498 1.762 0.542 ;
      RECT 1.478 0.088 1.546 0.132 ;
      RECT 1.478 0.498 1.546 0.542 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.198 0.79 0.242 ;
      RECT 0.614 0.198 0.682 0.242 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.384 0.142 0.428 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.79 0.428 1.006 0.472 ;
      RECT 0.79 0.068 1.114 0.112 ;
      RECT 1.37 0.158 1.438 0.472 ;
  END
END b15fpn000hn1n06x5

MACRO b15fpn000hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn000hn1n08x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.068 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.4645 2.086 0.5085 ;
        RECT 2.018 0.1205 2.086 0.1645 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.046 0.338 1.114 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.384 0.25 0.428 ;
        RECT 0.506 0.383 0.574 0.427 ;
        RECT 1.046 0.383 1.114 0.427 ;
        RECT 1.694 0.383 1.762 0.427 ;
        RECT 1.91 0.4645 1.978 0.5085 ;
        RECT 2.126 0.4645 2.194 0.5085 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.694 -0.022 1.762 0.292 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.198 0.574 0.242 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.694 0.203 1.762 0.247 ;
        RECT 1.91 0.1205 1.978 0.1645 ;
        RECT 2.126 0.1205 2.194 0.1645 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.338 1.256 0.382 ;
      RECT 0.04 0.158 1.348 0.202 ;
      RECT 1.336 0.338 1.996 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.154 0.428 1.37 0.472 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.262 0.158 1.33 0.382 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.91 0.248 1.978 0.382 ;
    LAYER v1 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.158 0.894 0.202 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.1205 1.87 0.1645 ;
      RECT 1.802 0.4645 1.87 0.5085 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.088 1.546 0.132 ;
      RECT 1.478 0.498 1.546 0.542 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.198 0.79 0.242 ;
      RECT 0.614 0.198 0.682 0.242 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.384 0.142 0.428 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.79 0.428 1.006 0.472 ;
      RECT 0.79 0.068 1.114 0.112 ;
      RECT 1.37 0.158 1.438 0.472 ;
  END
END b15fpn000hn1n08x5

MACRO b15fpn000hn1n08x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn000hn1n08x7 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.06625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.06625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.473 0.574 0.517 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.068 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.465 2.302 0.509 ;
        RECT 2.234 0.1205 2.302 0.1645 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.384 0.25 0.428 ;
        RECT 0.614 0.473 0.682 0.517 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 2.126 0.465 2.194 0.509 ;
        RECT 2.342 0.465 2.41 0.509 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.154 0.158 1.438 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.614 0.198 0.682 0.242 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.91 0.203 1.978 0.247 ;
        RECT 2.126 0.1205 2.194 0.1645 ;
        RECT 2.342 0.1205 2.41 0.1645 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 1.58 0.382 ;
      RECT 0.04 0.158 1.672 0.202 ;
      RECT 1.66 0.338 2.212 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 1.154 0.248 1.37 0.292 ;
      RECT 1.478 0.428 1.694 0.472 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 1.478 0.068 1.546 0.382 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 2.126 0.248 2.194 0.382 ;
    LAYER v1 ;
      RECT 2.13 0.338 2.19 0.382 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.59 0.158 1.65 0.202 ;
      RECT 1.482 0.338 1.542 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.158 0.894 0.202 ;
      RECT 0.402 0.338 0.462 0.382 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 2.126 0.293 2.194 0.337 ;
      RECT 2.018 0.203 2.086 0.247 ;
      RECT 2.018 0.383 2.086 0.427 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.203 1.762 0.247 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.383 1.438 0.427 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.046 0.198 1.114 0.242 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.722 0.198 0.79 0.242 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.384 0.466 0.428 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.384 0.142 0.428 ;
    LAYER m1 ;
      RECT 0.83 0.428 1.046 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 0.898 0.068 1.33 0.112 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.546 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.562 ;
  END
END b15fpn000hn1n08x7

MACRO b15fpn000hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn000hn1n12x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.06625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.06625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
        RECT 2.342 0.248 2.626 0.292 ;
        RECT 2.342 0.068 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.465 2.41 0.509 ;
        RECT 2.342 0.1175 2.41 0.1615 ;
        RECT 2.558 0.465 2.626 0.509 ;
        RECT 2.558 0.1175 2.626 0.1615 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.338 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.384 0.25 0.428 ;
        RECT 0.614 0.383 0.682 0.427 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 2.018 0.465 2.086 0.509 ;
        RECT 2.234 0.465 2.302 0.509 ;
        RECT 2.45 0.465 2.518 0.509 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.292 ;
        RECT 1.154 0.158 1.438 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.614 0.198 0.682 0.242 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 2.018 0.203 2.086 0.247 ;
        RECT 2.234 0.1175 2.302 0.1615 ;
        RECT 2.45 0.1175 2.518 0.1615 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 1.58 0.382 ;
      RECT 0.04 0.158 1.672 0.202 ;
      RECT 1.66 0.338 2.32 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 1.154 0.248 1.37 0.292 ;
      RECT 1.478 0.428 1.694 0.472 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 1.478 0.068 1.546 0.382 ;
      RECT 1.91 0.068 1.978 0.382 ;
      RECT 2.234 0.248 2.302 0.382 ;
    LAYER v1 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.59 0.158 1.65 0.202 ;
      RECT 1.482 0.338 1.542 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.158 0.894 0.202 ;
      RECT 0.402 0.338 0.462 0.382 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.126 0.203 2.194 0.247 ;
      RECT 2.126 0.465 2.194 0.509 ;
      RECT 1.91 0.088 1.978 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.203 1.762 0.247 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.383 1.438 0.427 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.046 0.198 1.114 0.242 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.722 0.198 0.79 0.242 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.384 0.466 0.428 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.384 0.142 0.428 ;
    LAYER m1 ;
      RECT 0.83 0.428 1.046 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 0.898 0.068 1.33 0.112 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.546 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.978 0.338 2.126 0.382 ;
      RECT 2.126 0.158 2.194 0.562 ;
  END
END b15fpn000hn1n12x5

MACRO b15fpn000hn1n12x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn000hn1n12x7 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.4385715 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.67833325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.562 ;
        RECT 2.666 0.248 2.95 0.292 ;
        RECT 2.666 0.068 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.666 0.138 2.734 0.182 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 2.882 0.138 2.95 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.586 0.338 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.384 0.25 0.428 ;
        RECT 0.722 0.403 0.79 0.447 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.4055 1.654 0.4495 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 1.78 0.382 ;
      RECT 0.04 0.158 1.996 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.046 0.248 1.114 0.382 ;
      RECT 0.938 0.428 1.154 0.472 ;
      RECT 1.262 0.158 1.33 0.382 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 1.478 0.068 1.546 0.472 ;
      RECT 1.91 0.158 1.978 0.382 ;
      RECT 1.802 0.428 2.018 0.472 ;
      RECT 2.45 0.068 2.518 0.562 ;
    LAYER v1 ;
      RECT 1.914 0.158 1.974 0.202 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.942 0.158 1.002 0.202 ;
      RECT 0.402 0.338 0.462 0.382 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.126 0.293 2.194 0.337 ;
      RECT 2.018 0.202 2.086 0.246 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.497 1.762 0.541 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.478 0.4055 1.546 0.4495 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.138 1.222 0.182 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.83 0.403 0.898 0.447 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.614 0.403 0.682 0.447 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.384 0.466 0.428 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.384 0.142 0.428 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.154 0.068 1.222 0.472 ;
      RECT 1.222 0.428 1.37 0.472 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.762 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.382 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 2.086 0.428 2.234 0.472 ;
      RECT 2.234 0.248 2.302 0.472 ;
  END
END b15fpn000hn1n12x7

MACRO b15fpn000hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn000hn1n16x5 0 0 ;
  SIZE 3.24 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.4385715 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.67833325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.068 3.058 0.562 ;
        RECT 2.774 0.338 3.058 0.382 ;
        RECT 2.774 0.068 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 2.99 0.138 3.058 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.274 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.586 0.338 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.384 0.25 0.428 ;
        RECT 0.722 0.403 0.79 0.447 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.4055 1.654 0.4495 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.45 0.538 2.518 0.582 ;
        RECT 2.666 0.538 2.734 0.582 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.274 0.022 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.292 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.234 0.202 2.302 0.246 ;
        RECT 2.45 0.1215 2.518 0.1655 ;
        RECT 2.666 0.138 2.734 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.098 0.138 3.166 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 1.78 0.382 ;
      RECT 0.04 0.158 1.996 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.046 0.248 1.114 0.382 ;
      RECT 0.938 0.428 1.154 0.472 ;
      RECT 1.262 0.158 1.33 0.382 ;
      RECT 1.802 0.428 2.018 0.472 ;
      RECT 1.478 0.068 1.546 0.472 ;
      RECT 1.91 0.158 1.978 0.382 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 2.342 0.248 2.41 0.472 ;
    LAYER v1 ;
      RECT 1.914 0.158 1.974 0.202 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.942 0.158 1.002 0.202 ;
      RECT 0.402 0.338 0.462 0.382 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.126 0.293 2.194 0.337 ;
      RECT 2.018 0.202 2.086 0.246 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.497 1.762 0.541 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.478 0.4055 1.546 0.4495 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.138 1.222 0.182 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.83 0.403 0.898 0.447 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.614 0.403 0.682 0.447 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.384 0.466 0.428 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.384 0.142 0.428 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.154 0.068 1.222 0.472 ;
      RECT 1.222 0.428 1.37 0.472 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 1.762 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.382 ;
      RECT 2.41 0.428 2.666 0.472 ;
      RECT 2.666 0.248 2.734 0.472 ;
  END
END b15fpn000hn1n16x5

MACRO b15fpn000hn1n16x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn000hn1n16x7 0 0 ;
  SIZE 3.564 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.9025 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.9025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.068 3.382 0.562 ;
        RECT 3.098 0.248 3.382 0.292 ;
        RECT 3.098 0.068 3.166 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.098 0.138 3.166 0.182 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.314 0.138 3.382 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.598 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.802 0.408 1.87 0.452 ;
        RECT 2.776 0.538 2.84 0.582 ;
        RECT 2.992 0.538 3.056 0.582 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.422 0.448 3.49 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.598 0.022 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 2.99 0.138 3.058 0.182 ;
        RECT 3.206 0.138 3.274 0.182 ;
        RECT 3.422 0.138 3.49 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.248 2.428 0.292 ;
      RECT 0.04 0.338 2.644 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.29 0.248 0.358 0.382 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.046 0.068 1.262 0.112 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.478 0.248 1.546 0.382 ;
      RECT 1.694 0.068 1.762 0.472 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.234 0.338 2.302 0.472 ;
      RECT 2.342 0.248 2.41 0.382 ;
      RECT 2.774 0.248 2.842 0.472 ;
      RECT 2.558 0.248 2.626 0.382 ;
    LAYER v1 ;
      RECT 2.562 0.338 2.622 0.382 ;
      RECT 2.346 0.248 2.406 0.292 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 1.482 0.248 1.542 0.292 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 0.942 0.248 1.002 0.292 ;
      RECT 0.402 0.248 0.462 0.292 ;
      RECT 0.294 0.338 0.354 0.382 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 2.99 0.293 3.058 0.337 ;
      RECT 2.882 0.428 2.95 0.472 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.558 0.293 2.626 0.337 ;
      RECT 2.45 0.202 2.518 0.246 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.342 0.518 2.41 0.562 ;
      RECT 2.234 0.202 2.302 0.246 ;
      RECT 2.234 0.408 2.302 0.452 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.694 0.138 1.762 0.182 ;
      RECT 1.694 0.408 1.762 0.452 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.178 1.438 0.222 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.83 0.088 0.898 0.132 ;
      RECT 0.83 0.498 0.898 0.542 ;
      RECT 0.614 0.088 0.682 0.132 ;
      RECT 0.614 0.498 0.682 0.542 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.4375 0.466 0.4815 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.562 ;
      RECT 0.898 0.158 1.154 0.202 ;
      RECT 1.154 0.158 1.222 0.382 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.114 0.428 1.37 0.472 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.762 0.248 1.91 0.292 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 1.978 0.248 2.126 0.292 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.086 0.518 2.45 0.562 ;
      RECT 2.302 0.068 2.45 0.112 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 2.842 0.428 2.99 0.472 ;
      RECT 2.99 0.248 3.058 0.472 ;
  END
END b15fpn000hn1n16x7

MACRO b15fpn010hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn010hn1n02x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.293 1.87 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.138 2.194 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 2.018 0.428 2.086 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.018 0.138 2.086 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.338 1.78 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 1.91 0.068 1.978 0.562 ;
    LAYER v1 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.482 0.338 1.542 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.473 1.762 0.517 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.264 0.498 1.328 0.542 ;
      RECT 1.154 0.3155 1.222 0.3595 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.338 0.25 0.382 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.33 0.428 1.37 0.472 ;
      RECT 1.37 0.068 1.438 0.472 ;
  END
END b15fpn010hn1n02x5

MACRO b15fpn010hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn010hn1n03x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.293 1.87 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.4235 2.194 0.4675 ;
        RECT 2.126 0.138 2.194 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 2.018 0.4235 2.086 0.4675 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.018 0.138 2.086 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.338 1.78 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 1.91 0.068 1.978 0.562 ;
    LAYER v1 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.482 0.338 1.542 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.4235 1.978 0.4675 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.473 1.762 0.517 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.264 0.498 1.328 0.542 ;
      RECT 1.154 0.3155 1.222 0.3595 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.338 0.25 0.382 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.33 0.428 1.37 0.472 ;
      RECT 1.37 0.068 1.438 0.472 ;
  END
END b15fpn010hn1n03x5

MACRO b15fpn010hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn010hn1n04x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.293 1.87 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.4235 2.194 0.4675 ;
        RECT 2.126 0.138 2.194 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 2.018 0.4235 2.086 0.4675 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.018 0.138 2.086 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.338 1.78 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 1.91 0.068 1.978 0.562 ;
    LAYER v1 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.482 0.338 1.542 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.4235 1.978 0.4675 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.473 1.762 0.517 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.264 0.498 1.328 0.542 ;
      RECT 1.154 0.3155 1.222 0.3595 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.338 0.25 0.382 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.33 0.428 1.37 0.472 ;
      RECT 1.37 0.068 1.438 0.472 ;
  END
END b15fpn010hn1n04x5

MACRO b15fpn010hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn010hn1n06x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.472 ;
      LAYER v0 ;
        RECT 2.018 0.248 2.086 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.397 2.41 0.441 ;
        RECT 2.342 0.138 2.41 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.234 0.397 2.302 0.441 ;
        RECT 2.45 0.397 2.518 0.441 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 1.154 0.192 1.222 0.236 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.248 1.996 0.292 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.694 0.158 1.762 0.382 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.126 0.068 2.194 0.472 ;
    LAYER v1 ;
      RECT 1.914 0.248 1.974 0.292 ;
      RECT 1.698 0.248 1.758 0.292 ;
      RECT 1.374 0.248 1.434 0.292 ;
      RECT 0.834 0.248 0.894 0.292 ;
      RECT 0.51 0.248 0.57 0.292 ;
    LAYER v0 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.397 2.194 0.441 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.192 1.33 0.236 ;
      RECT 1.262 0.448 1.33 0.492 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.155 0.79 0.199 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.614 0.155 0.682 0.199 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.074 0.248 0.142 0.292 ;
      RECT 0.074 0.4415 0.142 0.4855 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.142 0.158 0.398 0.202 ;
      RECT 0.398 0.068 0.466 0.202 ;
      RECT 0.466 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 1.006 0.338 1.262 0.382 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.546 0.338 1.586 0.382 ;
      RECT 1.586 0.068 1.654 0.382 ;
  END
END b15fpn010hn1n06x5

MACRO b15fpn010hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn010hn1n08x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.248 2.518 0.472 ;
      LAYER v0 ;
        RECT 2.45 0.293 2.518 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.4505 2.626 0.4945 ;
        RECT 2.558 0.113 2.626 0.157 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.29 0.473 0.358 0.517 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 2.018 0.473 2.086 0.517 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.666 0.4505 2.734 0.4945 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.1135 0.898 0.1575 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 2.018 0.113 2.086 0.157 ;
        RECT 2.45 0.113 2.518 0.157 ;
        RECT 2.666 0.113 2.734 0.157 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 2.32 0.382 ;
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 0.722 0.248 1.154 0.292 ;
      RECT 0.918 0.338 1.114 0.382 ;
      RECT 1.026 0.158 1.37 0.202 ;
      RECT 1.586 0.248 1.654 0.382 ;
      RECT 1.478 0.518 1.802 0.562 ;
      RECT 2.126 0.338 2.342 0.382 ;
      RECT 1.91 0.248 1.978 0.382 ;
    LAYER v1 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 2.342 0.113 2.41 0.157 ;
      RECT 2.342 0.4505 2.41 0.4945 ;
      RECT 1.91 0.2705 1.978 0.3145 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.694 0.2705 1.762 0.3145 ;
      RECT 1.586 0.2705 1.654 0.3145 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 1.48 0.178 1.544 0.222 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.38 0.574 0.424 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.473 0.25 0.517 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.248 0.466 0.562 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.466 0.518 0.702 0.562 ;
      RECT 0.682 0.428 1.006 0.472 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 1.222 0.248 1.478 0.292 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.438 0.068 1.694 0.112 ;
      RECT 1.694 0.068 1.762 0.382 ;
      RECT 1.802 0.158 1.87 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
  END
END b15fpn010hn1n08x5

MACRO b15fpn010hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn010hn1n12x5 0 0 ;
  SIZE 3.132 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5544445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.299 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.292 ;
      LAYER v0 ;
        RECT 2.342 0.113 2.41 0.157 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.068 3.058 0.562 ;
        RECT 2.774 0.338 3.058 0.382 ;
        RECT 2.774 0.068 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.774 0.113 2.842 0.157 ;
        RECT 2.99 0.428 3.058 0.472 ;
        RECT 2.99 0.113 3.058 0.157 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 2.126 0.538 2.194 0.582 ;
        RECT 2.45 0.538 2.518 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.166 0.022 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
        RECT 0.29 0.113 0.358 0.157 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 2.126 0.113 2.194 0.157 ;
        RECT 2.45 0.113 2.518 0.157 ;
        RECT 2.666 0.113 2.734 0.157 ;
        RECT 2.882 0.113 2.95 0.157 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 2.644 0.382 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.722 0.158 0.79 0.562 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.938 0.338 1.222 0.382 ;
      RECT 1.586 0.248 1.654 0.382 ;
      RECT 1.026 0.248 1.262 0.292 ;
      RECT 2.234 0.068 2.302 0.382 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 1.694 0.068 1.762 0.292 ;
      RECT 2.558 0.068 2.626 0.382 ;
    LAYER v1 ;
      RECT 2.562 0.338 2.622 0.382 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.558 0.113 2.626 0.157 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.234 0.113 2.302 0.157 ;
      RECT 2.126 0.2705 2.194 0.3145 ;
      RECT 2.018 0.2705 2.086 0.3145 ;
      RECT 1.91 0.178 1.978 0.222 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.178 1.762 0.222 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.586 0.2705 1.654 0.3145 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.448 1.33 0.492 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.218 0.79 0.262 ;
      RECT 0.506 0.197 0.574 0.241 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.398 0.197 0.466 0.241 ;
      RECT 0.182 0.113 0.25 0.157 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.682 0.562 ;
      RECT 0.79 0.518 1.114 0.562 ;
      RECT 0.466 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 0.898 0.158 1.37 0.202 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.438 0.068 1.654 0.112 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.33 0.248 1.478 0.292 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.546 0.428 1.802 0.472 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 2.302 0.338 2.43 0.382 ;
      RECT 1.478 0.518 1.91 0.562 ;
      RECT 1.762 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 1.978 0.428 2.126 0.472 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.194 0.428 2.666 0.472 ;
      RECT 2.666 0.248 2.734 0.472 ;
  END
END b15fpn010hn1n12x5

MACRO b15fpn010hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn010hn1n16x5 0 0 ;
  SIZE 3.78 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.7655555 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.7655555 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.292 ;
      LAYER v0 ;
        RECT 2.882 0.2035 2.95 0.2475 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.598 0.562 ;
        RECT 3.314 0.338 3.598 0.382 ;
        RECT 3.314 0.068 3.382 0.562 ;
      LAYER v0 ;
        RECT 3.314 0.428 3.382 0.472 ;
        RECT 3.314 0.113 3.382 0.157 ;
        RECT 3.53 0.428 3.598 0.472 ;
        RECT 3.53 0.203 3.598 0.247 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.814 0.652 ;
        RECT 3.638 0.518 3.706 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 3.206 0.518 3.274 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.99 0.538 3.058 0.582 ;
        RECT 3.206 0.538 3.274 0.582 ;
        RECT 3.424 0.538 3.488 0.582 ;
        RECT 3.64 0.538 3.704 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.814 0.022 ;
        RECT 3.638 -0.022 3.706 0.202 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.938 -0.022 1.006 0.292 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.262 0.129 1.33 0.173 ;
        RECT 1.478 0.129 1.546 0.173 ;
        RECT 1.694 0.129 1.762 0.173 ;
        RECT 2.666 0.1135 2.734 0.1575 ;
        RECT 2.99 0.1135 3.058 0.1575 ;
        RECT 3.206 0.113 3.274 0.157 ;
        RECT 3.422 0.113 3.49 0.157 ;
        RECT 3.638 0.113 3.706 0.157 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 3.184 0.382 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 1.046 0.248 1.114 0.382 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 2.774 0.068 2.842 0.382 ;
      RECT 2.558 0.248 2.626 0.382 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 3.098 0.158 3.166 0.382 ;
    LAYER v1 ;
      RECT 3.102 0.338 3.162 0.382 ;
      RECT 2.562 0.338 2.622 0.382 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.402 0.338 0.462 0.382 ;
    LAYER v0 ;
      RECT 3.206 0.313 3.274 0.357 ;
      RECT 3.098 0.203 3.166 0.247 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.774 0.1135 2.842 0.1575 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.558 0.293 2.626 0.337 ;
      RECT 2.45 0.1805 2.518 0.2245 ;
      RECT 2.342 0.1805 2.41 0.2245 ;
      RECT 2.342 0.518 2.41 0.562 ;
      RECT 2.234 0.1805 2.302 0.2245 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.1805 2.194 0.2245 ;
      RECT 2.126 0.518 2.194 0.562 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.616 0.448 0.68 0.492 ;
      RECT 0.398 0.268 0.466 0.312 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.29 0.472 ;
      RECT 0.074 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.338 0.722 0.382 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 0.682 0.518 1.114 0.562 ;
      RECT 0.898 0.428 1.154 0.472 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.222 0.248 1.91 0.292 ;
      RECT 1.91 0.068 1.978 0.292 ;
      RECT 1.978 0.068 2.194 0.112 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.472 ;
      RECT 1.87 0.428 2.126 0.472 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 2.194 0.428 2.342 0.472 ;
      RECT 2.342 0.158 2.41 0.472 ;
      RECT 2.842 0.338 3.058 0.382 ;
      RECT 2.018 0.518 2.45 0.562 ;
      RECT 2.302 0.068 2.45 0.112 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 2.518 0.428 2.666 0.472 ;
      RECT 2.666 0.248 2.734 0.472 ;
      RECT 2.734 0.428 3.206 0.472 ;
      RECT 3.206 0.248 3.274 0.472 ;
  END
END b15fpn010hn1n16x5

MACRO b15fpn040hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn040hn1n02x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.158 2.626 0.382 ;
      LAYER v0 ;
        RECT 2.558 0.248 2.626 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83901225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.068889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.381 2.95 0.425 ;
        RECT 2.882 0.1675 2.95 0.2115 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.774 0.381 2.842 0.425 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 0.722 0.248 1.222 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.722 0.158 0.79 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.724 0.178 0.788 0.222 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.694 0.114 1.762 0.158 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.774 0.1675 2.842 0.2115 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.812 0.518 2.752 0.562 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 1.37 0.068 1.438 0.472 ;
      RECT 1.674 0.248 1.802 0.292 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 1.802 0.518 2.126 0.562 ;
      RECT 2.666 0.068 2.734 0.562 ;
    LAYER v1 ;
      RECT 2.67 0.518 2.73 0.562 ;
      RECT 0.834 0.518 0.894 0.562 ;
    LAYER v0 ;
      RECT 2.666 0.1675 2.734 0.2115 ;
      RECT 2.666 0.381 2.734 0.425 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.018 0.3685 2.086 0.4125 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.802 0.114 1.87 0.158 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.386 1.438 0.43 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.3785 0.466 0.4225 ;
      RECT 0.29 0.518 0.358 0.562 ;
    LAYER m1 ;
      RECT 0.27 0.518 0.614 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.574 0.068 1.026 0.112 ;
      RECT 1.438 0.068 1.566 0.112 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.006 0.338 1.262 0.382 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.518 1.478 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.546 0.338 1.91 0.382 ;
      RECT 1.91 0.158 1.978 0.382 ;
      RECT 2.086 0.248 2.126 0.292 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.194 0.338 2.234 0.382 ;
      RECT 2.234 0.158 2.302 0.382 ;
      RECT 2.302 0.338 2.45 0.382 ;
      RECT 2.45 0.068 2.518 0.562 ;
  END
END b15fpn040hn1n02x5

MACRO b15fpn040hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn040hn1n03x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.158 2.626 0.382 ;
      LAYER v0 ;
        RECT 2.558 0.248 2.626 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83901225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.068889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.472 ;
      LAYER v0 ;
        RECT 2.882 0.383 2.95 0.427 ;
        RECT 2.882 0.1675 2.95 0.2115 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.774 0.383 2.842 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 0.722 0.248 1.222 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.722 0.158 0.79 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.724 0.178 0.788 0.222 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.694 0.114 1.762 0.158 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.774 0.1675 2.842 0.2115 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.812 0.518 2.752 0.562 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 1.37 0.068 1.438 0.472 ;
      RECT 1.674 0.248 1.802 0.292 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 1.802 0.518 2.126 0.562 ;
      RECT 2.666 0.068 2.734 0.562 ;
    LAYER v1 ;
      RECT 2.67 0.518 2.73 0.562 ;
      RECT 0.834 0.518 0.894 0.562 ;
    LAYER v0 ;
      RECT 2.666 0.1675 2.734 0.2115 ;
      RECT 2.666 0.383 2.734 0.427 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.018 0.3685 2.086 0.4125 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.802 0.114 1.87 0.158 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.386 1.438 0.43 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.3785 0.466 0.4225 ;
      RECT 0.29 0.518 0.358 0.562 ;
    LAYER m1 ;
      RECT 0.27 0.518 0.614 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.574 0.068 1.026 0.112 ;
      RECT 1.438 0.068 1.566 0.112 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.006 0.338 1.262 0.382 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.518 1.478 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.546 0.338 1.91 0.382 ;
      RECT 1.91 0.158 1.978 0.382 ;
      RECT 2.086 0.248 2.126 0.292 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.194 0.338 2.234 0.382 ;
      RECT 2.234 0.158 2.302 0.382 ;
      RECT 2.302 0.338 2.45 0.382 ;
      RECT 2.45 0.068 2.518 0.562 ;
  END
END b15fpn040hn1n03x5

MACRO b15fpn040hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn040hn1n04x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.158 2.626 0.382 ;
      LAYER v0 ;
        RECT 2.558 0.248 2.626 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83901225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.068889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.43 2.95 0.474 ;
        RECT 2.882 0.1675 2.95 0.2115 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.774 0.43 2.842 0.474 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 0.722 0.248 1.222 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.722 0.158 0.79 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.724 0.178 0.788 0.222 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.694 0.114 1.762 0.158 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.774 0.1675 2.842 0.2115 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.812 0.518 2.752 0.562 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 1.37 0.068 1.438 0.472 ;
      RECT 1.674 0.248 1.802 0.292 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 1.802 0.518 2.126 0.562 ;
      RECT 2.666 0.068 2.734 0.562 ;
    LAYER v1 ;
      RECT 2.67 0.518 2.73 0.562 ;
      RECT 0.834 0.518 0.894 0.562 ;
    LAYER v0 ;
      RECT 2.666 0.1675 2.734 0.2115 ;
      RECT 2.666 0.43 2.734 0.474 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.018 0.3685 2.086 0.4125 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.802 0.114 1.87 0.158 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.386 1.438 0.43 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.3785 0.466 0.4225 ;
      RECT 0.29 0.518 0.358 0.562 ;
    LAYER m1 ;
      RECT 0.27 0.518 0.614 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.574 0.068 1.026 0.112 ;
      RECT 1.438 0.068 1.566 0.112 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.006 0.338 1.262 0.382 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.518 1.478 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.546 0.338 1.91 0.382 ;
      RECT 1.91 0.158 1.978 0.382 ;
      RECT 2.086 0.248 2.126 0.292 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.194 0.338 2.234 0.382 ;
      RECT 2.234 0.158 2.302 0.382 ;
      RECT 2.302 0.338 2.45 0.382 ;
      RECT 2.45 0.068 2.518 0.562 ;
  END
END b15fpn040hn1n04x5

MACRO b15fpn040hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn040hn1n06x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.158 2.842 0.382 ;
      LAYER v0 ;
        RECT 2.774 0.248 2.842 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.068 3.166 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.098 0.138 3.166 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 1.586 0.428 1.998 0.472 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.403 0.25 0.447 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.206 0.448 3.274 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.183 0.25 0.227 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.694 0.114 1.762 0.158 ;
        RECT 1.91 0.114 1.978 0.158 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.99 0.138 3.058 0.182 ;
        RECT 3.206 0.138 3.274 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.812 0.518 2.968 0.562 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 1.37 0.068 1.438 0.472 ;
      RECT 1.674 0.248 1.802 0.292 ;
      RECT 0.938 0.068 1.006 0.562 ;
      RECT 2.214 0.428 2.342 0.472 ;
      RECT 1.782 0.518 2.45 0.562 ;
      RECT 2.882 0.068 2.95 0.562 ;
    LAYER v1 ;
      RECT 2.886 0.518 2.946 0.562 ;
      RECT 0.834 0.518 0.894 0.562 ;
    LAYER v0 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.882 0.448 2.95 0.492 ;
      RECT 2.666 0.138 2.734 0.182 ;
      RECT 2.666 0.448 2.734 0.492 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.342 0.1425 2.41 0.1865 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 1.802 0.114 1.87 0.158 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.386 1.438 0.43 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 0.938 0.138 1.006 0.182 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.83 0.358 0.898 0.402 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.398 0.384 0.466 0.428 ;
      RECT 0.398 0.518 0.466 0.562 ;
    LAYER m1 ;
      RECT 0.29 0.518 0.506 0.562 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 1.438 0.068 1.566 0.112 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.87 0.248 2.126 0.292 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 1.006 0.338 1.262 0.382 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.518 1.478 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.546 0.338 2.234 0.382 ;
      RECT 2.234 0.068 2.302 0.382 ;
      RECT 2.342 0.068 2.41 0.472 ;
      RECT 2.45 0.158 2.518 0.562 ;
      RECT 2.518 0.338 2.666 0.382 ;
      RECT 2.666 0.068 2.734 0.562 ;
  END
END b15fpn040hn1n06x5

MACRO b15fpn040hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn040hn1n08x5 0 0 ;
  SIZE 3.672 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.068 3.166 0.292 ;
      LAYER v0 ;
        RECT 3.098 0.088 3.166 0.132 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.736 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.81 0.112 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 0.722 0.068 0.79 0.112 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.158 3.49 0.562 ;
      LAYER v0 ;
        RECT 3.422 0.472 3.49 0.516 ;
        RECT 3.422 0.1885 3.49 0.2325 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.706 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 1.91 0.428 2.322 0.472 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 3.314 0.472 3.382 0.516 ;
        RECT 3.53 0.472 3.598 0.516 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.706 0.022 ;
        RECT 3.53 -0.022 3.598 0.292 ;
        RECT 3.314 -0.022 3.382 0.292 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.262 -0.022 1.33 0.292 ;
        RECT 0.702 0.248 1.114 0.292 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.262 0.2035 1.33 0.2475 ;
        RECT 2.018 0.114 2.086 0.158 ;
        RECT 2.234 0.114 2.302 0.158 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.314 0.1885 3.382 0.2325 ;
        RECT 3.53 0.1885 3.598 0.2325 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.518 0.7 0.562 ;
      RECT 1.028 0.518 3.076 0.562 ;
    LAYER m1 ;
      RECT 0.378 0.518 0.506 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.83 0.518 1.114 0.562 ;
      RECT 1.694 0.068 1.762 0.472 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.998 0.248 2.126 0.292 ;
      RECT 1.026 0.428 1.262 0.472 ;
      RECT 2.106 0.518 2.666 0.562 ;
      RECT 2.43 0.428 2.558 0.472 ;
      RECT 2.882 0.518 3.186 0.562 ;
    LAYER v1 ;
      RECT 2.994 0.518 3.054 0.562 ;
      RECT 1.05 0.518 1.11 0.562 ;
      RECT 0.618 0.518 0.678 0.562 ;
      RECT 0.186 0.518 0.246 0.562 ;
    LAYER v0 ;
      RECT 3.206 0.338 3.274 0.382 ;
      RECT 3.098 0.518 3.166 0.562 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.558 0.1535 2.626 0.1975 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.342 0.114 2.41 0.158 ;
      RECT 2.126 0.114 2.194 0.158 ;
      RECT 2.126 0.518 2.194 0.562 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.386 1.762 0.43 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.1885 1.546 0.2325 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.154 0.088 1.222 0.132 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.398 0.194 0.466 0.238 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.428 0.25 0.562 ;
      RECT 0.25 0.428 0.398 0.472 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.918 0.202 ;
      RECT 0.682 0.338 1.154 0.382 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.762 0.068 1.89 0.112 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.194 0.248 2.342 0.292 ;
      RECT 2.342 0.068 2.41 0.292 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.33 0.338 1.37 0.382 ;
      RECT 1.37 0.068 1.438 0.382 ;
      RECT 1.438 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.654 0.518 1.802 0.562 ;
      RECT 1.802 0.158 1.87 0.562 ;
      RECT 1.87 0.338 2.45 0.382 ;
      RECT 2.45 0.158 2.518 0.382 ;
      RECT 2.666 0.158 2.734 0.562 ;
      RECT 2.734 0.338 2.882 0.382 ;
      RECT 2.882 0.338 2.95 0.472 ;
      RECT 2.95 0.428 3.078 0.472 ;
      RECT 2.558 0.068 2.626 0.472 ;
      RECT 2.626 0.068 2.774 0.112 ;
      RECT 2.774 0.068 2.842 0.292 ;
      RECT 2.842 0.248 2.99 0.292 ;
      RECT 2.99 0.248 3.058 0.382 ;
      RECT 3.058 0.338 3.382 0.382 ;
  END
END b15fpn040hn1n08x5

MACRO b15fpn040hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn040hn1n12x5 0 0 ;
  SIZE 4.32 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.6044445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.805 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.338 3.814 0.382 ;
        RECT 3.746 0.068 3.814 0.382 ;
      LAYER v0 ;
        RECT 3.638 0.338 3.706 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.1046155 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.918 0.112 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.068 0.898 0.112 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.158 4.246 0.562 ;
        RECT 3.962 0.338 4.246 0.382 ;
        RECT 3.962 0.158 4.03 0.562 ;
      LAYER v0 ;
        RECT 3.962 0.472 4.03 0.516 ;
        RECT 3.962 0.203 4.03 0.247 ;
        RECT 4.178 0.472 4.246 0.516 ;
        RECT 4.178 0.203 4.246 0.247 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.354 0.652 ;
        RECT 4.07 0.428 4.138 0.652 ;
        RECT 3.854 0.428 3.922 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 3.854 0.472 3.922 0.516 ;
        RECT 4.07 0.472 4.138 0.516 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.354 0.022 ;
        RECT 4.07 -0.022 4.138 0.202 ;
        RECT 3.854 -0.022 3.922 0.202 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.702 0.248 1.222 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.154 0.1645 1.222 0.2085 ;
        RECT 1.478 0.114 1.546 0.158 ;
        RECT 2.234 0.114 2.302 0.158 ;
        RECT 2.45 0.114 2.518 0.158 ;
        RECT 3.424 0.048 3.488 0.092 ;
        RECT 3.854 0.113 3.922 0.157 ;
        RECT 4.07 0.113 4.138 0.157 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.518 0.824 0.562 ;
      RECT 0.904 0.518 3.832 0.562 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.83 0.518 1.026 0.562 ;
      RECT 1.35 0.248 1.802 0.292 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.026 0.338 1.586 0.382 ;
      RECT 2.214 0.248 2.342 0.292 ;
      RECT 2.646 0.518 3.206 0.562 ;
      RECT 2.754 0.428 3.098 0.472 ;
      RECT 3.746 0.428 3.814 0.562 ;
    LAYER v1 ;
      RECT 3.75 0.518 3.81 0.562 ;
      RECT 0.942 0.518 1.002 0.562 ;
      RECT 0.618 0.518 0.678 0.562 ;
      RECT 0.402 0.518 0.462 0.562 ;
    LAYER v0 ;
      RECT 3.746 0.472 3.814 0.516 ;
      RECT 3.64 0.088 3.704 0.132 ;
      RECT 3.53 0.248 3.598 0.292 ;
      RECT 3.422 0.448 3.49 0.492 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 3.098 0.15 3.166 0.194 ;
      RECT 2.99 0.15 3.058 0.194 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.884 0.318 2.948 0.362 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.342 0.114 2.41 0.158 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.018 0.361 2.086 0.405 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.802 0.3605 1.87 0.4045 ;
      RECT 1.696 0.138 1.76 0.182 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.506 0.49 0.574 0.534 ;
      RECT 0.398 0.194 0.466 0.238 ;
      RECT 0.29 0.428 0.358 0.472 ;
    LAYER m1 ;
      RECT 0.27 0.428 0.398 0.472 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.574 0.158 0.918 0.202 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.026 0.472 ;
      RECT 1.802 0.248 1.87 0.472 ;
      RECT 1.762 0.068 2.018 0.112 ;
      RECT 2.018 0.068 2.086 0.472 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.654 0.518 1.91 0.562 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 1.978 0.518 2.126 0.562 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.194 0.338 2.754 0.382 ;
      RECT 2.342 0.068 2.41 0.292 ;
      RECT 2.41 0.248 2.882 0.292 ;
      RECT 2.882 0.248 2.95 0.382 ;
      RECT 2.95 0.248 2.99 0.292 ;
      RECT 2.99 0.068 3.058 0.292 ;
      RECT 3.206 0.158 3.274 0.562 ;
      RECT 3.274 0.338 3.422 0.382 ;
      RECT 3.422 0.248 3.49 0.562 ;
      RECT 3.49 0.248 3.618 0.292 ;
      RECT 3.098 0.068 3.166 0.472 ;
      RECT 3.166 0.068 3.314 0.112 ;
      RECT 3.314 0.068 3.382 0.202 ;
      RECT 3.382 0.158 3.638 0.202 ;
      RECT 3.638 0.068 3.706 0.202 ;
  END
END b15fpn040hn1n12x5

MACRO b15fpn040hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn040hn1n16x5 0 0 ;
  SIZE 5.076 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33234575 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.338 4.462 0.382 ;
        RECT 4.394 0.158 4.462 0.382 ;
      LAYER v0 ;
        RECT 4.286 0.338 4.354 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53079375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 1.222 0.112 ;
        RECT 0.506 0.068 0.574 0.382 ;
        RECT 0.182 0.158 0.574 0.202 ;
        RECT 0.182 0.068 0.25 0.202 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 1.046 0.068 1.114 0.112 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.826 0.158 4.894 0.562 ;
        RECT 4.61 0.338 4.894 0.382 ;
        RECT 4.61 0.158 4.678 0.562 ;
      LAYER v0 ;
        RECT 4.61 0.472 4.678 0.516 ;
        RECT 4.61 0.1885 4.678 0.2325 ;
        RECT 4.826 0.472 4.894 0.516 ;
        RECT 4.826 0.1885 4.894 0.2325 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.11 0.652 ;
        RECT 4.934 0.428 5.002 0.652 ;
        RECT 4.718 0.428 4.786 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 2.97 0.428 3.294 0.472 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.478 0.471 1.546 0.515 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.99 0.428 3.058 0.472 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.962 0.448 4.03 0.492 ;
        RECT 4.178 0.448 4.246 0.492 ;
        RECT 4.502 0.472 4.57 0.516 ;
        RECT 4.718 0.472 4.786 0.516 ;
        RECT 4.934 0.472 5.002 0.516 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.11 0.022 ;
        RECT 4.934 -0.022 5.002 0.292 ;
        RECT 4.718 -0.022 4.786 0.292 ;
        RECT 4.502 -0.022 4.57 0.292 ;
        RECT 4.07 -0.022 4.138 0.112 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 1.478 0.248 1.89 0.292 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 0.918 0.158 1.33 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.478 0.1655 1.546 0.2095 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.99 0.1285 3.058 0.1725 ;
        RECT 3.206 0.1285 3.274 0.1725 ;
        RECT 4.072 0.048 4.136 0.092 ;
        RECT 4.502 0.1885 4.57 0.2325 ;
        RECT 4.718 0.1885 4.786 0.2325 ;
        RECT 4.934 0.1885 5.002 0.2325 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.518 1.04 0.562 ;
      RECT 1.12 0.518 4.48 0.562 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.722 0.248 0.79 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 1.046 0.518 1.242 0.562 ;
      RECT 1.674 0.158 2.018 0.202 ;
      RECT 2.214 0.338 2.342 0.382 ;
      RECT 1.35 0.338 1.91 0.382 ;
      RECT 2.774 0.338 3.422 0.382 ;
      RECT 3.206 0.518 3.854 0.562 ;
      RECT 3.53 0.068 3.598 0.292 ;
      RECT 4.394 0.428 4.462 0.562 ;
    LAYER v1 ;
      RECT 4.398 0.518 4.458 0.562 ;
      RECT 1.158 0.518 1.218 0.562 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.618 0.518 0.678 0.562 ;
      RECT 0.078 0.518 0.138 0.562 ;
    LAYER v0 ;
      RECT 4.394 0.472 4.462 0.516 ;
      RECT 4.288 0.088 4.352 0.132 ;
      RECT 4.178 0.248 4.246 0.292 ;
      RECT 4.07 0.448 4.138 0.492 ;
      RECT 3.854 0.248 3.922 0.292 ;
      RECT 3.748 0.138 3.812 0.182 ;
      RECT 3.638 0.223 3.706 0.267 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.53 0.338 3.598 0.382 ;
      RECT 3.532 0.138 3.596 0.182 ;
      RECT 3.422 0.223 3.49 0.267 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 3.314 0.1285 3.382 0.1725 ;
      RECT 3.314 0.518 3.382 0.562 ;
      RECT 3.098 0.338 3.166 0.382 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.452 0.178 2.516 0.222 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.02 0.358 2.084 0.402 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.156 0.318 1.22 0.362 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.49 0.79 0.534 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.158 0.81 0.202 ;
      RECT 0.79 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.472 ;
      RECT 1.114 0.428 1.438 0.472 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 2.086 0.158 2.214 0.202 ;
      RECT 2.086 0.428 2.43 0.472 ;
      RECT 1.998 0.068 2.342 0.112 ;
      RECT 2.342 0.068 2.41 0.382 ;
      RECT 2.41 0.338 2.538 0.382 ;
      RECT 2.41 0.068 2.558 0.112 ;
      RECT 2.558 0.068 2.626 0.202 ;
      RECT 2.626 0.158 2.862 0.202 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 2.45 0.158 2.518 0.292 ;
      RECT 1.978 0.518 2.666 0.562 ;
      RECT 2.518 0.248 2.666 0.292 ;
      RECT 2.666 0.248 2.734 0.562 ;
      RECT 2.734 0.248 3.314 0.292 ;
      RECT 3.314 0.068 3.382 0.292 ;
      RECT 3.422 0.158 3.49 0.382 ;
      RECT 3.49 0.338 3.638 0.382 ;
      RECT 3.638 0.158 3.706 0.382 ;
      RECT 3.854 0.158 3.922 0.562 ;
      RECT 3.922 0.338 4.07 0.382 ;
      RECT 4.07 0.248 4.138 0.562 ;
      RECT 4.138 0.248 4.266 0.292 ;
      RECT 3.402 0.428 3.746 0.472 ;
      RECT 3.598 0.068 3.746 0.112 ;
      RECT 3.746 0.068 3.814 0.472 ;
      RECT 3.814 0.068 3.962 0.112 ;
      RECT 3.962 0.068 4.03 0.202 ;
      RECT 4.03 0.158 4.286 0.202 ;
      RECT 4.286 0.068 4.354 0.202 ;
  END
END b15fpn040hn1n16x5

MACRO b15fpn080hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn080hn1n02x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.068 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.293 1.762 0.337 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.068 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.018 0.178 2.086 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.91 0.178 1.978 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 1.564 0.382 ;
      RECT 0.164 0.158 1.996 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 1.046 0.518 1.262 0.562 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.068 1.87 0.562 ;
    LAYER v1 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.158 0.246 0.202 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.2705 1.438 0.3145 ;
      RECT 1.262 0.1535 1.33 0.1975 ;
      RECT 1.154 0.3155 1.222 0.3595 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.83 0.3155 0.898 0.3595 ;
      RECT 0.722 0.3155 0.79 0.3595 ;
      RECT 0.614 0.1575 0.682 0.2015 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.248 0.25 0.292 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 1.262 0.068 1.33 0.562 ;
  END
END b15fpn080hn1n02x5

MACRO b15fpn080hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn080hn1n03x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.976 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.976 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.068 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.293 1.762 0.337 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.068 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.018 0.178 2.086 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.91 0.178 1.978 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 1.564 0.382 ;
      RECT 0.164 0.158 1.996 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 1.046 0.518 1.262 0.562 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.802 0.068 1.87 0.562 ;
    LAYER v1 ;
      RECT 1.806 0.158 1.866 0.202 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.158 0.246 0.202 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.2705 1.438 0.3145 ;
      RECT 1.262 0.1535 1.33 0.1975 ;
      RECT 1.154 0.3155 1.222 0.3595 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.83 0.3155 0.898 0.3595 ;
      RECT 0.722 0.3155 0.79 0.3595 ;
      RECT 0.614 0.1575 0.682 0.2015 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.248 0.25 0.292 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 1.262 0.068 1.33 0.562 ;
  END
END b15fpn080hn1n03x5

MACRO b15fpn080hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn080hn1n04x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.018 0.178 2.086 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.91 0.178 1.978 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.158 1.672 0.202 ;
      RECT 0.488 0.338 1.78 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 1.046 0.518 1.262 0.562 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.802 0.158 1.87 0.562 ;
    LAYER v1 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.59 0.158 1.65 0.202 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.694 0.178 1.762 0.222 ;
      RECT 1.586 0.3155 1.654 0.3595 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.1535 1.33 0.1975 ;
      RECT 1.154 0.3155 1.222 0.3595 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.83 0.3155 0.898 0.3595 ;
      RECT 0.722 0.3155 0.79 0.3595 ;
      RECT 0.614 0.1575 0.682 0.2015 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.074 0.133 0.142 0.177 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 1.262 0.068 1.33 0.562 ;
  END
END b15fpn080hn1n04x5

MACRO b15fpn080hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn080hn1n06x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.068 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.4645 2.086 0.5085 ;
        RECT 2.018 0.1205 2.086 0.1645 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.046 0.338 1.114 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 0.506 0.4645 0.574 0.5085 ;
        RECT 1.046 0.383 1.114 0.427 ;
        RECT 1.694 0.383 1.762 0.427 ;
        RECT 1.91 0.4645 1.978 0.5085 ;
        RECT 2.126 0.4645 2.194 0.5085 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.694 -0.022 1.762 0.292 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.116 0.25 0.16 ;
        RECT 0.506 0.116 0.574 0.16 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.694 0.203 1.762 0.247 ;
        RECT 1.91 0.1205 1.978 0.1645 ;
        RECT 2.126 0.1205 2.194 0.1645 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.338 1.256 0.382 ;
      RECT 0.04 0.158 1.348 0.202 ;
      RECT 1.336 0.338 1.996 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.154 0.428 1.37 0.472 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.91 0.248 1.978 0.382 ;
    LAYER v1 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.158 0.894 0.202 ;
      RECT 0.294 0.158 0.354 0.202 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.1205 1.87 0.1645 ;
      RECT 1.802 0.4645 1.87 0.5085 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.088 1.546 0.132 ;
      RECT 1.478 0.498 1.546 0.542 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.203 0.79 0.247 ;
      RECT 0.614 0.116 0.682 0.16 ;
      RECT 0.614 0.4645 0.682 0.5085 ;
      RECT 0.29 0.116 0.358 0.16 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.79 0.428 1.006 0.472 ;
      RECT 0.79 0.068 1.114 0.112 ;
      RECT 1.37 0.158 1.438 0.472 ;
  END
END b15fpn080hn1n06x5

MACRO b15fpn080hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn080hn1n08x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.068 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.4645 2.086 0.5085 ;
        RECT 2.018 0.1205 2.086 0.1645 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.046 0.338 1.114 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 0.506 0.4645 0.574 0.5085 ;
        RECT 1.046 0.383 1.114 0.427 ;
        RECT 1.694 0.383 1.762 0.427 ;
        RECT 1.91 0.4645 1.978 0.5085 ;
        RECT 2.126 0.4645 2.194 0.5085 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.694 -0.022 1.762 0.292 ;
        RECT 0.938 0.158 1.222 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.116 0.25 0.16 ;
        RECT 0.506 0.116 0.574 0.16 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.694 0.203 1.762 0.247 ;
        RECT 1.91 0.1205 1.978 0.1645 ;
        RECT 2.126 0.1205 2.194 0.1645 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.338 1.256 0.382 ;
      RECT 0.04 0.158 1.348 0.202 ;
      RECT 1.336 0.338 1.996 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.154 0.428 1.37 0.472 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.91 0.248 1.978 0.382 ;
    LAYER v1 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.158 0.894 0.202 ;
      RECT 0.294 0.158 0.354 0.202 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.1205 1.87 0.1645 ;
      RECT 1.802 0.4645 1.87 0.5085 ;
      RECT 1.586 0.088 1.654 0.132 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.088 1.546 0.132 ;
      RECT 1.478 0.498 1.546 0.542 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.203 0.79 0.247 ;
      RECT 0.614 0.116 0.682 0.16 ;
      RECT 0.614 0.4645 0.682 0.5085 ;
      RECT 0.29 0.116 0.358 0.16 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.79 0.428 1.006 0.472 ;
      RECT 0.79 0.068 1.114 0.112 ;
      RECT 1.37 0.158 1.438 0.472 ;
  END
END b15fpn080hn1n08x5

MACRO b15fpn080hn1n08x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn080hn1n08x7 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.06625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.06625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.473 0.574 0.517 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.068 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.465 2.302 0.509 ;
        RECT 2.234 0.1205 2.302 0.1645 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.384 0.25 0.428 ;
        RECT 0.614 0.473 0.682 0.517 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 2.126 0.465 2.194 0.509 ;
        RECT 2.342 0.465 2.41 0.509 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.154 0.158 1.438 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.614 0.198 0.682 0.242 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.91 0.203 1.978 0.247 ;
        RECT 2.126 0.1205 2.194 0.1645 ;
        RECT 2.342 0.1205 2.41 0.1645 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 1.58 0.382 ;
      RECT 0.04 0.158 1.672 0.202 ;
      RECT 1.66 0.338 2.212 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 1.154 0.248 1.37 0.292 ;
      RECT 1.478 0.428 1.694 0.472 ;
      RECT 1.478 0.248 1.546 0.382 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 2.126 0.248 2.194 0.382 ;
    LAYER v1 ;
      RECT 2.13 0.338 2.19 0.382 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.482 0.158 1.542 0.202 ;
      RECT 1.482 0.338 1.542 0.382 ;
      RECT 0.942 0.158 1.002 0.202 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.402 0.338 0.462 0.382 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 2.126 0.293 2.194 0.337 ;
      RECT 2.018 0.203 2.086 0.247 ;
      RECT 2.018 0.383 2.086 0.427 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.203 1.762 0.247 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.383 1.438 0.427 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.046 0.203 1.114 0.247 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.722 0.198 0.79 0.242 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.384 0.466 0.428 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.384 0.142 0.428 ;
    LAYER m1 ;
      RECT 0.83 0.428 1.046 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 0.898 0.068 1.33 0.112 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.546 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.562 ;
  END
END b15fpn080hn1n08x7

MACRO b15fpn080hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn080hn1n12x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.06625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.06625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
        RECT 2.342 0.248 2.626 0.292 ;
        RECT 2.342 0.068 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.465 2.41 0.509 ;
        RECT 2.342 0.1175 2.41 0.1615 ;
        RECT 2.558 0.465 2.626 0.509 ;
        RECT 2.558 0.1175 2.626 0.1615 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.338 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.384 0.25 0.428 ;
        RECT 0.614 0.383 0.682 0.427 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 2.018 0.465 2.086 0.509 ;
        RECT 2.234 0.465 2.302 0.509 ;
        RECT 2.45 0.465 2.518 0.509 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.292 ;
        RECT 1.154 0.158 1.438 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.614 0.198 0.682 0.242 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 2.018 0.203 2.086 0.247 ;
        RECT 2.234 0.1175 2.302 0.1615 ;
        RECT 2.45 0.1175 2.518 0.1615 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 1.58 0.382 ;
      RECT 0.04 0.158 1.672 0.202 ;
      RECT 1.66 0.338 2.32 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 1.154 0.248 1.37 0.292 ;
      RECT 1.478 0.428 1.694 0.472 ;
      RECT 1.478 0.248 1.546 0.382 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 1.91 0.068 1.978 0.382 ;
      RECT 2.234 0.248 2.302 0.382 ;
    LAYER v1 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.482 0.158 1.542 0.202 ;
      RECT 1.482 0.338 1.542 0.382 ;
      RECT 0.942 0.158 1.002 0.202 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.402 0.338 0.462 0.382 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.126 0.203 2.194 0.247 ;
      RECT 2.126 0.465 2.194 0.509 ;
      RECT 1.91 0.088 1.978 0.132 ;
      RECT 1.802 0.498 1.87 0.542 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.203 1.762 0.247 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.383 1.438 0.427 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.048 0.2005 1.112 0.2445 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.722 0.198 0.79 0.242 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.384 0.466 0.428 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.384 0.142 0.428 ;
    LAYER m1 ;
      RECT 0.83 0.518 1.046 0.562 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 0.898 0.068 1.33 0.112 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.546 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.978 0.338 2.126 0.382 ;
      RECT 2.126 0.158 2.194 0.562 ;
  END
END b15fpn080hn1n12x5

MACRO b15fpn080hn1n12x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn080hn1n12x7 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 3.07166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 3.07166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.428 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.448 2.302 0.492 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.562 ;
        RECT 2.666 0.338 2.95 0.382 ;
        RECT 2.666 0.068 2.734 0.382 ;
      LAYER v0 ;
        RECT 2.666 0.1525 2.734 0.1965 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 2.882 0.1525 2.95 0.1965 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.91 0.473 1.978 0.517 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.558 -0.022 2.626 0.292 ;
        RECT 2.342 -0.022 2.41 0.292 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.91 0.138 1.978 0.182 ;
        RECT 2.342 0.1525 2.41 0.1965 ;
        RECT 2.558 0.1525 2.626 0.1965 ;
        RECT 2.774 0.1525 2.842 0.1965 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.428 1.996 0.472 ;
    LAYER m1 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.722 0.518 0.938 0.562 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.586 0.158 1.654 0.562 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.694 0.248 1.762 0.562 ;
      RECT 1.802 0.338 2.45 0.382 ;
    LAYER v1 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.402 0.428 0.462 0.472 ;
    LAYER v0 ;
      RECT 2.45 0.1525 2.518 0.1965 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.234 0.1525 2.302 0.1965 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.43 1.654 0.474 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.37 0.138 1.438 0.182 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.154 0.138 1.222 0.182 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.466 0.338 0.79 0.382 ;
      RECT 0.614 0.158 0.938 0.202 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.006 0.338 1.33 0.382 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.654 0.158 1.802 0.202 ;
      RECT 1.802 0.158 1.87 0.292 ;
      RECT 1.87 0.248 2.234 0.292 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.45 0.068 2.518 0.562 ;
  END
END b15fpn080hn1n12x7

MACRO b15fpn080hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn080hn1n16x5 0 0 ;
  SIZE 3.24 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.4385715 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.67833325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.068 3.058 0.562 ;
        RECT 2.774 0.338 3.058 0.382 ;
        RECT 2.774 0.068 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 2.99 0.138 3.058 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.274 0.652 ;
        RECT 3.098 0.338 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.586 0.338 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.384 0.25 0.428 ;
        RECT 0.722 0.403 0.79 0.447 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.4055 1.654 0.4495 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.45 0.538 2.518 0.582 ;
        RECT 2.666 0.538 2.734 0.582 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.274 0.022 ;
        RECT 3.098 -0.022 3.166 0.292 ;
        RECT 2.882 -0.022 2.95 0.292 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.292 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.234 0.202 2.302 0.246 ;
        RECT 2.45 0.1215 2.518 0.1655 ;
        RECT 2.666 0.138 2.734 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.098 0.138 3.166 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 1.78 0.382 ;
      RECT 0.164 0.158 2.104 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.046 0.248 1.114 0.382 ;
      RECT 0.938 0.428 1.154 0.472 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.802 0.428 2.018 0.472 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.91 0.158 1.978 0.382 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 2.342 0.248 2.41 0.472 ;
    LAYER v1 ;
      RECT 1.914 0.158 1.974 0.202 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.942 0.158 1.002 0.202 ;
      RECT 0.402 0.158 0.462 0.202 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.126 0.293 2.194 0.337 ;
      RECT 2.018 0.202 2.086 0.246 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.497 1.762 0.541 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.478 0.4055 1.546 0.4495 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.138 1.222 0.182 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.83 0.403 0.898 0.447 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.614 0.403 0.682 0.447 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.384 0.466 0.428 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.384 0.142 0.428 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.562 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.154 0.068 1.222 0.472 ;
      RECT 1.222 0.428 1.37 0.472 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 1.762 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.382 ;
      RECT 2.41 0.428 2.666 0.472 ;
      RECT 2.666 0.248 2.734 0.472 ;
  END
END b15fpn080hn1n16x5

MACRO b15fpn080hn1n16x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpn080hn1n16x7 0 0 ;
  SIZE 3.564 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.9025 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.9025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.068 3.382 0.562 ;
        RECT 3.098 0.248 3.382 0.292 ;
        RECT 3.098 0.068 3.166 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.098 0.138 3.166 0.182 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.314 0.138 3.382 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.598 0.652 ;
        RECT 3.422 0.338 3.49 0.652 ;
        RECT 3.206 0.338 3.274 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.776 0.538 2.84 0.582 ;
        RECT 2.992 0.538 3.056 0.582 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.422 0.448 3.49 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.598 0.022 ;
        RECT 3.422 -0.022 3.49 0.292 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.722 0.088 0.79 0.132 ;
        RECT 1.586 0.135 1.654 0.179 ;
        RECT 1.802 0.135 1.87 0.179 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 2.99 0.138 3.058 0.182 ;
        RECT 3.206 0.138 3.274 0.182 ;
        RECT 3.422 0.138 3.49 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 2.644 0.382 ;
      RECT 0.38 0.158 2.752 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 2.018 0.068 2.086 0.202 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.342 0.248 2.41 0.472 ;
      RECT 2.774 0.248 2.842 0.472 ;
      RECT 2.558 0.068 2.626 0.382 ;
    LAYER v1 ;
      RECT 2.562 0.158 2.622 0.202 ;
      RECT 2.346 0.338 2.406 0.382 ;
      RECT 2.022 0.158 2.082 0.202 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 0.942 0.158 1.002 0.202 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.402 0.158 0.462 0.202 ;
      RECT 0.294 0.338 0.354 0.382 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 2.99 0.293 3.058 0.337 ;
      RECT 2.882 0.428 2.95 0.472 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.558 0.293 2.626 0.337 ;
      RECT 2.45 0.202 2.518 0.246 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.342 0.518 2.41 0.562 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 2.018 0.135 2.086 0.179 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.135 1.978 0.179 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.694 0.135 1.762 0.179 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.586 0.3155 1.654 0.3595 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.313 1.438 0.357 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.938 0.088 1.006 0.132 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.83 0.088 0.898 0.132 ;
      RECT 0.83 0.498 0.898 0.542 ;
      RECT 0.614 0.088 0.682 0.132 ;
      RECT 0.614 0.498 0.682 0.542 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.4375 0.466 0.4815 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.562 ;
      RECT 0.898 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.046 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.518 1.478 0.562 ;
      RECT 1.478 0.428 1.546 0.562 ;
      RECT 1.33 0.158 1.546 0.202 ;
      RECT 1.546 0.428 1.586 0.472 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.978 0.248 2.126 0.292 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.086 0.518 2.45 0.562 ;
      RECT 2.302 0.068 2.45 0.112 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 2.842 0.428 2.99 0.472 ;
      RECT 2.99 0.248 3.058 0.472 ;
  END
END b15fpn080hn1n16x7

MACRO b15fpy000hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy000hn1n02x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.338 2.302 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.158 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.558 0.2085 2.626 0.2525 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.478 0.408 1.546 0.452 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.45 0.2085 2.518 0.2525 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.428 1.996 0.472 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.37 0.248 1.586 0.292 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.586 0.518 1.802 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.91 0.158 1.978 0.472 ;
      RECT 2.342 0.158 2.41 0.562 ;
    LAYER v1 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 0.942 0.428 1.002 0.472 ;
    LAYER v0 ;
      RECT 2.342 0.2085 2.41 0.2525 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.802 0.1535 1.87 0.1975 ;
      RECT 1.694 0.3155 1.762 0.3595 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.1575 1.222 0.2015 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.1575 1.114 0.2015 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.508 0.231 0.572 0.275 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.978 0.338 2.126 0.382 ;
      RECT 2.126 0.068 2.194 0.562 ;
  END
END b15fpy000hn1n02x5

MACRO b15fpy000hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy000hn1n03x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.338 2.302 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.158 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.558 0.2085 2.626 0.2525 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.478 0.408 1.546 0.452 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.45 0.2085 2.518 0.2525 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.428 1.996 0.472 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.37 0.248 1.586 0.292 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.586 0.518 1.802 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.91 0.158 1.978 0.472 ;
      RECT 2.342 0.158 2.41 0.562 ;
    LAYER v1 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 0.942 0.428 1.002 0.472 ;
    LAYER v0 ;
      RECT 2.342 0.2085 2.41 0.2525 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.802 0.1535 1.87 0.1975 ;
      RECT 1.694 0.3155 1.762 0.3595 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.1575 1.222 0.2015 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.1575 1.114 0.2015 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.508 0.231 0.572 0.275 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.978 0.338 2.126 0.382 ;
      RECT 2.126 0.068 2.194 0.562 ;
  END
END b15fpy000hn1n03x5

MACRO b15fpy000hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy000hn1n04x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.338 2.302 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.4285 2.626 0.4725 ;
        RECT 2.558 0.1585 2.626 0.2025 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.478 0.408 1.546 0.452 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.45 0.4285 2.518 0.4725 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.45 0.1585 2.518 0.2025 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.428 1.996 0.472 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.37 0.248 1.586 0.292 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.586 0.518 1.802 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.91 0.158 1.978 0.472 ;
      RECT 2.342 0.068 2.41 0.562 ;
    LAYER v1 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 0.942 0.428 1.002 0.472 ;
    LAYER v0 ;
      RECT 2.342 0.1585 2.41 0.2025 ;
      RECT 2.342 0.4285 2.41 0.4725 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.802 0.1535 1.87 0.1975 ;
      RECT 1.694 0.3155 1.762 0.3595 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.1575 1.222 0.2015 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.1575 1.114 0.2015 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.508 0.231 0.572 0.275 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.978 0.338 2.126 0.382 ;
      RECT 2.126 0.068 2.194 0.562 ;
  END
END b15fpy000hn1n04x5

MACRO b15fpy000hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy000hn1n06x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.248 2.41 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.3155 2.41 0.3595 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.406 2.734 0.45 ;
        RECT 2.666 0.1805 2.734 0.2245 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.126 0.338 2.194 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.452 0.25 0.496 ;
        RECT 0.722 0.452 0.79 0.496 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.558 0.406 2.626 0.45 ;
        RECT 2.774 0.406 2.842 0.45 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.558 -0.022 2.626 0.292 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1975 0.25 0.2415 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.558 0.1805 2.626 0.2245 ;
        RECT 2.774 0.1805 2.842 0.2245 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.428 2.32 0.472 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.802 0.158 1.87 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.45 0.068 2.518 0.562 ;
    LAYER v1 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 0.942 0.428 1.002 0.472 ;
    LAYER v0 ;
      RECT 2.45 0.1805 2.518 0.2245 ;
      RECT 2.45 0.406 2.518 0.45 ;
      RECT 2.234 0.138 2.302 0.182 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.2705 2.086 0.3145 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.1575 1.222 0.2015 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.1575 1.114 0.2015 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.508 0.2345 0.572 0.2785 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.87 0.158 2.086 0.202 ;
  END
END b15fpy000hn1n06x5

MACRO b15fpy000hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy000hn1n08x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.248 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.338 2.41 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.158 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.424 2.734 0.468 ;
        RECT 2.666 0.178 2.734 0.222 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.126 0.338 2.194 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.452 0.25 0.496 ;
        RECT 0.722 0.452 0.79 0.496 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.558 0.424 2.626 0.468 ;
        RECT 2.774 0.424 2.842 0.468 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.558 -0.022 2.626 0.292 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1975 0.25 0.2415 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.558 0.178 2.626 0.222 ;
        RECT 2.774 0.178 2.842 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.428 2.32 0.472 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.802 0.158 1.87 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.45 0.158 2.518 0.562 ;
    LAYER v1 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 0.942 0.428 1.002 0.472 ;
    LAYER v0 ;
      RECT 2.45 0.178 2.518 0.222 ;
      RECT 2.45 0.424 2.518 0.468 ;
      RECT 2.234 0.138 2.302 0.182 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.2705 2.086 0.3145 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.1575 1.222 0.2015 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.1575 1.114 0.2015 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.508 0.2345 0.572 0.2785 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.87 0.158 2.086 0.202 ;
  END
END b15fpy000hn1n08x5

MACRO b15fpy000hn1n08x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy000hn1n08x7 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.338 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.4665 2.842 0.5105 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.825679 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.81 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.068 3.166 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.4665 3.166 0.5105 ;
        RECT 3.098 0.158 3.166 0.202 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.61777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.452 0.25 0.496 ;
        RECT 0.722 0.473 0.79 0.517 ;
        RECT 1.478 0.472 1.546 0.516 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.558 0.4665 2.626 0.5105 ;
        RECT 2.99 0.4665 3.058 0.5105 ;
        RECT 3.206 0.4665 3.274 0.5105 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 3.206 -0.022 3.274 0.292 ;
        RECT 2.99 -0.022 3.058 0.292 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.37 0.158 1.566 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.702 0.158 0.898 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1975 0.25 0.2415 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.206 0.158 3.274 0.202 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.028 0.428 2.32 0.472 ;
    LAYER m1 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.35 0.338 1.694 0.382 ;
      RECT 1.37 0.248 1.91 0.292 ;
      RECT 2.234 0.338 2.302 0.472 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 2.126 0.158 2.194 0.562 ;
      RECT 2.882 0.068 2.95 0.562 ;
    LAYER v1 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.05 0.428 1.11 0.472 ;
    LAYER v0 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.882 0.4665 2.95 0.5105 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.666 0.4665 2.734 0.5105 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.43 2.194 0.474 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.1785 1.222 0.2225 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.439 1.006 0.483 ;
      RECT 0.94 0.178 1.004 0.222 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.248 0.938 0.292 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.006 0.518 1.242 0.562 ;
      RECT 1.222 0.428 1.438 0.472 ;
      RECT 1.694 0.338 1.762 0.472 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.302 0.338 2.666 0.382 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.194 0.158 2.342 0.202 ;
      RECT 2.342 0.158 2.41 0.292 ;
      RECT 2.41 0.248 2.774 0.292 ;
      RECT 2.774 0.068 2.842 0.292 ;
  END
END b15fpy000hn1n08x7

MACRO b15fpy000hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy000hn1n12x5 0 0 ;
  SIZE 3.564 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.338 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.4665 2.842 0.5105 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.825679 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.81 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.068 3.49 0.562 ;
        RECT 3.206 0.338 3.49 0.382 ;
        RECT 3.206 0.068 3.274 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.4665 3.274 0.5105 ;
        RECT 3.206 0.158 3.274 0.202 ;
        RECT 3.422 0.4665 3.49 0.5105 ;
        RECT 3.422 0.158 3.49 0.202 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.61777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.452 0.25 0.496 ;
        RECT 0.722 0.473 0.79 0.517 ;
        RECT 1.478 0.472 1.546 0.516 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.558 0.4665 2.626 0.5105 ;
        RECT 2.882 0.4665 2.95 0.5105 ;
        RECT 3.098 0.4665 3.166 0.5105 ;
        RECT 3.314 0.4665 3.382 0.5105 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.598 0.022 ;
        RECT 3.314 -0.022 3.382 0.292 ;
        RECT 3.098 -0.022 3.166 0.292 ;
        RECT 2.882 -0.022 2.95 0.292 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.37 0.158 1.566 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.702 0.158 0.898 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1975 0.25 0.2415 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.882 0.158 2.95 0.202 ;
        RECT 3.098 0.158 3.166 0.202 ;
        RECT 3.314 0.158 3.382 0.202 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.028 0.428 2.32 0.472 ;
    LAYER m1 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.35 0.338 1.694 0.382 ;
      RECT 1.37 0.248 1.91 0.292 ;
      RECT 2.234 0.338 2.302 0.472 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 2.126 0.158 2.194 0.562 ;
      RECT 2.99 0.068 3.058 0.562 ;
    LAYER v1 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.05 0.428 1.11 0.472 ;
    LAYER v0 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.99 0.4665 3.058 0.5105 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.666 0.4665 2.734 0.5105 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.43 2.194 0.474 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.1785 1.222 0.2225 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.439 1.006 0.483 ;
      RECT 0.94 0.178 1.004 0.222 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.248 0.938 0.292 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.006 0.518 1.242 0.562 ;
      RECT 1.222 0.428 1.438 0.472 ;
      RECT 1.694 0.338 1.762 0.472 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.302 0.338 2.666 0.382 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.194 0.158 2.342 0.202 ;
      RECT 2.342 0.158 2.41 0.292 ;
      RECT 2.41 0.248 2.774 0.292 ;
      RECT 2.774 0.068 2.842 0.292 ;
  END
END b15fpy000hn1n12x5

MACRO b15fpy000hn1n12x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy000hn1n12x7 0 0 ;
  SIZE 3.996 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.248 3.274 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.2705 3.274 0.3145 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.222 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.068 3.922 0.562 ;
        RECT 3.638 0.338 3.922 0.382 ;
        RECT 3.638 0.068 3.706 0.562 ;
      LAYER v0 ;
        RECT 3.638 0.448 3.706 0.492 ;
        RECT 3.638 0.1525 3.706 0.1965 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 3.854 0.1525 3.922 0.1965 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.13925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.338 3.382 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.472 0.25 0.516 ;
        RECT 0.722 0.4725 0.79 0.5165 ;
        RECT 1.154 0.4725 1.222 0.5165 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 3.746 0.448 3.814 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.03 0.022 ;
        RECT 3.746 -0.022 3.814 0.292 ;
        RECT 3.314 0.248 3.598 0.292 ;
        RECT 3.53 -0.022 3.598 0.292 ;
        RECT 3.314 0.158 3.382 0.292 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.702 0.158 0.898 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1905 0.25 0.2345 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.882 0.048 2.95 0.092 ;
        RECT 3.316 0.178 3.38 0.222 ;
        RECT 3.53 0.1525 3.598 0.1965 ;
        RECT 3.746 0.1525 3.814 0.1965 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.352 0.428 2.86 0.472 ;
    LAYER m1 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.694 0.518 1.91 0.562 ;
      RECT 1.802 0.248 1.87 0.472 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.774 0.248 2.842 0.472 ;
      RECT 2.45 0.248 2.518 0.472 ;
      RECT 2.558 0.158 2.626 0.562 ;
    LAYER v1 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.454 0.428 2.514 0.472 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.374 0.428 1.434 0.472 ;
    LAYER v0 ;
      RECT 3.206 0.068 3.274 0.112 ;
      RECT 3.098 0.406 3.166 0.45 ;
      RECT 3.1 0.178 3.164 0.222 ;
      RECT 2.774 0.338 2.842 0.382 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.558 0.43 2.626 0.474 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 1.802 0.3155 1.87 0.3595 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.408 1.762 0.452 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.248 1.694 0.292 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.566 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 1.978 0.338 2.302 0.382 ;
      RECT 2.194 0.248 2.342 0.292 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.842 0.248 3.098 0.292 ;
      RECT 3.098 0.158 3.166 0.472 ;
      RECT 2.626 0.158 2.99 0.202 ;
      RECT 2.99 0.068 3.058 0.202 ;
      RECT 3.058 0.068 3.382 0.112 ;
  END
END b15fpy000hn1n12x7

MACRO b15fpy000hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy000hn1n16x5 0 0 ;
  SIZE 4.212 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.248 3.166 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.2705 3.166 0.3145 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.222 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.158 4.03 0.562 ;
        RECT 3.746 0.338 4.03 0.382 ;
        RECT 3.746 0.158 3.814 0.562 ;
      LAYER v0 ;
        RECT 3.746 0.448 3.814 0.492 ;
        RECT 3.746 0.178 3.814 0.222 ;
        RECT 3.962 0.448 4.03 0.492 ;
        RECT 3.962 0.178 4.03 0.222 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.13925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.246 0.652 ;
        RECT 4.07 0.428 4.138 0.652 ;
        RECT 3.854 0.428 3.922 0.652 ;
        RECT 3.638 0.428 3.706 0.652 ;
        RECT 3.422 0.338 3.49 0.652 ;
        RECT 2.99 0.338 3.058 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.472 0.25 0.516 ;
        RECT 0.722 0.4725 0.79 0.5165 ;
        RECT 1.154 0.4725 1.222 0.5165 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.99 0.428 3.058 0.472 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.638 0.448 3.706 0.492 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 4.07 0.448 4.138 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.246 0.022 ;
        RECT 4.07 -0.022 4.138 0.292 ;
        RECT 3.854 -0.022 3.922 0.292 ;
        RECT 3.638 -0.022 3.706 0.292 ;
        RECT 3.422 -0.022 3.49 0.292 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.342 -0.022 2.41 0.292 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.702 0.158 0.898 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1905 0.25 0.2345 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 2.126 0.143 2.194 0.187 ;
        RECT 2.342 0.143 2.41 0.187 ;
        RECT 2.99 0.048 3.058 0.092 ;
        RECT 3.422 0.178 3.49 0.222 ;
        RECT 3.638 0.178 3.706 0.222 ;
        RECT 3.854 0.178 3.922 0.222 ;
        RECT 4.07 0.178 4.138 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.352 0.428 3.292 0.472 ;
    LAYER m1 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 2.018 0.158 2.086 0.382 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 2.666 0.158 2.734 0.562 ;
      RECT 2.558 0.248 2.626 0.472 ;
      RECT 2.882 0.248 2.95 0.472 ;
      RECT 3.206 0.158 3.274 0.472 ;
      RECT 3.53 0.158 3.598 0.562 ;
    LAYER v1 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.374 0.428 1.434 0.472 ;
    LAYER v0 ;
      RECT 3.53 0.178 3.598 0.222 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.314 0.178 3.382 0.222 ;
      RECT 3.206 0.178 3.274 0.222 ;
      RECT 3.206 0.406 3.274 0.45 ;
      RECT 2.882 0.3155 2.95 0.3595 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.666 0.43 2.734 0.474 ;
      RECT 2.558 0.338 2.626 0.382 ;
      RECT 2.45 0.143 2.518 0.187 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.234 0.143 2.302 0.187 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.802 0.157 1.87 0.201 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.694 0.157 1.762 0.201 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.248 1.262 0.292 ;
      RECT 1.262 0.068 1.33 0.292 ;
      RECT 1.33 0.068 1.694 0.112 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 2.086 0.338 2.234 0.382 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.302 0.338 2.45 0.382 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 2.734 0.158 3.098 0.202 ;
      RECT 3.098 0.068 3.166 0.202 ;
      RECT 3.166 0.068 3.314 0.112 ;
      RECT 3.314 0.068 3.382 0.292 ;
  END
END b15fpy000hn1n16x5

MACRO b15fpy000hn1n16x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy000hn1n16x7 0 0 ;
  SIZE 5.076 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.30375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.30375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.158 4.138 0.472 ;
      LAYER v0 ;
        RECT 4.07 0.408 4.138 0.452 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.242 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.826 0.068 4.894 0.562 ;
        RECT 4.61 0.248 4.894 0.292 ;
        RECT 4.61 0.068 4.678 0.562 ;
      LAYER v0 ;
        RECT 4.61 0.43 4.678 0.474 ;
        RECT 4.61 0.138 4.678 0.182 ;
        RECT 4.826 0.43 4.894 0.474 ;
        RECT 4.826 0.138 4.894 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 2.4594445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.11 0.652 ;
        RECT 4.934 0.338 5.002 0.652 ;
        RECT 4.718 0.338 4.786 0.652 ;
        RECT 4.502 0.338 4.57 0.652 ;
        RECT 4.286 0.338 4.354 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.472 0.25 0.516 ;
        RECT 0.722 0.4725 0.79 0.5165 ;
        RECT 1.154 0.4725 1.222 0.5165 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 3.422 0.478 3.49 0.522 ;
        RECT 3.746 0.448 3.814 0.492 ;
        RECT 4.286 0.43 4.354 0.474 ;
        RECT 4.502 0.43 4.57 0.474 ;
        RECT 4.718 0.43 4.786 0.474 ;
        RECT 4.934 0.43 5.002 0.474 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.11 0.022 ;
        RECT 4.934 -0.022 5.002 0.202 ;
        RECT 4.718 -0.022 4.786 0.202 ;
        RECT 4.502 -0.022 4.57 0.292 ;
        RECT 4.286 -0.022 4.354 0.202 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.046 0.158 1.242 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.702 0.158 0.898 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1905 0.25 0.2345 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 3.424 0.138 3.488 0.182 ;
        RECT 3.748 0.048 3.812 0.092 ;
        RECT 4.286 0.138 4.354 0.182 ;
        RECT 4.502 0.138 4.57 0.182 ;
        RECT 4.718 0.138 4.786 0.182 ;
        RECT 4.934 0.138 5.002 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.46 0.428 4.048 0.472 ;
    LAYER m1 ;
      RECT 1.478 0.068 1.546 0.472 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.774 0.248 2.842 0.472 ;
      RECT 2.666 0.158 2.882 0.202 ;
      RECT 3.206 0.248 3.274 0.472 ;
      RECT 3.53 0.428 3.598 0.562 ;
      RECT 3.962 0.158 4.03 0.472 ;
      RECT 3.402 0.338 3.854 0.382 ;
    LAYER v1 ;
      RECT 3.966 0.428 4.026 0.472 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
    LAYER v0 ;
      RECT 4.394 0.138 4.462 0.182 ;
      RECT 4.394 0.43 4.462 0.474 ;
      RECT 4.07 0.068 4.138 0.112 ;
      RECT 3.962 0.178 4.03 0.222 ;
      RECT 3.962 0.408 4.03 0.452 ;
      RECT 3.53 0.478 3.598 0.522 ;
      RECT 3.422 0.338 3.49 0.382 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.206 0.338 3.274 0.382 ;
      RECT 3.098 0.498 3.166 0.542 ;
      RECT 2.99 0.178 3.058 0.222 ;
      RECT 2.99 0.408 3.058 0.452 ;
      RECT 2.882 0.408 2.95 0.452 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.3155 2.842 0.3595 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.4385 1.978 0.4825 ;
      RECT 1.694 0.4135 1.762 0.4575 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.586 0.3135 1.654 0.3575 ;
      RECT 1.37 0.422 1.438 0.466 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.438 0.518 1.694 0.562 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.546 0.068 1.762 0.112 ;
      RECT 1.654 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 1.978 0.158 2.234 0.202 ;
      RECT 2.234 0.158 2.302 0.382 ;
      RECT 2.302 0.338 2.538 0.382 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.194 0.428 2.666 0.472 ;
      RECT 2.518 0.248 2.666 0.292 ;
      RECT 2.666 0.248 2.734 0.562 ;
      RECT 2.734 0.518 2.99 0.562 ;
      RECT 2.99 0.158 3.058 0.562 ;
      RECT 2.882 0.068 2.95 0.472 ;
      RECT 2.95 0.068 3.098 0.112 ;
      RECT 3.098 0.068 3.166 0.562 ;
      RECT 3.166 0.158 3.314 0.202 ;
      RECT 3.314 0.158 3.382 0.292 ;
      RECT 3.382 0.248 3.854 0.292 ;
      RECT 3.854 0.068 3.922 0.292 ;
      RECT 3.922 0.068 4.246 0.112 ;
      RECT 3.854 0.338 3.922 0.562 ;
      RECT 3.922 0.518 4.178 0.562 ;
      RECT 4.178 0.248 4.246 0.562 ;
      RECT 4.246 0.248 4.394 0.292 ;
      RECT 4.394 0.068 4.462 0.562 ;
  END
END b15fpy000hn1n16x7

MACRO b15fpy010hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy010hn1n02x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.248 2.41 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.138 2.734 0.182 ;
    END
  END o1
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.558 0.428 2.626 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.074 0.158 0.27 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.338 2.32 0.382 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.694 0.518 1.91 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.45 0.068 2.518 0.562 ;
    LAYER v1 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
    LAYER v0 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.138 2.302 0.182 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.223 1.654 0.267 ;
      RECT 1.586 0.469 1.654 0.513 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.155 1.222 0.199 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 1.046 0.155 1.114 0.199 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.508 0.228 0.572 0.272 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.378 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.654 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.91 0.068 1.978 0.562 ;
  END
END b15fpy010hn1n02x5

MACRO b15fpy010hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy010hn1n03x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.248 2.41 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.138 2.734 0.182 ;
    END
  END o1
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.558 0.428 2.626 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.074 0.158 0.27 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.338 2.32 0.382 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.694 0.518 1.91 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.45 0.068 2.518 0.562 ;
    LAYER v1 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
    LAYER v0 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.138 2.302 0.182 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.223 1.654 0.267 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.155 1.222 0.199 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 1.046 0.155 1.114 0.199 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.508 0.228 0.572 0.272 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.378 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.654 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.91 0.068 1.978 0.562 ;
  END
END b15fpy010hn1n03x5

MACRO b15fpy010hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy010hn1n04x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.248 2.41 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.4085 2.734 0.4525 ;
        RECT 2.666 0.138 2.734 0.182 ;
    END
  END o1
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.558 0.4085 2.626 0.4525 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.074 0.158 0.27 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.338 2.32 0.382 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.694 0.518 1.91 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.45 0.068 2.518 0.562 ;
    LAYER v1 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
    LAYER v0 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.4085 2.518 0.4525 ;
      RECT 2.234 0.138 2.302 0.182 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.223 1.654 0.267 ;
      RECT 1.586 0.469 1.654 0.513 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.155 1.222 0.199 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 1.046 0.155 1.114 0.199 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.508 0.228 0.572 0.272 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.378 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.654 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.91 0.068 1.978 0.562 ;
  END
END b15fpy010hn1n04x5

MACRO b15fpy010hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy010hn1n06x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.158 2.518 0.472 ;
      LAYER v0 ;
        RECT 2.45 0.338 2.518 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.068 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.774 0.138 2.842 0.182 ;
    END
  END o1
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.882 0.448 2.95 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.223 0.25 0.267 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.586 0.192 1.654 0.236 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.666 0.138 2.734 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.338 2.428 0.382 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.802 0.248 1.87 0.472 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.558 0.068 2.626 0.562 ;
    LAYER v1 ;
      RECT 2.346 0.338 2.406 0.382 ;
      RECT 2.13 0.338 2.19 0.382 ;
      RECT 1.806 0.338 1.866 0.382 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
    LAYER v0 ;
      RECT 2.558 0.138 2.626 0.182 ;
      RECT 2.558 0.448 2.626 0.492 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.694 0.192 1.762 0.236 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.155 1.222 0.199 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 1.046 0.155 1.114 0.199 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.508 0.228 0.572 0.272 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.378 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.438 0.338 1.694 0.382 ;
      RECT 1.694 0.158 1.762 0.562 ;
      RECT 1.978 0.338 2.018 0.382 ;
      RECT 2.018 0.068 2.086 0.382 ;
  END
END b15fpy010hn1n06x5

MACRO b15fpy010hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy010hn1n08x5 0 0 ;
  SIZE 3.564 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 5.561111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 5.561111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.382 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER m2 ;
        RECT 0.04 0.338 0.592 0.382 ;
      LAYER v1 ;
        RECT 0.186 0.338 0.246 0.382 ;
        RECT 0.51 0.338 0.57 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END ssb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.158 3.382 0.382 ;
        RECT 3.206 0.158 3.382 0.202 ;
        RECT 3.206 0.068 3.274 0.202 ;
      LAYER v0 ;
        RECT 3.314 0.2705 3.382 0.3145 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.338 3.274 0.562 ;
        RECT 2.99 0.338 3.274 0.382 ;
        RECT 2.99 0.068 3.058 0.562 ;
      LAYER v0 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 2.99 0.113 3.058 0.157 ;
        RECT 3.206 0.448 3.274 0.492 ;
    END
  END o1
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END si
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.4285 0.358 0.4725 ;
        RECT 0.83 0.4285 0.898 0.4725 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.314 0.448 3.382 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.598 0.022 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.159 0.358 0.203 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.478 0.113 1.546 0.157 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.666 0.113 2.734 0.157 ;
        RECT 3.098 0.113 3.166 0.157 ;
        RECT 3.314 0.048 3.382 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.136 0.338 3.524 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.182 0.158 0.25 0.382 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 1.154 0.338 1.222 0.472 ;
      RECT 1.262 0.068 1.33 0.472 ;
      RECT 1.37 0.248 1.802 0.292 ;
      RECT 1.478 0.338 1.762 0.382 ;
      RECT 1.586 0.158 2.018 0.202 ;
      RECT 2.234 0.248 2.302 0.382 ;
      RECT 2.126 0.518 2.45 0.562 ;
      RECT 2.558 0.248 2.626 0.382 ;
      RECT 2.774 0.068 2.842 0.562 ;
      RECT 3.422 0.068 3.49 0.562 ;
    LAYER v1 ;
      RECT 3.426 0.338 3.486 0.382 ;
      RECT 2.562 0.338 2.622 0.382 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
    LAYER v0 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.422 0.448 3.49 0.492 ;
      RECT 2.774 0.113 2.842 0.157 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.558 0.2705 2.626 0.3145 ;
      RECT 2.45 0.178 2.518 0.222 ;
      RECT 2.342 0.2705 2.41 0.3145 ;
      RECT 2.234 0.2705 2.302 0.3145 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.126 0.383 2.194 0.427 ;
      RECT 2.128 0.178 2.192 0.222 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.138 1.33 0.182 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.154 0.138 1.222 0.182 ;
      RECT 1.154 0.38 1.222 0.424 ;
      RECT 0.614 0.4295 0.682 0.4735 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.074 0.159 0.142 0.203 ;
      RECT 0.074 0.4285 0.142 0.4725 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.158 0.938 0.202 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.248 1.046 0.292 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.114 0.518 1.35 0.562 ;
      RECT 1.33 0.428 1.654 0.472 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.87 0.248 2.126 0.292 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 2.018 0.068 2.086 0.202 ;
      RECT 2.086 0.068 2.342 0.112 ;
      RECT 2.342 0.068 2.41 0.382 ;
      RECT 2.45 0.158 2.518 0.562 ;
  END
END b15fpy010hn1n08x5

MACRO b15fpy010hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy010hn1n12x5 0 0 ;
  SIZE 4.212 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 8.845 LAYER m1 ;
      ANTENNAMAXAREACAR 13.076111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0153 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 5.561111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.382 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER m2 ;
        RECT 0.164 0.338 1.024 0.382 ;
      LAYER v1 ;
        RECT 0.186 0.338 0.246 0.382 ;
        RECT 0.51 0.338 0.57 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END ssb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5544445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.299 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.068 3.49 0.292 ;
      LAYER v0 ;
        RECT 3.422 0.113 3.49 0.157 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.07166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.63285725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 1.33 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.154 0.248 1.222 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.068 4.138 0.562 ;
        RECT 3.854 0.248 4.138 0.292 ;
        RECT 3.854 0.068 3.922 0.562 ;
      LAYER v0 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 3.854 0.113 3.922 0.157 ;
        RECT 4.07 0.448 4.138 0.492 ;
        RECT 4.07 0.113 4.138 0.157 ;
    END
  END o1
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END si
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.246 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.206 0.518 3.274 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.4285 0.358 0.4725 ;
        RECT 0.83 0.468 0.898 0.512 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 3.206 0.538 3.274 0.582 ;
        RECT 3.53 0.538 3.598 0.582 ;
        RECT 3.746 0.538 3.814 0.582 ;
        RECT 3.962 0.448 4.03 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.246 0.022 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.53 -0.022 3.598 0.292 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.159 0.358 0.203 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.262 0.1135 1.33 0.1575 ;
        RECT 1.91 0.138 1.978 0.182 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 3.206 0.113 3.274 0.157 ;
        RECT 3.53 0.228 3.598 0.272 ;
        RECT 3.746 0.113 3.814 0.157 ;
        RECT 3.962 0.113 4.03 0.157 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.46 0.338 3.724 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.182 0.158 0.25 0.382 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 1.478 0.248 1.546 0.382 ;
      RECT 1.694 0.158 1.762 0.562 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.91 0.338 2.194 0.382 ;
      RECT 2.558 0.248 2.626 0.382 ;
      RECT 2.234 0.248 2.302 0.562 ;
      RECT 3.314 0.068 3.382 0.382 ;
      RECT 3.098 0.248 3.166 0.382 ;
      RECT 2.774 0.068 2.842 0.292 ;
      RECT 3.638 0.068 3.706 0.382 ;
    LAYER v1 ;
      RECT 3.642 0.338 3.702 0.382 ;
      RECT 3.102 0.338 3.162 0.382 ;
      RECT 2.562 0.338 2.622 0.382 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.482 0.338 1.542 0.382 ;
    LAYER v0 ;
      RECT 3.746 0.293 3.814 0.337 ;
      RECT 3.638 0.113 3.706 0.157 ;
      RECT 3.422 0.338 3.49 0.382 ;
      RECT 3.314 0.113 3.382 0.157 ;
      RECT 3.206 0.2705 3.274 0.3145 ;
      RECT 3.098 0.2705 3.166 0.3145 ;
      RECT 2.99 0.1805 3.058 0.2245 ;
      RECT 2.882 0.1805 2.95 0.2245 ;
      RECT 2.882 0.518 2.95 0.562 ;
      RECT 2.774 0.1805 2.842 0.2245 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.1805 2.734 0.2245 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.558 0.2705 2.626 0.3145 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.56 0.088 2.624 0.132 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.694 0.178 1.762 0.222 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.37 0.197 1.438 0.241 ;
      RECT 1.046 0.4335 1.114 0.4775 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.074 0.159 0.142 0.203 ;
      RECT 0.074 0.4285 0.142 0.4725 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.518 1.654 0.562 ;
      RECT 1.762 0.518 2.086 0.562 ;
      RECT 1.438 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.472 ;
      RECT 1.87 0.248 2.126 0.292 ;
      RECT 2.126 0.158 2.194 0.292 ;
      RECT 2.194 0.158 2.558 0.202 ;
      RECT 2.558 0.068 2.626 0.202 ;
      RECT 2.302 0.248 2.45 0.292 ;
      RECT 2.45 0.248 2.518 0.472 ;
      RECT 2.518 0.428 2.666 0.472 ;
      RECT 2.666 0.158 2.734 0.472 ;
      RECT 2.734 0.428 2.882 0.472 ;
      RECT 2.882 0.158 2.95 0.472 ;
      RECT 3.382 0.338 3.598 0.382 ;
      RECT 2.558 0.518 2.99 0.562 ;
      RECT 2.842 0.068 2.99 0.112 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.058 0.428 3.206 0.472 ;
      RECT 3.206 0.248 3.274 0.472 ;
      RECT 3.274 0.428 3.746 0.472 ;
      RECT 3.746 0.248 3.814 0.472 ;
  END
END b15fpy010hn1n12x5

MACRO b15fpy010hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy010hn1n16x5 0 0 ;
  SIZE 4.86 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 6.565 LAYER m1 ;
      ANTENNAMAXAREACAR 10.796111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
      ANTENNAMAXAREACAR 5.561111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.382 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER m2 ;
        RECT 0.164 0.248 0.592 0.292 ;
      LAYER v1 ;
        RECT 0.186 0.248 0.246 0.292 ;
        RECT 0.51 0.248 0.57 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END ssb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.13222225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.919 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.068 4.03 0.382 ;
      LAYER v0 ;
        RECT 3.962 0.088 4.03 0.132 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.318125 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.318125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.202 ;
      LAYER v0 ;
        RECT 1.046 0.133 1.114 0.177 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.068 4.678 0.562 ;
        RECT 4.394 0.338 4.678 0.382 ;
        RECT 4.394 0.068 4.462 0.562 ;
      LAYER v0 ;
        RECT 4.394 0.428 4.462 0.472 ;
        RECT 4.394 0.138 4.462 0.182 ;
        RECT 4.61 0.428 4.678 0.472 ;
        RECT 4.61 0.138 4.678 0.182 ;
    END
  END o1
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END si
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.894 0.652 ;
        RECT 4.718 0.518 4.786 0.652 ;
        RECT 4.502 0.518 4.57 0.652 ;
        RECT 4.286 0.518 4.354 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.4285 0.358 0.4725 ;
        RECT 1.154 0.538 1.222 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 4.07 0.538 4.138 0.582 ;
        RECT 4.286 0.538 4.354 0.582 ;
        RECT 4.504 0.538 4.568 0.582 ;
        RECT 4.72 0.538 4.784 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.894 0.022 ;
        RECT 4.718 -0.022 4.786 0.202 ;
        RECT 4.502 -0.022 4.57 0.202 ;
        RECT 4.286 -0.022 4.354 0.202 ;
        RECT 4.07 -0.022 4.138 0.292 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.159 0.358 0.203 ;
        RECT 1.154 0.133 1.222 0.177 ;
        RECT 1.37 0.133 1.438 0.177 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 3.746 0.138 3.814 0.182 ;
        RECT 4.07 0.223 4.138 0.267 ;
        RECT 4.286 0.138 4.354 0.182 ;
        RECT 4.502 0.138 4.57 0.182 ;
        RECT 4.718 0.138 4.786 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.46 0.248 4.264 0.292 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.182 0.158 0.25 0.382 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.398 0.158 0.614 0.202 ;
      RECT 0.722 0.428 1.438 0.472 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 2.126 0.248 2.194 0.382 ;
      RECT 3.098 0.248 3.166 0.382 ;
      RECT 2.342 0.338 2.882 0.382 ;
      RECT 3.314 0.068 3.382 0.292 ;
      RECT 3.638 0.248 3.706 0.382 ;
      RECT 4.178 0.068 4.246 0.382 ;
    LAYER v1 ;
      RECT 4.182 0.248 4.242 0.292 ;
      RECT 3.642 0.248 3.702 0.292 ;
      RECT 3.102 0.248 3.162 0.292 ;
      RECT 2.13 0.248 2.19 0.292 ;
      RECT 1.482 0.248 1.542 0.292 ;
    LAYER v0 ;
      RECT 4.286 0.293 4.354 0.337 ;
      RECT 4.178 0.138 4.246 0.182 ;
      RECT 3.746 0.293 3.814 0.337 ;
      RECT 3.638 0.293 3.706 0.337 ;
      RECT 3.53 0.178 3.598 0.222 ;
      RECT 3.422 0.178 3.49 0.222 ;
      RECT 3.422 0.518 3.49 0.562 ;
      RECT 3.314 0.178 3.382 0.222 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 3.206 0.178 3.274 0.222 ;
      RECT 3.206 0.518 3.274 0.562 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 3.098 0.293 3.166 0.337 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.882 0.248 2.95 0.292 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.126 0.293 2.194 0.337 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.133 1.87 0.177 ;
      RECT 1.694 0.133 1.762 0.177 ;
      RECT 1.588 0.448 1.652 0.492 ;
      RECT 1.478 0.133 1.546 0.177 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.262 0.133 1.33 0.177 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.139 0.898 0.183 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.074 0.159 0.142 0.203 ;
      RECT 0.074 0.4285 0.142 0.4725 ;
    LAYER m1 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 0.898 0.248 1.262 0.292 ;
      RECT 1.262 0.068 1.33 0.292 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.338 1.694 0.382 ;
      RECT 1.694 0.068 1.762 0.382 ;
      RECT 1.654 0.518 1.802 0.562 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.87 0.518 2.194 0.562 ;
      RECT 1.978 0.428 2.234 0.472 ;
      RECT 2.234 0.248 2.302 0.472 ;
      RECT 2.302 0.248 2.99 0.292 ;
      RECT 2.99 0.068 3.058 0.292 ;
      RECT 3.058 0.068 3.274 0.112 ;
      RECT 2.882 0.338 2.95 0.472 ;
      RECT 2.95 0.428 3.206 0.472 ;
      RECT 3.206 0.158 3.274 0.472 ;
      RECT 3.274 0.428 3.422 0.472 ;
      RECT 3.422 0.158 3.49 0.472 ;
      RECT 3.098 0.518 3.53 0.562 ;
      RECT 3.382 0.068 3.53 0.112 ;
      RECT 3.53 0.068 3.598 0.562 ;
      RECT 3.598 0.428 3.746 0.472 ;
      RECT 3.746 0.248 3.814 0.472 ;
      RECT 3.814 0.428 4.286 0.472 ;
      RECT 4.286 0.248 4.354 0.472 ;
  END
END b15fpy010hn1n16x5

MACRO b15fpy040hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy040hn1n02x5 0 0 ;
  SIZE 3.78 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.158 3.382 0.382 ;
      LAYER v0 ;
        RECT 3.314 0.248 3.382 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.088 0.79 0.132 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.068 3.706 0.472 ;
      LAYER v0 ;
        RECT 3.638 0.383 3.706 0.427 ;
        RECT 3.638 0.1675 3.706 0.2115 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.814 0.652 ;
        RECT 3.53 0.338 3.598 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.83 0.428 1.026 0.472 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.53 0.383 3.598 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.814 0.022 ;
        RECT 3.53 -0.022 3.598 0.292 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 1.782 0.248 1.978 0.292 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.938 0.1135 1.006 0.1575 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.45 0.114 2.518 0.158 ;
        RECT 3.098 0.138 3.166 0.182 ;
        RECT 3.53 0.1675 3.598 0.2115 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.518 1.472 0.562 ;
      RECT 1.552 0.518 3.508 0.562 ;
    LAYER m1 ;
      RECT 1.026 0.518 1.262 0.562 ;
      RECT 0.506 0.518 0.722 0.562 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 2.126 0.068 2.194 0.472 ;
      RECT 2.43 0.248 2.558 0.292 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 2.774 0.248 2.842 0.472 ;
      RECT 2.558 0.518 2.882 0.562 ;
      RECT 3.422 0.068 3.49 0.562 ;
    LAYER v1 ;
      RECT 3.426 0.518 3.486 0.562 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 0.294 0.518 0.354 0.562 ;
    LAYER v0 ;
      RECT 3.422 0.1675 3.49 0.2115 ;
      RECT 3.422 0.383 3.49 0.427 ;
      RECT 3.206 0.138 3.274 0.182 ;
      RECT 3.206 0.448 3.274 0.492 ;
      RECT 2.99 0.248 3.058 0.292 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.774 0.3685 2.842 0.4125 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.558 0.114 2.626 0.158 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.386 2.194 0.43 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.156 0.408 1.22 0.452 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.228 0.574 0.272 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.338 1.154 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.222 0.158 1.438 0.202 ;
      RECT 1.438 0.248 1.586 0.292 ;
      RECT 1.586 0.068 1.654 0.292 ;
      RECT 1.654 0.068 1.782 0.112 ;
      RECT 2.194 0.068 2.322 0.112 ;
      RECT 2.558 0.068 2.626 0.292 ;
      RECT 1.762 0.338 2.018 0.382 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 2.086 0.518 2.234 0.562 ;
      RECT 2.234 0.158 2.302 0.562 ;
      RECT 2.302 0.338 2.666 0.382 ;
      RECT 2.666 0.158 2.734 0.382 ;
      RECT 2.842 0.248 2.882 0.292 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 2.95 0.338 2.99 0.382 ;
      RECT 2.99 0.158 3.058 0.382 ;
      RECT 3.058 0.338 3.206 0.382 ;
      RECT 3.206 0.068 3.274 0.562 ;
  END
END b15fpy040hn1n02x5

MACRO b15fpy040hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy040hn1n03x5 0 0 ;
  SIZE 3.78 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.158 3.382 0.382 ;
      LAYER v0 ;
        RECT 3.314 0.248 3.382 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.088 0.79 0.132 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.068 3.706 0.472 ;
      LAYER v0 ;
        RECT 3.638 0.383 3.706 0.427 ;
        RECT 3.638 0.1675 3.706 0.2115 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.814 0.652 ;
        RECT 3.53 0.338 3.598 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.83 0.428 1.026 0.472 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.53 0.383 3.598 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.814 0.022 ;
        RECT 3.53 -0.022 3.598 0.292 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 1.782 0.248 1.978 0.292 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.938 0.1135 1.006 0.1575 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.45 0.114 2.518 0.158 ;
        RECT 3.098 0.138 3.166 0.182 ;
        RECT 3.53 0.1675 3.598 0.2115 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.518 1.472 0.562 ;
      RECT 1.552 0.518 3.508 0.562 ;
    LAYER m1 ;
      RECT 1.026 0.518 1.262 0.562 ;
      RECT 0.506 0.518 0.722 0.562 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 2.126 0.068 2.194 0.472 ;
      RECT 2.43 0.248 2.558 0.292 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 2.774 0.248 2.842 0.472 ;
      RECT 2.558 0.518 2.882 0.562 ;
      RECT 3.422 0.068 3.49 0.562 ;
    LAYER v1 ;
      RECT 3.426 0.518 3.486 0.562 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 0.294 0.518 0.354 0.562 ;
    LAYER v0 ;
      RECT 3.422 0.1675 3.49 0.2115 ;
      RECT 3.422 0.383 3.49 0.427 ;
      RECT 3.206 0.138 3.274 0.182 ;
      RECT 3.206 0.448 3.274 0.492 ;
      RECT 2.99 0.248 3.058 0.292 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.774 0.3685 2.842 0.4125 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.558 0.114 2.626 0.158 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.386 2.194 0.43 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.156 0.408 1.22 0.452 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.228 0.574 0.272 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.338 1.154 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.222 0.158 1.438 0.202 ;
      RECT 1.438 0.248 1.586 0.292 ;
      RECT 1.586 0.068 1.654 0.292 ;
      RECT 1.654 0.068 1.782 0.112 ;
      RECT 2.194 0.068 2.322 0.112 ;
      RECT 2.558 0.068 2.626 0.292 ;
      RECT 1.762 0.338 2.018 0.382 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 2.086 0.518 2.234 0.562 ;
      RECT 2.234 0.158 2.302 0.562 ;
      RECT 2.302 0.338 2.666 0.382 ;
      RECT 2.666 0.158 2.734 0.382 ;
      RECT 2.842 0.248 2.882 0.292 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 2.95 0.338 2.99 0.382 ;
      RECT 2.99 0.158 3.058 0.382 ;
      RECT 3.058 0.338 3.206 0.382 ;
      RECT 3.206 0.068 3.274 0.562 ;
  END
END b15fpy040hn1n03x5

MACRO b15fpy040hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy040hn1n04x5 0 0 ;
  SIZE 3.78 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.158 3.382 0.382 ;
      LAYER v0 ;
        RECT 3.314 0.248 3.382 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.088 0.79 0.132 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.068 3.706 0.472 ;
      LAYER v0 ;
        RECT 3.638 0.383 3.706 0.427 ;
        RECT 3.638 0.1675 3.706 0.2115 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.814 0.652 ;
        RECT 3.53 0.338 3.598 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.83 0.428 1.026 0.472 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.53 0.383 3.598 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.814 0.022 ;
        RECT 3.53 -0.022 3.598 0.292 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 1.782 0.248 1.978 0.292 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.938 0.1135 1.006 0.1575 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.45 0.114 2.518 0.158 ;
        RECT 3.098 0.138 3.166 0.182 ;
        RECT 3.53 0.1675 3.598 0.2115 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.518 1.472 0.562 ;
      RECT 1.552 0.518 3.508 0.562 ;
    LAYER m1 ;
      RECT 1.026 0.518 1.262 0.562 ;
      RECT 0.506 0.518 0.722 0.562 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 2.126 0.068 2.194 0.472 ;
      RECT 2.43 0.248 2.558 0.292 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 2.774 0.248 2.842 0.472 ;
      RECT 2.558 0.518 2.882 0.562 ;
      RECT 3.422 0.068 3.49 0.562 ;
    LAYER v1 ;
      RECT 3.426 0.518 3.486 0.562 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 0.294 0.518 0.354 0.562 ;
    LAYER v0 ;
      RECT 3.422 0.1675 3.49 0.2115 ;
      RECT 3.422 0.383 3.49 0.427 ;
      RECT 3.206 0.138 3.274 0.182 ;
      RECT 3.206 0.448 3.274 0.492 ;
      RECT 2.99 0.248 3.058 0.292 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.774 0.3685 2.842 0.4125 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.558 0.114 2.626 0.158 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.386 2.194 0.43 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.156 0.408 1.22 0.452 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.228 0.574 0.272 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.338 1.154 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.222 0.158 1.438 0.202 ;
      RECT 1.438 0.248 1.586 0.292 ;
      RECT 1.586 0.068 1.654 0.292 ;
      RECT 1.654 0.068 1.782 0.112 ;
      RECT 2.194 0.068 2.322 0.112 ;
      RECT 2.558 0.068 2.626 0.292 ;
      RECT 1.762 0.338 2.018 0.382 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 2.086 0.518 2.234 0.562 ;
      RECT 2.234 0.158 2.302 0.562 ;
      RECT 2.302 0.338 2.666 0.382 ;
      RECT 2.666 0.158 2.734 0.382 ;
      RECT 2.842 0.248 2.882 0.292 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 2.95 0.338 2.99 0.382 ;
      RECT 2.99 0.158 3.058 0.382 ;
      RECT 3.058 0.338 3.206 0.382 ;
      RECT 3.206 0.068 3.274 0.562 ;
  END
END b15fpy040hn1n04x5

MACRO b15fpy040hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy040hn1n06x5 0 0 ;
  SIZE 4.104 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.158 3.598 0.382 ;
      LAYER v0 ;
        RECT 3.53 0.248 3.598 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.088 0.79 0.132 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.068 3.922 0.562 ;
      LAYER v0 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 3.854 0.138 3.922 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.138 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.342 0.428 2.754 0.472 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.83 0.428 1.026 0.472 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.746 0.448 3.814 0.492 ;
        RECT 3.962 0.448 4.03 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.138 0.022 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.938 0.114 1.006 0.158 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.45 0.114 2.518 0.158 ;
        RECT 2.666 0.114 2.734 0.158 ;
        RECT 3.314 0.138 3.382 0.182 ;
        RECT 3.746 0.138 3.814 0.182 ;
        RECT 3.962 0.138 4.03 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.518 1.472 0.562 ;
      RECT 1.552 0.518 3.724 0.562 ;
    LAYER m1 ;
      RECT 1.026 0.518 1.262 0.562 ;
      RECT 0.506 0.518 0.722 0.562 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 2.126 0.068 2.194 0.472 ;
      RECT 2.43 0.248 2.558 0.292 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 2.97 0.428 3.098 0.472 ;
      RECT 2.538 0.518 3.206 0.562 ;
      RECT 3.638 0.068 3.706 0.562 ;
    LAYER v1 ;
      RECT 3.642 0.518 3.702 0.562 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 0.294 0.518 0.354 0.562 ;
    LAYER v0 ;
      RECT 3.638 0.138 3.706 0.182 ;
      RECT 3.638 0.448 3.706 0.492 ;
      RECT 3.422 0.138 3.49 0.182 ;
      RECT 3.422 0.448 3.49 0.492 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 3.098 0.1425 3.166 0.1865 ;
      RECT 2.99 0.248 3.058 0.292 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.558 0.114 2.626 0.158 ;
      RECT 2.558 0.518 2.626 0.562 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.386 2.194 0.43 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.694 0.138 1.762 0.182 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.358 1.654 0.402 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.156 0.408 1.22 0.452 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.228 0.574 0.272 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.338 1.154 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.222 0.158 1.438 0.202 ;
      RECT 1.438 0.248 1.586 0.292 ;
      RECT 1.586 0.068 1.654 0.292 ;
      RECT 2.194 0.068 2.322 0.112 ;
      RECT 2.558 0.068 2.626 0.292 ;
      RECT 2.626 0.248 2.882 0.292 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 1.762 0.338 2.018 0.382 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 2.086 0.518 2.234 0.562 ;
      RECT 2.234 0.158 2.302 0.562 ;
      RECT 2.302 0.338 2.99 0.382 ;
      RECT 2.99 0.068 3.058 0.382 ;
      RECT 3.098 0.068 3.166 0.472 ;
      RECT 3.206 0.158 3.274 0.562 ;
      RECT 3.274 0.338 3.422 0.382 ;
      RECT 3.422 0.068 3.49 0.562 ;
  END
END b15fpy040hn1n06x5

MACRO b15fpy040hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy040hn1n08x5 0 0 ;
  SIZE 4.428 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.068 3.922 0.292 ;
      LAYER v0 ;
        RECT 3.854 0.088 3.922 0.132 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 2.22571425 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.1045 0.79 0.1485 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.736 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.566 0.112 ;
        RECT 1.046 0.068 1.114 0.292 ;
      LAYER v0 ;
        RECT 1.262 0.068 1.33 0.112 ;
        RECT 1.478 0.068 1.546 0.112 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.158 4.246 0.562 ;
      LAYER v0 ;
        RECT 4.178 0.472 4.246 0.516 ;
        RECT 4.178 0.1885 4.246 0.2325 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.116 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.462 0.652 ;
        RECT 4.286 0.428 4.354 0.652 ;
        RECT 4.07 0.428 4.138 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 2.666 0.428 3.078 0.472 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.99 0.428 3.058 0.472 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 4.07 0.472 4.138 0.516 ;
        RECT 4.286 0.472 4.354 0.516 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.462 0.022 ;
        RECT 4.286 -0.022 4.354 0.292 ;
        RECT 4.07 -0.022 4.138 0.292 ;
        RECT 3.638 -0.022 3.706 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.018 -0.022 2.086 0.292 ;
        RECT 1.458 0.248 1.87 0.292 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.83 0.1975 0.898 0.2415 ;
        RECT 1.478 0.248 1.546 0.292 ;
        RECT 2.018 0.2035 2.086 0.2475 ;
        RECT 2.774 0.114 2.842 0.158 ;
        RECT 2.99 0.114 3.058 0.158 ;
        RECT 3.638 0.138 3.706 0.182 ;
        RECT 4.07 0.1885 4.138 0.2325 ;
        RECT 4.286 0.1885 4.354 0.2325 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.518 1.456 0.562 ;
      RECT 1.784 0.518 3.832 0.562 ;
    LAYER m1 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 1.046 0.518 1.262 0.562 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.586 0.518 1.87 0.562 ;
      RECT 2.45 0.068 2.518 0.472 ;
      RECT 2.234 0.158 2.302 0.562 ;
      RECT 2.754 0.248 2.882 0.292 ;
      RECT 1.782 0.428 2.018 0.472 ;
      RECT 2.862 0.518 3.422 0.562 ;
      RECT 3.186 0.428 3.314 0.472 ;
      RECT 3.638 0.518 3.942 0.562 ;
    LAYER v1 ;
      RECT 3.75 0.518 3.81 0.562 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 0.51 0.518 0.57 0.562 ;
    LAYER v0 ;
      RECT 3.962 0.338 4.03 0.382 ;
      RECT 3.854 0.518 3.922 0.562 ;
      RECT 3.746 0.428 3.814 0.472 ;
      RECT 3.422 0.248 3.49 0.292 ;
      RECT 3.314 0.1535 3.382 0.1975 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.114 3.166 0.158 ;
      RECT 2.882 0.114 2.95 0.158 ;
      RECT 2.882 0.518 2.95 0.562 ;
      RECT 2.774 0.248 2.842 0.292 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.45 0.386 2.518 0.43 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.234 0.1885 2.302 0.2325 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 1.91 0.088 1.978 0.132 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.154 0.194 1.222 0.238 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.048 0.408 1.112 0.452 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.506 0.228 0.574 0.272 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.378 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.79 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.472 ;
      RECT 1.114 0.338 1.154 0.382 ;
      RECT 1.154 0.158 1.222 0.382 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.674 0.202 ;
      RECT 1.438 0.338 1.91 0.382 ;
      RECT 1.91 0.068 1.978 0.382 ;
      RECT 2.518 0.068 2.646 0.112 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 2.95 0.248 3.098 0.292 ;
      RECT 3.098 0.068 3.166 0.292 ;
      RECT 2.018 0.338 2.086 0.472 ;
      RECT 2.086 0.338 2.126 0.382 ;
      RECT 2.126 0.068 2.194 0.382 ;
      RECT 2.194 0.068 2.342 0.112 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.41 0.518 2.558 0.562 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 2.626 0.338 3.206 0.382 ;
      RECT 3.206 0.158 3.274 0.382 ;
      RECT 3.422 0.158 3.49 0.562 ;
      RECT 3.49 0.338 3.638 0.382 ;
      RECT 3.638 0.338 3.706 0.472 ;
      RECT 3.706 0.428 3.834 0.472 ;
      RECT 3.314 0.068 3.382 0.472 ;
      RECT 3.382 0.068 3.53 0.112 ;
      RECT 3.53 0.068 3.598 0.292 ;
      RECT 3.598 0.248 3.746 0.292 ;
      RECT 3.746 0.248 3.814 0.382 ;
      RECT 3.814 0.338 4.138 0.382 ;
  END
END b15fpy040hn1n08x5

MACRO b15fpy040hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy040hn1n12x5 0 0 ;
  SIZE 5.076 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.6044445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.805 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.338 4.57 0.382 ;
        RECT 4.502 0.068 4.57 0.382 ;
      LAYER v0 ;
        RECT 4.394 0.338 4.462 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.1046155 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.674 0.112 ;
        RECT 1.046 0.068 1.114 0.292 ;
      LAYER v0 ;
        RECT 1.586 0.068 1.654 0.112 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.934 0.068 5.002 0.562 ;
        RECT 4.718 0.338 5.002 0.382 ;
        RECT 4.718 0.068 4.786 0.562 ;
      LAYER v0 ;
        RECT 4.718 0.472 4.786 0.516 ;
        RECT 4.718 0.138 4.786 0.182 ;
        RECT 4.934 0.472 5.002 0.516 ;
        RECT 4.934 0.138 5.002 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.4225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.398 0.068 0.79 0.112 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.722 0.186 0.79 0.23 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.11 0.652 ;
        RECT 4.826 0.428 4.894 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 4.286 0.428 4.354 0.652 ;
        RECT 4.07 0.428 4.138 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 4.07 0.448 4.138 0.492 ;
        RECT 4.286 0.448 4.354 0.492 ;
        RECT 4.61 0.472 4.678 0.516 ;
        RECT 4.826 0.472 4.894 0.516 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.11 0.022 ;
        RECT 4.826 -0.022 4.894 0.202 ;
        RECT 4.61 -0.022 4.678 0.202 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.458 0.248 1.978 0.292 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.197 0.25 0.241 ;
        RECT 0.83 0.186 0.898 0.23 ;
        RECT 1.478 0.248 1.546 0.292 ;
        RECT 1.91 0.1645 1.978 0.2085 ;
        RECT 2.234 0.114 2.302 0.158 ;
        RECT 2.99 0.114 3.058 0.158 ;
        RECT 3.206 0.114 3.274 0.158 ;
        RECT 4.18 0.048 4.244 0.092 ;
        RECT 4.61 0.138 4.678 0.182 ;
        RECT 4.826 0.138 4.894 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.704 0.518 1.58 0.562 ;
      RECT 1.66 0.518 4.588 0.562 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.586 0.518 1.782 0.562 ;
      RECT 2.106 0.248 2.558 0.292 ;
      RECT 2.45 0.068 2.518 0.202 ;
      RECT 1.782 0.338 2.342 0.382 ;
      RECT 2.97 0.248 3.098 0.292 ;
      RECT 3.402 0.518 3.962 0.562 ;
      RECT 3.51 0.428 3.854 0.472 ;
      RECT 4.502 0.428 4.57 0.562 ;
    LAYER v1 ;
      RECT 4.506 0.518 4.566 0.562 ;
      RECT 1.698 0.518 1.758 0.562 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 0.726 0.518 0.786 0.562 ;
    LAYER v0 ;
      RECT 4.502 0.472 4.57 0.516 ;
      RECT 4.396 0.088 4.46 0.132 ;
      RECT 4.286 0.248 4.354 0.292 ;
      RECT 4.178 0.448 4.246 0.492 ;
      RECT 3.962 0.248 4.03 0.292 ;
      RECT 3.854 0.15 3.922 0.194 ;
      RECT 3.746 0.15 3.814 0.194 ;
      RECT 3.746 0.428 3.814 0.472 ;
      RECT 3.64 0.318 3.704 0.362 ;
      RECT 3.53 0.428 3.598 0.472 ;
      RECT 3.422 0.338 3.49 0.382 ;
      RECT 3.422 0.518 3.49 0.562 ;
      RECT 3.314 0.248 3.382 0.292 ;
      RECT 3.098 0.114 3.166 0.158 ;
      RECT 2.99 0.248 3.058 0.292 ;
      RECT 2.774 0.361 2.842 0.405 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.558 0.3605 2.626 0.4045 ;
      RECT 2.452 0.138 2.516 0.182 ;
      RECT 2.342 0.248 2.41 0.292 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.262 0.49 1.33 0.534 ;
      RECT 1.154 0.194 1.222 0.238 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.614 0.186 0.682 0.23 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.186 0.574 0.23 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.378 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.154 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.33 0.158 1.674 0.202 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.338 1.654 0.472 ;
      RECT 1.654 0.428 1.782 0.472 ;
      RECT 2.558 0.248 2.626 0.472 ;
      RECT 2.518 0.068 2.774 0.112 ;
      RECT 2.774 0.068 2.842 0.472 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.41 0.518 2.666 0.562 ;
      RECT 2.666 0.158 2.734 0.562 ;
      RECT 2.734 0.518 2.882 0.562 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 2.95 0.338 3.51 0.382 ;
      RECT 3.098 0.068 3.166 0.292 ;
      RECT 3.166 0.248 3.638 0.292 ;
      RECT 3.638 0.248 3.706 0.382 ;
      RECT 3.706 0.248 3.746 0.292 ;
      RECT 3.746 0.068 3.814 0.292 ;
      RECT 3.962 0.158 4.03 0.562 ;
      RECT 4.03 0.338 4.178 0.382 ;
      RECT 4.178 0.248 4.246 0.562 ;
      RECT 4.246 0.248 4.374 0.292 ;
      RECT 3.854 0.068 3.922 0.472 ;
      RECT 3.922 0.068 4.07 0.112 ;
      RECT 4.07 0.068 4.138 0.202 ;
      RECT 4.138 0.158 4.394 0.202 ;
      RECT 4.394 0.068 4.462 0.202 ;
  END
END b15fpy040hn1n12x5

MACRO b15fpy040hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy040hn1n16x5 0 0 ;
  SIZE 5.94 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33234575 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.042 0.338 5.326 0.382 ;
        RECT 5.258 0.158 5.326 0.382 ;
      LAYER v0 ;
        RECT 5.15 0.338 5.218 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 1.242 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 2.086 0.112 ;
        RECT 1.37 0.068 1.438 0.382 ;
        RECT 1.046 0.158 1.438 0.202 ;
        RECT 1.046 0.068 1.114 0.202 ;
        RECT 0.83 0.068 1.114 0.112 ;
        RECT 0.83 0.068 0.898 0.202 ;
      LAYER v0 ;
        RECT 0.832 0.138 0.896 0.182 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.91 0.068 1.978 0.112 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.69 0.158 5.758 0.562 ;
        RECT 5.474 0.338 5.758 0.382 ;
        RECT 5.474 0.158 5.542 0.562 ;
      LAYER v0 ;
        RECT 5.474 0.472 5.542 0.516 ;
        RECT 5.474 0.1885 5.542 0.2325 ;
        RECT 5.69 0.472 5.758 0.516 ;
        RECT 5.69 0.1885 5.758 0.2325 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.974 0.652 ;
        RECT 5.798 0.428 5.866 0.652 ;
        RECT 5.582 0.428 5.65 0.652 ;
        RECT 5.366 0.428 5.434 0.652 ;
        RECT 5.042 0.428 5.11 0.652 ;
        RECT 4.826 0.428 4.894 0.652 ;
        RECT 3.834 0.428 4.158 0.472 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.638 0.428 3.706 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.342 0.471 2.41 0.515 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 3.638 0.448 3.706 0.492 ;
        RECT 3.854 0.428 3.922 0.472 ;
        RECT 4.07 0.428 4.138 0.472 ;
        RECT 4.826 0.448 4.894 0.492 ;
        RECT 5.042 0.448 5.11 0.492 ;
        RECT 5.366 0.472 5.434 0.516 ;
        RECT 5.582 0.472 5.65 0.516 ;
        RECT 5.798 0.472 5.866 0.516 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.974 0.022 ;
        RECT 5.798 -0.022 5.866 0.292 ;
        RECT 5.582 -0.022 5.65 0.292 ;
        RECT 5.366 -0.022 5.434 0.292 ;
        RECT 4.934 -0.022 5.002 0.112 ;
        RECT 4.07 -0.022 4.138 0.202 ;
        RECT 3.854 -0.022 3.922 0.202 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 2.342 0.248 2.754 0.292 ;
        RECT 2.342 -0.022 2.41 0.292 ;
        RECT 1.782 0.158 2.194 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.197 0.25 0.241 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.342 0.1655 2.41 0.2095 ;
        RECT 2.666 0.248 2.734 0.292 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.854 0.1285 3.922 0.1725 ;
        RECT 4.07 0.1285 4.138 0.1725 ;
        RECT 4.936 0.048 5 0.092 ;
        RECT 5.366 0.1885 5.434 0.2325 ;
        RECT 5.582 0.1885 5.65 0.2325 ;
        RECT 5.798 0.1885 5.866 0.2325 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.704 0.518 1.904 0.562 ;
      RECT 1.984 0.518 5.344 0.562 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 1.586 0.248 1.654 0.562 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.91 0.518 2.106 0.562 ;
      RECT 2.538 0.158 2.882 0.202 ;
      RECT 3.078 0.338 3.206 0.382 ;
      RECT 2.214 0.338 2.774 0.382 ;
      RECT 3.638 0.338 4.286 0.382 ;
      RECT 4.07 0.518 4.718 0.562 ;
      RECT 4.394 0.068 4.462 0.292 ;
      RECT 5.258 0.428 5.326 0.562 ;
    LAYER v1 ;
      RECT 5.262 0.518 5.322 0.562 ;
      RECT 2.022 0.518 2.082 0.562 ;
      RECT 1.698 0.518 1.758 0.562 ;
      RECT 0.726 0.518 0.786 0.562 ;
    LAYER v0 ;
      RECT 5.258 0.472 5.326 0.516 ;
      RECT 5.152 0.088 5.216 0.132 ;
      RECT 5.042 0.248 5.11 0.292 ;
      RECT 4.934 0.448 5.002 0.492 ;
      RECT 4.718 0.248 4.786 0.292 ;
      RECT 4.612 0.138 4.676 0.182 ;
      RECT 4.502 0.223 4.57 0.267 ;
      RECT 4.502 0.428 4.57 0.472 ;
      RECT 4.394 0.338 4.462 0.382 ;
      RECT 4.396 0.138 4.46 0.182 ;
      RECT 4.286 0.223 4.354 0.267 ;
      RECT 4.286 0.428 4.354 0.472 ;
      RECT 4.178 0.1285 4.246 0.1725 ;
      RECT 4.178 0.518 4.246 0.562 ;
      RECT 3.962 0.338 4.03 0.382 ;
      RECT 3.746 0.338 3.814 0.382 ;
      RECT 3.638 0.158 3.706 0.202 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 3.316 0.178 3.38 0.222 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 3.098 0.338 3.166 0.382 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.884 0.358 2.948 0.402 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 2.02 0.318 2.084 0.362 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.49 1.654 0.534 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.614 0.202 0.682 0.246 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.202 0.574 0.246 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.378 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.338 1.114 0.472 ;
      RECT 1.114 0.338 1.262 0.382 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.33 0.428 1.478 0.472 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.546 0.158 1.674 0.202 ;
      RECT 1.654 0.248 2.018 0.292 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 1.762 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.472 ;
      RECT 1.978 0.428 2.302 0.472 ;
      RECT 2.882 0.158 2.95 0.472 ;
      RECT 2.95 0.158 3.078 0.202 ;
      RECT 2.95 0.428 3.294 0.472 ;
      RECT 2.862 0.068 3.206 0.112 ;
      RECT 3.206 0.068 3.274 0.382 ;
      RECT 3.274 0.338 3.402 0.382 ;
      RECT 3.274 0.068 3.422 0.112 ;
      RECT 3.422 0.068 3.49 0.202 ;
      RECT 3.49 0.158 3.726 0.202 ;
      RECT 2.774 0.338 2.842 0.562 ;
      RECT 3.314 0.158 3.382 0.292 ;
      RECT 2.842 0.518 3.53 0.562 ;
      RECT 3.382 0.248 3.53 0.292 ;
      RECT 3.53 0.248 3.598 0.562 ;
      RECT 3.598 0.248 4.178 0.292 ;
      RECT 4.178 0.068 4.246 0.292 ;
      RECT 4.286 0.158 4.354 0.382 ;
      RECT 4.354 0.338 4.502 0.382 ;
      RECT 4.502 0.158 4.57 0.382 ;
      RECT 4.718 0.158 4.786 0.562 ;
      RECT 4.786 0.338 4.934 0.382 ;
      RECT 4.934 0.248 5.002 0.562 ;
      RECT 5.002 0.248 5.13 0.292 ;
      RECT 4.266 0.428 4.61 0.472 ;
      RECT 4.462 0.068 4.61 0.112 ;
      RECT 4.61 0.068 4.678 0.472 ;
      RECT 4.678 0.068 4.826 0.112 ;
      RECT 4.826 0.068 4.894 0.202 ;
      RECT 4.894 0.158 5.15 0.202 ;
      RECT 5.15 0.068 5.218 0.202 ;
  END
END b15fpy040hn1n16x5

MACRO b15fpy080hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy080hn1n02x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.338 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.448 2.302 0.492 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.558 0.113 2.626 0.157 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.84 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.42 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.79 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.614 0.068 0.682 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.478 0.473 1.546 0.517 ;
        RECT 2.018 0.383 2.086 0.427 ;
        RECT 2.45 0.448 2.518 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.478 0.113 1.546 0.157 ;
        RECT 2.018 0.113 2.086 0.157 ;
        RECT 2.45 0.113 2.518 0.157 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.518 2.428 0.562 ;
      RECT 1.568 0.068 2.428 0.112 ;
    LAYER m1 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.938 0.068 1.262 0.112 ;
      RECT 1.37 0.248 1.586 0.292 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.694 0.248 1.762 0.562 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
    LAYER v1 ;
      RECT 2.346 0.518 2.406 0.562 ;
      RECT 2.238 0.068 2.298 0.112 ;
      RECT 1.914 0.518 1.974 0.562 ;
      RECT 1.698 0.068 1.758 0.112 ;
      RECT 1.698 0.518 1.758 0.562 ;
      RECT 0.942 0.518 1.002 0.562 ;
    LAYER v0 ;
      RECT 2.342 0.113 2.41 0.157 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.234 0.113 2.302 0.157 ;
      RECT 1.91 0.383 1.978 0.427 ;
      RECT 1.802 0.473 1.87 0.517 ;
      RECT 1.694 0.113 1.762 0.157 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.113 1.654 0.157 ;
      RECT 1.586 0.473 1.654 0.517 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.2435 1.222 0.2875 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.046 0.2435 1.114 0.2875 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.508 0.231 0.572 0.275 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.518 1.33 0.562 ;
      RECT 1.222 0.428 1.438 0.472 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.33 0.338 1.546 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.87 0.248 2.234 0.292 ;
      RECT 2.234 0.068 2.302 0.292 ;
  END
END b15fpy080hn1n02x5

MACRO b15fpy080hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy080hn1n03x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.338 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.448 2.302 0.492 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.558 0.113 2.626 0.157 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.84 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.42 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.79 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.614 0.068 0.682 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.478 0.473 1.546 0.517 ;
        RECT 2.018 0.383 2.086 0.427 ;
        RECT 2.45 0.448 2.518 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.478 0.113 1.546 0.157 ;
        RECT 2.018 0.113 2.086 0.157 ;
        RECT 2.45 0.113 2.518 0.157 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.518 2.428 0.562 ;
      RECT 1.568 0.068 2.428 0.112 ;
    LAYER m1 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.938 0.068 1.262 0.112 ;
      RECT 1.37 0.248 1.586 0.292 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.694 0.248 1.762 0.562 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
    LAYER v1 ;
      RECT 2.346 0.518 2.406 0.562 ;
      RECT 2.238 0.068 2.298 0.112 ;
      RECT 1.914 0.518 1.974 0.562 ;
      RECT 1.698 0.068 1.758 0.112 ;
      RECT 1.698 0.518 1.758 0.562 ;
      RECT 0.942 0.518 1.002 0.562 ;
    LAYER v0 ;
      RECT 2.342 0.113 2.41 0.157 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.234 0.113 2.302 0.157 ;
      RECT 1.91 0.383 1.978 0.427 ;
      RECT 1.802 0.473 1.87 0.517 ;
      RECT 1.694 0.113 1.762 0.157 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.113 1.654 0.157 ;
      RECT 1.586 0.473 1.654 0.517 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.2435 1.222 0.2875 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.046 0.2435 1.114 0.2875 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.508 0.231 0.572 0.275 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.518 1.33 0.562 ;
      RECT 1.222 0.428 1.438 0.472 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.33 0.338 1.546 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.87 0.248 2.234 0.292 ;
      RECT 2.234 0.068 2.302 0.292 ;
  END
END b15fpy080hn1n03x5

MACRO b15fpy080hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy080hn1n04x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.6075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.6075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.428 1.006 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.448 1.006 0.492 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.4285 2.626 0.4725 ;
        RECT 2.558 0.1585 2.626 0.2025 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.478 0.408 1.546 0.452 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.45 0.4285 2.518 0.4725 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.018 -0.022 2.086 0.292 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.45 0.1585 2.518 0.2025 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.704 0.248 2.32 0.292 ;
      RECT 0.812 0.158 2.32 0.202 ;
    LAYER m1 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.37 0.248 1.586 0.292 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.262 0.068 1.33 0.472 ;
      RECT 1.586 0.518 1.802 0.562 ;
      RECT 1.694 0.068 1.762 0.472 ;
      RECT 1.91 0.068 1.978 0.472 ;
      RECT 2.126 0.068 2.194 0.562 ;
      RECT 2.234 0.158 2.302 0.382 ;
      RECT 2.342 0.068 2.41 0.562 ;
    LAYER v1 ;
      RECT 2.238 0.248 2.298 0.292 ;
      RECT 2.13 0.158 2.19 0.202 ;
      RECT 1.914 0.158 1.974 0.202 ;
      RECT 1.698 0.158 1.758 0.202 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 0.942 0.158 1.002 0.202 ;
      RECT 0.834 0.248 0.894 0.292 ;
    LAYER v0 ;
      RECT 2.342 0.1585 2.41 0.2025 ;
      RECT 2.342 0.4285 2.41 0.4725 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.802 0.1535 1.87 0.1975 ;
      RECT 1.694 0.3155 1.762 0.3595 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.1575 1.222 0.2015 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 1.046 0.1575 1.114 0.2015 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.508 0.231 0.572 0.275 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.802 0.068 1.87 0.562 ;
  END
END b15fpy080hn1n04x5

MACRO b15fpy080hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy080hn1n06x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.292 ;
      LAYER v0 ;
        RECT 2.342 0.088 2.41 0.132 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.158 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.666 0.203 2.734 0.247 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.452 0.25 0.496 ;
        RECT 0.722 0.452 0.79 0.496 ;
        RECT 1.478 0.472 1.546 0.516 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.558 -0.022 2.626 0.292 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1975 0.25 0.2415 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.478 0.048 1.546 0.092 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.558 0.203 2.626 0.247 ;
        RECT 2.774 0.203 2.842 0.247 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.812 0.428 2.536 0.472 ;
    LAYER m1 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.37 0.248 1.586 0.292 ;
      RECT 0.83 0.068 1.262 0.112 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 1.694 0.518 2.018 0.562 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.45 0.068 2.518 0.562 ;
    LAYER v1 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 0.942 0.428 1.002 0.472 ;
    LAYER v0 ;
      RECT 2.45 0.203 2.518 0.247 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.472 1.654 0.516 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.2435 1.222 0.2875 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.2435 1.114 0.2875 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.508 0.2345 0.572 0.2785 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.518 1.33 0.562 ;
      RECT 1.222 0.428 1.438 0.472 ;
      RECT 1.586 0.248 1.654 0.562 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.33 0.338 1.546 0.382 ;
      RECT 1.33 0.158 1.694 0.202 ;
      RECT 1.694 0.068 1.762 0.472 ;
      RECT 1.762 0.068 1.978 0.112 ;
      RECT 1.802 0.158 2.018 0.202 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 2.086 0.338 2.342 0.382 ;
      RECT 2.342 0.338 2.41 0.562 ;
  END
END b15fpy080hn1n06x5

MACRO b15fpy080hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy080hn1n08x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.292 ;
      LAYER v0 ;
        RECT 2.342 0.088 2.41 0.132 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.158 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.666 0.203 2.734 0.247 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.452 0.25 0.496 ;
        RECT 0.722 0.452 0.79 0.496 ;
        RECT 1.478 0.472 1.546 0.516 ;
        RECT 2.126 0.473 2.194 0.517 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.558 -0.022 2.626 0.292 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1975 0.25 0.2415 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.478 0.048 1.546 0.092 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.558 0.203 2.626 0.247 ;
        RECT 2.774 0.203 2.842 0.247 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.812 0.428 2.536 0.472 ;
    LAYER m1 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.37 0.248 1.586 0.292 ;
      RECT 0.83 0.068 1.262 0.112 ;
      RECT 1.91 0.248 1.978 0.562 ;
      RECT 1.802 0.158 1.87 0.562 ;
      RECT 2.018 0.338 2.45 0.382 ;
      RECT 2.234 0.428 2.302 0.562 ;
    LAYER v1 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 0.942 0.428 1.002 0.472 ;
    LAYER v0 ;
      RECT 2.45 0.203 2.518 0.247 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.234 0.473 2.302 0.517 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.472 1.654 0.516 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.2435 1.222 0.2875 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.2435 1.114 0.2875 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.508 0.2345 0.572 0.2785 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.518 1.33 0.562 ;
      RECT 1.222 0.428 1.438 0.472 ;
      RECT 1.586 0.248 1.654 0.562 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.33 0.338 1.546 0.382 ;
      RECT 1.33 0.158 1.694 0.202 ;
      RECT 1.694 0.068 1.762 0.472 ;
      RECT 1.762 0.068 1.978 0.112 ;
      RECT 1.87 0.158 2.086 0.202 ;
      RECT 2.45 0.068 2.518 0.562 ;
  END
END b15fpy080hn1n08x5

MACRO b15fpy080hn1n08x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy080hn1n08x7 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.428 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.4665 2.842 0.5105 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.09777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.898 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.068 3.166 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.4665 3.166 0.5105 ;
        RECT 3.098 0.158 3.166 0.202 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.61777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.452 0.25 0.496 ;
        RECT 0.722 0.473 0.79 0.517 ;
        RECT 1.478 0.472 1.546 0.516 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.558 0.4665 2.626 0.5105 ;
        RECT 2.99 0.4665 3.058 0.5105 ;
        RECT 3.206 0.4665 3.274 0.5105 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 3.206 -0.022 3.274 0.292 ;
        RECT 2.99 -0.022 3.058 0.292 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.37 0.158 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.702 0.158 0.898 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1975 0.25 0.2415 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.206 0.158 3.274 0.202 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.028 0.428 2.32 0.472 ;
    LAYER m1 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.37 0.248 1.91 0.292 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 2.126 0.158 2.194 0.562 ;
      RECT 2.018 0.248 2.086 0.562 ;
      RECT 2.234 0.248 2.302 0.562 ;
      RECT 2.342 0.338 2.882 0.382 ;
    LAYER v1 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 1.05 0.428 1.11 0.472 ;
    LAYER v0 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.882 0.4665 2.95 0.5105 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.126 0.43 2.194 0.474 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.154 0.1785 1.222 0.2225 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.439 1.006 0.483 ;
      RECT 0.94 0.178 1.004 0.222 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.068 0.574 0.472 ;
      RECT 0.574 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.562 ;
      RECT 1.222 0.518 1.438 0.562 ;
      RECT 1.33 0.338 1.546 0.382 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.194 0.158 2.342 0.202 ;
      RECT 2.342 0.158 2.41 0.292 ;
      RECT 2.41 0.248 2.774 0.292 ;
      RECT 2.774 0.068 2.842 0.292 ;
      RECT 2.882 0.068 2.95 0.562 ;
  END
END b15fpy080hn1n08x7

MACRO b15fpy080hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy080hn1n12x5 0 0 ;
  SIZE 3.564 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 5.28833325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 5.28833325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.338 2.842 0.472 ;
      LAYER v0 ;
        RECT 2.774 0.3825 2.842 0.4265 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.825679 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.81 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.068 3.49 0.562 ;
        RECT 3.206 0.338 3.49 0.382 ;
        RECT 3.206 0.068 3.274 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.4665 3.274 0.5105 ;
        RECT 3.206 0.113 3.274 0.157 ;
        RECT 3.422 0.4665 3.49 0.5105 ;
        RECT 3.422 0.113 3.49 0.157 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.61777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.452 0.25 0.496 ;
        RECT 0.722 0.473 0.79 0.517 ;
        RECT 1.478 0.472 1.546 0.516 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.558 0.4665 2.626 0.5105 ;
        RECT 2.882 0.4665 2.95 0.5105 ;
        RECT 3.098 0.4665 3.166 0.5105 ;
        RECT 3.314 0.4665 3.382 0.5105 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.598 0.022 ;
        RECT 3.314 -0.022 3.382 0.292 ;
        RECT 3.098 -0.022 3.166 0.292 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.614 0.158 0.898 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1975 0.25 0.2415 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.478 0.114 1.546 0.158 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.45 0.048 2.518 0.092 ;
        RECT 2.882 0.113 2.95 0.157 ;
        RECT 3.098 0.113 3.166 0.157 ;
        RECT 3.314 0.113 3.382 0.157 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.028 0.428 2.212 0.472 ;
    LAYER m1 ;
      RECT 1.154 0.068 1.222 0.562 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.37 0.248 1.586 0.292 ;
      RECT 1.694 0.428 1.762 0.562 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.234 0.338 2.666 0.382 ;
      RECT 1.694 0.068 1.762 0.292 ;
      RECT 2.342 0.248 2.99 0.292 ;
    LAYER v1 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 1.05 0.428 1.11 0.472 ;
    LAYER v0 ;
      RECT 2.99 0.113 3.058 0.157 ;
      RECT 2.99 0.3825 3.058 0.4265 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.666 0.4665 2.734 0.5105 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.694 0.138 1.762 0.182 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.154 0.1785 1.222 0.2225 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.439 1.006 0.483 ;
      RECT 0.94 0.178 1.004 0.222 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.068 0.574 0.472 ;
      RECT 0.574 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.562 ;
      RECT 1.222 0.518 1.438 0.562 ;
      RECT 1.33 0.338 1.546 0.382 ;
      RECT 1.586 0.248 1.654 0.382 ;
      RECT 1.654 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 2.086 0.158 2.302 0.202 ;
      RECT 2.086 0.518 2.41 0.562 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 1.762 0.248 1.91 0.292 ;
      RECT 1.91 0.068 1.978 0.292 ;
      RECT 1.978 0.068 2.342 0.112 ;
      RECT 2.342 0.068 2.41 0.202 ;
      RECT 2.41 0.158 2.842 0.202 ;
      RECT 2.99 0.068 3.058 0.472 ;
  END
END b15fpy080hn1n12x5

MACRO b15fpy080hn1n12x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy080hn1n12x7 0 0 ;
  SIZE 3.996 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 3.07166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 3.07166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.428 3.274 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.448 3.274 0.492 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.222 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.068 3.922 0.562 ;
        RECT 3.638 0.338 3.922 0.382 ;
        RECT 3.638 0.068 3.706 0.382 ;
      LAYER v0 ;
        RECT 3.638 0.1525 3.706 0.1965 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 3.854 0.1525 3.922 0.1965 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.13925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.472 0.25 0.516 ;
        RECT 0.722 0.4725 0.79 0.5165 ;
        RECT 1.154 0.4725 1.222 0.5165 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.882 0.473 2.95 0.517 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 3.746 0.448 3.814 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.03 0.022 ;
        RECT 3.746 -0.022 3.814 0.292 ;
        RECT 3.53 -0.022 3.598 0.292 ;
        RECT 3.314 -0.022 3.382 0.292 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.702 0.158 0.898 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1905 0.25 0.2345 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.314 0.1525 3.382 0.1965 ;
        RECT 3.53 0.1525 3.598 0.1965 ;
        RECT 3.746 0.1525 3.814 0.1965 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.244 0.428 2.86 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 1.694 0.518 1.91 0.562 ;
      RECT 1.802 0.248 1.87 0.472 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 2.45 0.248 2.518 0.472 ;
      RECT 2.666 0.248 2.734 0.472 ;
      RECT 2.774 0.338 3.422 0.382 ;
    LAYER v1 ;
      RECT 2.67 0.428 2.73 0.472 ;
      RECT 2.454 0.428 2.514 0.472 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
    LAYER v0 ;
      RECT 3.422 0.1525 3.49 0.1965 ;
      RECT 3.422 0.448 3.49 0.492 ;
      RECT 3.206 0.1525 3.274 0.1965 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.558 0.43 2.626 0.474 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 1.802 0.3155 1.87 0.3595 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.408 1.762 0.452 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.262 0.4725 1.33 0.5165 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.33 0.338 1.654 0.382 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.248 1.694 0.292 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.566 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 1.978 0.338 2.302 0.382 ;
      RECT 2.194 0.248 2.342 0.292 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.626 0.158 2.774 0.202 ;
      RECT 2.774 0.158 2.842 0.292 ;
      RECT 2.842 0.248 3.206 0.292 ;
      RECT 3.206 0.068 3.274 0.292 ;
      RECT 3.422 0.068 3.49 0.562 ;
  END
END b15fpy080hn1n12x7

MACRO b15fpy080hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy080hn1n16x5 0 0 ;
  SIZE 4.212 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.248 3.166 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.2705 3.166 0.3145 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.222 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.068 4.03 0.562 ;
        RECT 3.746 0.338 4.03 0.382 ;
        RECT 3.746 0.068 3.814 0.562 ;
      LAYER v0 ;
        RECT 3.746 0.448 3.814 0.492 ;
        RECT 3.746 0.178 3.814 0.222 ;
        RECT 3.962 0.448 4.03 0.492 ;
        RECT 3.962 0.178 4.03 0.222 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.13925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.246 0.652 ;
        RECT 4.07 0.338 4.138 0.652 ;
        RECT 3.854 0.428 3.922 0.652 ;
        RECT 3.638 0.338 3.706 0.652 ;
        RECT 3.422 0.338 3.49 0.652 ;
        RECT 2.99 0.338 3.058 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.472 0.25 0.516 ;
        RECT 0.722 0.4725 0.79 0.5165 ;
        RECT 1.154 0.4725 1.222 0.5165 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.99 0.428 3.058 0.472 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.638 0.448 3.706 0.492 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 4.07 0.448 4.138 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.246 0.022 ;
        RECT 4.07 -0.022 4.138 0.292 ;
        RECT 3.854 -0.022 3.922 0.292 ;
        RECT 3.638 -0.022 3.706 0.292 ;
        RECT 3.422 -0.022 3.49 0.292 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.342 -0.022 2.41 0.292 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.702 0.158 0.898 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1905 0.25 0.2345 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 2.126 0.143 2.194 0.187 ;
        RECT 2.342 0.143 2.41 0.187 ;
        RECT 2.99 0.048 3.058 0.092 ;
        RECT 3.422 0.178 3.49 0.222 ;
        RECT 3.638 0.178 3.706 0.222 ;
        RECT 3.854 0.178 3.922 0.222 ;
        RECT 4.07 0.178 4.138 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.136 0.428 3.292 0.472 ;
      RECT 1.244 0.158 3.4 0.202 ;
    LAYER m1 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 2.018 0.158 2.086 0.382 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 2.666 0.158 2.734 0.562 ;
      RECT 2.558 0.248 2.626 0.472 ;
      RECT 2.882 0.248 2.95 0.472 ;
      RECT 3.206 0.158 3.274 0.562 ;
      RECT 3.53 0.068 3.598 0.562 ;
    LAYER v1 ;
      RECT 3.21 0.158 3.27 0.202 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.374 0.158 1.434 0.202 ;
      RECT 1.266 0.428 1.326 0.472 ;
    LAYER v0 ;
      RECT 3.53 0.178 3.598 0.222 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.314 0.178 3.382 0.222 ;
      RECT 3.206 0.178 3.274 0.222 ;
      RECT 3.206 0.406 3.274 0.45 ;
      RECT 2.882 0.3155 2.95 0.3595 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.666 0.43 2.734 0.474 ;
      RECT 2.558 0.338 2.626 0.382 ;
      RECT 2.45 0.143 2.518 0.187 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.234 0.143 2.302 0.187 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.802 0.157 1.87 0.201 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.694 0.157 1.762 0.201 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.4725 1.33 0.5165 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.068 0.574 0.472 ;
      RECT 0.574 0.248 1.262 0.292 ;
      RECT 1.262 0.068 1.33 0.292 ;
      RECT 1.33 0.068 1.694 0.112 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 2.086 0.338 2.234 0.382 ;
      RECT 2.234 0.068 2.302 0.562 ;
      RECT 2.302 0.338 2.45 0.382 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 2.734 0.158 3.098 0.202 ;
      RECT 3.098 0.068 3.166 0.202 ;
      RECT 3.166 0.068 3.314 0.112 ;
      RECT 3.314 0.068 3.382 0.292 ;
  END
END b15fpy080hn1n16x5

MACRO b15fpy080hn1n16x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy080hn1n16x7 0 0 ;
  SIZE 5.076 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.30375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.30375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.158 4.138 0.472 ;
      LAYER v0 ;
        RECT 4.07 0.408 4.138 0.452 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.242 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.826 0.068 4.894 0.562 ;
        RECT 4.61 0.248 4.894 0.292 ;
        RECT 4.61 0.068 4.678 0.562 ;
      LAYER v0 ;
        RECT 4.61 0.43 4.678 0.474 ;
        RECT 4.61 0.138 4.678 0.182 ;
        RECT 4.826 0.43 4.894 0.474 ;
        RECT 4.826 0.138 4.894 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 2.4594445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.11 0.652 ;
        RECT 4.934 0.338 5.002 0.652 ;
        RECT 4.718 0.338 4.786 0.652 ;
        RECT 4.502 0.338 4.57 0.652 ;
        RECT 4.286 0.338 4.354 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.472 0.25 0.516 ;
        RECT 0.722 0.4725 0.79 0.5165 ;
        RECT 1.154 0.4725 1.222 0.5165 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 3.422 0.478 3.49 0.522 ;
        RECT 3.746 0.448 3.814 0.492 ;
        RECT 4.286 0.43 4.354 0.474 ;
        RECT 4.502 0.43 4.57 0.474 ;
        RECT 4.718 0.43 4.786 0.474 ;
        RECT 4.934 0.43 5.002 0.474 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.11 0.022 ;
        RECT 4.934 -0.022 5.002 0.292 ;
        RECT 4.718 -0.022 4.786 0.202 ;
        RECT 4.502 -0.022 4.57 0.292 ;
        RECT 4.286 -0.022 4.354 0.202 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.292 ;
        RECT 1.046 0.158 1.242 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.702 0.158 0.898 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.1905 0.25 0.2345 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 3.424 0.138 3.488 0.182 ;
        RECT 3.746 0.138 3.814 0.182 ;
        RECT 4.286 0.138 4.354 0.182 ;
        RECT 4.502 0.138 4.57 0.182 ;
        RECT 4.718 0.138 4.786 0.182 ;
        RECT 4.934 0.138 5.002 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.46 0.428 3.616 0.472 ;
      RECT 1.676 0.248 4.156 0.292 ;
    LAYER m1 ;
      RECT 1.478 0.068 1.546 0.472 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.774 0.248 2.842 0.472 ;
      RECT 2.666 0.158 2.882 0.202 ;
      RECT 3.206 0.248 3.274 0.472 ;
      RECT 3.53 0.428 3.598 0.562 ;
      RECT 3.962 0.158 4.03 0.472 ;
      RECT 3.402 0.338 3.854 0.382 ;
    LAYER v1 ;
      RECT 3.966 0.248 4.026 0.292 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.806 0.248 1.866 0.292 ;
      RECT 1.482 0.428 1.542 0.472 ;
    LAYER v0 ;
      RECT 4.394 0.138 4.462 0.182 ;
      RECT 4.394 0.43 4.462 0.474 ;
      RECT 4.07 0.068 4.138 0.112 ;
      RECT 3.962 0.178 4.03 0.222 ;
      RECT 3.962 0.408 4.03 0.452 ;
      RECT 3.53 0.478 3.598 0.522 ;
      RECT 3.422 0.338 3.49 0.382 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.206 0.338 3.274 0.382 ;
      RECT 3.098 0.498 3.166 0.542 ;
      RECT 2.99 0.178 3.058 0.222 ;
      RECT 2.99 0.408 3.058 0.452 ;
      RECT 2.882 0.408 2.95 0.452 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.3155 2.842 0.3595 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.4385 1.978 0.4825 ;
      RECT 1.802 0.4385 1.87 0.4825 ;
      RECT 1.694 0.3135 1.762 0.3575 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.586 0.3135 1.654 0.3575 ;
      RECT 1.37 0.422 1.438 0.466 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.068 0.574 0.472 ;
      RECT 0.574 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.438 0.518 1.694 0.562 ;
      RECT 1.694 0.248 1.762 0.562 ;
      RECT 1.546 0.068 1.762 0.112 ;
      RECT 1.654 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 1.978 0.158 2.234 0.202 ;
      RECT 2.234 0.158 2.302 0.382 ;
      RECT 2.302 0.338 2.538 0.382 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 2.194 0.428 2.666 0.472 ;
      RECT 2.518 0.248 2.666 0.292 ;
      RECT 2.666 0.248 2.734 0.562 ;
      RECT 2.734 0.518 2.99 0.562 ;
      RECT 2.99 0.158 3.058 0.562 ;
      RECT 2.882 0.068 2.95 0.472 ;
      RECT 2.95 0.068 3.098 0.112 ;
      RECT 3.098 0.068 3.166 0.562 ;
      RECT 3.166 0.158 3.314 0.202 ;
      RECT 3.314 0.158 3.382 0.292 ;
      RECT 3.382 0.248 3.854 0.292 ;
      RECT 3.854 0.068 3.922 0.292 ;
      RECT 3.922 0.068 4.246 0.112 ;
      RECT 3.854 0.338 3.922 0.562 ;
      RECT 3.922 0.518 4.178 0.562 ;
      RECT 4.178 0.248 4.246 0.562 ;
      RECT 4.246 0.248 4.394 0.292 ;
      RECT 4.394 0.068 4.462 0.562 ;
  END
END b15fpy080hn1n16x7

MACRO b15fpy200hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy200hn1n02x5 0 0 ;
  SIZE 4.752 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.472 ;
      LAYER v0 ;
        RECT 2.018 0.338 2.086 0.382 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.158 2.95 0.472 ;
      LAYER v0 ;
        RECT 2.882 0.338 2.95 0.382 ;
    END
  END d2
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.068 4.678 0.562 ;
      LAYER v0 ;
        RECT 4.61 0.448 4.678 0.492 ;
        RECT 4.61 0.138 4.678 0.182 ;
    END
  END o2
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.292 ;
      LAYER v0 ;
        RECT 2.342 0.088 2.41 0.132 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.292 ;
      LAYER v0 ;
        RECT 2.558 0.088 2.626 0.132 ;
    END
  END si2
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 5.51 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.95 0.112 ;
        RECT 2.234 0.338 2.734 0.382 ;
        RECT 2.666 0.068 2.734 0.382 ;
        RECT 2.234 0.068 2.302 0.382 ;
        RECT 2.018 0.068 2.302 0.112 ;
      LAYER v0 ;
        RECT 2.126 0.068 2.194 0.112 ;
        RECT 2.342 0.338 2.41 0.382 ;
        RECT 2.558 0.338 2.626 0.382 ;
        RECT 2.774 0.068 2.842 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.786 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.638 0.428 3.706 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.638 0.473 3.706 0.517 ;
        RECT 4.178 0.448 4.246 0.492 ;
        RECT 4.502 0.448 4.57 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.786 0.022 ;
        RECT 4.502 -0.022 4.57 0.112 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.638 -0.022 3.706 0.202 ;
        RECT 2.99 -0.022 3.058 0.292 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.262 0.113 1.33 0.157 ;
        RECT 1.91 0.138 1.978 0.182 ;
        RECT 2.45 0.222 2.518 0.266 ;
        RECT 2.99 0.183 3.058 0.227 ;
        RECT 3.638 0.138 3.706 0.182 ;
        RECT 4.178 0.138 4.246 0.182 ;
        RECT 4.502 0.048 4.57 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.338 1.024 0.382 ;
      RECT 1.568 0.338 2.212 0.382 ;
      RECT 2.756 0.338 3.4 0.382 ;
      RECT 0.488 0.428 4.156 0.472 ;
      RECT 1.784 0.518 4.372 0.562 ;
      RECT 3.944 0.338 4.588 0.382 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.382 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 0.938 0.068 1.006 0.562 ;
      RECT 1.242 0.338 1.478 0.382 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 2.558 0.428 2.774 0.472 ;
      RECT 3.098 0.338 3.166 0.472 ;
      RECT 3.206 0.428 3.274 0.562 ;
      RECT 3.314 0.068 3.382 0.562 ;
      RECT 3.422 0.068 3.49 0.562 ;
      RECT 3.53 0.158 3.598 0.562 ;
      RECT 3.746 0.068 3.814 0.562 ;
      RECT 3.854 0.248 3.922 0.472 ;
      RECT 3.962 0.068 4.03 0.562 ;
      RECT 4.07 0.158 4.138 0.472 ;
      RECT 4.286 0.068 4.354 0.562 ;
      RECT 4.394 0.068 4.462 0.562 ;
      RECT 4.502 0.158 4.57 0.382 ;
    LAYER v1 ;
      RECT 4.506 0.338 4.566 0.382 ;
      RECT 4.29 0.518 4.35 0.562 ;
      RECT 4.074 0.428 4.134 0.472 ;
      RECT 3.966 0.338 4.026 0.382 ;
      RECT 3.858 0.428 3.918 0.472 ;
      RECT 3.534 0.518 3.594 0.562 ;
      RECT 3.318 0.338 3.378 0.382 ;
      RECT 3.21 0.518 3.27 0.562 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.778 0.338 2.838 0.382 ;
      RECT 2.13 0.338 2.19 0.382 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 4.502 0.248 4.57 0.292 ;
      RECT 4.394 0.138 4.462 0.182 ;
      RECT 4.394 0.448 4.462 0.492 ;
      RECT 4.286 0.138 4.354 0.182 ;
      RECT 4.286 0.448 4.354 0.492 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 3.962 0.138 4.03 0.182 ;
      RECT 3.962 0.448 4.03 0.492 ;
      RECT 3.854 0.338 3.922 0.382 ;
      RECT 3.746 0.138 3.814 0.182 ;
      RECT 3.746 0.473 3.814 0.517 ;
      RECT 3.53 0.248 3.598 0.292 ;
      RECT 3.422 0.1515 3.49 0.1955 ;
      RECT 3.422 0.47 3.49 0.514 ;
      RECT 3.314 0.1515 3.382 0.1955 ;
      RECT 3.314 0.47 3.382 0.514 ;
      RECT 3.206 0.47 3.274 0.514 ;
      RECT 3.208 0.268 3.272 0.312 ;
      RECT 2.774 0.203 2.842 0.247 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.203 2.194 0.247 ;
      RECT 1.802 0.138 1.87 0.182 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.694 0.292 1.762 0.336 ;
      RECT 1.586 0.1515 1.654 0.1955 ;
      RECT 1.586 0.453 1.654 0.497 ;
      RECT 1.478 0.1515 1.546 0.1955 ;
      RECT 1.478 0.453 1.546 0.497 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.113 1.222 0.157 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.113 1.006 0.157 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.29 0.448 0.358 0.492 ;
      RECT 0.182 0.293 0.25 0.337 ;
    LAYER m1 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.248 1.35 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 2.194 0.428 2.41 0.472 ;
      RECT 2.774 0.158 2.842 0.472 ;
      RECT 3.166 0.338 3.206 0.382 ;
      RECT 3.206 0.248 3.274 0.382 ;
  END
END b15fpy200hn1n02x5

MACRO b15fpy200hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy200hn1n03x5 0 0 ;
  SIZE 4.752 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.472 ;
      LAYER v0 ;
        RECT 2.018 0.338 2.086 0.382 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.158 2.95 0.472 ;
      LAYER v0 ;
        RECT 2.882 0.338 2.95 0.382 ;
    END
  END d2
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.068 4.678 0.562 ;
      LAYER v0 ;
        RECT 4.61 0.448 4.678 0.492 ;
        RECT 4.61 0.138 4.678 0.182 ;
    END
  END o2
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.292 ;
      LAYER v0 ;
        RECT 2.342 0.088 2.41 0.132 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.292 ;
      LAYER v0 ;
        RECT 2.558 0.088 2.626 0.132 ;
    END
  END si2
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 5.51 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.95 0.112 ;
        RECT 2.234 0.338 2.734 0.382 ;
        RECT 2.666 0.068 2.734 0.382 ;
        RECT 2.234 0.068 2.302 0.382 ;
        RECT 2.018 0.068 2.302 0.112 ;
      LAYER v0 ;
        RECT 2.126 0.068 2.194 0.112 ;
        RECT 2.342 0.338 2.41 0.382 ;
        RECT 2.558 0.338 2.626 0.382 ;
        RECT 2.774 0.068 2.842 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.786 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.638 0.428 3.706 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.638 0.473 3.706 0.517 ;
        RECT 4.178 0.448 4.246 0.492 ;
        RECT 4.502 0.448 4.57 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.786 0.022 ;
        RECT 4.502 -0.022 4.57 0.112 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.638 -0.022 3.706 0.202 ;
        RECT 2.99 -0.022 3.058 0.292 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.262 0.113 1.33 0.157 ;
        RECT 1.91 0.138 1.978 0.182 ;
        RECT 2.45 0.222 2.518 0.266 ;
        RECT 2.99 0.183 3.058 0.227 ;
        RECT 3.638 0.138 3.706 0.182 ;
        RECT 4.178 0.138 4.246 0.182 ;
        RECT 4.502 0.048 4.57 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.338 1.024 0.382 ;
      RECT 1.568 0.338 2.212 0.382 ;
      RECT 2.756 0.338 3.4 0.382 ;
      RECT 0.488 0.428 4.156 0.472 ;
      RECT 1.784 0.518 4.372 0.562 ;
      RECT 3.944 0.338 4.588 0.382 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.382 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 0.938 0.068 1.006 0.562 ;
      RECT 1.242 0.338 1.478 0.382 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 2.558 0.428 2.774 0.472 ;
      RECT 3.098 0.338 3.166 0.472 ;
      RECT 3.206 0.428 3.274 0.562 ;
      RECT 3.314 0.068 3.382 0.562 ;
      RECT 3.422 0.068 3.49 0.562 ;
      RECT 3.53 0.158 3.598 0.562 ;
      RECT 3.746 0.068 3.814 0.562 ;
      RECT 3.854 0.248 3.922 0.472 ;
      RECT 3.962 0.068 4.03 0.562 ;
      RECT 4.07 0.158 4.138 0.472 ;
      RECT 4.286 0.068 4.354 0.562 ;
      RECT 4.394 0.068 4.462 0.562 ;
      RECT 4.502 0.158 4.57 0.382 ;
    LAYER v1 ;
      RECT 4.506 0.338 4.566 0.382 ;
      RECT 4.29 0.518 4.35 0.562 ;
      RECT 4.074 0.428 4.134 0.472 ;
      RECT 3.966 0.338 4.026 0.382 ;
      RECT 3.858 0.428 3.918 0.472 ;
      RECT 3.534 0.518 3.594 0.562 ;
      RECT 3.318 0.338 3.378 0.382 ;
      RECT 3.21 0.518 3.27 0.562 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.778 0.338 2.838 0.382 ;
      RECT 2.13 0.338 2.19 0.382 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 4.502 0.248 4.57 0.292 ;
      RECT 4.394 0.138 4.462 0.182 ;
      RECT 4.394 0.448 4.462 0.492 ;
      RECT 4.286 0.138 4.354 0.182 ;
      RECT 4.286 0.448 4.354 0.492 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 3.962 0.138 4.03 0.182 ;
      RECT 3.962 0.448 4.03 0.492 ;
      RECT 3.854 0.338 3.922 0.382 ;
      RECT 3.746 0.138 3.814 0.182 ;
      RECT 3.746 0.473 3.814 0.517 ;
      RECT 3.53 0.248 3.598 0.292 ;
      RECT 3.422 0.1515 3.49 0.1955 ;
      RECT 3.422 0.47 3.49 0.514 ;
      RECT 3.314 0.1515 3.382 0.1955 ;
      RECT 3.314 0.47 3.382 0.514 ;
      RECT 3.206 0.47 3.274 0.514 ;
      RECT 3.208 0.268 3.272 0.312 ;
      RECT 2.774 0.203 2.842 0.247 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.203 2.194 0.247 ;
      RECT 1.802 0.138 1.87 0.182 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.694 0.292 1.762 0.336 ;
      RECT 1.586 0.1515 1.654 0.1955 ;
      RECT 1.586 0.453 1.654 0.497 ;
      RECT 1.478 0.1515 1.546 0.1955 ;
      RECT 1.478 0.453 1.546 0.497 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.113 1.222 0.157 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.113 1.006 0.157 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.29 0.448 0.358 0.492 ;
      RECT 0.182 0.293 0.25 0.337 ;
    LAYER m1 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.248 1.35 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 2.194 0.428 2.41 0.472 ;
      RECT 2.774 0.158 2.842 0.472 ;
      RECT 3.166 0.338 3.206 0.382 ;
      RECT 3.206 0.248 3.274 0.382 ;
  END
END b15fpy200hn1n03x5

MACRO b15fpy200hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy200hn1n04x5 0 0 ;
  SIZE 4.752 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.472 ;
      LAYER v0 ;
        RECT 2.018 0.338 2.086 0.382 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.158 2.95 0.472 ;
      LAYER v0 ;
        RECT 2.882 0.338 2.95 0.382 ;
    END
  END d2
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.068 4.678 0.562 ;
      LAYER v0 ;
        RECT 4.61 0.448 4.678 0.492 ;
        RECT 4.61 0.138 4.678 0.182 ;
    END
  END o2
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.292 ;
      LAYER v0 ;
        RECT 2.342 0.088 2.41 0.132 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.292 ;
      LAYER v0 ;
        RECT 2.558 0.088 2.626 0.132 ;
    END
  END si2
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 5.51 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.95 0.112 ;
        RECT 2.234 0.338 2.734 0.382 ;
        RECT 2.666 0.068 2.734 0.382 ;
        RECT 2.234 0.068 2.302 0.382 ;
        RECT 2.018 0.068 2.302 0.112 ;
      LAYER v0 ;
        RECT 2.126 0.068 2.194 0.112 ;
        RECT 2.342 0.338 2.41 0.382 ;
        RECT 2.558 0.338 2.626 0.382 ;
        RECT 2.774 0.068 2.842 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.786 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.638 0.428 3.706 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.638 0.473 3.706 0.517 ;
        RECT 4.178 0.448 4.246 0.492 ;
        RECT 4.502 0.448 4.57 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.786 0.022 ;
        RECT 4.502 -0.022 4.57 0.112 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.638 -0.022 3.706 0.202 ;
        RECT 2.99 -0.022 3.058 0.292 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.262 0.113 1.33 0.157 ;
        RECT 1.91 0.138 1.978 0.182 ;
        RECT 2.45 0.222 2.518 0.266 ;
        RECT 2.99 0.183 3.058 0.227 ;
        RECT 3.638 0.138 3.706 0.182 ;
        RECT 4.178 0.138 4.246 0.182 ;
        RECT 4.504 0.048 4.568 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.338 1.024 0.382 ;
      RECT 1.568 0.338 2.212 0.382 ;
      RECT 2.756 0.338 3.4 0.382 ;
      RECT 0.488 0.428 4.156 0.472 ;
      RECT 1.784 0.518 4.372 0.562 ;
      RECT 3.944 0.338 4.588 0.382 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.382 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 0.938 0.068 1.006 0.562 ;
      RECT 1.242 0.338 1.478 0.382 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 2.558 0.428 2.774 0.472 ;
      RECT 3.098 0.338 3.166 0.472 ;
      RECT 3.206 0.428 3.274 0.562 ;
      RECT 3.314 0.068 3.382 0.562 ;
      RECT 3.422 0.068 3.49 0.562 ;
      RECT 3.53 0.158 3.598 0.562 ;
      RECT 3.746 0.068 3.814 0.562 ;
      RECT 3.854 0.248 3.922 0.472 ;
      RECT 3.962 0.068 4.03 0.562 ;
      RECT 4.07 0.158 4.138 0.472 ;
      RECT 4.286 0.068 4.354 0.562 ;
      RECT 4.394 0.068 4.462 0.562 ;
      RECT 4.502 0.158 4.57 0.382 ;
    LAYER v1 ;
      RECT 4.506 0.338 4.566 0.382 ;
      RECT 4.29 0.518 4.35 0.562 ;
      RECT 4.074 0.428 4.134 0.472 ;
      RECT 3.966 0.338 4.026 0.382 ;
      RECT 3.858 0.428 3.918 0.472 ;
      RECT 3.534 0.518 3.594 0.562 ;
      RECT 3.318 0.338 3.378 0.382 ;
      RECT 3.21 0.518 3.27 0.562 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.778 0.338 2.838 0.382 ;
      RECT 2.13 0.338 2.19 0.382 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 4.502 0.248 4.57 0.292 ;
      RECT 4.394 0.138 4.462 0.182 ;
      RECT 4.394 0.448 4.462 0.492 ;
      RECT 4.286 0.138 4.354 0.182 ;
      RECT 4.286 0.448 4.354 0.492 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 3.962 0.138 4.03 0.182 ;
      RECT 3.962 0.448 4.03 0.492 ;
      RECT 3.854 0.338 3.922 0.382 ;
      RECT 3.746 0.138 3.814 0.182 ;
      RECT 3.746 0.473 3.814 0.517 ;
      RECT 3.53 0.248 3.598 0.292 ;
      RECT 3.422 0.1515 3.49 0.1955 ;
      RECT 3.422 0.47 3.49 0.514 ;
      RECT 3.314 0.1515 3.382 0.1955 ;
      RECT 3.314 0.47 3.382 0.514 ;
      RECT 3.206 0.47 3.274 0.514 ;
      RECT 3.208 0.268 3.272 0.312 ;
      RECT 2.774 0.203 2.842 0.247 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.203 2.194 0.247 ;
      RECT 1.802 0.138 1.87 0.182 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.694 0.292 1.762 0.336 ;
      RECT 1.586 0.1515 1.654 0.1955 ;
      RECT 1.586 0.453 1.654 0.497 ;
      RECT 1.478 0.1515 1.546 0.1955 ;
      RECT 1.478 0.453 1.546 0.497 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.113 1.222 0.157 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.113 1.006 0.157 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.29 0.448 0.358 0.492 ;
      RECT 0.182 0.293 0.25 0.337 ;
    LAYER m1 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.248 1.35 0.292 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 2.194 0.428 2.41 0.472 ;
      RECT 2.774 0.158 2.842 0.472 ;
      RECT 3.166 0.338 3.206 0.382 ;
      RECT 3.206 0.248 3.274 0.382 ;
  END
END b15fpy200hn1n04x5

MACRO b15fpy200hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy200hn1n08x5 0 0 ;
  SIZE 5.832 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.068 2.086 0.382 ;
      LAYER v0 ;
        RECT 2.018 0.3155 2.086 0.3595 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.068 3.814 0.382 ;
      LAYER v0 ;
        RECT 3.746 0.3155 3.814 0.3595 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.068 2.302 0.382 ;
      LAYER v0 ;
        RECT 2.234 0.3155 2.302 0.3595 ;
    END
  END d2
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.582 0.068 5.65 0.562 ;
      LAYER v0 ;
        RECT 5.582 0.448 5.65 0.492 ;
        RECT 5.582 0.138 5.65 0.182 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o2
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.078 0.248 3.274 0.292 ;
        RECT 3.206 0.068 3.274 0.292 ;
      LAYER v0 ;
        RECT 3.098 0.248 3.166 0.292 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.248 2.862 0.292 ;
        RECT 2.666 0.068 2.734 0.292 ;
      LAYER v0 ;
        RECT 2.774 0.248 2.842 0.292 ;
    END
  END si2
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.598 0.382 ;
        RECT 3.314 0.068 3.598 0.112 ;
        RECT 2.558 0.338 3.382 0.382 ;
        RECT 3.314 0.068 3.382 0.382 ;
        RECT 2.558 0.068 2.626 0.382 ;
        RECT 2.342 0.068 2.626 0.112 ;
        RECT 2.342 0.068 2.41 0.382 ;
      LAYER v0 ;
        RECT 2.342 0.3155 2.41 0.3595 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 2.99 0.338 3.058 0.382 ;
        RECT 3.206 0.338 3.274 0.382 ;
        RECT 3.53 0.3155 3.598 0.3595 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.866 0.652 ;
        RECT 5.69 0.428 5.758 0.652 ;
        RECT 5.474 0.428 5.542 0.652 ;
        RECT 5.258 0.428 5.326 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 2.126 0.538 2.194 0.582 ;
        RECT 2.774 0.452 2.842 0.496 ;
        RECT 3.098 0.452 3.166 0.496 ;
        RECT 3.746 0.538 3.814 0.582 ;
        RECT 4.61 0.448 4.678 0.492 ;
        RECT 5.258 0.448 5.326 0.492 ;
        RECT 5.474 0.448 5.542 0.492 ;
        RECT 5.69 0.448 5.758 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.866 0.022 ;
        RECT 5.69 -0.022 5.758 0.202 ;
        RECT 5.474 -0.022 5.542 0.202 ;
        RECT 5.258 -0.022 5.326 0.202 ;
        RECT 4.61 -0.022 4.678 0.202 ;
        RECT 3.854 -0.022 3.922 0.202 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.774 0.114 2.842 0.158 ;
        RECT 3.098 0.114 3.166 0.158 ;
        RECT 3.854 0.138 3.922 0.182 ;
        RECT 4.61 0.138 4.678 0.182 ;
        RECT 5.258 0.138 5.326 0.182 ;
        RECT 5.474 0.138 5.542 0.182 ;
        RECT 5.69 0.138 5.758 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.596 0.338 5.236 0.382 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.248 0.682 0.382 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.694 0.248 1.762 0.382 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.91 0.068 1.978 0.472 ;
      RECT 3.294 0.428 3.422 0.472 ;
      RECT 3.854 0.248 3.922 0.382 ;
      RECT 3.962 0.068 4.03 0.472 ;
      RECT 4.07 0.158 4.138 0.382 ;
      RECT 4.502 0.158 4.57 0.382 ;
      RECT 4.286 0.068 4.354 0.562 ;
      RECT 4.394 0.248 4.462 0.472 ;
      RECT 4.826 0.518 5.042 0.562 ;
      RECT 4.826 0.248 4.894 0.472 ;
      RECT 5.15 0.248 5.218 0.382 ;
      RECT 5.366 0.068 5.434 0.562 ;
    LAYER v1 ;
      RECT 5.154 0.338 5.214 0.382 ;
      RECT 4.83 0.338 4.89 0.382 ;
      RECT 4.398 0.338 4.458 0.382 ;
      RECT 4.074 0.338 4.134 0.382 ;
      RECT 3.858 0.338 3.918 0.382 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.618 0.338 0.678 0.382 ;
    LAYER v0 ;
      RECT 5.366 0.138 5.434 0.182 ;
      RECT 5.366 0.448 5.434 0.492 ;
      RECT 5.15 0.293 5.218 0.337 ;
      RECT 5.042 0.1505 5.11 0.1945 ;
      RECT 4.934 0.518 5.002 0.562 ;
      RECT 4.826 0.338 4.894 0.382 ;
      RECT 4.718 0.138 4.786 0.182 ;
      RECT 4.718 0.448 4.786 0.492 ;
      RECT 4.502 0.248 4.57 0.292 ;
      RECT 4.394 0.338 4.462 0.382 ;
      RECT 4.286 0.1575 4.354 0.2015 ;
      RECT 4.286 0.428 4.354 0.472 ;
      RECT 4.178 0.1575 4.246 0.2015 ;
      RECT 4.178 0.428 4.246 0.472 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 3.962 0.138 4.03 0.182 ;
      RECT 3.962 0.408 4.03 0.452 ;
      RECT 3.854 0.3155 3.922 0.3595 ;
      RECT 3.422 0.178 3.49 0.222 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.45 0.178 2.518 0.222 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.3155 1.762 0.3595 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.1605 0.79 0.2045 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.79 0.518 1.006 0.562 ;
      RECT 1.114 0.338 1.262 0.382 ;
      RECT 1.262 0.158 1.33 0.382 ;
      RECT 1.546 0.158 1.762 0.202 ;
      RECT 1.654 0.518 1.802 0.562 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.87 0.518 2.018 0.562 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 2.086 0.428 2.45 0.472 ;
      RECT 2.45 0.158 2.518 0.472 ;
      RECT 2.518 0.428 2.646 0.472 ;
      RECT 3.422 0.158 3.49 0.472 ;
      RECT 3.49 0.428 3.854 0.472 ;
      RECT 3.854 0.428 3.922 0.562 ;
      RECT 3.922 0.518 4.178 0.562 ;
      RECT 4.178 0.068 4.246 0.562 ;
      RECT 4.57 0.338 4.718 0.382 ;
      RECT 4.718 0.068 4.786 0.562 ;
      RECT 5.042 0.068 5.11 0.562 ;
  END
END b15fpy200hn1n08x5

MACRO b15fpy400hn1d02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy400hn1d02x5 0 0 ;
  SIZE 4.536 BY 1.26 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.338 1.762 0.382 ;
        RECT 1.478 0.158 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.248 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.338 2.734 0.382 ;
    END
  END d2
  PIN d3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.788 2.734 1.102 ;
      LAYER v0 ;
        RECT 2.666 0.878 2.734 0.922 ;
    END
  END d3
  PIN d4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.788 1.87 1.102 ;
      LAYER v0 ;
        RECT 1.802 0.878 1.87 0.922 ;
    END
  END d4
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.068 4.462 0.562 ;
      LAYER v0 ;
        RECT 4.394 0.453 4.462 0.497 ;
        RECT 4.394 0.138 4.462 0.182 ;
    END
  END o2
  PIN o3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.698 4.462 1.192 ;
      LAYER v0 ;
        RECT 4.394 1.103 4.462 1.147 ;
        RECT 4.394 0.768 4.462 0.812 ;
    END
  END o3
  PIN o4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.698 0.142 1.192 ;
      LAYER v0 ;
        RECT 0.074 1.078 0.142 1.122 ;
        RECT 0.074 0.768 0.142 0.812 ;
    END
  END o4
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.292 ;
      LAYER v0 ;
        RECT 2.126 0.088 2.194 0.132 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.292 ;
      LAYER v0 ;
        RECT 2.342 0.088 2.41 0.132 ;
    END
  END si2
  PIN si3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.968 2.41 1.192 ;
      LAYER v0 ;
        RECT 2.342 1.013 2.41 1.057 ;
    END
  END si3
  PIN si4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.968 2.194 1.192 ;
      LAYER v0 ;
        RECT 2.126 1.013 2.194 1.057 ;
    END
  END si4
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 11.2538385 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 9.54822225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.734 0.112 ;
        RECT 1.91 0.518 2.518 0.562 ;
        RECT 2.018 0.338 2.518 0.382 ;
        RECT 2.45 0.068 2.518 0.382 ;
        RECT 2.234 0.338 2.302 0.562 ;
        RECT 2.018 0.068 2.086 0.382 ;
        RECT 1.802 0.068 2.086 0.112 ;
        RECT 2.45 1.148 2.734 1.192 ;
        RECT 2.45 0.878 2.518 1.192 ;
        RECT 2.018 0.878 2.518 0.922 ;
        RECT 1.802 1.148 2.086 1.192 ;
        RECT 2.018 0.878 2.086 1.192 ;
      LAYER v0 ;
        RECT 1.91 1.148 1.978 1.192 ;
        RECT 1.91 0.068 1.978 0.112 ;
        RECT 2.126 0.878 2.194 0.922 ;
        RECT 2.126 0.518 2.194 0.562 ;
        RECT 2.342 0.878 2.41 0.922 ;
        RECT 2.342 0.518 2.41 0.562 ;
        RECT 2.558 1.148 2.626 1.192 ;
        RECT 2.558 0.068 2.626 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.57 0.652 ;
        RECT 4.286 0.518 4.354 0.742 ;
        RECT 3.962 0.518 4.03 0.832 ;
        RECT 3.422 0.428 3.49 0.832 ;
        RECT 1.694 0.428 1.762 0.832 ;
        RECT 1.046 0.428 1.114 0.832 ;
        RECT 0.506 0.428 0.574 0.832 ;
        RECT 0.182 0.518 0.25 0.742 ;
      LAYER v0 ;
        RECT 0.182 0.678 0.25 0.722 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.506 0.724 0.574 0.768 ;
        RECT 0.506 0.493 0.574 0.537 ;
        RECT 1.046 0.743 1.114 0.787 ;
        RECT 1.046 0.473 1.114 0.517 ;
        RECT 1.694 0.763 1.762 0.807 ;
        RECT 1.694 0.498 1.762 0.542 ;
        RECT 2.234 0.608 2.302 0.652 ;
        RECT 2.774 0.608 2.842 0.652 ;
        RECT 3.422 0.743 3.49 0.787 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 3.962 0.768 4.03 0.812 ;
        RECT 4.286 0.678 4.354 0.722 ;
        RECT 4.286 0.538 4.354 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.57 0.022 ;
        RECT 4.286 -0.022 4.354 0.202 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.234 -0.022 2.302 0.292 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
        RECT -0.034 1.238 4.57 1.282 ;
        RECT 4.286 1.058 4.354 1.282 ;
        RECT 3.962 1.058 4.03 1.282 ;
        RECT 3.422 1.058 3.49 1.282 ;
        RECT 2.774 1.058 2.842 1.282 ;
        RECT 2.234 1.148 2.302 1.282 ;
        RECT 1.694 0.968 1.762 1.282 ;
        RECT 1.046 1.058 1.114 1.282 ;
        RECT 0.506 1.058 0.574 1.282 ;
        RECT 0.182 1.058 0.25 1.282 ;
      LAYER v0 ;
        RECT 0.182 1.078 0.25 1.122 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.506 1.078 0.574 1.122 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.046 1.103 1.114 1.147 ;
        RECT 1.046 0.113 1.114 0.157 ;
        RECT 1.694 1.033 1.762 1.077 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 2.236 1.168 2.3 1.212 ;
        RECT 2.234 0.222 2.302 0.266 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.774 1.078 2.842 1.122 ;
        RECT 3.422 1.078 3.49 1.122 ;
        RECT 3.422 0.048 3.49 0.092 ;
        RECT 3.962 1.103 4.03 1.147 ;
        RECT 3.962 0.138 4.03 0.182 ;
        RECT 4.286 1.103 4.354 1.147 ;
        RECT 4.286 0.138 4.354 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.878 0.808 0.922 ;
      RECT 0.164 0.428 0.824 0.472 ;
      RECT 1.352 0.878 1.996 0.922 ;
      RECT 2.54 0.878 3.184 0.922 ;
      RECT 0.904 0.428 3.74 0.472 ;
      RECT 0.596 0.788 3.94 0.832 ;
      RECT 0.38 0.698 4.156 0.742 ;
      RECT 3.728 0.878 4.372 0.922 ;
      RECT 3.82 0.428 4.372 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.878 0.25 1.012 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.29 0.698 0.358 1.192 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.398 0.698 0.466 1.192 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.788 0.682 1.102 ;
      RECT 0.722 0.698 0.79 1.192 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.83 0.698 0.898 1.012 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 1.026 0.878 1.262 0.922 ;
      RECT 0.938 0.338 1.262 0.382 ;
      RECT 1.91 0.788 1.978 1.102 ;
      RECT 1.37 0.698 1.438 1.192 ;
      RECT 1.478 0.698 1.546 0.832 ;
      RECT 1.586 0.698 1.654 1.102 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 2.342 0.788 2.558 0.832 ;
      RECT 1.802 0.698 2.774 0.742 ;
      RECT 2.882 0.788 2.95 0.922 ;
      RECT 2.342 0.428 2.558 0.472 ;
      RECT 2.99 0.698 3.058 0.832 ;
      RECT 2.99 0.248 3.058 0.472 ;
      RECT 3.098 0.698 3.166 1.192 ;
      RECT 3.422 0.158 3.49 0.382 ;
      RECT 3.206 0.698 3.274 1.192 ;
      RECT 3.206 0.068 3.274 0.562 ;
      RECT 3.314 0.698 3.382 1.102 ;
      RECT 3.314 0.248 3.382 0.472 ;
      RECT 3.53 0.698 3.598 1.192 ;
      RECT 3.746 0.068 3.814 0.562 ;
      RECT 3.638 0.788 3.706 1.012 ;
      RECT 3.638 0.248 3.706 0.472 ;
      RECT 3.746 0.698 3.814 1.192 ;
      RECT 3.854 0.788 3.922 1.102 ;
      RECT 4.07 0.698 4.138 1.192 ;
      RECT 4.07 0.068 4.138 0.472 ;
      RECT 4.178 0.698 4.246 1.192 ;
      RECT 4.178 0.068 4.246 0.562 ;
      RECT 4.286 0.788 4.354 1.012 ;
      RECT 4.286 0.248 4.354 0.472 ;
    LAYER v1 ;
      RECT 4.29 0.428 4.35 0.472 ;
      RECT 4.29 0.878 4.35 0.922 ;
      RECT 4.074 0.698 4.134 0.742 ;
      RECT 3.858 0.428 3.918 0.472 ;
      RECT 3.858 0.788 3.918 0.832 ;
      RECT 3.75 0.878 3.81 0.922 ;
      RECT 3.642 0.428 3.702 0.472 ;
      RECT 3.642 0.788 3.702 0.832 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 3.318 0.698 3.378 0.742 ;
      RECT 3.102 0.878 3.162 0.922 ;
      RECT 2.994 0.428 3.054 0.472 ;
      RECT 2.994 0.698 3.054 0.742 ;
      RECT 2.886 0.788 2.946 0.832 ;
      RECT 2.562 0.878 2.622 0.922 ;
      RECT 1.914 0.878 1.974 0.922 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.59 0.698 1.65 0.742 ;
      RECT 1.482 0.788 1.542 0.832 ;
      RECT 1.374 0.878 1.434 0.922 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.726 0.428 0.786 0.472 ;
      RECT 0.726 0.878 0.786 0.922 ;
      RECT 0.618 0.788 0.678 0.832 ;
      RECT 0.402 0.698 0.462 0.742 ;
      RECT 0.186 0.428 0.246 0.472 ;
      RECT 0.186 0.878 0.246 0.922 ;
    LAYER v0 ;
      RECT 4.286 0.3605 4.354 0.4045 ;
      RECT 4.286 0.878 4.354 0.922 ;
      RECT 4.178 0.138 4.246 0.182 ;
      RECT 4.178 0.453 4.246 0.497 ;
      RECT 4.178 0.768 4.246 0.812 ;
      RECT 4.178 1.103 4.246 1.147 ;
      RECT 4.07 0.138 4.138 0.182 ;
      RECT 4.07 0.3695 4.138 0.4135 ;
      RECT 4.07 0.768 4.138 0.812 ;
      RECT 4.07 1.103 4.138 1.147 ;
      RECT 3.854 0.968 3.922 1.012 ;
      RECT 3.746 0.138 3.814 0.182 ;
      RECT 3.746 0.768 3.814 0.812 ;
      RECT 3.746 1.078 3.814 1.122 ;
      RECT 3.748 0.498 3.812 0.542 ;
      RECT 3.638 0.338 3.706 0.382 ;
      RECT 3.638 0.878 3.706 0.922 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.53 0.743 3.598 0.787 ;
      RECT 3.53 1.078 3.598 1.122 ;
      RECT 3.422 0.248 3.49 0.292 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 3.314 0.968 3.382 1.012 ;
      RECT 3.206 0.1515 3.274 0.1955 ;
      RECT 3.206 0.47 3.274 0.514 ;
      RECT 3.206 0.746 3.274 0.79 ;
      RECT 3.206 1.0645 3.274 1.1085 ;
      RECT 3.098 0.1515 3.166 0.1955 ;
      RECT 3.098 0.47 3.166 0.514 ;
      RECT 3.098 0.746 3.166 0.79 ;
      RECT 3.098 1.0645 3.166 1.1085 ;
      RECT 2.99 0.293 3.058 0.337 ;
      RECT 2.99 0.746 3.058 0.79 ;
      RECT 2.992 0.948 3.056 0.992 ;
      RECT 2.882 1.078 2.95 1.122 ;
      RECT 2.558 1.013 2.626 1.057 ;
      RECT 2.56 0.228 2.624 0.272 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.45 0.698 2.518 0.742 ;
      RECT 2.45 0.788 2.518 0.832 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 2.018 0.788 2.086 0.832 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.91 0.698 1.978 0.742 ;
      RECT 1.91 1.013 1.978 1.057 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.586 0.763 1.654 0.807 ;
      RECT 1.586 1.033 1.654 1.077 ;
      RECT 1.478 0.763 1.546 0.807 ;
      RECT 1.37 0.1515 1.438 0.1955 ;
      RECT 1.37 0.453 1.438 0.497 ;
      RECT 1.37 0.763 1.438 0.807 ;
      RECT 1.37 1.0645 1.438 1.1085 ;
      RECT 1.262 0.1515 1.33 0.1955 ;
      RECT 1.262 0.453 1.33 0.497 ;
      RECT 1.262 0.763 1.33 0.807 ;
      RECT 1.262 1.0645 1.33 1.1085 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 1.046 0.878 1.114 0.922 ;
      RECT 1.046 0.968 1.114 1.012 ;
      RECT 0.938 0.113 1.006 0.157 ;
      RECT 0.938 1.103 1.006 1.147 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.83 0.763 0.898 0.807 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.408 0.79 0.452 ;
      RECT 0.722 0.763 0.79 0.807 ;
      RECT 0.722 1.078 0.79 1.122 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.614 0.923 0.682 0.967 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.493 0.466 0.537 ;
      RECT 0.398 0.724 0.466 0.768 ;
      RECT 0.398 1.078 0.466 1.122 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.29 0.3855 0.358 0.4295 ;
      RECT 0.29 0.8305 0.358 0.8745 ;
      RECT 0.29 1.078 0.358 1.122 ;
      RECT 0.182 0.293 0.25 0.337 ;
      RECT 0.182 0.923 0.25 0.967 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.898 0.968 0.938 1.012 ;
      RECT 0.938 0.968 1.006 1.192 ;
      RECT 1.006 0.968 1.134 1.012 ;
      RECT 0.898 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.006 0.248 1.134 0.292 ;
      RECT 1.262 0.698 1.33 1.192 ;
      RECT 1.262 0.068 1.33 0.562 ;
      RECT 1.978 0.788 2.194 0.832 ;
      RECT 1.438 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.202 ;
      RECT 1.654 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.472 ;
      RECT 1.978 0.428 2.194 0.472 ;
      RECT 2.558 0.788 2.626 1.102 ;
      RECT 2.774 0.698 2.842 1.012 ;
      RECT 2.842 0.968 2.882 1.012 ;
      RECT 2.882 0.968 2.95 1.192 ;
      RECT 2.95 0.878 2.99 0.922 ;
      RECT 2.99 0.878 3.058 1.012 ;
      RECT 2.558 0.158 2.626 0.472 ;
      RECT 2.626 0.158 2.882 0.202 ;
      RECT 2.882 0.068 2.95 0.202 ;
      RECT 2.95 0.068 3.098 0.112 ;
      RECT 3.098 0.068 3.166 0.562 ;
      RECT 3.49 0.338 3.53 0.382 ;
      RECT 3.53 0.338 3.598 0.562 ;
      RECT 3.814 0.428 4.03 0.472 ;
  END
END b15fpy400hn1d02x5

MACRO b15fpy400hn1d03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy400hn1d03x5 0 0 ;
  SIZE 4.536 BY 1.26 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.338 1.762 0.382 ;
        RECT 1.478 0.158 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.248 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.338 2.734 0.382 ;
    END
  END d2
  PIN d3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.788 2.734 1.102 ;
      LAYER v0 ;
        RECT 2.666 0.878 2.734 0.922 ;
    END
  END d3
  PIN d4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.788 1.87 1.102 ;
      LAYER v0 ;
        RECT 1.802 0.878 1.87 0.922 ;
    END
  END d4
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.068 4.462 0.562 ;
      LAYER v0 ;
        RECT 4.394 0.453 4.462 0.497 ;
        RECT 4.394 0.138 4.462 0.182 ;
    END
  END o2
  PIN o3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.698 4.462 1.192 ;
      LAYER v0 ;
        RECT 4.394 1.103 4.462 1.147 ;
        RECT 4.394 0.768 4.462 0.812 ;
    END
  END o3
  PIN o4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.698 0.142 1.192 ;
      LAYER v0 ;
        RECT 0.074 1.078 0.142 1.122 ;
        RECT 0.074 0.768 0.142 0.812 ;
    END
  END o4
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.292 ;
      LAYER v0 ;
        RECT 2.126 0.088 2.194 0.132 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.292 ;
      LAYER v0 ;
        RECT 2.342 0.088 2.41 0.132 ;
    END
  END si2
  PIN si3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.968 2.41 1.192 ;
      LAYER v0 ;
        RECT 2.342 1.013 2.41 1.057 ;
    END
  END si3
  PIN si4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.968 2.194 1.192 ;
      LAYER v0 ;
        RECT 2.126 1.013 2.194 1.057 ;
    END
  END si4
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 11.2538385 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 9.54822225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.734 0.112 ;
        RECT 1.91 0.518 2.518 0.562 ;
        RECT 2.018 0.338 2.518 0.382 ;
        RECT 2.45 0.068 2.518 0.382 ;
        RECT 2.234 0.338 2.302 0.562 ;
        RECT 2.018 0.068 2.086 0.382 ;
        RECT 1.802 0.068 2.086 0.112 ;
        RECT 2.45 1.148 2.734 1.192 ;
        RECT 2.45 0.878 2.518 1.192 ;
        RECT 2.018 0.878 2.518 0.922 ;
        RECT 1.802 1.148 2.086 1.192 ;
        RECT 2.018 0.878 2.086 1.192 ;
      LAYER v0 ;
        RECT 1.91 1.148 1.978 1.192 ;
        RECT 1.91 0.068 1.978 0.112 ;
        RECT 2.126 0.878 2.194 0.922 ;
        RECT 2.126 0.518 2.194 0.562 ;
        RECT 2.342 0.878 2.41 0.922 ;
        RECT 2.342 0.518 2.41 0.562 ;
        RECT 2.558 1.148 2.626 1.192 ;
        RECT 2.558 0.068 2.626 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.57 0.652 ;
        RECT 4.286 0.518 4.354 0.742 ;
        RECT 3.962 0.518 4.03 0.832 ;
        RECT 3.422 0.428 3.49 0.832 ;
        RECT 1.694 0.428 1.762 0.832 ;
        RECT 1.046 0.428 1.114 0.832 ;
        RECT 0.506 0.428 0.574 0.832 ;
        RECT 0.182 0.518 0.25 0.742 ;
      LAYER v0 ;
        RECT 0.182 0.678 0.25 0.722 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.506 0.724 0.574 0.768 ;
        RECT 0.506 0.493 0.574 0.537 ;
        RECT 1.046 0.743 1.114 0.787 ;
        RECT 1.046 0.473 1.114 0.517 ;
        RECT 1.694 0.763 1.762 0.807 ;
        RECT 1.694 0.498 1.762 0.542 ;
        RECT 2.234 0.608 2.302 0.652 ;
        RECT 2.774 0.608 2.842 0.652 ;
        RECT 3.422 0.743 3.49 0.787 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 3.962 0.768 4.03 0.812 ;
        RECT 4.286 0.678 4.354 0.722 ;
        RECT 4.286 0.538 4.354 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.57 0.022 ;
        RECT 4.286 -0.022 4.354 0.202 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.234 -0.022 2.302 0.292 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
        RECT -0.034 1.238 4.57 1.282 ;
        RECT 4.286 1.058 4.354 1.282 ;
        RECT 3.962 1.058 4.03 1.282 ;
        RECT 3.422 1.058 3.49 1.282 ;
        RECT 2.774 1.058 2.842 1.282 ;
        RECT 2.234 1.148 2.302 1.282 ;
        RECT 1.694 0.968 1.762 1.282 ;
        RECT 1.046 1.058 1.114 1.282 ;
        RECT 0.506 1.058 0.574 1.282 ;
        RECT 0.182 1.058 0.25 1.282 ;
      LAYER v0 ;
        RECT 0.182 1.078 0.25 1.122 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.506 1.078 0.574 1.122 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.046 1.103 1.114 1.147 ;
        RECT 1.046 0.113 1.114 0.157 ;
        RECT 1.694 1.033 1.762 1.077 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 2.236 1.168 2.3 1.212 ;
        RECT 2.234 0.222 2.302 0.266 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.774 1.078 2.842 1.122 ;
        RECT 3.422 1.078 3.49 1.122 ;
        RECT 3.422 0.048 3.49 0.092 ;
        RECT 3.962 1.103 4.03 1.147 ;
        RECT 3.962 0.138 4.03 0.182 ;
        RECT 4.286 1.103 4.354 1.147 ;
        RECT 4.286 0.138 4.354 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.878 0.808 0.922 ;
      RECT 0.164 0.428 0.824 0.472 ;
      RECT 1.352 0.878 1.996 0.922 ;
      RECT 2.54 0.878 3.184 0.922 ;
      RECT 0.904 0.428 3.74 0.472 ;
      RECT 0.596 0.788 3.94 0.832 ;
      RECT 0.38 0.698 4.156 0.742 ;
      RECT 3.728 0.878 4.372 0.922 ;
      RECT 3.82 0.428 4.372 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.878 0.25 1.012 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.29 0.698 0.358 1.192 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.398 0.698 0.466 1.192 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.788 0.682 1.102 ;
      RECT 0.722 0.698 0.79 1.192 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.83 0.698 0.898 1.012 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 1.026 0.878 1.262 0.922 ;
      RECT 0.938 0.338 1.262 0.382 ;
      RECT 1.91 0.788 1.978 1.102 ;
      RECT 1.37 0.698 1.438 1.192 ;
      RECT 1.478 0.698 1.546 0.832 ;
      RECT 1.586 0.698 1.654 1.102 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 2.342 0.788 2.558 0.832 ;
      RECT 1.802 0.698 2.774 0.742 ;
      RECT 2.882 0.788 2.95 0.922 ;
      RECT 2.342 0.428 2.558 0.472 ;
      RECT 2.99 0.698 3.058 0.832 ;
      RECT 2.99 0.248 3.058 0.472 ;
      RECT 3.098 0.698 3.166 1.192 ;
      RECT 3.422 0.158 3.49 0.382 ;
      RECT 3.206 0.698 3.274 1.192 ;
      RECT 3.206 0.068 3.274 0.562 ;
      RECT 3.314 0.698 3.382 1.102 ;
      RECT 3.314 0.248 3.382 0.472 ;
      RECT 3.53 0.698 3.598 1.192 ;
      RECT 3.746 0.068 3.814 0.562 ;
      RECT 3.638 0.788 3.706 1.012 ;
      RECT 3.638 0.248 3.706 0.472 ;
      RECT 3.746 0.698 3.814 1.192 ;
      RECT 3.854 0.788 3.922 1.102 ;
      RECT 4.07 0.698 4.138 1.192 ;
      RECT 4.07 0.068 4.138 0.472 ;
      RECT 4.178 0.698 4.246 1.192 ;
      RECT 4.178 0.068 4.246 0.562 ;
      RECT 4.286 0.788 4.354 1.012 ;
      RECT 4.286 0.248 4.354 0.472 ;
    LAYER v1 ;
      RECT 4.29 0.428 4.35 0.472 ;
      RECT 4.29 0.878 4.35 0.922 ;
      RECT 4.074 0.698 4.134 0.742 ;
      RECT 3.858 0.428 3.918 0.472 ;
      RECT 3.858 0.788 3.918 0.832 ;
      RECT 3.75 0.878 3.81 0.922 ;
      RECT 3.642 0.428 3.702 0.472 ;
      RECT 3.642 0.788 3.702 0.832 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 3.318 0.698 3.378 0.742 ;
      RECT 3.102 0.878 3.162 0.922 ;
      RECT 2.994 0.428 3.054 0.472 ;
      RECT 2.994 0.698 3.054 0.742 ;
      RECT 2.886 0.788 2.946 0.832 ;
      RECT 2.562 0.878 2.622 0.922 ;
      RECT 1.914 0.878 1.974 0.922 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.59 0.698 1.65 0.742 ;
      RECT 1.482 0.788 1.542 0.832 ;
      RECT 1.374 0.878 1.434 0.922 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.726 0.428 0.786 0.472 ;
      RECT 0.726 0.878 0.786 0.922 ;
      RECT 0.618 0.788 0.678 0.832 ;
      RECT 0.402 0.698 0.462 0.742 ;
      RECT 0.186 0.428 0.246 0.472 ;
      RECT 0.186 0.878 0.246 0.922 ;
    LAYER v0 ;
      RECT 4.286 0.338 4.354 0.382 ;
      RECT 4.286 0.878 4.354 0.922 ;
      RECT 4.178 0.138 4.246 0.182 ;
      RECT 4.178 0.453 4.246 0.497 ;
      RECT 4.178 0.768 4.246 0.812 ;
      RECT 4.178 1.103 4.246 1.147 ;
      RECT 4.07 0.138 4.138 0.182 ;
      RECT 4.07 0.3695 4.138 0.4135 ;
      RECT 4.07 0.768 4.138 0.812 ;
      RECT 4.07 1.103 4.138 1.147 ;
      RECT 3.854 0.968 3.922 1.012 ;
      RECT 3.746 0.138 3.814 0.182 ;
      RECT 3.746 0.768 3.814 0.812 ;
      RECT 3.746 1.078 3.814 1.122 ;
      RECT 3.748 0.498 3.812 0.542 ;
      RECT 3.638 0.338 3.706 0.382 ;
      RECT 3.638 0.878 3.706 0.922 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.53 0.743 3.598 0.787 ;
      RECT 3.53 1.078 3.598 1.122 ;
      RECT 3.422 0.248 3.49 0.292 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 3.314 0.968 3.382 1.012 ;
      RECT 3.206 0.1515 3.274 0.1955 ;
      RECT 3.206 0.47 3.274 0.514 ;
      RECT 3.206 0.746 3.274 0.79 ;
      RECT 3.206 1.0645 3.274 1.1085 ;
      RECT 3.098 0.1515 3.166 0.1955 ;
      RECT 3.098 0.47 3.166 0.514 ;
      RECT 3.098 0.746 3.166 0.79 ;
      RECT 3.098 1.0645 3.166 1.1085 ;
      RECT 2.99 0.293 3.058 0.337 ;
      RECT 2.99 0.746 3.058 0.79 ;
      RECT 2.992 0.948 3.056 0.992 ;
      RECT 2.882 1.078 2.95 1.122 ;
      RECT 2.558 1.013 2.626 1.057 ;
      RECT 2.56 0.228 2.624 0.272 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.45 0.698 2.518 0.742 ;
      RECT 2.45 0.788 2.518 0.832 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 2.018 0.788 2.086 0.832 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.91 0.698 1.978 0.742 ;
      RECT 1.91 1.013 1.978 1.057 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.586 0.763 1.654 0.807 ;
      RECT 1.586 1.033 1.654 1.077 ;
      RECT 1.478 0.763 1.546 0.807 ;
      RECT 1.37 0.1515 1.438 0.1955 ;
      RECT 1.37 0.453 1.438 0.497 ;
      RECT 1.37 0.763 1.438 0.807 ;
      RECT 1.37 1.0645 1.438 1.1085 ;
      RECT 1.262 0.1515 1.33 0.1955 ;
      RECT 1.262 0.453 1.33 0.497 ;
      RECT 1.262 0.763 1.33 0.807 ;
      RECT 1.262 1.0645 1.33 1.1085 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 1.046 0.878 1.114 0.922 ;
      RECT 1.046 0.968 1.114 1.012 ;
      RECT 0.938 0.113 1.006 0.157 ;
      RECT 0.938 1.103 1.006 1.147 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.83 0.763 0.898 0.807 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.408 0.79 0.452 ;
      RECT 0.722 0.763 0.79 0.807 ;
      RECT 0.722 1.078 0.79 1.122 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.614 0.923 0.682 0.967 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.493 0.466 0.537 ;
      RECT 0.398 0.724 0.466 0.768 ;
      RECT 0.398 1.078 0.466 1.122 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.29 0.3855 0.358 0.4295 ;
      RECT 0.29 0.8305 0.358 0.8745 ;
      RECT 0.29 1.078 0.358 1.122 ;
      RECT 0.182 0.293 0.25 0.337 ;
      RECT 0.182 0.923 0.25 0.967 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.898 0.968 0.938 1.012 ;
      RECT 0.938 0.968 1.006 1.192 ;
      RECT 1.006 0.968 1.134 1.012 ;
      RECT 0.898 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.006 0.248 1.134 0.292 ;
      RECT 1.262 0.698 1.33 1.192 ;
      RECT 1.262 0.068 1.33 0.562 ;
      RECT 1.978 0.788 2.194 0.832 ;
      RECT 1.438 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.202 ;
      RECT 1.654 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.472 ;
      RECT 1.978 0.428 2.194 0.472 ;
      RECT 2.558 0.788 2.626 1.102 ;
      RECT 2.774 0.698 2.842 1.012 ;
      RECT 2.842 0.968 2.882 1.012 ;
      RECT 2.882 0.968 2.95 1.192 ;
      RECT 2.95 0.878 2.99 0.922 ;
      RECT 2.99 0.878 3.058 1.012 ;
      RECT 2.558 0.158 2.626 0.472 ;
      RECT 2.626 0.158 2.882 0.202 ;
      RECT 2.882 0.068 2.95 0.202 ;
      RECT 2.95 0.068 3.098 0.112 ;
      RECT 3.098 0.068 3.166 0.562 ;
      RECT 3.49 0.338 3.53 0.382 ;
      RECT 3.53 0.338 3.598 0.562 ;
      RECT 3.814 0.428 4.03 0.472 ;
  END
END b15fpy400hn1d03x5

MACRO b15fpy400hn1d04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy400hn1d04x5 0 0 ;
  SIZE 4.536 BY 1.26 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.338 1.762 0.382 ;
        RECT 1.478 0.158 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.248 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.338 2.734 0.382 ;
    END
  END d2
  PIN d3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.788 2.734 1.102 ;
      LAYER v0 ;
        RECT 2.666 0.878 2.734 0.922 ;
    END
  END d3
  PIN d4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.788 1.87 1.102 ;
      LAYER v0 ;
        RECT 1.802 0.878 1.87 0.922 ;
    END
  END d4
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.068 4.462 0.562 ;
      LAYER v0 ;
        RECT 4.394 0.453 4.462 0.497 ;
        RECT 4.394 0.138 4.462 0.182 ;
    END
  END o2
  PIN o3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.698 4.462 1.192 ;
      LAYER v0 ;
        RECT 4.394 1.103 4.462 1.147 ;
        RECT 4.394 0.768 4.462 0.812 ;
    END
  END o3
  PIN o4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.698 0.142 1.192 ;
      LAYER v0 ;
        RECT 0.074 1.078 0.142 1.122 ;
        RECT 0.074 0.768 0.142 0.812 ;
    END
  END o4
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.292 ;
      LAYER v0 ;
        RECT 2.126 0.088 2.194 0.132 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.292 ;
      LAYER v0 ;
        RECT 2.342 0.088 2.41 0.132 ;
    END
  END si2
  PIN si3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.968 2.41 1.192 ;
      LAYER v0 ;
        RECT 2.342 1.013 2.41 1.057 ;
    END
  END si3
  PIN si4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.968 2.194 1.192 ;
      LAYER v0 ;
        RECT 2.126 1.013 2.194 1.057 ;
    END
  END si4
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 11.2538385 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 9.54822225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.734 0.112 ;
        RECT 1.91 0.518 2.518 0.562 ;
        RECT 2.018 0.338 2.518 0.382 ;
        RECT 2.45 0.068 2.518 0.382 ;
        RECT 2.234 0.338 2.302 0.562 ;
        RECT 2.018 0.068 2.086 0.382 ;
        RECT 1.802 0.068 2.086 0.112 ;
        RECT 2.45 1.148 2.734 1.192 ;
        RECT 2.45 0.878 2.518 1.192 ;
        RECT 2.018 0.878 2.518 0.922 ;
        RECT 1.802 1.148 2.086 1.192 ;
        RECT 2.018 0.878 2.086 1.192 ;
      LAYER v0 ;
        RECT 1.91 1.148 1.978 1.192 ;
        RECT 1.91 0.068 1.978 0.112 ;
        RECT 2.126 0.878 2.194 0.922 ;
        RECT 2.126 0.518 2.194 0.562 ;
        RECT 2.342 0.878 2.41 0.922 ;
        RECT 2.342 0.518 2.41 0.562 ;
        RECT 2.558 1.148 2.626 1.192 ;
        RECT 2.558 0.068 2.626 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.57 0.652 ;
        RECT 4.286 0.518 4.354 0.742 ;
        RECT 3.962 0.518 4.03 0.832 ;
        RECT 3.422 0.428 3.49 0.832 ;
        RECT 1.694 0.428 1.762 0.832 ;
        RECT 1.046 0.428 1.114 0.832 ;
        RECT 0.506 0.428 0.574 0.832 ;
        RECT 0.182 0.518 0.25 0.742 ;
      LAYER v0 ;
        RECT 0.182 0.678 0.25 0.722 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.506 0.724 0.574 0.768 ;
        RECT 0.506 0.493 0.574 0.537 ;
        RECT 1.046 0.743 1.114 0.787 ;
        RECT 1.046 0.473 1.114 0.517 ;
        RECT 1.694 0.763 1.762 0.807 ;
        RECT 1.694 0.498 1.762 0.542 ;
        RECT 2.234 0.608 2.302 0.652 ;
        RECT 2.774 0.608 2.842 0.652 ;
        RECT 3.422 0.743 3.49 0.787 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 3.962 0.768 4.03 0.812 ;
        RECT 4.288 0.678 4.352 0.722 ;
        RECT 4.288 0.538 4.352 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.57 0.022 ;
        RECT 4.286 -0.022 4.354 0.202 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.234 -0.022 2.302 0.292 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
        RECT -0.034 1.238 4.57 1.282 ;
        RECT 4.286 1.058 4.354 1.282 ;
        RECT 3.962 1.058 4.03 1.282 ;
        RECT 3.422 1.058 3.49 1.282 ;
        RECT 2.774 1.058 2.842 1.282 ;
        RECT 2.234 1.148 2.302 1.282 ;
        RECT 1.694 0.968 1.762 1.282 ;
        RECT 1.046 1.058 1.114 1.282 ;
        RECT 0.506 1.058 0.574 1.282 ;
        RECT 0.182 1.058 0.25 1.282 ;
      LAYER v0 ;
        RECT 0.182 1.078 0.25 1.122 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.506 1.078 0.574 1.122 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.046 1.103 1.114 1.147 ;
        RECT 1.046 0.113 1.114 0.157 ;
        RECT 1.694 1.033 1.762 1.077 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 2.236 1.168 2.3 1.212 ;
        RECT 2.234 0.222 2.302 0.266 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.774 1.078 2.842 1.122 ;
        RECT 3.422 1.078 3.49 1.122 ;
        RECT 3.422 0.048 3.49 0.092 ;
        RECT 3.962 1.103 4.03 1.147 ;
        RECT 3.962 0.138 4.03 0.182 ;
        RECT 4.286 1.103 4.354 1.147 ;
        RECT 4.286 0.138 4.354 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.878 0.808 0.922 ;
      RECT 0.164 0.428 0.824 0.472 ;
      RECT 1.352 0.878 1.996 0.922 ;
      RECT 2.54 0.878 3.184 0.922 ;
      RECT 0.904 0.428 3.74 0.472 ;
      RECT 0.596 0.788 3.94 0.832 ;
      RECT 0.38 0.698 4.156 0.742 ;
      RECT 3.728 0.878 4.372 0.922 ;
      RECT 3.82 0.428 4.372 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.878 0.25 1.012 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.29 0.698 0.358 1.192 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.398 0.698 0.466 1.192 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.788 0.682 1.102 ;
      RECT 0.722 0.698 0.79 1.192 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.83 0.698 0.898 1.012 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 1.026 0.878 1.262 0.922 ;
      RECT 0.938 0.338 1.262 0.382 ;
      RECT 1.91 0.788 1.978 1.102 ;
      RECT 1.37 0.698 1.438 1.192 ;
      RECT 1.478 0.698 1.546 0.832 ;
      RECT 1.586 0.698 1.654 1.102 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 2.342 0.788 2.558 0.832 ;
      RECT 1.802 0.698 2.774 0.742 ;
      RECT 2.882 0.788 2.95 0.922 ;
      RECT 2.342 0.428 2.558 0.472 ;
      RECT 2.99 0.698 3.058 0.832 ;
      RECT 2.99 0.248 3.058 0.472 ;
      RECT 3.098 0.698 3.166 1.192 ;
      RECT 3.422 0.158 3.49 0.382 ;
      RECT 3.206 0.698 3.274 1.192 ;
      RECT 3.206 0.068 3.274 0.562 ;
      RECT 3.314 0.698 3.382 1.102 ;
      RECT 3.314 0.248 3.382 0.472 ;
      RECT 3.53 0.698 3.598 1.192 ;
      RECT 3.746 0.068 3.814 0.562 ;
      RECT 3.638 0.788 3.706 1.012 ;
      RECT 3.638 0.248 3.706 0.472 ;
      RECT 3.746 0.698 3.814 1.192 ;
      RECT 3.854 0.788 3.922 1.102 ;
      RECT 4.07 0.698 4.138 1.192 ;
      RECT 4.07 0.068 4.138 0.472 ;
      RECT 4.178 0.698 4.246 1.192 ;
      RECT 4.178 0.068 4.246 0.562 ;
      RECT 4.286 0.788 4.354 1.012 ;
      RECT 4.286 0.248 4.354 0.472 ;
    LAYER v1 ;
      RECT 4.29 0.428 4.35 0.472 ;
      RECT 4.29 0.878 4.35 0.922 ;
      RECT 4.074 0.698 4.134 0.742 ;
      RECT 3.858 0.428 3.918 0.472 ;
      RECT 3.858 0.788 3.918 0.832 ;
      RECT 3.75 0.878 3.81 0.922 ;
      RECT 3.642 0.428 3.702 0.472 ;
      RECT 3.642 0.788 3.702 0.832 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 3.318 0.698 3.378 0.742 ;
      RECT 3.102 0.878 3.162 0.922 ;
      RECT 2.994 0.428 3.054 0.472 ;
      RECT 2.994 0.698 3.054 0.742 ;
      RECT 2.886 0.788 2.946 0.832 ;
      RECT 2.562 0.878 2.622 0.922 ;
      RECT 1.914 0.878 1.974 0.922 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.59 0.698 1.65 0.742 ;
      RECT 1.482 0.788 1.542 0.832 ;
      RECT 1.374 0.878 1.434 0.922 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.726 0.428 0.786 0.472 ;
      RECT 0.726 0.878 0.786 0.922 ;
      RECT 0.618 0.788 0.678 0.832 ;
      RECT 0.402 0.698 0.462 0.742 ;
      RECT 0.186 0.428 0.246 0.472 ;
      RECT 0.186 0.878 0.246 0.922 ;
    LAYER v0 ;
      RECT 4.286 0.338 4.354 0.382 ;
      RECT 4.286 0.878 4.354 0.922 ;
      RECT 4.178 0.138 4.246 0.182 ;
      RECT 4.178 0.453 4.246 0.497 ;
      RECT 4.178 0.768 4.246 0.812 ;
      RECT 4.178 1.103 4.246 1.147 ;
      RECT 4.07 0.138 4.138 0.182 ;
      RECT 4.07 0.3695 4.138 0.4135 ;
      RECT 4.07 0.768 4.138 0.812 ;
      RECT 4.07 1.103 4.138 1.147 ;
      RECT 3.854 0.968 3.922 1.012 ;
      RECT 3.746 0.138 3.814 0.182 ;
      RECT 3.746 0.768 3.814 0.812 ;
      RECT 3.746 1.078 3.814 1.122 ;
      RECT 3.748 0.498 3.812 0.542 ;
      RECT 3.638 0.338 3.706 0.382 ;
      RECT 3.638 0.878 3.706 0.922 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.53 0.743 3.598 0.787 ;
      RECT 3.53 1.078 3.598 1.122 ;
      RECT 3.422 0.248 3.49 0.292 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 3.314 0.968 3.382 1.012 ;
      RECT 3.206 0.1515 3.274 0.1955 ;
      RECT 3.206 0.47 3.274 0.514 ;
      RECT 3.206 0.746 3.274 0.79 ;
      RECT 3.206 1.0645 3.274 1.1085 ;
      RECT 3.098 0.1515 3.166 0.1955 ;
      RECT 3.098 0.47 3.166 0.514 ;
      RECT 3.098 0.746 3.166 0.79 ;
      RECT 3.098 1.0645 3.166 1.1085 ;
      RECT 2.99 0.293 3.058 0.337 ;
      RECT 2.99 0.746 3.058 0.79 ;
      RECT 2.992 0.948 3.056 0.992 ;
      RECT 2.882 1.078 2.95 1.122 ;
      RECT 2.558 1.013 2.626 1.057 ;
      RECT 2.56 0.228 2.624 0.272 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.45 0.698 2.518 0.742 ;
      RECT 2.45 0.788 2.518 0.832 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 2.018 0.788 2.086 0.832 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.91 0.698 1.978 0.742 ;
      RECT 1.91 1.013 1.978 1.057 ;
      RECT 1.586 0.498 1.654 0.542 ;
      RECT 1.586 0.763 1.654 0.807 ;
      RECT 1.586 1.033 1.654 1.077 ;
      RECT 1.478 0.763 1.546 0.807 ;
      RECT 1.37 0.1515 1.438 0.1955 ;
      RECT 1.37 0.453 1.438 0.497 ;
      RECT 1.37 0.763 1.438 0.807 ;
      RECT 1.37 1.0645 1.438 1.1085 ;
      RECT 1.262 0.1515 1.33 0.1955 ;
      RECT 1.262 0.453 1.33 0.497 ;
      RECT 1.262 0.763 1.33 0.807 ;
      RECT 1.262 1.0645 1.33 1.1085 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 1.046 0.878 1.114 0.922 ;
      RECT 1.046 0.968 1.114 1.012 ;
      RECT 0.938 0.113 1.006 0.157 ;
      RECT 0.938 1.103 1.006 1.147 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.83 0.763 0.898 0.807 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.408 0.79 0.452 ;
      RECT 0.722 0.763 0.79 0.807 ;
      RECT 0.722 1.078 0.79 1.122 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.614 0.923 0.682 0.967 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.493 0.466 0.537 ;
      RECT 0.398 0.724 0.466 0.768 ;
      RECT 0.398 1.078 0.466 1.122 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.29 0.3855 0.358 0.4295 ;
      RECT 0.29 0.8305 0.358 0.8745 ;
      RECT 0.29 1.078 0.358 1.122 ;
      RECT 0.182 0.293 0.25 0.337 ;
      RECT 0.182 0.923 0.25 0.967 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.898 0.968 0.938 1.012 ;
      RECT 0.938 0.968 1.006 1.192 ;
      RECT 1.006 0.968 1.134 1.012 ;
      RECT 0.898 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.006 0.248 1.134 0.292 ;
      RECT 1.262 0.698 1.33 1.192 ;
      RECT 1.262 0.068 1.33 0.562 ;
      RECT 1.978 0.788 2.194 0.832 ;
      RECT 1.438 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.202 ;
      RECT 1.654 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.472 ;
      RECT 1.978 0.428 2.194 0.472 ;
      RECT 2.558 0.788 2.626 1.102 ;
      RECT 2.774 0.698 2.842 1.012 ;
      RECT 2.842 0.968 2.882 1.012 ;
      RECT 2.882 0.968 2.95 1.192 ;
      RECT 2.95 0.878 2.99 0.922 ;
      RECT 2.99 0.878 3.058 1.012 ;
      RECT 2.558 0.158 2.626 0.472 ;
      RECT 2.626 0.158 2.882 0.202 ;
      RECT 2.882 0.068 2.95 0.202 ;
      RECT 2.95 0.068 3.098 0.112 ;
      RECT 3.098 0.068 3.166 0.562 ;
      RECT 3.49 0.338 3.53 0.382 ;
      RECT 3.53 0.338 3.598 0.562 ;
      RECT 3.814 0.428 4.03 0.472 ;
  END
END b15fpy400hn1d04x5

MACRO b15fpy400hn1d08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fpy400hn1d08x5 0 0 ;
  SIZE 5.94 BY 1.26 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 9.22027775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 9.22027775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.248 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.248 3.922 0.562 ;
      LAYER v0 ;
        RECT 3.854 0.293 3.922 0.337 ;
    END
  END d2
  PIN d3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.788 2.41 1.192 ;
      LAYER v0 ;
        RECT 2.342 0.878 2.41 0.922 ;
    END
  END d3
  PIN d4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.788 3.814 1.012 ;
      LAYER v0 ;
        RECT 3.746 0.923 3.814 0.967 ;
    END
  END d4
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.425 0.25 0.469 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.69 0.068 5.758 0.562 ;
      LAYER v0 ;
        RECT 5.69 0.448 5.758 0.492 ;
        RECT 5.69 0.138 5.758 0.182 ;
    END
  END o2
  PIN o3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.698 0.25 1.192 ;
      LAYER v0 ;
        RECT 0.182 1.078 0.25 1.122 ;
        RECT 0.182 0.7905 0.25 0.8345 ;
    END
  END o3
  PIN o4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.69 0.698 5.758 1.192 ;
      LAYER v0 ;
        RECT 5.69 1.078 5.758 1.122 ;
        RECT 5.69 0.768 5.758 0.812 ;
    END
  END o4
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.068 2.842 0.382 ;
      LAYER v0 ;
        RECT 2.774 0.2705 2.842 0.3145 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.068 3.382 0.382 ;
      LAYER v0 ;
        RECT 3.314 0.2705 3.382 0.3145 ;
    END
  END si2
  PIN si3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.878 2.842 1.192 ;
      LAYER v0 ;
        RECT 2.774 0.9455 2.842 0.9895 ;
    END
  END si3
  PIN si4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.878 3.382 1.192 ;
      LAYER v0 ;
        RECT 3.314 0.9455 3.382 0.9895 ;
    END
  END si4
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0252 LAYER m1 ;
      ANTENNAMAXAREACAR 6.22047625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0252 LAYER m1 ;
      ANTENNAMAXAREACAR 18.1090475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.518 3.598 0.562 ;
        RECT 3.53 0.248 3.598 0.562 ;
        RECT 3.53 0.698 3.598 1.012 ;
        RECT 3.206 0.698 3.598 0.742 ;
        RECT 2.558 0.518 2.95 0.562 ;
        RECT 2.558 0.248 2.626 0.562 ;
        RECT 2.558 0.698 2.95 0.742 ;
        RECT 2.558 0.698 2.626 1.012 ;
      LAYER v0 ;
        RECT 2.558 0.9005 2.626 0.9445 ;
        RECT 2.558 0.293 2.626 0.337 ;
        RECT 2.774 0.698 2.842 0.742 ;
        RECT 2.774 0.518 2.842 0.562 ;
        RECT 3.314 0.698 3.382 0.742 ;
        RECT 3.314 0.518 3.382 0.562 ;
        RECT 3.53 0.923 3.598 0.967 ;
        RECT 3.53 0.293 3.598 0.337 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.974 0.652 ;
        RECT 5.798 0.428 5.866 0.832 ;
        RECT 5.582 0.248 5.65 1.012 ;
        RECT 5.042 0.788 5.65 0.832 ;
        RECT 5.042 0.428 5.65 0.472 ;
        RECT 5.366 0.788 5.434 1.012 ;
        RECT 5.366 0.248 5.434 0.472 ;
        RECT 4.502 0.338 4.57 0.832 ;
        RECT 2.774 0.788 3.382 0.832 ;
        RECT 2.774 0.428 3.382 0.472 ;
        RECT 2.99 0.428 3.058 0.832 ;
        RECT 1.478 0.338 1.546 0.922 ;
        RECT 0.29 0.338 0.358 1.012 ;
        RECT 0.074 0.338 0.142 0.922 ;
      LAYER v0 ;
        RECT 0.074 0.7905 0.142 0.8345 ;
        RECT 0.074 0.425 0.142 0.469 ;
        RECT 0.29 0.7905 0.358 0.8345 ;
        RECT 0.29 0.425 0.358 0.469 ;
        RECT 0.506 0.608 0.574 0.652 ;
        RECT 0.83 0.608 0.898 0.652 ;
        RECT 1.478 0.788 1.546 0.832 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 2.234 0.608 2.302 0.652 ;
        RECT 2.882 0.788 2.95 0.832 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 3.206 0.788 3.274 0.832 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.746 0.608 3.814 0.652 ;
        RECT 4.502 0.744 4.57 0.788 ;
        RECT 4.502 0.408 4.57 0.452 ;
        RECT 5.15 0.788 5.218 0.832 ;
        RECT 5.15 0.428 5.218 0.472 ;
        RECT 5.366 0.878 5.434 0.922 ;
        RECT 5.366 0.338 5.434 0.382 ;
        RECT 5.582 0.878 5.65 0.922 ;
        RECT 5.582 0.338 5.65 0.382 ;
        RECT 5.798 0.768 5.866 0.812 ;
        RECT 5.798 0.448 5.866 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.974 0.022 ;
        RECT 5.798 -0.022 5.866 0.202 ;
        RECT 5.582 -0.022 5.65 0.202 ;
        RECT 5.366 -0.022 5.434 0.202 ;
        RECT 5.15 -0.022 5.218 0.202 ;
        RECT 4.394 -0.022 4.462 0.202 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
        RECT -0.034 1.238 5.974 1.282 ;
        RECT 5.798 1.058 5.866 1.282 ;
        RECT 5.582 1.058 5.65 1.282 ;
        RECT 5.366 1.058 5.434 1.282 ;
        RECT 5.15 1.058 5.218 1.282 ;
        RECT 4.502 1.058 4.57 1.282 ;
        RECT 3.746 1.058 3.814 1.282 ;
        RECT 3.206 1.058 3.274 1.282 ;
        RECT 2.882 1.058 2.95 1.282 ;
        RECT 2.234 1.058 2.302 1.282 ;
        RECT 1.478 1.058 1.546 1.282 ;
        RECT 0.83 1.058 0.898 1.282 ;
        RECT 0.506 1.058 0.574 1.282 ;
        RECT 0.29 1.058 0.358 1.282 ;
        RECT 0.074 1.058 0.142 1.282 ;
      LAYER v0 ;
        RECT 0.074 1.078 0.142 1.122 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 1.078 0.358 1.122 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 1.078 0.574 1.122 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.83 1.078 0.898 1.122 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.478 1.078 1.546 1.122 ;
        RECT 1.478 0.113 1.546 0.157 ;
        RECT 2.234 1.078 2.302 1.122 ;
        RECT 2.342 0.048 2.41 0.092 ;
        RECT 2.882 1.078 2.95 1.122 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.206 1.078 3.274 1.122 ;
        RECT 3.206 0.138 3.274 0.182 ;
        RECT 3.746 1.078 3.814 1.122 ;
        RECT 3.746 0.048 3.814 0.092 ;
        RECT 4.394 0.138 4.462 0.182 ;
        RECT 4.502 1.078 4.57 1.122 ;
        RECT 5.15 1.078 5.218 1.122 ;
        RECT 5.15 0.138 5.218 0.182 ;
        RECT 5.366 1.078 5.434 1.122 ;
        RECT 5.366 0.138 5.434 0.182 ;
        RECT 5.582 1.078 5.65 1.122 ;
        RECT 5.582 0.138 5.65 0.182 ;
        RECT 5.798 1.078 5.866 1.122 ;
        RECT 5.798 0.138 5.866 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.704 0.968 5.128 1.012 ;
      RECT 0.812 0.338 5.128 0.382 ;
    LAYER m1 ;
      RECT 0.398 0.698 0.466 1.192 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.722 0.788 0.79 1.192 ;
      RECT 0.938 0.878 1.006 1.012 ;
      RECT 0.506 0.698 0.574 1.012 ;
      RECT 1.262 0.788 1.33 1.012 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 1.37 0.698 1.438 1.192 ;
      RECT 1.262 0.248 1.33 0.382 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.586 1.058 1.802 1.102 ;
      RECT 1.694 0.788 1.762 1.012 ;
      RECT 1.586 0.158 1.802 0.202 ;
      RECT 1.91 0.698 1.978 1.192 ;
      RECT 2.018 0.788 2.086 1.192 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 2.126 0.788 2.194 1.012 ;
      RECT 2.126 0.158 2.194 0.562 ;
      RECT 2.234 0.248 2.302 0.382 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 3.422 0.788 3.49 1.102 ;
      RECT 3.098 0.068 3.166 0.382 ;
      RECT 3.854 0.788 3.922 1.192 ;
      RECT 3.962 0.878 4.03 1.102 ;
      RECT 3.962 0.248 4.03 0.382 ;
      RECT 3.422 0.158 3.49 0.472 ;
      RECT 3.962 0.068 4.178 0.112 ;
      RECT 4.178 0.698 4.246 1.192 ;
      RECT 4.286 0.788 4.354 1.012 ;
      RECT 4.286 0.248 4.354 0.472 ;
      RECT 4.482 0.878 4.61 0.922 ;
      RECT 4.394 0.248 4.61 0.292 ;
      RECT 4.718 0.698 4.934 0.742 ;
      RECT 4.718 0.788 4.786 1.012 ;
      RECT 4.718 0.248 4.786 0.472 ;
      RECT 5.042 0.878 5.11 1.012 ;
      RECT 5.042 0.248 5.11 0.382 ;
      RECT 4.61 0.518 4.934 0.562 ;
    LAYER v1 ;
      RECT 5.046 0.338 5.106 0.382 ;
      RECT 5.046 0.968 5.106 1.012 ;
      RECT 4.722 0.338 4.782 0.382 ;
      RECT 4.722 0.968 4.782 1.012 ;
      RECT 4.29 0.338 4.35 0.382 ;
      RECT 4.29 0.968 4.35 1.012 ;
      RECT 3.966 0.338 4.026 0.382 ;
      RECT 3.966 0.968 4.026 1.012 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 2.13 0.968 2.19 1.012 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.698 0.968 1.758 1.012 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 1.266 0.968 1.326 1.012 ;
      RECT 0.942 0.968 1.002 1.012 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.726 0.968 0.786 1.012 ;
    LAYER v0 ;
      RECT 5.258 0.518 5.326 0.562 ;
      RECT 5.258 0.698 5.326 0.742 ;
      RECT 5.042 0.2705 5.11 0.3145 ;
      RECT 5.042 0.9455 5.11 0.9895 ;
      RECT 4.934 0.1535 5.002 0.1975 ;
      RECT 4.934 1.0625 5.002 1.1065 ;
      RECT 4.826 0.698 4.894 0.742 ;
      RECT 4.718 0.3155 4.786 0.3595 ;
      RECT 4.718 0.518 4.786 0.562 ;
      RECT 4.718 0.9005 4.786 0.9445 ;
      RECT 4.61 0.138 4.678 0.182 ;
      RECT 4.61 0.408 4.678 0.452 ;
      RECT 4.61 0.744 4.678 0.788 ;
      RECT 4.61 1.078 4.678 1.122 ;
      RECT 4.502 0.248 4.57 0.292 ;
      RECT 4.502 0.878 4.57 0.922 ;
      RECT 4.286 0.338 4.354 0.382 ;
      RECT 4.286 0.698 4.354 0.742 ;
      RECT 4.286 0.878 4.354 0.922 ;
      RECT 4.178 0.428 4.246 0.472 ;
      RECT 4.178 1.058 4.246 1.102 ;
      RECT 4.07 0.068 4.138 0.112 ;
      RECT 4.07 0.428 4.138 0.472 ;
      RECT 4.07 0.788 4.138 0.832 ;
      RECT 4.07 1.058 4.138 1.102 ;
      RECT 3.962 0.158 4.03 0.202 ;
      RECT 3.962 0.293 4.03 0.337 ;
      RECT 3.962 0.923 4.03 0.967 ;
      RECT 3.854 0.808 3.922 0.852 ;
      RECT 3.854 1.078 3.922 1.122 ;
      RECT 3.53 0.158 3.598 0.202 ;
      RECT 3.53 1.058 3.598 1.102 ;
      RECT 3.422 0.408 3.49 0.452 ;
      RECT 3.422 0.808 3.49 0.852 ;
      RECT 3.098 0.138 3.166 0.182 ;
      RECT 3.098 0.318 3.166 0.362 ;
      RECT 2.666 0.408 2.734 0.452 ;
      RECT 2.666 0.808 2.734 0.852 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.558 1.058 2.626 1.102 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.126 0.178 2.194 0.222 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.126 0.878 2.194 0.922 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 2.018 0.878 2.086 0.922 ;
      RECT 2.018 1.078 2.086 1.122 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.4375 1.978 0.4815 ;
      RECT 1.91 0.788 1.978 0.832 ;
      RECT 1.91 1.078 1.978 1.122 ;
      RECT 1.802 0.4375 1.87 0.4815 ;
      RECT 1.802 0.788 1.87 0.832 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.878 1.762 0.922 ;
      RECT 1.694 1.058 1.762 1.102 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.586 0.878 1.654 0.922 ;
      RECT 1.37 0.113 1.438 0.157 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.37 0.788 1.438 0.832 ;
      RECT 1.37 1.078 1.438 1.122 ;
      RECT 1.262 0.3155 1.33 0.3595 ;
      RECT 1.262 0.9005 1.33 0.9445 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.154 0.698 1.222 0.742 ;
      RECT 1.046 0.1535 1.114 0.1975 ;
      RECT 1.046 1.0625 1.114 1.1065 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.9455 1.006 0.9895 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.808 0.79 0.852 ;
      RECT 0.722 1.078 0.79 1.122 ;
      RECT 0.724 0.408 0.788 0.452 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.506 0.923 0.574 0.967 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.425 0.466 0.469 ;
      RECT 0.398 0.7905 0.466 0.8345 ;
      RECT 0.398 1.078 0.466 1.122 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.79 0.338 0.938 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 0.574 0.698 1.046 0.742 ;
      RECT 1.046 0.698 1.114 1.192 ;
      RECT 1.114 0.698 1.33 0.742 ;
      RECT 0.574 0.518 1.046 0.562 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.114 0.518 1.33 0.562 ;
      RECT 1.438 0.968 1.586 1.012 ;
      RECT 1.586 0.788 1.654 1.012 ;
      RECT 1.438 0.248 1.586 0.292 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.802 0.698 1.87 1.102 ;
      RECT 1.802 0.158 1.87 0.562 ;
      RECT 1.978 0.698 2.45 0.742 ;
      RECT 2.45 0.698 2.518 1.102 ;
      RECT 2.518 1.058 2.666 1.102 ;
      RECT 2.666 0.788 2.734 1.102 ;
      RECT 1.978 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.202 ;
      RECT 2.302 0.158 2.666 0.202 ;
      RECT 2.666 0.158 2.734 0.472 ;
      RECT 3.49 1.058 3.638 1.102 ;
      RECT 3.638 0.698 3.706 1.102 ;
      RECT 3.706 0.698 4.07 0.742 ;
      RECT 4.07 0.698 4.138 1.192 ;
      RECT 3.49 0.158 4.07 0.202 ;
      RECT 4.07 0.158 4.138 0.562 ;
      RECT 4.178 0.068 4.246 0.562 ;
      RECT 4.246 0.698 4.374 0.742 ;
      RECT 4.61 0.698 4.678 1.192 ;
      RECT 4.61 0.068 4.678 0.472 ;
      RECT 4.934 0.698 5.002 1.192 ;
      RECT 5.002 0.698 5.434 0.742 ;
      RECT 4.934 0.068 5.002 0.562 ;
      RECT 5.002 0.518 5.434 0.562 ;
  END
END b15fpy400hn1d08x5

MACRO b15fqn003hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn003hn1n02x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.428 1.222 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
      LAYER m2 ;
        RECT 0.38 0.518 1.24 0.562 ;
      LAYER v1 ;
        RECT 0.402 0.518 0.462 0.562 ;
        RECT 1.158 0.518 1.218 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.498 0.466 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.292 ;
        RECT 1.998 0.068 2.194 0.112 ;
      LAYER v0 ;
        RECT 2.018 0.068 2.086 0.112 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.248 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.498 1.978 0.542 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.403 0.25 0.447 ;
        RECT 0.182 0.1915 0.25 0.2355 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 1.046 0.338 1.114 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.506 0.403 0.574 0.447 ;
        RECT 1.046 0.402 1.114 0.446 ;
        RECT 1.37 0.403 1.438 0.447 ;
        RECT 1.802 0.393 1.87 0.437 ;
        RECT 2.234 0.377 2.302 0.421 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.234 -0.022 2.302 0.292 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.046 0.158 1.33 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.398 0.088 0.466 0.132 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.234 0.208 2.302 0.252 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 0.824 0.382 ;
      RECT 0.904 0.338 1.688 0.382 ;
      RECT 1.568 0.518 2.212 0.562 ;
      RECT 0.812 0.428 2.444 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.382 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.83 0.248 1.262 0.292 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.37 0.158 1.586 0.202 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.478 0.518 1.694 0.562 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.342 0.158 2.41 0.472 ;
    LAYER v1 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.13 0.518 2.19 0.562 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 2.342 0.208 2.41 0.252 ;
      RECT 2.342 0.377 2.41 0.421 ;
      RECT 2.126 0.377 2.194 0.421 ;
      RECT 2.018 0.498 2.086 0.542 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.586 0.3835 1.654 0.4275 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.403 1.33 0.447 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.498 0.898 0.542 ;
      RECT 0.722 0.363 0.79 0.407 ;
      RECT 0.614 0.498 0.682 0.542 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.79 0.158 1.006 0.202 ;
      RECT 0.682 0.068 1.006 0.112 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.478 0.068 1.694 0.112 ;
      RECT 1.694 0.068 1.762 0.562 ;
  END
END b15fqn003hn1n02x5

MACRO b15fqn003hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn003hn1n03x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 4.948889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 4.948889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.428 1.33 0.562 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.518 1.348 0.562 ;
      LAYER v1 ;
        RECT 0.51 0.518 0.57 0.562 ;
        RECT 1.266 0.518 1.326 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 1.262 0.498 1.33 0.542 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.068 2.302 0.292 ;
        RECT 2.106 0.068 2.302 0.112 ;
      LAYER v0 ;
        RECT 2.126 0.068 2.194 0.112 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.248 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.498 2.086 0.542 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.403 0.142 0.447 ;
        RECT 0.074 0.183 0.142 0.227 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.614 0.338 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.403 0.25 0.447 ;
        RECT 0.614 0.383 0.682 0.427 ;
        RECT 1.154 0.383 1.222 0.427 ;
        RECT 1.478 0.403 1.546 0.447 ;
        RECT 1.91 0.393 1.978 0.437 ;
        RECT 2.342 0.377 2.41 0.421 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.342 -0.022 2.41 0.292 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.183 0.25 0.227 ;
        RECT 0.506 0.203 0.574 0.247 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.91 0.138 1.978 0.182 ;
        RECT 2.342 0.208 2.41 0.252 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 0.932 0.382 ;
      RECT 1.012 0.338 1.796 0.382 ;
      RECT 1.676 0.518 2.32 0.562 ;
      RECT 0.92 0.428 2.552 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 0.938 0.248 1.37 0.292 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.478 0.158 1.694 0.202 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.586 0.518 1.802 0.562 ;
      RECT 2.126 0.428 2.194 0.562 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 2.45 0.158 2.518 0.472 ;
    LAYER v1 ;
      RECT 2.454 0.428 2.514 0.472 ;
      RECT 2.238 0.518 2.298 0.562 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.698 0.518 1.758 0.562 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.402 0.338 0.462 0.382 ;
    LAYER v0 ;
      RECT 2.45 0.208 2.518 0.252 ;
      RECT 2.45 0.377 2.518 0.421 ;
      RECT 2.234 0.377 2.302 0.421 ;
      RECT 2.126 0.498 2.194 0.542 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.3835 1.762 0.4275 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.37 0.403 1.438 0.447 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.498 1.114 0.542 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.398 0.403 0.466 0.447 ;
      RECT 0.29 0.183 0.358 0.227 ;
      RECT 0.29 0.403 0.358 0.447 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.79 0.068 1.006 0.112 ;
      RECT 0.898 0.158 1.114 0.202 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.674 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.562 ;
  END
END b15fqn003hn1n03x5

MACRO b15fqn003hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn003hn1n04x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 6.748611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 6.748611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.438 0.382 ;
        RECT 1.154 0.338 1.222 0.562 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.518 1.24 0.562 ;
      LAYER v1 ;
        RECT 0.51 0.518 0.57 0.562 ;
        RECT 1.158 0.518 1.218 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.292 ;
        RECT 2.214 0.068 2.41 0.112 ;
      LAYER v0 ;
        RECT 2.234 0.068 2.302 0.112 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.248 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.498 2.194 0.542 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.403 0.142 0.447 ;
        RECT 0.074 0.178 0.142 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.586 0.338 1.654 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.338 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.403 0.25 0.447 ;
        RECT 0.614 0.363 0.682 0.407 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.586 0.403 1.654 0.447 ;
        RECT 2.018 0.393 2.086 0.437 ;
        RECT 2.45 0.377 2.518 0.421 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.178 0.25 0.222 ;
        RECT 0.506 0.222 0.574 0.266 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.45 0.208 2.518 0.252 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 0.932 0.382 ;
      RECT 1.012 0.338 1.904 0.382 ;
      RECT 1.784 0.518 2.428 0.562 ;
      RECT 0.92 0.428 2.66 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.046 0.248 1.478 0.292 ;
      RECT 1.586 0.158 1.802 0.202 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.558 0.158 2.626 0.472 ;
    LAYER v1 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.346 0.518 2.406 0.562 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 1.806 0.338 1.866 0.382 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.402 0.338 0.462 0.382 ;
    LAYER v0 ;
      RECT 2.558 0.208 2.626 0.252 ;
      RECT 2.558 0.377 2.626 0.421 ;
      RECT 2.342 0.377 2.41 0.421 ;
      RECT 2.234 0.498 2.302 0.542 ;
      RECT 1.802 0.3835 1.87 0.4275 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.478 0.403 1.546 0.447 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.395 0.898 0.439 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.398 0.403 0.466 0.447 ;
      RECT 0.29 0.178 0.358 0.222 ;
      RECT 0.29 0.403 0.358 0.447 ;
    LAYER m1 ;
      RECT 0.83 0.518 1.046 0.562 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 0.898 0.158 1.114 0.202 ;
      RECT 1.222 0.338 1.438 0.382 ;
      RECT 1.478 0.248 1.546 0.562 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 0.79 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 1.694 0.518 1.91 0.562 ;
      RECT 1.546 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.562 ;
  END
END b15fqn003hn1n04x5

MACRO b15fqn003hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn003hn1n06x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    ANTENNADIFFAREA 0.03672 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.428 0.484 0.472 ;
      LAYER v1 ;
        RECT 0.078 0.428 0.138 0.472 ;
        RECT 0.294 0.428 0.354 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.179 0.142 0.223 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAGATEAREA 0.0117 LAYER m2 ;
      ANTENNAMAXAREACAR 0.3144445 LAYER m1 ;
      ANTENNAMAXAREACAR 4.950889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.2515555 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.3930555 LAYER m1 ;
      ANTENNAMAXAREACAR 6.188611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.338 1.654 0.562 ;
        RECT 1.458 0.338 1.654 0.382 ;
        RECT 0.398 0.428 0.466 0.562 ;
      LAYER m2 ;
        RECT 0.38 0.518 1.672 0.562 ;
      LAYER v1 ;
        RECT 0.402 0.518 0.462 0.562 ;
        RECT 1.59 0.518 1.65 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.498 0.466 0.542 ;
        RECT 1.478 0.338 1.546 0.382 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.292 ;
        RECT 2.342 0.068 2.626 0.112 ;
      LAYER v0 ;
        RECT 2.45 0.068 2.518 0.112 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 2.926 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 2.926 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.248 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.498 2.518 0.542 ;
    END
  END d
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.498 0.25 0.542 ;
        RECT 0.614 0.467 0.682 0.511 ;
        RECT 1.262 0.503 1.33 0.547 ;
        RECT 1.802 0.403 1.87 0.447 ;
        RECT 2.234 0.393 2.302 0.437 ;
        RECT 2.666 0.377 2.734 0.421 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.088 0.25 0.132 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.666 0.208 2.734 0.252 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.338 0.916 0.382 ;
      RECT 1.244 0.338 2.104 0.382 ;
      RECT 2 0.518 2.644 0.562 ;
      RECT 0.812 0.428 2.876 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.182 0.248 0.25 0.382 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.398 0.338 0.682 0.382 ;
      RECT 0.83 0.158 0.898 0.562 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.458 0.338 1.586 0.382 ;
      RECT 1.154 0.338 1.35 0.382 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.802 0.158 2.018 0.202 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 2.342 0.158 2.41 0.472 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 2.774 0.158 2.842 0.472 ;
    LAYER v1 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.562 0.518 2.622 0.562 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 2.022 0.518 2.082 0.562 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 2.774 0.208 2.842 0.252 ;
      RECT 2.774 0.377 2.842 0.421 ;
      RECT 2.558 0.377 2.626 0.421 ;
      RECT 2.342 0.223 2.41 0.267 ;
      RECT 2.342 0.393 2.41 0.437 ;
      RECT 2.018 0.3835 2.086 0.4275 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.694 0.403 1.762 0.447 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 1.046 0.467 1.114 0.511 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.467 0.898 0.511 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.088 0.682 0.132 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.182 0.293 0.25 0.337 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.898 0.158 1.114 0.202 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.114 0.248 1.694 0.292 ;
      RECT 1.694 0.248 1.762 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 0.79 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.438 0.158 1.694 0.202 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.91 0.518 2.126 0.562 ;
      RECT 1.762 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.562 ;
  END
END b15fqn003hn1n06x5

MACRO b15fqn003hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn003hn1n08x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 7.788889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 7.788889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.338 1.762 0.382 ;
        RECT 1.37 0.518 1.546 0.562 ;
        RECT 1.478 0.338 1.546 0.562 ;
        RECT 0.506 0.248 0.574 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.518 1.472 0.562 ;
      LAYER v1 ;
        RECT 0.51 0.518 0.57 0.562 ;
        RECT 1.374 0.518 1.434 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.068 3.294 0.112 ;
        RECT 3.098 0.068 3.166 0.292 ;
      LAYER v0 ;
        RECT 3.206 0.068 3.274 0.112 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.43833325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.43833325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.338 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.498 2.842 0.542 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 2.99 0.338 3.058 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.694 0.472 1.762 0.516 ;
        RECT 1.91 0.472 1.978 0.516 ;
        RECT 2.558 0.393 2.626 0.437 ;
        RECT 2.99 0.377 3.058 0.421 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 2.99 -0.022 3.058 0.292 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.614 0.1245 0.682 0.1685 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.91 0.048 1.978 0.092 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.99 0.208 3.058 0.252 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.596 0.248 1.04 0.292 ;
      RECT 1.552 0.518 2.32 0.562 ;
      RECT 1.46 0.068 2.752 0.112 ;
      RECT 1.12 0.248 3.308 0.292 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.37 0.518 1.478 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.242 0.158 1.978 0.202 ;
      RECT 2.018 0.158 2.234 0.202 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.666 0.068 2.882 0.112 ;
      RECT 2.342 0.068 2.41 0.472 ;
      RECT 3.206 0.158 3.274 0.472 ;
    LAYER v1 ;
      RECT 3.21 0.248 3.27 0.292 ;
      RECT 2.67 0.068 2.73 0.112 ;
      RECT 2.346 0.068 2.406 0.112 ;
      RECT 2.238 0.518 2.298 0.562 ;
      RECT 2.13 0.248 2.19 0.292 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.482 0.068 1.542 0.112 ;
      RECT 1.158 0.248 1.218 0.292 ;
      RECT 0.942 0.248 1.002 0.292 ;
      RECT 0.618 0.248 0.678 0.292 ;
    LAYER v0 ;
      RECT 3.206 0.208 3.274 0.252 ;
      RECT 3.206 0.377 3.274 0.421 ;
      RECT 2.882 0.208 2.95 0.252 ;
      RECT 2.882 0.377 2.95 0.421 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.344 0.088 2.408 0.132 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.472 1.87 0.516 ;
      RECT 1.586 0.472 1.654 0.516 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.154 0.473 1.222 0.517 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.006 0.158 1.134 0.202 ;
      RECT 1.114 0.248 1.33 0.292 ;
      RECT 0.898 0.068 1.654 0.112 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.546 0.338 1.762 0.382 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.248 1.438 0.382 ;
      RECT 1.438 0.248 1.802 0.292 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.87 0.248 2.018 0.292 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 2.234 0.158 2.302 0.562 ;
      RECT 2.882 0.068 2.95 0.472 ;
  END
END b15fqn003hn1n08x5

MACRO b15fqn003hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn003hn1n12x5 0 0 ;
  SIZE 3.996 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0207 LAYER m2 ;
      ANTENNAMAXAREACAR 0.61185175 LAYER m1 ;
      ANTENNAMAXAREACAR 4.05925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 0.61185175 LAYER m1 ;
      ANTENNAMAXAREACAR 4.05925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.338 1.978 0.382 ;
        RECT 1.694 0.338 1.762 0.472 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER m2 ;
        RECT 0.596 0.428 1.796 0.472 ;
      LAYER v1 ;
        RECT 0.618 0.428 0.678 0.472 ;
        RECT 1.698 0.428 1.758 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.068 3.814 0.382 ;
      LAYER v0 ;
        RECT 3.746 0.293 3.814 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.158 3.382 0.382 ;
      LAYER v0 ;
        RECT 3.314 0.293 3.382 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.03 0.652 ;
        RECT 3.638 0.338 3.706 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 2.126 0.338 2.194 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.83 0.4485 0.898 0.4925 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 1.802 0.473 1.87 0.517 ;
        RECT 2.126 0.473 2.194 0.517 ;
        RECT 2.342 0.473 2.41 0.517 ;
        RECT 2.99 0.538 3.058 0.582 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.638 0.377 3.706 0.421 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.03 0.022 ;
        RECT 3.638 -0.022 3.706 0.292 ;
        RECT 3.206 -0.022 3.274 0.292 ;
        RECT 2.99 -0.022 3.058 0.292 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.722 0.1245 0.79 0.1685 ;
        RECT 2.126 0.048 2.194 0.092 ;
        RECT 2.99 0.178 3.058 0.222 ;
        RECT 3.206 0.178 3.274 0.222 ;
        RECT 3.638 0.158 3.706 0.202 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.704 0.338 1.148 0.382 ;
      RECT 1.876 0.428 2.66 0.472 ;
      RECT 2.74 0.428 3.184 0.472 ;
      RECT 1.568 0.068 3.616 0.112 ;
      RECT 1.228 0.338 3.956 0.382 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 1.154 0.338 1.438 0.382 ;
      RECT 0.938 0.068 1.006 0.472 ;
      RECT 1.694 0.338 1.762 0.472 ;
      RECT 1.91 0.428 1.978 0.562 ;
      RECT 1.154 0.248 1.478 0.292 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 1.566 0.158 2.41 0.202 ;
      RECT 2.45 0.248 2.518 0.472 ;
      RECT 2.666 0.158 2.734 0.382 ;
      RECT 2.342 0.068 2.774 0.112 ;
      RECT 3.314 0.518 3.53 0.562 ;
      RECT 2.882 0.158 2.95 0.562 ;
      RECT 3.098 0.158 3.166 0.562 ;
      RECT 3.53 0.068 3.598 0.292 ;
      RECT 3.854 0.158 3.922 0.472 ;
    LAYER v1 ;
      RECT 3.858 0.338 3.918 0.382 ;
      RECT 3.534 0.068 3.594 0.112 ;
      RECT 3.534 0.338 3.594 0.382 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 2.778 0.068 2.838 0.112 ;
      RECT 2.67 0.338 2.73 0.382 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.454 0.338 2.514 0.382 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.59 0.068 1.65 0.112 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
    LAYER v0 ;
      RECT 3.854 0.178 3.922 0.222 ;
      RECT 3.854 0.408 3.922 0.452 ;
      RECT 3.53 0.158 3.598 0.202 ;
      RECT 3.422 0.518 3.49 0.562 ;
      RECT 3.098 0.178 3.166 0.222 ;
      RECT 3.098 0.448 3.166 0.492 ;
      RECT 2.882 0.178 2.95 0.222 ;
      RECT 2.882 0.4185 2.95 0.4625 ;
      RECT 2.774 0.338 2.842 0.382 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.473 2.302 0.517 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 2.018 0.473 2.086 0.517 ;
      RECT 1.91 0.473 1.978 0.517 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.3485 1.546 0.3925 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.048 0.498 1.112 0.542 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.722 0.4485 0.79 0.4925 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.448 0.574 0.492 ;
    LAYER m1 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.428 1.35 0.472 ;
      RECT 1.114 0.158 1.458 0.202 ;
      RECT 1.006 0.068 1.654 0.112 ;
      RECT 1.762 0.338 1.978 0.382 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.546 0.248 2.018 0.292 ;
      RECT 2.018 0.248 2.086 0.562 ;
      RECT 2.086 0.248 2.234 0.292 ;
      RECT 2.234 0.248 2.302 0.562 ;
      RECT 2.626 0.518 2.842 0.562 ;
      RECT 2.774 0.068 2.842 0.472 ;
      RECT 3.53 0.338 3.598 0.562 ;
  END
END b15fqn003hn1n12x5

MACRO b15fqn003hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn003hn1n16x5 0 0 ;
  SIZE 4.752 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 5.1925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0342 LAYER m2 ;
      ANTENNAMAXAREACAR 5.1925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.338 2.518 0.382 ;
        RECT 2.018 0.338 2.086 0.562 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER m2 ;
        RECT 0.704 0.518 2.228 0.562 ;
      LAYER v1 ;
        RECT 0.726 0.518 0.786 0.562 ;
        RECT 2.022 0.518 2.082 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.3155 0.79 0.3595 ;
        RECT 2.342 0.338 2.41 0.382 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.502 0.068 4.57 0.382 ;
      LAYER v0 ;
        RECT 4.502 0.293 4.57 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.338 4.246 0.562 ;
      LAYER v0 ;
        RECT 4.178 0.498 4.246 0.542 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.786 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.91 0.473 1.978 0.517 ;
        RECT 2.126 0.473 2.194 0.517 ;
        RECT 2.45 0.473 2.518 0.517 ;
        RECT 2.666 0.473 2.734 0.517 ;
        RECT 2.99 0.473 3.058 0.517 ;
        RECT 3.746 0.473 3.814 0.517 ;
        RECT 3.962 0.473 4.03 0.517 ;
        RECT 4.502 0.493 4.57 0.537 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.786 0.022 ;
        RECT 4.394 -0.022 4.462 0.202 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.746 -0.022 3.814 0.292 ;
        RECT 2.342 0.158 3.078 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.746 0.228 3.814 0.272 ;
        RECT 3.962 0.138 4.03 0.182 ;
        RECT 4.394 0.138 4.462 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.812 0.338 1.256 0.382 ;
      RECT 2.308 0.518 3.616 0.562 ;
      RECT 1.46 0.068 4.372 0.112 ;
      RECT 1.336 0.338 4.712 0.382 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.248 0.79 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 1.262 0.338 1.762 0.382 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 1.89 0.158 2.214 0.202 ;
      RECT 2.342 0.428 2.41 0.562 ;
      RECT 1.37 0.518 1.802 0.562 ;
      RECT 3.186 0.158 3.314 0.202 ;
      RECT 3.206 0.248 3.274 0.472 ;
      RECT 2.99 0.068 3.638 0.112 ;
      RECT 3.53 0.428 3.598 0.562 ;
      RECT 3.422 0.248 3.49 0.562 ;
      RECT 4.07 0.068 4.138 0.472 ;
      RECT 4.286 0.068 4.354 0.472 ;
      RECT 4.394 0.248 4.462 0.382 ;
      RECT 4.61 0.158 4.678 0.472 ;
    LAYER v1 ;
      RECT 4.614 0.338 4.674 0.382 ;
      RECT 4.398 0.338 4.458 0.382 ;
      RECT 4.29 0.068 4.35 0.112 ;
      RECT 3.642 0.068 3.702 0.112 ;
      RECT 3.534 0.518 3.594 0.562 ;
      RECT 3.318 0.518 3.378 0.562 ;
      RECT 3.21 0.338 3.27 0.382 ;
      RECT 3.102 0.068 3.162 0.112 ;
      RECT 2.346 0.518 2.406 0.562 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.482 0.068 1.542 0.112 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.834 0.338 0.894 0.382 ;
    LAYER v0 ;
      RECT 4.61 0.178 4.678 0.222 ;
      RECT 4.61 0.408 4.678 0.452 ;
      RECT 4.394 0.293 4.462 0.337 ;
      RECT 4.286 0.138 4.354 0.182 ;
      RECT 4.286 0.408 4.354 0.452 ;
      RECT 4.07 0.138 4.138 0.182 ;
      RECT 4.07 0.338 4.138 0.382 ;
      RECT 3.854 0.228 3.922 0.272 ;
      RECT 3.854 0.473 3.922 0.517 ;
      RECT 3.64 0.138 3.704 0.182 ;
      RECT 3.53 0.248 3.598 0.292 ;
      RECT 3.53 0.498 3.598 0.542 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.422 0.498 3.49 0.542 ;
      RECT 3.314 0.498 3.382 0.542 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.206 0.293 3.274 0.337 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 2.99 0.338 3.058 0.382 ;
      RECT 2.774 0.473 2.842 0.517 ;
      RECT 2.558 0.473 2.626 0.517 ;
      RECT 2.342 0.473 2.41 0.517 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.3455 1.87 0.3895 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.156 0.498 1.22 0.542 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.614 0.448 0.682 0.492 ;
    LAYER m1 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 1.222 0.428 1.674 0.472 ;
      RECT 1.222 0.158 1.782 0.202 ;
      RECT 1.114 0.068 1.782 0.112 ;
      RECT 2.086 0.338 2.518 0.382 ;
      RECT 1.478 0.248 1.802 0.292 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.87 0.248 2.558 0.292 ;
      RECT 2.558 0.248 2.626 0.562 ;
      RECT 2.626 0.248 2.774 0.292 ;
      RECT 2.774 0.248 2.842 0.562 ;
      RECT 2.842 0.338 3.078 0.382 ;
      RECT 3.314 0.158 3.382 0.562 ;
      RECT 3.382 0.158 3.51 0.202 ;
      RECT 3.638 0.068 3.706 0.202 ;
      RECT 3.49 0.248 3.638 0.292 ;
      RECT 3.638 0.248 3.706 0.382 ;
      RECT 3.706 0.338 3.854 0.382 ;
      RECT 3.854 0.158 3.922 0.562 ;
  END
END b15fqn003hn1n16x5

MACRO b15fqn00chn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00chn1n02x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.498 2.626 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.068 2.302 0.292 ;
      LAYER v0 ;
        RECT 2.234 0.203 2.302 0.247 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 6.08 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.472 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.574 0.112 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.068 0.466 0.112 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.366 2.518 0.41 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.566 0.158 1.978 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 0.486 0.158 0.682 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.126 0.203 2.194 0.247 ;
        RECT 2.45 0.203 2.518 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 1.242 0.248 1.91 0.292 ;
      RECT 0.81 0.518 1.046 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
    LAYER v0 ;
      RECT 2.342 0.203 2.41 0.247 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.018 0.203 2.086 0.247 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.2705 1.114 0.3145 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.83 0.2705 0.898 0.3145 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.398 0.363 0.466 0.407 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.702 0.292 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.428 0.938 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 0.898 0.068 1.782 0.112 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.33 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 2.126 0.562 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.194 0.338 2.342 0.382 ;
      RECT 2.342 0.158 2.41 0.562 ;
  END
END b15fqn00chn1n02x5

MACRO b15fqn00chn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00chn1n03x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.498 2.626 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.068 2.302 0.292 ;
      LAYER v0 ;
        RECT 2.234 0.203 2.302 0.247 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 6.08 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.472 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.574 0.112 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.068 0.466 0.112 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.366 2.518 0.41 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.566 0.158 1.978 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 0.486 0.158 0.682 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.126 0.203 2.194 0.247 ;
        RECT 2.45 0.203 2.518 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 1.242 0.248 1.91 0.292 ;
      RECT 0.81 0.518 1.046 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
    LAYER v0 ;
      RECT 2.342 0.203 2.41 0.247 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.018 0.203 2.086 0.247 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.2705 1.114 0.3145 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.83 0.2705 0.898 0.3145 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.398 0.363 0.466 0.407 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.702 0.292 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.428 0.938 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 0.898 0.068 1.782 0.112 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.33 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 2.126 0.562 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.194 0.338 2.342 0.382 ;
      RECT 2.342 0.158 2.41 0.562 ;
  END
END b15fqn00chn1n03x5

MACRO b15fqn00chn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00chn1n04x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.498 2.626 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.068 2.302 0.292 ;
      LAYER v0 ;
        RECT 2.234 0.203 2.302 0.247 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 6.08 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.472 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.574 0.112 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.068 0.466 0.112 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.366 2.518 0.41 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.566 0.158 1.978 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 0.486 0.158 0.682 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.126 0.203 2.194 0.247 ;
        RECT 2.45 0.203 2.518 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 1.242 0.248 1.91 0.292 ;
      RECT 0.81 0.518 1.046 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
    LAYER v0 ;
      RECT 2.342 0.203 2.41 0.247 ;
      RECT 2.342 0.448 2.41 0.492 ;
      RECT 2.018 0.203 2.086 0.247 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.2705 1.114 0.3145 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.83 0.2705 0.898 0.3145 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.398 0.363 0.466 0.407 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.702 0.292 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.428 0.938 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 0.898 0.068 1.782 0.112 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.33 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 2.126 0.562 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.194 0.338 2.342 0.382 ;
      RECT 2.342 0.158 2.41 0.562 ;
  END
END b15fqn00chn1n04x5

MACRO b15fqn00chn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00chn1n06x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.338 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.498 2.842 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 2.3614285 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.518 0.292 ;
      LAYER v0 ;
        RECT 2.45 0.203 2.518 0.247 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.182 0.186 0.25 0.23 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.016 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.29 0.3905 0.358 0.4345 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.666 0.366 2.734 0.41 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 2.342 -0.022 2.41 0.292 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 0.594 0.158 0.79 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.186 0.142 0.23 ;
        RECT 0.29 0.186 0.358 0.23 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 2.342 0.203 2.41 0.247 ;
        RECT 2.666 0.203 2.734 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.154 0.248 1.782 0.292 ;
      RECT 1.458 0.338 1.91 0.382 ;
      RECT 0.918 0.518 1.154 0.562 ;
      RECT 2.234 0.158 2.302 0.472 ;
    LAYER v0 ;
      RECT 2.558 0.203 2.626 0.247 ;
      RECT 2.558 0.448 2.626 0.492 ;
      RECT 2.234 0.203 2.302 0.247 ;
      RECT 2.234 0.408 2.302 0.452 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 2.018 0.3155 2.086 0.3595 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.358 1.222 0.402 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.938 0.2705 1.006 0.3145 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.363 0.574 0.407 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.248 0.81 0.292 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.006 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.158 1.802 0.202 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 1.87 0.068 1.998 0.112 ;
      RECT 1.91 0.158 1.978 0.382 ;
      RECT 1.978 0.158 2.126 0.202 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.518 1.37 0.562 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.438 0.428 2.018 0.472 ;
      RECT 2.018 0.248 2.086 0.562 ;
      RECT 2.086 0.518 2.342 0.562 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.41 0.338 2.558 0.382 ;
      RECT 2.558 0.158 2.626 0.562 ;
  END
END b15fqn00chn1n06x5

MACRO b15fqn00chn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00chn1n08x5 0 0 ;
  SIZE 3.24 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.158 3.166 0.472 ;
      LAYER v0 ;
        RECT 3.098 0.293 3.166 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.248 2.842 0.472 ;
      LAYER v0 ;
        RECT 2.774 0.293 2.842 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.87666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.274 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.882 0.4605 2.95 0.5045 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.274 0.022 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 1.566 0.158 2.214 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 0.594 0.158 0.79 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.884 0.048 2.948 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.458 0.338 2.018 0.382 ;
      RECT 0.918 0.518 1.154 0.562 ;
      RECT 2.558 0.068 2.774 0.112 ;
    LAYER v0 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 3.098 0.518 3.166 0.562 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.558 0.384 2.626 0.428 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.938 0.2705 1.006 0.3145 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.363 0.574 0.407 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.248 0.81 0.292 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.33 0.248 1.89 0.292 ;
      RECT 1.006 0.068 1.89 0.112 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 2.086 0.248 2.342 0.292 ;
      RECT 2.342 0.158 2.41 0.292 ;
      RECT 2.41 0.158 2.558 0.202 ;
      RECT 2.558 0.158 2.626 0.472 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.518 1.37 0.562 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.438 0.428 2.126 0.472 ;
      RECT 2.126 0.338 2.194 0.472 ;
      RECT 2.194 0.338 2.45 0.382 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.518 0.518 2.842 0.562 ;
      RECT 2.774 0.068 2.842 0.202 ;
      RECT 2.842 0.158 2.99 0.202 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.058 0.518 3.186 0.562 ;
      RECT 3.058 0.068 3.186 0.112 ;
  END
END b15fqn00chn1n08x5

MACRO b15fqn00chn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00chn1n12x5 0 0 ;
  SIZE 3.672 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.428 3.166 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.453 3.166 0.497 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.248 3.598 0.472 ;
      LAYER v0 ;
        RECT 3.53 0.3155 3.598 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.408 0.142 0.452 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.408 0.358 0.452 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 3.9425 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 3.154 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.706 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.398 0.493 0.466 0.537 ;
        RECT 0.614 0.493 0.682 0.537 ;
        RECT 0.938 0.383 1.006 0.427 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.018 0.538 2.086 0.582 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 3.314 0.453 3.382 0.497 ;
        RECT 3.53 0.538 3.598 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.706 0.022 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 1.89 0.158 2.626 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 3.314 0.138 3.382 0.182 ;
        RECT 3.53 0.048 3.598 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.782 0.338 2.882 0.382 ;
      RECT 1.134 0.518 1.478 0.562 ;
      RECT 2.99 0.338 3.058 0.562 ;
    LAYER v0 ;
      RECT 3.422 0.223 3.49 0.267 ;
      RECT 3.422 0.453 3.49 0.497 ;
      RECT 2.99 0.248 3.058 0.292 ;
      RECT 2.99 0.453 3.058 0.497 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.882 0.453 2.95 0.497 ;
      RECT 2.774 0.338 2.842 0.382 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.342 0.248 2.41 0.292 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.586 0.268 1.654 0.312 ;
      RECT 1.478 0.4055 1.546 0.4495 ;
      RECT 1.37 0.178 1.438 0.222 ;
      RECT 1.262 0.2705 1.33 0.3145 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.493 0.79 0.537 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.508 0.408 0.572 0.452 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.472 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.898 0.248 1.046 0.292 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.114 0.428 1.37 0.472 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 1.654 0.428 2.302 0.472 ;
      RECT 1.33 0.068 2.322 0.112 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.546 0.158 1.694 0.202 ;
      RECT 1.694 0.158 1.762 0.292 ;
      RECT 1.762 0.248 3.078 0.292 ;
      RECT 3.058 0.338 3.206 0.382 ;
      RECT 2.862 0.158 3.206 0.202 ;
      RECT 3.206 0.158 3.274 0.382 ;
      RECT 3.274 0.338 3.422 0.382 ;
      RECT 3.422 0.158 3.49 0.562 ;
  END
END b15fqn00chn1n12x5

MACRO b15fqn00chn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00chn1n16x5 0 0 ;
  SIZE 4.644 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0198 LAYER m2 ;
      ANTENNAMAXAREACAR 1.497037 LAYER m1 ;
      ANTENNAMAXAREACAR 5.734074 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 1.497037 LAYER m1 ;
      ANTENNAMAXAREACAR 5.734074 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.214 0.338 2.734 0.382 ;
        RECT 0.83 0.338 0.898 0.562 ;
      LAYER m2 ;
        RECT 0.812 0.338 2.32 0.382 ;
      LAYER v1 ;
        RECT 0.834 0.338 0.894 0.382 ;
        RECT 2.238 0.338 2.298 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 2.234 0.338 2.302 0.382 ;
        RECT 2.558 0.338 2.626 0.382 ;
    END
  END psb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.63625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.63625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.338 4.246 0.562 ;
      LAYER v0 ;
        RECT 4.178 0.453 4.246 0.497 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.502 0.248 4.57 0.472 ;
      LAYER v0 ;
        RECT 4.502 0.3155 4.57 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.4495 0.25 0.4935 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.398 0.4495 0.466 0.4935 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.678 0.652 ;
        RECT 4.502 0.518 4.57 0.652 ;
        RECT 4.286 0.518 4.354 0.652 ;
        RECT 3.854 0.428 3.922 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.666 0.4505 2.734 0.4945 ;
        RECT 3.854 0.473 3.922 0.517 ;
        RECT 4.288 0.538 4.352 0.582 ;
        RECT 4.504 0.538 4.568 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.678 0.022 ;
        RECT 4.502 -0.022 4.57 0.112 ;
        RECT 4.286 -0.022 4.354 0.202 ;
        RECT 3.854 -0.022 3.922 0.202 ;
        RECT 2.214 0.158 3.166 0.202 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
        RECT 0.29 0.113 0.358 0.157 ;
        RECT 0.506 0.113 0.574 0.157 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.882 0.158 2.95 0.202 ;
        RECT 3.854 0.138 3.922 0.182 ;
        RECT 4.286 0.138 4.354 0.182 ;
        RECT 4.502 0.048 4.57 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 1.37 0.068 1.438 0.382 ;
      RECT 1.91 0.428 2.538 0.472 ;
      RECT 2.214 0.338 2.734 0.382 ;
      RECT 1.242 0.518 1.802 0.562 ;
      RECT 2.774 0.338 2.842 0.472 ;
      RECT 3.402 0.518 3.746 0.562 ;
    LAYER v0 ;
      RECT 4.394 0.138 4.462 0.182 ;
      RECT 4.394 0.408 4.462 0.452 ;
      RECT 3.53 0.428 3.598 0.472 ;
      RECT 3.422 0.248 3.49 0.292 ;
      RECT 3.422 0.338 3.49 0.382 ;
      RECT 3.422 0.518 3.49 0.562 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 2.99 0.338 3.058 0.382 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.776 0.358 2.84 0.402 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.614 0.223 0.682 0.267 ;
      RECT 0.614 0.4495 0.682 0.4935 ;
    LAYER m1 ;
      RECT 0.938 0.248 1.006 0.562 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.222 0.428 1.478 0.472 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.546 0.428 1.674 0.472 ;
      RECT 1.546 0.158 1.89 0.202 ;
      RECT 1.438 0.068 2.97 0.112 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.87 0.248 2.882 0.292 ;
      RECT 2.882 0.248 2.95 0.382 ;
      RECT 2.95 0.338 3.51 0.382 ;
      RECT 2.842 0.428 3.638 0.472 ;
      RECT 3.098 0.248 3.638 0.292 ;
      RECT 3.638 0.248 3.706 0.472 ;
      RECT 3.294 0.158 3.746 0.202 ;
      RECT 3.746 0.158 3.814 0.562 ;
      RECT 3.814 0.248 4.394 0.292 ;
      RECT 4.394 0.068 4.462 0.472 ;
  END
END b15fqn00chn1n16x5

MACRO b15fqn00fhn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00fhn1n02x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 8.348889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 8.348889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.158 3.058 0.562 ;
        RECT 1.37 0.518 1.654 0.562 ;
      LAYER m2 ;
        RECT 1.46 0.518 3.076 0.562 ;
      LAYER v1 ;
        RECT 1.482 0.518 1.542 0.562 ;
        RECT 2.994 0.518 3.054 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.518 1.546 0.562 ;
        RECT 2.99 0.248 3.058 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.382 ;
        RECT 1.91 0.338 2.194 0.382 ;
      LAYER m2 ;
        RECT 1.984 0.338 2.644 0.382 ;
      LAYER v1 ;
        RECT 2.13 0.338 2.19 0.382 ;
        RECT 2.562 0.338 2.622 0.382 ;
      LAYER v0 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.558 0.088 2.626 0.132 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.37 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.37 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.068 3.274 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.206 0.138 3.274 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.408 0.358 0.452 ;
        RECT 0.722 0.47 0.79 0.514 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.1 0.538 3.164 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 1.262 0.158 1.978 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.666 0.203 2.734 0.247 ;
        RECT 3.098 0.138 3.166 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 0.824 0.382 ;
      RECT 0.164 0.518 1.024 0.562 ;
      RECT 0.904 0.338 1.904 0.382 ;
      RECT 0.596 0.428 2.228 0.472 ;
      RECT 2.308 0.428 3.184 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.722 0.248 0.79 0.382 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 0.83 0.518 1.114 0.562 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.37 0.518 1.654 0.562 ;
      RECT 1.694 0.248 1.762 0.382 ;
      RECT 1.91 0.338 2.194 0.382 ;
      RECT 2.126 0.428 2.234 0.472 ;
      RECT 2.126 0.158 2.342 0.202 ;
      RECT 1.478 0.068 2.45 0.112 ;
      RECT 2.774 0.248 2.842 0.562 ;
      RECT 2.558 0.068 2.626 0.382 ;
      RECT 2.666 0.428 2.734 0.562 ;
      RECT 2.99 0.158 3.058 0.562 ;
      RECT 3.098 0.248 3.166 0.472 ;
    LAYER v1 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.67 0.428 2.73 0.472 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.942 0.518 1.002 0.562 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.402 0.518 0.462 0.562 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 3.098 0.338 3.166 0.382 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.774 0.448 2.842 0.492 ;
      RECT 2.666 0.448 2.734 0.492 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.938 0.3835 1.006 0.4275 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.83 0.3835 0.898 0.4275 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.408 0.142 0.452 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.006 0.158 1.222 0.202 ;
      RECT 1.33 0.428 1.802 0.472 ;
      RECT 1.802 0.248 1.87 0.472 ;
      RECT 1.87 0.248 2.194 0.292 ;
      RECT 2.234 0.248 2.302 0.472 ;
      RECT 2.342 0.158 2.41 0.562 ;
      RECT 2.45 0.068 2.518 0.472 ;
      RECT 2.842 0.248 2.882 0.292 ;
      RECT 2.882 0.068 2.95 0.292 ;
  END
END b15fqn00fhn1n02x5

MACRO b15fqn00fhn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00fhn1n03x5 0 0 ;
  SIZE 3.564 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 6.679111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 6.679111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.158 3.274 0.562 ;
        RECT 1.37 0.518 1.654 0.562 ;
      LAYER m2 ;
        RECT 1.46 0.518 3.292 0.562 ;
      LAYER v1 ;
        RECT 1.482 0.518 1.542 0.562 ;
        RECT 3.21 0.518 3.27 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.518 1.546 0.562 ;
        RECT 3.206 0.248 3.274 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.068 2.842 0.382 ;
        RECT 2.214 0.338 2.41 0.382 ;
      LAYER m2 ;
        RECT 2.308 0.338 2.86 0.382 ;
      LAYER v1 ;
        RECT 2.346 0.338 2.406 0.382 ;
        RECT 2.778 0.338 2.838 0.382 ;
      LAYER v0 ;
        RECT 2.234 0.338 2.302 0.382 ;
        RECT 2.774 0.088 2.842 0.132 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.37 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.37 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.068 3.49 0.562 ;
      LAYER v0 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.422 0.138 3.49 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.408 0.358 0.452 ;
        RECT 0.722 0.47 0.79 0.514 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 2.126 0.538 2.194 0.582 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.316 0.538 3.38 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.598 0.022 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 2.882 -0.022 2.95 0.292 ;
        RECT 1.262 0.158 1.978 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.882 0.203 2.95 0.247 ;
        RECT 3.314 0.138 3.382 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 0.824 0.382 ;
      RECT 0.164 0.518 1.024 0.562 ;
      RECT 0.904 0.338 2.228 0.382 ;
      RECT 0.596 0.428 2.444 0.472 ;
      RECT 2.524 0.428 3.4 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.722 0.248 0.79 0.382 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 0.83 0.518 1.114 0.562 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.37 0.518 1.654 0.562 ;
      RECT 1.91 0.338 2.106 0.382 ;
      RECT 2.342 0.428 2.45 0.472 ;
      RECT 2.214 0.338 2.41 0.382 ;
      RECT 2.43 0.158 2.558 0.202 ;
      RECT 1.478 0.068 2.666 0.112 ;
      RECT 2.99 0.248 3.058 0.562 ;
      RECT 2.774 0.068 2.842 0.382 ;
      RECT 2.882 0.428 2.95 0.562 ;
      RECT 3.206 0.158 3.274 0.562 ;
      RECT 3.314 0.248 3.382 0.472 ;
    LAYER v1 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.942 0.518 1.002 0.562 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.402 0.518 0.462 0.562 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 3.098 0.138 3.166 0.182 ;
      RECT 2.99 0.448 3.058 0.492 ;
      RECT 2.882 0.448 2.95 0.492 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.938 0.3835 1.006 0.4275 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.83 0.3835 0.898 0.4275 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.408 0.142 0.452 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.006 0.158 1.222 0.202 ;
      RECT 1.33 0.428 1.802 0.472 ;
      RECT 1.802 0.248 1.87 0.472 ;
      RECT 1.87 0.428 1.998 0.472 ;
      RECT 1.87 0.248 2.322 0.292 ;
      RECT 2.45 0.248 2.518 0.472 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 2.666 0.068 2.734 0.472 ;
      RECT 3.058 0.248 3.098 0.292 ;
      RECT 3.098 0.068 3.166 0.292 ;
  END
END b15fqn00fhn1n03x5

MACRO b15fqn00fhn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00fhn1n04x5 0 0 ;
  SIZE 3.564 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 5.751111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 5.751111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.158 3.274 0.562 ;
        RECT 1.37 0.518 1.654 0.562 ;
      LAYER m2 ;
        RECT 1.46 0.518 3.292 0.562 ;
      LAYER v1 ;
        RECT 1.482 0.518 1.542 0.562 ;
        RECT 3.21 0.518 3.27 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.518 1.546 0.562 ;
        RECT 3.206 0.248 3.274 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.068 2.842 0.382 ;
        RECT 2.214 0.338 2.41 0.382 ;
      LAYER m2 ;
        RECT 2.308 0.338 2.86 0.382 ;
      LAYER v1 ;
        RECT 2.346 0.338 2.406 0.382 ;
        RECT 2.778 0.338 2.838 0.382 ;
      LAYER v0 ;
        RECT 2.234 0.338 2.302 0.382 ;
        RECT 2.774 0.088 2.842 0.132 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.37 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.37 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.068 3.49 0.562 ;
      LAYER v0 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.422 0.138 3.49 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.408 0.358 0.452 ;
        RECT 0.722 0.47 0.79 0.514 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 2.126 0.538 2.194 0.582 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.316 0.538 3.38 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.598 0.022 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 2.882 -0.022 2.95 0.292 ;
        RECT 1.262 0.158 1.978 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.882 0.203 2.95 0.247 ;
        RECT 3.314 0.138 3.382 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 0.824 0.382 ;
      RECT 0.164 0.518 1.024 0.562 ;
      RECT 0.904 0.338 2.228 0.382 ;
      RECT 0.596 0.428 2.444 0.472 ;
      RECT 2.524 0.428 3.4 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.722 0.248 0.79 0.382 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 0.83 0.518 1.114 0.562 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.37 0.518 1.654 0.562 ;
      RECT 1.91 0.338 2.106 0.382 ;
      RECT 2.342 0.428 2.45 0.472 ;
      RECT 2.214 0.338 2.41 0.382 ;
      RECT 2.43 0.158 2.558 0.202 ;
      RECT 1.478 0.068 2.666 0.112 ;
      RECT 2.99 0.248 3.058 0.562 ;
      RECT 2.774 0.068 2.842 0.382 ;
      RECT 2.882 0.428 2.95 0.562 ;
      RECT 3.206 0.158 3.274 0.562 ;
      RECT 3.314 0.248 3.382 0.472 ;
    LAYER v1 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.346 0.428 2.406 0.472 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.942 0.518 1.002 0.562 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.402 0.518 0.462 0.562 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 3.098 0.138 3.166 0.182 ;
      RECT 2.99 0.448 3.058 0.492 ;
      RECT 2.882 0.448 2.95 0.492 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.938 0.3835 1.006 0.4275 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.83 0.3835 0.898 0.4275 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.408 0.142 0.452 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.006 0.158 1.222 0.202 ;
      RECT 1.33 0.428 1.478 0.472 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.546 0.428 1.998 0.472 ;
      RECT 1.546 0.248 2.322 0.292 ;
      RECT 2.45 0.248 2.518 0.472 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 2.666 0.068 2.734 0.472 ;
      RECT 3.058 0.248 3.098 0.292 ;
      RECT 3.098 0.068 3.166 0.292 ;
  END
END b15fqn00fhn1n04x5

MACRO b15fqn00fhn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00fhn1n06x5 0 0 ;
  SIZE 3.888 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 6.679111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 6.679111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.158 3.49 0.562 ;
        RECT 1.37 0.518 1.654 0.562 ;
      LAYER m2 ;
        RECT 1.46 0.518 3.508 0.562 ;
      LAYER v1 ;
        RECT 1.482 0.518 1.542 0.562 ;
        RECT 3.426 0.518 3.486 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.518 1.546 0.562 ;
        RECT 3.422 0.248 3.49 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.068 3.058 0.382 ;
        RECT 2.43 0.338 2.626 0.382 ;
      LAYER m2 ;
        RECT 2.416 0.338 3.076 0.382 ;
      LAYER v1 ;
        RECT 2.454 0.338 2.514 0.382 ;
        RECT 2.994 0.338 3.054 0.382 ;
      LAYER v0 ;
        RECT 2.45 0.338 2.518 0.382 ;
        RECT 2.99 0.088 3.058 0.132 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.068 3.706 0.562 ;
      LAYER v0 ;
        RECT 3.638 0.448 3.706 0.492 ;
        RECT 3.638 0.138 3.706 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.922 0.652 ;
        RECT 3.746 0.338 3.814 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.389 0.358 0.433 ;
        RECT 0.722 0.47 0.79 0.514 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.532 0.538 3.596 0.582 ;
        RECT 3.746 0.448 3.814 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.922 0.022 ;
        RECT 3.746 -0.022 3.814 0.292 ;
        RECT 3.53 -0.022 3.598 0.202 ;
        RECT 3.098 -0.022 3.166 0.292 ;
        RECT 1.262 0.158 2.106 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 3.098 0.203 3.166 0.247 ;
        RECT 3.53 0.138 3.598 0.182 ;
        RECT 3.746 0.138 3.814 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 0.824 0.382 ;
      RECT 0.164 0.518 1.132 0.562 ;
      RECT 0.904 0.338 2.336 0.382 ;
      RECT 0.596 0.428 2.66 0.472 ;
      RECT 2.74 0.428 3.616 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.722 0.248 0.79 0.382 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.83 0.518 1.134 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.37 0.518 1.654 0.562 ;
      RECT 2.126 0.338 2.322 0.382 ;
      RECT 2.45 0.428 2.666 0.472 ;
      RECT 2.43 0.338 2.626 0.382 ;
      RECT 2.646 0.158 2.774 0.202 ;
      RECT 1.478 0.068 2.882 0.112 ;
      RECT 3.206 0.248 3.274 0.562 ;
      RECT 2.99 0.068 3.058 0.382 ;
      RECT 3.098 0.428 3.166 0.562 ;
      RECT 3.422 0.158 3.49 0.562 ;
      RECT 3.53 0.248 3.598 0.472 ;
    LAYER v1 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.238 0.338 2.298 0.382 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 1.05 0.518 1.11 0.562 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.402 0.518 0.462 0.562 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 3.53 0.338 3.598 0.382 ;
      RECT 3.314 0.138 3.382 0.182 ;
      RECT 3.206 0.448 3.274 0.492 ;
      RECT 3.098 0.448 3.166 0.492 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.3835 1.006 0.4275 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.83 0.3835 0.898 0.4275 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.498 0.466 0.542 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.389 0.142 0.433 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.006 0.158 1.222 0.202 ;
      RECT 1.33 0.428 1.478 0.472 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.546 0.248 2.018 0.292 ;
      RECT 2.018 0.248 2.086 0.562 ;
      RECT 2.086 0.248 2.538 0.292 ;
      RECT 2.666 0.248 2.734 0.472 ;
      RECT 2.774 0.158 2.842 0.562 ;
      RECT 2.882 0.068 2.95 0.472 ;
      RECT 3.274 0.248 3.314 0.292 ;
      RECT 3.314 0.068 3.382 0.292 ;
  END
END b15fqn00fhn1n06x5

MACRO b15fqn00fhn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00fhn1n08x5 0 0 ;
  SIZE 4.428 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 5.751111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 5.751111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.158 4.03 0.562 ;
        RECT 1.586 0.518 1.87 0.562 ;
      LAYER m2 ;
        RECT 1.676 0.518 4.048 0.562 ;
      LAYER v1 ;
        RECT 1.698 0.518 1.758 0.562 ;
        RECT 3.966 0.518 4.026 0.562 ;
      LAYER v0 ;
        RECT 1.694 0.518 1.762 0.562 ;
        RECT 3.962 0.248 4.03 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.598 0.382 ;
        RECT 2.862 0.338 3.166 0.382 ;
      LAYER m2 ;
        RECT 3.08 0.338 3.616 0.382 ;
      LAYER v1 ;
        RECT 3.102 0.338 3.162 0.382 ;
        RECT 3.534 0.338 3.594 0.382 ;
      LAYER v0 ;
        RECT 2.99 0.338 3.058 0.382 ;
        RECT 3.53 0.088 3.598 0.132 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.068 4.246 0.562 ;
      LAYER v0 ;
        RECT 4.178 0.448 4.246 0.492 ;
        RECT 4.178 0.138 4.246 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.462 0.652 ;
        RECT 4.286 0.428 4.354 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.854 0.428 3.922 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.126 0.338 2.194 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.408 0.358 0.452 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.91 0.3835 1.978 0.4275 ;
        RECT 2.128 0.428 2.192 0.472 ;
        RECT 2.882 0.538 2.95 0.582 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 4.072 0.538 4.136 0.582 ;
        RECT 4.286 0.448 4.354 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.462 0.022 ;
        RECT 4.286 -0.022 4.354 0.202 ;
        RECT 4.07 -0.022 4.138 0.202 ;
        RECT 3.638 -0.022 3.706 0.292 ;
        RECT 1.478 0.158 2.646 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 3.638 0.203 3.706 0.247 ;
        RECT 4.07 0.138 4.138 0.182 ;
        RECT 4.286 0.138 4.354 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 1.04 0.382 ;
      RECT 0.38 0.518 1.24 0.562 ;
      RECT 1.12 0.338 2.536 0.382 ;
      RECT 0.596 0.428 3.2 0.472 ;
      RECT 3.28 0.428 4.156 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.83 0.248 0.898 0.382 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.154 0.518 1.35 0.562 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.586 0.518 1.87 0.562 ;
      RECT 2.342 0.338 2.754 0.382 ;
      RECT 2.862 0.338 3.166 0.382 ;
      RECT 2.99 0.428 3.206 0.472 ;
      RECT 3.098 0.158 3.314 0.202 ;
      RECT 1.694 0.068 3.422 0.112 ;
      RECT 3.746 0.248 3.814 0.562 ;
      RECT 3.53 0.068 3.598 0.382 ;
      RECT 3.638 0.428 3.706 0.562 ;
      RECT 3.962 0.158 4.03 0.562 ;
      RECT 4.07 0.248 4.138 0.472 ;
    LAYER v1 ;
      RECT 4.074 0.428 4.134 0.472 ;
      RECT 3.642 0.428 3.702 0.472 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.454 0.338 2.514 0.382 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 1.158 0.518 1.218 0.562 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.402 0.518 0.462 0.562 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 4.07 0.338 4.138 0.382 ;
      RECT 3.854 0.138 3.922 0.182 ;
      RECT 3.746 0.448 3.814 0.492 ;
      RECT 3.638 0.448 3.706 0.492 ;
      RECT 3.422 0.338 3.49 0.382 ;
      RECT 3.314 0.068 3.382 0.112 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.206 0.338 3.274 0.382 ;
      RECT 2.99 0.248 3.058 0.292 ;
      RECT 2.774 0.248 2.842 0.292 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.154 0.3835 1.222 0.4275 ;
      RECT 1.048 0.088 1.112 0.132 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.4055 0.142 0.4495 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.466 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.158 1.046 0.202 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.222 0.158 1.438 0.202 ;
      RECT 1.546 0.428 1.802 0.472 ;
      RECT 1.802 0.248 1.87 0.472 ;
      RECT 1.87 0.248 2.234 0.292 ;
      RECT 2.234 0.248 2.302 0.472 ;
      RECT 2.302 0.428 2.95 0.472 ;
      RECT 2.302 0.248 3.166 0.292 ;
      RECT 3.206 0.248 3.274 0.472 ;
      RECT 3.314 0.158 3.382 0.562 ;
      RECT 3.422 0.068 3.49 0.472 ;
      RECT 3.814 0.248 3.854 0.292 ;
      RECT 3.854 0.068 3.922 0.292 ;
  END
END b15fqn00fhn1n08x5

MACRO b15fqn00fhn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00fhn1n12x5 0 0 ;
  SIZE 5.508 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 5.565926 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 5.565926 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.934 0.158 5.002 0.562 ;
        RECT 2.234 0.428 2.302 0.562 ;
      LAYER m2 ;
        RECT 2.216 0.518 5.02 0.562 ;
      LAYER v1 ;
        RECT 2.238 0.518 2.298 0.562 ;
        RECT 4.938 0.518 4.998 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.49 2.302 0.534 ;
        RECT 4.934 0.248 5.002 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAGATEAREA 0.0207 LAYER m2 ;
      ANTENNAMAXAREACAR 2.49714275 LAYER m1 ;
      ANTENNAMAXAREACAR 6.640635 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.89396825 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
      ANTENNAMAXAREACAR 7.7474075 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.248 4.786 0.292 ;
        RECT 4.718 0.068 4.786 0.292 ;
        RECT 4.61 0.248 4.678 0.382 ;
        RECT 3.53 0.338 3.726 0.382 ;
      LAYER m2 ;
        RECT 3.604 0.338 4.696 0.382 ;
      LAYER v1 ;
        RECT 3.642 0.338 3.702 0.382 ;
        RECT 4.614 0.338 4.674 0.382 ;
      LAYER v0 ;
        RECT 3.638 0.338 3.706 0.382 ;
        RECT 4.718 0.138 4.786 0.182 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.366 0.068 5.434 0.562 ;
        RECT 5.15 0.338 5.434 0.382 ;
        RECT 5.15 0.068 5.218 0.562 ;
      LAYER v0 ;
        RECT 5.15 0.448 5.218 0.492 ;
        RECT 5.15 0.138 5.218 0.182 ;
        RECT 5.366 0.448 5.434 0.492 ;
        RECT 5.366 0.138 5.434 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.542 0.652 ;
        RECT 5.258 0.428 5.326 0.652 ;
        RECT 5.042 0.518 5.11 0.652 ;
        RECT 4.826 0.428 4.894 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 3.638 0.518 3.706 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.154 0.4575 1.222 0.5015 ;
        RECT 1.91 0.538 1.978 0.582 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 3.64 0.538 3.704 0.582 ;
        RECT 4.502 0.448 4.57 0.492 ;
        RECT 4.826 0.448 4.894 0.492 ;
        RECT 5.044 0.538 5.108 0.582 ;
        RECT 5.258 0.448 5.326 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.542 0.022 ;
        RECT 5.258 -0.022 5.326 0.292 ;
        RECT 5.042 -0.022 5.11 0.202 ;
        RECT 4.61 -0.022 4.678 0.202 ;
        RECT 1.91 0.158 3.186 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.154 0.203 1.222 0.247 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.882 0.158 2.95 0.202 ;
        RECT 3.098 0.158 3.166 0.202 ;
        RECT 4.61 0.138 4.678 0.182 ;
        RECT 5.042 0.138 5.11 0.182 ;
        RECT 5.258 0.138 5.326 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 1.024 0.382 ;
      RECT 0.164 0.518 1.456 0.562 ;
      RECT 1.568 0.338 3.524 0.382 ;
      RECT 0.596 0.428 4.172 0.472 ;
      RECT 4.252 0.428 5.128 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 3.098 0.248 3.166 0.472 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 3.422 0.338 3.49 0.472 ;
      RECT 3.53 0.338 3.726 0.382 ;
      RECT 3.294 0.158 3.726 0.202 ;
      RECT 3.962 0.338 4.03 0.562 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 4.07 0.338 4.138 0.562 ;
      RECT 2.126 0.068 4.394 0.112 ;
      RECT 4.61 0.248 4.678 0.382 ;
      RECT 4.61 0.428 4.678 0.562 ;
      RECT 4.718 0.338 4.786 0.562 ;
      RECT 4.934 0.158 5.002 0.562 ;
      RECT 5.042 0.248 5.11 0.472 ;
    LAYER v1 ;
      RECT 5.046 0.428 5.106 0.472 ;
      RECT 4.614 0.428 4.674 0.472 ;
      RECT 4.29 0.428 4.35 0.472 ;
      RECT 3.966 0.428 4.026 0.472 ;
      RECT 3.426 0.338 3.486 0.382 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.402 0.518 0.462 0.562 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 5.042 0.338 5.11 0.382 ;
      RECT 4.826 0.138 4.894 0.182 ;
      RECT 4.718 0.448 4.786 0.492 ;
      RECT 4.61 0.448 4.678 0.492 ;
      RECT 4.394 0.338 4.462 0.382 ;
      RECT 4.288 0.448 4.352 0.492 ;
      RECT 4.178 0.158 4.246 0.202 ;
      RECT 4.178 0.3675 4.246 0.4115 ;
      RECT 4.07 0.068 4.138 0.112 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 4.072 0.448 4.136 0.492 ;
      RECT 3.962 0.158 4.03 0.202 ;
      RECT 3.962 0.3675 4.03 0.4115 ;
      RECT 3.746 0.248 3.814 0.292 ;
      RECT 3.746 0.428 3.814 0.472 ;
      RECT 3.638 0.158 3.706 0.202 ;
      RECT 3.53 0.248 3.598 0.292 ;
      RECT 3.422 0.3835 3.49 0.4275 ;
      RECT 3.422 0.518 3.49 0.562 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.098 0.383 3.166 0.427 ;
      RECT 2.882 0.428 2.95 0.472 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.478 0.203 1.546 0.247 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.4575 1.33 0.5015 ;
      RECT 1.046 0.203 1.114 0.247 ;
      RECT 1.046 0.4575 1.114 0.5015 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.338 1.262 0.382 ;
      RECT 1.262 0.068 1.33 0.562 ;
      RECT 1.33 0.068 1.478 0.112 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 1.546 0.338 1.586 0.382 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 1.654 0.158 1.87 0.202 ;
      RECT 3.098 0.518 3.53 0.562 ;
      RECT 3.53 0.428 3.598 0.562 ;
      RECT 3.598 0.428 3.854 0.472 ;
      RECT 3.166 0.248 3.854 0.292 ;
      RECT 3.854 0.248 3.922 0.472 ;
      RECT 3.922 0.248 4.178 0.292 ;
      RECT 4.178 0.248 4.246 0.472 ;
      RECT 1.978 0.428 2.126 0.472 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.194 0.248 2.882 0.292 ;
      RECT 2.882 0.248 2.95 0.562 ;
      RECT 2.95 0.518 3.098 0.562 ;
      RECT 2.95 0.248 3.098 0.292 ;
      RECT 4.138 0.518 4.286 0.562 ;
      RECT 3.942 0.158 4.286 0.202 ;
      RECT 4.286 0.158 4.354 0.562 ;
      RECT 4.394 0.068 4.462 0.472 ;
      RECT 4.678 0.248 4.718 0.292 ;
      RECT 4.718 0.068 4.786 0.292 ;
      RECT 4.786 0.338 4.826 0.382 ;
      RECT 4.826 0.068 4.894 0.382 ;
  END
END b15fqn00fhn1n12x5

MACRO b15fqn00fhn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn00fhn1n16x5 0 0 ;
  SIZE 6.372 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAGATEAREA 0.0135 LAYER m2 ;
      ANTENNAMAXAREACAR 0.711746 LAYER m1 ;
      ANTENNAMAXAREACAR 5.072381 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.89396825 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAGATEAREA 0.0135 LAYER m2 ;
      ANTENNAMAXAREACAR 0.711746 LAYER m1 ;
      ANTENNAMAXAREACAR 5.072381 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.89396825 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.69 0.158 5.758 0.562 ;
        RECT 2.45 0.428 2.518 0.562 ;
      LAYER m2 ;
        RECT 2.432 0.518 5.776 0.562 ;
      LAYER v1 ;
        RECT 2.454 0.518 2.514 0.562 ;
        RECT 5.694 0.518 5.754 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.49 2.518 0.534 ;
        RECT 5.69 0.248 5.758 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAGATEAREA 0.0279 LAYER m2 ;
      ANTENNAMAXAREACAR 2.49714275 LAYER m1 ;
      ANTENNAMAXAREACAR 6.640635 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.89396825 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0351 LAYER m2 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
      ANTENNAMAXAREACAR 7.7474075 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.258 0.248 5.434 0.292 ;
        RECT 5.366 0.068 5.434 0.292 ;
        RECT 5.258 0.248 5.326 0.382 ;
        RECT 4.07 0.338 4.266 0.382 ;
      LAYER m2 ;
        RECT 4.144 0.338 5.344 0.382 ;
      LAYER v1 ;
        RECT 4.182 0.338 4.242 0.382 ;
        RECT 5.262 0.338 5.322 0.382 ;
      LAYER v0 ;
        RECT 4.178 0.338 4.246 0.382 ;
        RECT 5.366 0.138 5.434 0.182 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 6.122 0.068 6.19 0.562 ;
        RECT 5.906 0.338 6.19 0.382 ;
        RECT 5.906 0.068 5.974 0.562 ;
      LAYER v0 ;
        RECT 5.906 0.448 5.974 0.492 ;
        RECT 5.906 0.138 5.974 0.182 ;
        RECT 6.122 0.448 6.19 0.492 ;
        RECT 6.122 0.138 6.19 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.406 0.652 ;
        RECT 6.23 0.428 6.298 0.652 ;
        RECT 6.014 0.428 6.082 0.652 ;
        RECT 5.798 0.518 5.866 0.652 ;
        RECT 5.474 0.428 5.542 0.652 ;
        RECT 5.15 0.428 5.218 0.652 ;
        RECT 4.394 0.518 4.462 0.652 ;
        RECT 4.178 0.518 4.246 0.652 ;
        RECT 3.098 0.338 3.166 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.154 0.4575 1.222 0.5015 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.666 0.403 2.734 0.447 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 3.098 0.428 3.166 0.472 ;
        RECT 4.18 0.538 4.244 0.582 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 5.15 0.448 5.218 0.492 ;
        RECT 5.474 0.448 5.542 0.492 ;
        RECT 5.8 0.538 5.864 0.582 ;
        RECT 6.014 0.448 6.082 0.492 ;
        RECT 6.23 0.448 6.298 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.406 0.022 ;
        RECT 6.23 -0.022 6.298 0.292 ;
        RECT 6.014 -0.022 6.082 0.292 ;
        RECT 5.798 -0.022 5.866 0.202 ;
        RECT 5.258 -0.022 5.326 0.202 ;
        RECT 1.91 0.158 3.834 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.154 0.203 1.222 0.247 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.882 0.158 2.95 0.202 ;
        RECT 3.098 0.158 3.166 0.202 ;
        RECT 3.314 0.158 3.382 0.202 ;
        RECT 3.53 0.158 3.598 0.202 ;
        RECT 3.746 0.158 3.814 0.202 ;
        RECT 5.258 0.138 5.326 0.182 ;
        RECT 5.798 0.138 5.866 0.182 ;
        RECT 6.014 0.138 6.082 0.182 ;
        RECT 6.23 0.138 6.298 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 1.024 0.382 ;
      RECT 0.164 0.518 1.348 0.562 ;
      RECT 1.784 0.338 4.064 0.382 ;
      RECT 0.596 0.428 4.712 0.472 ;
      RECT 4.792 0.428 5.884 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 3.53 0.338 3.598 0.562 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 2.45 0.428 2.518 0.562 ;
      RECT 3.962 0.338 4.03 0.472 ;
      RECT 4.07 0.338 4.266 0.382 ;
      RECT 3.942 0.158 4.482 0.202 ;
      RECT 4.502 0.338 4.57 0.562 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 4.718 0.338 4.786 0.562 ;
      RECT 2.106 0.068 5.042 0.112 ;
      RECT 5.258 0.248 5.326 0.382 ;
      RECT 5.258 0.428 5.326 0.562 ;
      RECT 5.366 0.338 5.434 0.562 ;
      RECT 5.69 0.158 5.758 0.562 ;
      RECT 5.798 0.248 5.866 0.472 ;
    LAYER v1 ;
      RECT 5.802 0.428 5.862 0.472 ;
      RECT 5.262 0.428 5.322 0.472 ;
      RECT 4.938 0.428 4.998 0.472 ;
      RECT 4.506 0.428 4.566 0.472 ;
      RECT 3.966 0.338 4.026 0.382 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.806 0.338 1.866 0.382 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.266 0.518 1.326 0.562 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.402 0.518 0.462 0.562 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 5.798 0.338 5.866 0.382 ;
      RECT 5.582 0.448 5.65 0.492 ;
      RECT 5.474 0.138 5.542 0.182 ;
      RECT 5.366 0.448 5.434 0.492 ;
      RECT 5.258 0.448 5.326 0.492 ;
      RECT 5.042 0.338 5.11 0.382 ;
      RECT 4.936 0.448 5 0.492 ;
      RECT 4.826 0.158 4.894 0.202 ;
      RECT 4.826 0.3675 4.894 0.4115 ;
      RECT 4.718 0.248 4.786 0.292 ;
      RECT 4.72 0.448 4.784 0.492 ;
      RECT 4.61 0.158 4.678 0.202 ;
      RECT 4.61 0.3675 4.678 0.4115 ;
      RECT 4.502 0.068 4.57 0.112 ;
      RECT 4.502 0.448 4.57 0.492 ;
      RECT 4.394 0.158 4.462 0.202 ;
      RECT 4.286 0.248 4.354 0.292 ;
      RECT 4.286 0.428 4.354 0.472 ;
      RECT 4.178 0.158 4.246 0.202 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 3.962 0.158 4.03 0.202 ;
      RECT 3.962 0.3835 4.03 0.4275 ;
      RECT 3.962 0.518 4.03 0.562 ;
      RECT 3.746 0.383 3.814 0.427 ;
      RECT 3.53 0.428 3.598 0.472 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.383 1.978 0.427 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.479 1.87 0.523 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.262 0.4575 1.33 0.5015 ;
      RECT 1.046 0.203 1.114 0.247 ;
      RECT 1.046 0.4575 1.114 0.5015 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.338 1.478 0.382 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.546 0.158 1.762 0.202 ;
      RECT 1.438 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 3.53 0.248 3.746 0.292 ;
      RECT 3.746 0.248 3.814 0.472 ;
      RECT 3.598 0.518 4.07 0.562 ;
      RECT 4.07 0.428 4.138 0.562 ;
      RECT 4.138 0.428 4.394 0.472 ;
      RECT 3.814 0.248 4.394 0.292 ;
      RECT 4.394 0.248 4.462 0.472 ;
      RECT 4.462 0.248 4.61 0.292 ;
      RECT 4.61 0.248 4.678 0.562 ;
      RECT 4.678 0.248 4.826 0.292 ;
      RECT 4.826 0.248 4.894 0.472 ;
      RECT 2.086 0.428 2.234 0.472 ;
      RECT 2.234 0.248 2.302 0.472 ;
      RECT 2.302 0.248 3.314 0.292 ;
      RECT 3.314 0.248 3.382 0.562 ;
      RECT 3.382 0.518 3.53 0.562 ;
      RECT 3.382 0.248 3.53 0.292 ;
      RECT 4.786 0.518 4.934 0.562 ;
      RECT 4.59 0.158 4.934 0.202 ;
      RECT 4.934 0.158 5.002 0.562 ;
      RECT 5.042 0.068 5.11 0.472 ;
      RECT 5.326 0.248 5.366 0.292 ;
      RECT 5.366 0.068 5.434 0.292 ;
      RECT 5.434 0.338 5.474 0.382 ;
      RECT 5.474 0.068 5.542 0.382 ;
      RECT 5.542 0.338 5.582 0.382 ;
      RECT 5.582 0.338 5.65 0.562 ;
  END
END b15fqn00fhn1n16x5

MACRO b15fqn043hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn043hn1n02x5 0 0 ;
  SIZE 3.564 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.338 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.498 2.518 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.248 3.382 0.472 ;
      LAYER v0 ;
        RECT 3.314 0.338 3.382 0.382 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 3.166 0.382 ;
        RECT 3.098 0.158 3.166 0.382 ;
      LAYER v0 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 2.882 0.338 2.95 0.382 ;
        RECT 3.098 0.248 3.166 0.292 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.182 0.203 0.25 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.9825 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.586 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.088 0.574 0.132 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.5235 0.142 0.5675 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 1.154 0.472 1.222 0.516 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 2.342 0.403 2.41 0.447 ;
        RECT 2.774 0.472 2.842 0.516 ;
        RECT 3.314 0.538 3.382 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.598 0.022 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.0915 0.142 0.1355 ;
        RECT 0.398 0.203 0.466 0.247 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 3.314 0.138 3.382 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.068 2.536 0.112 ;
      RECT 2.864 0.068 3.524 0.112 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.614 0.068 0.682 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 0.702 0.518 0.938 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 2.45 0.068 2.646 0.112 ;
      RECT 2.97 0.428 3.206 0.472 ;
      RECT 3.422 0.068 3.49 0.562 ;
    LAYER v1 ;
      RECT 3.426 0.068 3.486 0.112 ;
      RECT 2.886 0.068 2.946 0.112 ;
      RECT 2.454 0.068 2.514 0.112 ;
      RECT 0.618 0.068 0.678 0.112 ;
      RECT 0.294 0.068 0.354 0.112 ;
    LAYER v0 ;
      RECT 3.422 0.138 3.49 0.182 ;
      RECT 3.422 0.4185 3.49 0.4625 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.234 0.403 2.302 0.447 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.018 0.178 2.086 0.222 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.804 0.178 1.868 0.222 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.154 0.268 1.222 0.312 ;
      RECT 1.046 0.472 1.114 0.516 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.4 0.358 0.464 0.402 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.398 0.338 0.466 0.472 ;
      RECT 0.466 0.428 0.83 0.472 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.114 0.338 1.154 0.382 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.438 0.248 1.802 0.292 ;
      RECT 1.802 0.158 1.87 0.292 ;
      RECT 1.87 0.248 1.91 0.292 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 0.79 0.068 1.478 0.112 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 1.546 0.158 1.694 0.202 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.762 0.068 2.214 0.112 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.006 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.518 1.478 0.562 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.546 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 2.234 0.562 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 2.086 0.248 2.882 0.292 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 3.078 0.068 3.206 0.112 ;
      RECT 3.206 0.068 3.274 0.472 ;
  END
END b15fqn043hn1n02x5

MACRO b15fqn043hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn043hn1n03x5 0 0 ;
  SIZE 3.672 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.498 2.626 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.248 3.49 0.472 ;
      LAYER v0 ;
        RECT 3.422 0.338 3.49 0.382 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.338 3.274 0.382 ;
        RECT 3.206 0.158 3.274 0.382 ;
      LAYER v0 ;
        RECT 2.774 0.338 2.842 0.382 ;
        RECT 2.99 0.338 3.058 0.382 ;
        RECT 3.206 0.248 3.274 0.292 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.95875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.567 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.706 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.262 0.338 1.33 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 1.262 0.472 1.33 0.516 ;
        RECT 1.694 0.473 1.762 0.517 ;
        RECT 2.45 0.403 2.518 0.447 ;
        RECT 2.882 0.472 2.95 0.516 ;
        RECT 3.422 0.538 3.49 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.706 0.022 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.178 0.574 0.222 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.422 0.138 3.49 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.068 2.644 0.112 ;
      RECT 2.972 0.068 3.632 0.112 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 0.81 0.518 1.154 0.562 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 2.558 0.068 2.754 0.112 ;
      RECT 3.078 0.428 3.314 0.472 ;
      RECT 3.53 0.068 3.598 0.562 ;
    LAYER v1 ;
      RECT 3.534 0.068 3.594 0.112 ;
      RECT 2.994 0.068 3.054 0.112 ;
      RECT 2.562 0.068 2.622 0.112 ;
      RECT 0.726 0.068 0.786 0.112 ;
      RECT 0.294 0.068 0.354 0.112 ;
    LAYER v0 ;
      RECT 3.53 0.138 3.598 0.182 ;
      RECT 3.53 0.4185 3.598 0.4625 ;
      RECT 3.206 0.068 3.274 0.112 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.342 0.403 2.41 0.447 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.126 0.178 2.194 0.222 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.912 0.178 1.976 0.222 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.83 0.2705 0.898 0.3145 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.2705 0.79 0.3145 ;
      RECT 0.508 0.358 0.572 0.402 ;
      RECT 0.29 0.203 0.358 0.247 ;
      RECT 0.29 0.3905 0.358 0.4345 ;
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 0.574 0.428 0.938 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.114 0.158 1.35 0.202 ;
      RECT 1.546 0.248 1.91 0.292 ;
      RECT 1.91 0.158 1.978 0.292 ;
      RECT 1.978 0.248 2.018 0.292 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 0.898 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.202 ;
      RECT 1.654 0.158 1.802 0.202 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 1.87 0.068 2.322 0.112 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.438 0.518 1.586 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.654 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.978 0.518 2.342 0.562 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.194 0.248 2.99 0.292 ;
      RECT 2.99 0.068 3.058 0.292 ;
      RECT 3.186 0.068 3.314 0.112 ;
      RECT 3.314 0.068 3.382 0.472 ;
  END
END b15fqn043hn1n03x5

MACRO b15fqn043hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn043hn1n04x5 0 0 ;
  SIZE 3.672 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.498 2.626 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.248 3.49 0.472 ;
      LAYER v0 ;
        RECT 3.422 0.338 3.49 0.382 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.338 3.274 0.382 ;
        RECT 3.206 0.158 3.274 0.382 ;
      LAYER v0 ;
        RECT 2.774 0.338 2.842 0.382 ;
        RECT 2.99 0.338 3.058 0.382 ;
        RECT 3.206 0.248 3.274 0.292 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.25916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.706 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.674 0.428 1.87 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 2.45 0.403 2.518 0.447 ;
        RECT 2.882 0.472 2.95 0.516 ;
        RECT 3.422 0.538 3.49 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.706 0.022 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.198 0.574 0.242 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.422 0.138 3.49 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.068 2.644 0.112 ;
      RECT 2.972 0.068 3.632 0.112 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.89 0.158 2.018 0.202 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 0.81 0.518 1.046 0.562 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 2.558 0.068 2.754 0.112 ;
      RECT 3.078 0.428 3.314 0.472 ;
      RECT 3.53 0.068 3.598 0.562 ;
    LAYER v1 ;
      RECT 3.534 0.068 3.594 0.112 ;
      RECT 2.994 0.068 3.054 0.112 ;
      RECT 2.562 0.068 2.622 0.112 ;
      RECT 0.726 0.068 0.786 0.112 ;
      RECT 0.294 0.068 0.354 0.112 ;
    LAYER v0 ;
      RECT 3.53 0.138 3.598 0.182 ;
      RECT 3.53 0.4225 3.598 0.4665 ;
      RECT 3.206 0.068 3.274 0.112 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.342 0.403 2.41 0.447 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.126 0.178 2.194 0.222 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 1.046 0.33 1.114 0.374 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.508 0.358 0.572 0.402 ;
      RECT 0.29 0.203 0.358 0.247 ;
      RECT 0.29 0.3905 0.358 0.4345 ;
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 0.574 0.428 0.938 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.222 0.338 1.478 0.382 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.546 0.338 1.782 0.382 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 0.898 0.068 1.478 0.112 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 1.546 0.158 1.694 0.202 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.762 0.068 2.322 0.112 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.248 1.91 0.292 ;
      RECT 1.91 0.248 1.978 0.562 ;
      RECT 1.978 0.518 2.342 0.562 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.194 0.248 2.99 0.292 ;
      RECT 2.99 0.068 3.058 0.292 ;
      RECT 3.186 0.068 3.314 0.112 ;
      RECT 3.314 0.068 3.382 0.472 ;
  END
END b15fqn043hn1n04x5

MACRO b15fqn043hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn043hn1n06x5 0 0 ;
  SIZE 3.996 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.338 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.498 2.95 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.248 3.814 0.472 ;
      LAYER v0 ;
        RECT 3.746 0.338 3.814 0.382 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.338 3.598 0.382 ;
        RECT 3.53 0.158 3.598 0.382 ;
      LAYER v0 ;
        RECT 3.098 0.338 3.166 0.382 ;
        RECT 3.314 0.338 3.382 0.382 ;
        RECT 3.53 0.248 3.598 0.292 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.182 0.203 0.25 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.63916675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 3.274706 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.088 0.574 0.132 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.29 0.3905 0.358 0.4345 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.774 0.403 2.842 0.447 ;
        RECT 3.206 0.472 3.274 0.516 ;
        RECT 3.746 0.538 3.814 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.03 0.022 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 1.566 0.158 2.086 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.29 0.203 0.358 0.247 ;
        RECT 0.614 0.178 0.682 0.222 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 3.206 0.138 3.274 0.182 ;
        RECT 3.746 0.138 3.814 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.068 2.968 0.112 ;
      RECT 3.296 0.068 3.956 0.112 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.35 0.338 1.89 0.382 ;
      RECT 2.214 0.158 2.342 0.202 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 2.45 0.158 2.518 0.472 ;
      RECT 2.882 0.068 3.078 0.112 ;
      RECT 3.402 0.428 3.638 0.472 ;
      RECT 3.854 0.068 3.922 0.562 ;
    LAYER v1 ;
      RECT 3.858 0.068 3.918 0.112 ;
      RECT 3.318 0.068 3.378 0.112 ;
      RECT 2.886 0.068 2.946 0.112 ;
      RECT 0.834 0.068 0.894 0.112 ;
      RECT 0.402 0.068 0.462 0.112 ;
    LAYER v0 ;
      RECT 3.854 0.138 3.922 0.182 ;
      RECT 3.854 0.4185 3.922 0.4625 ;
      RECT 3.53 0.068 3.598 0.112 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 2.99 0.068 3.058 0.112 ;
      RECT 2.666 0.403 2.734 0.447 ;
      RECT 2.45 0.178 2.518 0.222 ;
      RECT 2.45 0.408 2.518 0.452 ;
      RECT 2.342 0.408 2.41 0.452 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.616 0.358 0.68 0.402 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.3905 0.466 0.4345 ;
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.472 ;
      RECT 0.682 0.428 1.046 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.006 0.068 1.89 0.112 ;
      RECT 2.342 0.158 2.41 0.472 ;
      RECT 1.222 0.158 1.37 0.202 ;
      RECT 1.37 0.158 1.438 0.292 ;
      RECT 1.438 0.248 2.234 0.292 ;
      RECT 2.234 0.248 2.302 0.562 ;
      RECT 2.302 0.518 2.666 0.562 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.518 0.248 3.314 0.292 ;
      RECT 3.314 0.068 3.382 0.292 ;
      RECT 3.51 0.068 3.638 0.112 ;
      RECT 3.638 0.068 3.706 0.472 ;
  END
END b15fqn043hn1n06x5

MACRO b15fqn043hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn043hn1n08x5 0 0 ;
  SIZE 4.212 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.862 0.518 3.058 0.562 ;
        RECT 2.99 0.338 3.058 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.518 2.95 0.562 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 1.06158725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.248 3.814 0.472 ;
      LAYER v0 ;
        RECT 3.746 0.338 3.814 0.382 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 1.95428575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.726 0.112 ;
        RECT 3.53 0.068 3.598 0.472 ;
        RECT 3.314 0.248 3.598 0.292 ;
        RECT 3.314 0.248 3.382 0.472 ;
      LAYER v0 ;
        RECT 3.314 0.338 3.382 0.382 ;
        RECT 3.53 0.338 3.598 0.382 ;
        RECT 3.638 0.068 3.706 0.112 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.1995 0.25 0.2435 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 4.001875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 3.2015 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.113 0.574 0.157 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.246 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.234 0.472 2.302 0.516 ;
        RECT 3.098 0.453 3.166 0.497 ;
        RECT 3.422 0.472 3.49 0.516 ;
        RECT 3.964 0.538 4.028 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.246 0.022 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 1.154 0.158 2.322 0.202 ;
        RECT 0.83 0.338 1.222 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
        RECT 0.83 -0.022 0.898 0.382 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.0975 0.142 0.1415 ;
        RECT 0.29 0.0975 0.358 0.1415 ;
        RECT 0.614 0.113 0.682 0.157 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.99 0.088 3.058 0.132 ;
        RECT 3.422 0.138 3.49 0.182 ;
        RECT 3.964 0.048 4.028 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.068 3.2 0.112 ;
      RECT 3.28 0.068 4.172 0.112 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 2.43 0.158 2.558 0.202 ;
      RECT 0.918 0.518 1.37 0.562 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 2.774 0.158 2.842 0.292 ;
      RECT 3.098 0.068 3.166 0.202 ;
      RECT 3.638 0.428 3.706 0.562 ;
      RECT 4.07 0.068 4.138 0.472 ;
    LAYER v1 ;
      RECT 4.074 0.068 4.134 0.112 ;
      RECT 3.318 0.068 3.378 0.112 ;
      RECT 3.102 0.068 3.162 0.112 ;
      RECT 0.726 0.068 0.786 0.112 ;
      RECT 0.402 0.068 0.462 0.112 ;
    LAYER v0 ;
      RECT 4.07 0.138 4.138 0.182 ;
      RECT 4.07 0.406 4.138 0.45 ;
      RECT 3.962 0.248 4.03 0.292 ;
      RECT 3.746 0.158 3.814 0.202 ;
      RECT 3.64 0.448 3.704 0.492 ;
      RECT 3.098 0.088 3.166 0.132 ;
      RECT 2.776 0.178 2.84 0.222 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.666 0.3155 2.734 0.3595 ;
      RECT 2.558 0.408 2.626 0.452 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.342 0.248 2.41 0.292 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.37 0.3605 1.438 0.4045 ;
      RECT 1.262 0.268 1.33 0.312 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.938 0.228 1.006 0.272 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.616 0.358 0.68 0.402 ;
      RECT 0.398 0.206 0.466 0.25 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.472 ;
      RECT 0.682 0.428 1.262 0.472 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.546 0.338 1.694 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.762 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.978 0.338 2.322 0.382 ;
      RECT 2.558 0.158 2.626 0.472 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.438 0.248 2.45 0.292 ;
      RECT 2.45 0.248 2.518 0.562 ;
      RECT 2.518 0.518 2.666 0.562 ;
      RECT 2.666 0.248 2.734 0.562 ;
      RECT 1.006 0.068 2.842 0.112 ;
      RECT 2.842 0.248 3.206 0.292 ;
      RECT 3.206 0.068 3.274 0.292 ;
      RECT 3.274 0.068 3.382 0.112 ;
      RECT 3.706 0.518 3.854 0.562 ;
      RECT 3.854 0.428 3.922 0.562 ;
      RECT 3.922 0.428 3.962 0.472 ;
      RECT 3.726 0.158 3.962 0.202 ;
      RECT 3.962 0.158 4.03 0.472 ;
  END
END b15fqn043hn1n08x5

MACRO b15fqn043hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn043hn1n12x5 0 0 ;
  SIZE 4.752 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0117 LAYER m2 ;
      ANTENNAMAXAREACAR 9.19365075 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0126 LAYER m2 ;
      ANTENNAMAXAREACAR 8.3505555 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.518 4.246 0.562 ;
        RECT 4.178 0.158 4.246 0.562 ;
        RECT 3.962 0.248 4.03 0.562 ;
        RECT 3.53 0.518 3.814 0.562 ;
        RECT 3.746 0.338 3.814 0.562 ;
      LAYER m2 ;
        RECT 3.728 0.428 4.156 0.472 ;
      LAYER v1 ;
        RECT 3.75 0.428 3.81 0.472 ;
        RECT 3.966 0.428 4.026 0.472 ;
      LAYER v0 ;
        RECT 3.638 0.518 3.706 0.562 ;
        RECT 3.962 0.293 4.03 0.337 ;
        RECT 4.178 0.248 4.246 0.292 ;
    END
  END den
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0207 LAYER m2 ;
      ANTENNAMAXAREACAR 2.82185175 LAYER m1 ;
      ANTENNAMAXAREACAR 4.418889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0279 LAYER m2 ;
      ANTENNAMAXAREACAR 2.82185175 LAYER m1 ;
      ANTENNAMAXAREACAR 4.418889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.428 2.43 0.472 ;
        RECT 0.594 0.428 0.79 0.472 ;
      LAYER m2 ;
        RECT 0.596 0.428 2.32 0.472 ;
      LAYER v1 ;
        RECT 0.618 0.428 0.678 0.472 ;
        RECT 2.238 0.428 2.298 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 2.342 0.428 2.41 0.472 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.158 3.49 0.382 ;
      LAYER v0 ;
        RECT 3.422 0.248 3.49 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.248 4.354 0.472 ;
      LAYER v0 ;
        RECT 4.286 0.338 4.354 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.562 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.1995 0.142 0.2435 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.29 0.1995 0.358 0.2435 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.786 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 4.394 0.518 4.462 0.652 ;
        RECT 3.854 0.338 3.922 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.83 0.338 0.898 0.472 ;
        RECT 0.398 0.338 0.898 0.382 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.832 0.408 0.896 0.452 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.666 0.538 2.734 0.582 ;
        RECT 3.422 0.538 3.49 0.582 ;
        RECT 3.854 0.4265 3.922 0.4705 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 4.61 0.453 4.678 0.497 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.786 0.022 ;
        RECT 4.61 -0.022 4.678 0.202 ;
        RECT 4.394 -0.022 4.462 0.112 ;
        RECT 3.854 -0.022 3.922 0.112 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 1.782 0.158 2.842 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.0975 0.25 0.1415 ;
        RECT 0.398 0.0975 0.466 0.1415 ;
        RECT 0.722 0.113 0.79 0.157 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.856 0.048 3.92 0.092 ;
        RECT 4.396 0.048 4.46 0.092 ;
        RECT 4.61 0.133 4.678 0.177 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 2.864 0.428 3.292 0.472 ;
      RECT 0.488 0.068 3.848 0.112 ;
      RECT 3.928 0.068 4.588 0.112 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.594 0.428 0.79 0.472 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 2.234 0.428 2.43 0.472 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 2.322 0.518 2.558 0.562 ;
      RECT 3.53 0.518 3.746 0.562 ;
      RECT 3.206 0.428 3.274 0.562 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 3.746 0.068 3.814 0.202 ;
      RECT 3.962 0.248 4.03 0.562 ;
      RECT 4.07 0.068 4.138 0.472 ;
      RECT 4.502 0.068 4.57 0.562 ;
    LAYER v1 ;
      RECT 4.506 0.068 4.566 0.112 ;
      RECT 3.966 0.068 4.026 0.112 ;
      RECT 3.75 0.068 3.81 0.112 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 0.942 0.068 1.002 0.112 ;
      RECT 0.51 0.068 0.57 0.112 ;
    LAYER v0 ;
      RECT 4.502 0.133 4.57 0.177 ;
      RECT 4.502 0.453 4.57 0.497 ;
      RECT 4.394 0.248 4.462 0.292 ;
      RECT 4.178 0.068 4.246 0.112 ;
      RECT 4.07 0.3985 4.138 0.4425 ;
      RECT 3.746 0.138 3.814 0.182 ;
      RECT 3.206 0.473 3.274 0.517 ;
      RECT 3.098 0.473 3.166 0.517 ;
      RECT 2.99 0.338 3.058 0.382 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.884 0.138 2.948 0.182 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.342 0.518 2.41 0.562 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.408 1.438 0.452 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 1.048 0.138 1.112 0.182 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.206 0.574 0.25 ;
    LAYER m1 ;
      RECT 0.702 0.518 1.046 0.562 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.248 1.262 0.292 ;
      RECT 1.262 0.158 1.33 0.472 ;
      RECT 1.33 0.158 1.458 0.202 ;
      RECT 1.114 0.068 2.538 0.112 ;
      RECT 1.222 0.518 1.478 0.562 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.546 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.338 2.754 0.382 ;
      RECT 1.438 0.248 2.882 0.292 ;
      RECT 2.882 0.248 2.95 0.472 ;
      RECT 2.558 0.428 2.626 0.562 ;
      RECT 2.626 0.428 2.774 0.472 ;
      RECT 2.774 0.428 2.842 0.562 ;
      RECT 2.882 0.068 2.95 0.202 ;
      RECT 2.842 0.518 2.99 0.562 ;
      RECT 2.99 0.248 3.058 0.562 ;
      RECT 3.058 0.248 3.098 0.292 ;
      RECT 2.95 0.068 3.098 0.112 ;
      RECT 3.098 0.068 3.166 0.292 ;
      RECT 3.746 0.338 3.814 0.562 ;
      RECT 3.166 0.338 3.314 0.382 ;
      RECT 3.314 0.338 3.382 0.472 ;
      RECT 3.382 0.428 3.638 0.472 ;
      RECT 3.638 0.248 3.706 0.472 ;
      RECT 3.706 0.248 3.854 0.292 ;
      RECT 3.854 0.158 3.922 0.292 ;
      RECT 3.922 0.158 3.962 0.202 ;
      RECT 3.962 0.068 4.03 0.202 ;
      RECT 4.03 0.518 4.178 0.562 ;
      RECT 4.178 0.158 4.246 0.562 ;
      RECT 4.138 0.068 4.286 0.112 ;
      RECT 4.286 0.068 4.354 0.202 ;
      RECT 4.354 0.158 4.394 0.202 ;
      RECT 4.394 0.158 4.462 0.382 ;
  END
END b15fqn043hn1n12x5

MACRO b15fqn043hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn043hn1n16x5 0 0 ;
  SIZE 5.832 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0297 LAYER m2 ;
      ANTENNAMAXAREACAR 4.05925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0342 LAYER m2 ;
      ANTENNAMAXAREACAR 4.05925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.042 0.248 5.11 0.472 ;
        RECT 4.07 0.338 4.138 0.472 ;
        RECT 3.51 0.338 4.138 0.382 ;
      LAYER m2 ;
        RECT 4.052 0.428 5.128 0.472 ;
      LAYER v1 ;
        RECT 4.074 0.428 4.134 0.472 ;
        RECT 5.046 0.428 5.106 0.472 ;
      LAYER v0 ;
        RECT 3.53 0.338 3.598 0.382 ;
        RECT 5.042 0.338 5.11 0.382 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.562 ;
      LAYER v0 ;
        RECT 1.802 0.448 1.87 0.492 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.262 0.068 1.33 0.472 ;
        RECT 0.81 0.068 1.33 0.112 ;
      LAYER v0 ;
        RECT 0.83 0.068 0.898 0.112 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.586 0.248 1.654 0.292 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.582 0.068 5.65 0.562 ;
        RECT 5.366 0.338 5.65 0.382 ;
        RECT 5.366 0.068 5.434 0.562 ;
      LAYER v0 ;
        RECT 5.366 0.448 5.434 0.492 ;
        RECT 5.366 0.158 5.434 0.202 ;
        RECT 5.582 0.448 5.65 0.492 ;
        RECT 5.582 0.158 5.65 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.866 0.652 ;
        RECT 5.69 0.428 5.758 0.652 ;
        RECT 5.474 0.428 5.542 0.652 ;
        RECT 5.258 0.428 5.326 0.652 ;
        RECT 4.826 0.338 4.894 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 3.206 0.518 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.4395 0.358 0.4835 ;
        RECT 0.506 0.4395 0.574 0.4835 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.99 0.457 3.058 0.501 ;
        RECT 3.208 0.538 3.272 0.582 ;
        RECT 3.424 0.538 3.488 0.582 ;
        RECT 3.746 0.457 3.814 0.501 ;
        RECT 3.962 0.448 4.03 0.492 ;
        RECT 4.826 0.4485 4.894 0.4925 ;
        RECT 5.258 0.448 5.326 0.492 ;
        RECT 5.474 0.448 5.542 0.492 ;
        RECT 5.69 0.448 5.758 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.866 0.022 ;
        RECT 5.69 -0.022 5.758 0.292 ;
        RECT 5.474 -0.022 5.542 0.292 ;
        RECT 5.258 -0.022 5.326 0.292 ;
        RECT 4.934 -0.022 5.002 0.292 ;
        RECT 2.774 0.158 3.51 0.202 ;
        RECT 2.126 0.248 2.842 0.292 ;
        RECT 2.774 0.158 2.842 0.292 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.206 0.158 3.274 0.202 ;
        RECT 3.422 0.158 3.49 0.202 ;
        RECT 4.934 0.158 5.002 0.202 ;
        RECT 5.258 0.158 5.326 0.202 ;
        RECT 5.474 0.158 5.542 0.202 ;
        RECT 5.69 0.158 5.758 0.202 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.518 0.7 0.562 ;
      RECT 0.164 0.068 0.7 0.112 ;
      RECT 1.028 0.518 1.904 0.562 ;
      RECT 0.38 0.428 2.66 0.472 ;
      RECT 2.74 0.428 3.616 0.472 ;
      RECT 1.984 0.518 4.264 0.562 ;
      RECT 4.592 0.518 5.02 0.562 ;
      RECT 1.46 0.068 5.236 0.112 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.182 0.068 0.25 0.202 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.614 0.338 1.046 0.382 ;
      RECT 0.506 0.248 1.154 0.292 ;
      RECT 2.43 0.338 2.774 0.382 ;
      RECT 1.478 0.068 1.546 0.382 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 2.018 0.068 2.086 0.562 ;
      RECT 2.558 0.428 2.626 0.562 ;
      RECT 3.51 0.338 4.07 0.382 ;
      RECT 2.882 0.248 2.95 0.562 ;
      RECT 3.422 0.428 3.618 0.472 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 4.178 0.338 4.246 0.562 ;
      RECT 4.394 0.428 4.462 0.562 ;
      RECT 2.342 0.068 2.41 0.202 ;
      RECT 4.934 0.338 5.002 0.562 ;
      RECT 5.042 0.248 5.11 0.472 ;
      RECT 5.15 0.068 5.218 0.562 ;
    LAYER v1 ;
      RECT 5.154 0.068 5.214 0.112 ;
      RECT 4.938 0.518 4.998 0.562 ;
      RECT 4.614 0.518 4.674 0.562 ;
      RECT 4.182 0.518 4.242 0.562 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 2.886 0.518 2.946 0.562 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.022 0.518 2.082 0.562 ;
      RECT 1.698 0.518 1.758 0.562 ;
      RECT 1.482 0.068 1.542 0.112 ;
      RECT 1.05 0.518 1.11 0.562 ;
      RECT 0.618 0.068 0.678 0.112 ;
      RECT 0.618 0.518 0.678 0.562 ;
      RECT 0.402 0.428 0.462 0.472 ;
      RECT 0.186 0.068 0.246 0.112 ;
      RECT 0.186 0.518 0.246 0.562 ;
    LAYER v0 ;
      RECT 5.15 0.158 5.218 0.202 ;
      RECT 5.15 0.448 5.218 0.492 ;
      RECT 4.934 0.4485 5.002 0.4925 ;
      RECT 4.718 0.338 4.786 0.382 ;
      RECT 4.612 0.448 4.676 0.492 ;
      RECT 4.502 0.158 4.57 0.202 ;
      RECT 4.502 0.3685 4.57 0.4125 ;
      RECT 4.396 0.448 4.46 0.492 ;
      RECT 4.286 0.248 4.354 0.292 ;
      RECT 4.178 0.068 4.246 0.112 ;
      RECT 4.178 0.158 4.246 0.202 ;
      RECT 4.178 0.3685 4.246 0.4125 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 3.854 0.248 3.922 0.292 ;
      RECT 3.638 0.248 3.706 0.292 ;
      RECT 3.53 0.428 3.598 0.472 ;
      RECT 3.314 0.457 3.382 0.501 ;
      RECT 3.098 0.457 3.166 0.501 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.558 0.448 2.626 0.492 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.344 0.138 2.408 0.182 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.694 0.138 1.762 0.182 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.154 0.4855 1.222 0.5295 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.832 0.448 0.896 0.492 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.398 0.4395 0.466 0.4835 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.4395 0.25 0.4835 ;
    LAYER m1 ;
      RECT 0.614 0.518 0.83 0.562 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.682 0.158 0.918 0.202 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 2.774 0.338 2.842 0.472 ;
      RECT 4.07 0.338 4.138 0.472 ;
      RECT 3.166 0.338 3.314 0.382 ;
      RECT 3.314 0.248 3.382 0.562 ;
      RECT 3.382 0.248 4.502 0.292 ;
      RECT 4.502 0.248 4.57 0.472 ;
      RECT 4.462 0.518 4.61 0.562 ;
      RECT 4.158 0.158 4.61 0.202 ;
      RECT 4.61 0.158 4.678 0.562 ;
      RECT 2.41 0.068 4.718 0.112 ;
      RECT 4.718 0.068 4.786 0.562 ;
  END
END b15fqn043hn1n16x5

MACRO b15fqn08fhn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn08fhn1n02x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 5.32 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 5.32 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.518 0.292 ;
      LAYER v0 ;
        RECT 2.45 0.228 2.518 0.272 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.248 3.166 0.472 ;
      LAYER v0 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.4 0.142 0.444 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.15375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.15375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.398 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.496 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.566 0.202 ;
        RECT 1.046 0.068 1.114 0.202 ;
        RECT 0.83 0.068 1.114 0.112 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.383 0.466 0.427 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.234 0.358 2.302 0.402 ;
        RECT 2.558 0.473 2.626 0.517 ;
        RECT 3.1 0.538 3.164 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.782 0.158 2.41 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 3.098 0.138 3.166 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.428 1.148 0.472 ;
      RECT 1.228 0.428 2.968 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 1.046 0.338 1.262 0.382 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.91 0.338 2.126 0.382 ;
      RECT 1.674 0.248 1.998 0.292 ;
      RECT 2.126 0.428 2.194 0.562 ;
      RECT 1.242 0.068 2.214 0.112 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.206 0.068 3.274 0.562 ;
    LAYER v1 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 2.67 0.428 2.73 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.186 0.428 0.246 0.472 ;
    LAYER v0 ;
      RECT 3.206 0.138 3.274 0.182 ;
      RECT 3.206 0.453 3.274 0.497 ;
      RECT 2.99 0.138 3.058 0.182 ;
      RECT 2.99 0.4575 3.058 0.5015 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.882 0.358 2.95 0.402 ;
      RECT 2.774 0.472 2.842 0.516 ;
      RECT 2.666 0.383 2.734 0.427 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.182 0.293 0.25 0.337 ;
    LAYER m1 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.358 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.574 0.338 0.938 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.114 0.518 1.37 0.562 ;
      RECT 1.242 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 1.998 0.562 ;
      RECT 2.126 0.248 2.194 0.382 ;
      RECT 2.194 0.248 2.342 0.292 ;
      RECT 2.342 0.248 2.41 0.382 ;
      RECT 2.41 0.338 2.558 0.382 ;
      RECT 2.558 0.248 2.626 0.382 ;
      RECT 2.626 0.248 2.774 0.292 ;
      RECT 2.774 0.248 2.842 0.562 ;
      RECT 2.842 0.248 2.882 0.292 ;
      RECT 2.882 0.068 2.95 0.292 ;
  END
END b15fqn08fhn1n02x5

MACRO b15fqn08fhn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn08fhn1n04x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 5.32 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 5.32 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.518 0.292 ;
      LAYER v0 ;
        RECT 2.45 0.228 2.518 0.272 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.248 3.166 0.472 ;
      LAYER v0 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.4 0.142 0.444 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 4.123 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 4.123 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.398 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 2.49714275 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.566 0.202 ;
        RECT 1.046 0.068 1.114 0.202 ;
        RECT 0.83 0.068 1.114 0.112 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.383 0.466 0.427 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.234 0.358 2.302 0.402 ;
        RECT 2.558 0.473 2.626 0.517 ;
        RECT 3.1 0.538 3.164 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.782 0.158 2.41 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 3.098 0.138 3.166 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.428 1.148 0.472 ;
      RECT 1.228 0.428 2.984 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 1.046 0.338 1.262 0.382 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.91 0.338 2.126 0.382 ;
      RECT 1.674 0.248 1.998 0.292 ;
      RECT 2.126 0.428 2.194 0.562 ;
      RECT 1.242 0.068 2.214 0.112 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.206 0.068 3.274 0.562 ;
    LAYER v1 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 2.67 0.428 2.73 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.186 0.428 0.246 0.472 ;
    LAYER v0 ;
      RECT 3.206 0.138 3.274 0.182 ;
      RECT 3.206 0.4575 3.274 0.5015 ;
      RECT 2.99 0.138 3.058 0.182 ;
      RECT 2.99 0.4575 3.058 0.5015 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.882 0.358 2.95 0.402 ;
      RECT 2.774 0.472 2.842 0.516 ;
      RECT 2.666 0.383 2.734 0.427 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.182 0.293 0.25 0.337 ;
    LAYER m1 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.358 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.574 0.338 0.938 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.114 0.518 1.37 0.562 ;
      RECT 1.242 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 1.998 0.562 ;
      RECT 2.126 0.248 2.194 0.382 ;
      RECT 2.194 0.248 2.342 0.292 ;
      RECT 2.342 0.248 2.41 0.382 ;
      RECT 2.41 0.338 2.558 0.382 ;
      RECT 2.558 0.248 2.626 0.382 ;
      RECT 2.626 0.248 2.774 0.292 ;
      RECT 2.774 0.248 2.842 0.562 ;
      RECT 2.842 0.248 2.882 0.292 ;
      RECT 2.882 0.068 2.95 0.292 ;
  END
END b15fqn08fhn1n04x5

MACRO b15fqn08fhn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn08fhn1n08x5 0 0 ;
  SIZE 4.32 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.158 3.274 0.382 ;
        RECT 2.99 0.248 3.274 0.292 ;
      LAYER v0 ;
        RECT 3.098 0.248 3.166 0.292 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.248 4.138 0.472 ;
      LAYER v0 ;
        RECT 4.07 0.338 4.138 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.4 0.25 0.444 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 4.123 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 4.123 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.614 0.068 0.682 0.112 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.59916675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 1.199375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 2.214 0.112 ;
        RECT 0.938 0.068 1.006 0.292 ;
      LAYER v0 ;
        RECT 1.046 0.068 1.114 0.112 ;
        RECT 2.126 0.068 2.194 0.112 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.354 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.493 0.142 0.537 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.383 0.574 0.427 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 4.072 0.538 4.136 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.354 0.022 ;
        RECT 4.07 -0.022 4.138 0.202 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.99 0.048 3.058 0.092 ;
        RECT 3.422 0.138 3.49 0.182 ;
        RECT 4.07 0.138 4.138 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.428 1.24 0.472 ;
      RECT 1.784 0.428 2.66 0.472 ;
      RECT 2.74 0.428 3.848 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 2.558 0.428 2.626 0.562 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 1.89 0.158 2.754 0.202 ;
      RECT 1.458 0.338 3.098 0.382 ;
      RECT 2.666 0.428 2.862 0.472 ;
      RECT 3.638 0.338 3.706 0.562 ;
      RECT 1.262 0.248 2.882 0.292 ;
      RECT 3.962 0.158 4.03 0.562 ;
      RECT 4.178 0.068 4.246 0.562 ;
    LAYER v1 ;
      RECT 3.642 0.428 3.702 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.158 0.428 1.218 0.472 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.294 0.428 0.354 0.472 ;
    LAYER v0 ;
      RECT 4.178 0.138 4.246 0.182 ;
      RECT 4.178 0.4285 4.246 0.4725 ;
      RECT 3.962 0.2185 4.03 0.2625 ;
      RECT 3.962 0.4575 4.03 0.5015 ;
      RECT 3.854 0.338 3.922 0.382 ;
      RECT 3.746 0.178 3.814 0.222 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.53 0.338 3.598 0.382 ;
      RECT 3.314 0.333 3.382 0.377 ;
      RECT 3.098 0.448 3.166 0.492 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.774 0.518 2.842 0.562 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.56 0.448 2.624 0.492 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.588 0.448 1.652 0.492 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.614 0.498 0.682 0.542 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.29 0.293 0.358 0.337 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.158 0.574 0.292 ;
      RECT 0.574 0.248 0.614 0.292 ;
      RECT 0.614 0.248 0.682 0.382 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.158 1.114 0.382 ;
      RECT 1.222 0.158 1.458 0.202 ;
      RECT 1.222 0.518 1.586 0.562 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 2.626 0.518 2.862 0.562 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 3.706 0.338 3.746 0.382 ;
      RECT 3.746 0.158 3.814 0.382 ;
      RECT 2.882 0.158 2.95 0.292 ;
      RECT 2.95 0.158 3.098 0.202 ;
      RECT 3.098 0.068 3.166 0.202 ;
      RECT 3.166 0.068 3.314 0.112 ;
      RECT 3.314 0.068 3.382 0.472 ;
      RECT 3.382 0.248 3.53 0.292 ;
      RECT 3.53 0.068 3.598 0.472 ;
      RECT 3.598 0.068 3.854 0.112 ;
      RECT 3.854 0.068 3.922 0.472 ;
  END
END b15fqn08fhn1n08x5

MACRO b15fqn08fhn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqn08fhn1n16x5 0 0 ;
  SIZE 5.94 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.158 4.462 0.382 ;
        RECT 4.158 0.248 4.462 0.292 ;
      LAYER v0 ;
        RECT 4.178 0.248 4.246 0.292 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.366 0.248 5.434 0.562 ;
      LAYER v0 ;
        RECT 5.366 0.49 5.434 0.534 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.408 0.466 0.452 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0135 LAYER m1 ;
      ANTENNAMAXAREACAR 5.4014285 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0135 LAYER m1 ;
      ANTENNAMAXAREACAR 2.52066675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.3155 0.898 0.3595 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.027 LAYER m1 ;
      ANTENNAMAXAREACAR 3.04 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0342 LAYER m1 ;
      ANTENNAMAXAREACAR 3.04 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 2.322 0.112 ;
        RECT 1.37 0.068 1.438 0.292 ;
      LAYER v0 ;
        RECT 1.478 0.068 1.546 0.112 ;
        RECT 2.234 0.068 2.302 0.112 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.974 0.652 ;
        RECT 5.798 0.518 5.866 0.652 ;
        RECT 5.582 0.428 5.65 0.652 ;
        RECT 4.718 0.428 4.786 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.493 0.358 0.537 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 4.178 0.448 4.246 0.492 ;
        RECT 4.718 0.456 4.786 0.5 ;
        RECT 5.582 0.456 5.65 0.5 ;
        RECT 5.798 0.538 5.866 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.974 0.022 ;
        RECT 5.798 -0.022 5.866 0.202 ;
        RECT 5.582 -0.022 5.65 0.202 ;
        RECT 4.61 -0.022 4.678 0.292 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.316 0.048 3.38 0.092 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.748 0.048 3.812 0.092 ;
        RECT 4.18 0.048 4.244 0.092 ;
        RECT 4.61 0.1715 4.678 0.2155 ;
        RECT 5.582 0.13 5.65 0.174 ;
        RECT 5.798 0.13 5.866 0.174 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.428 1.564 0.472 ;
      RECT 2.216 0.428 3.848 0.472 ;
      RECT 3.928 0.428 5.36 0.472 ;
      RECT 5.44 0.428 5.9 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.472 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 1.046 0.338 1.114 0.472 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 3.746 0.428 3.814 0.562 ;
      RECT 1.89 0.428 2.322 0.472 ;
      RECT 2.558 0.428 2.626 0.562 ;
      RECT 2.774 0.428 2.842 0.562 ;
      RECT 3.53 0.428 3.598 0.562 ;
      RECT 2.43 0.158 3.854 0.202 ;
      RECT 3.854 0.428 4.05 0.472 ;
      RECT 1.586 0.338 1.654 0.472 ;
      RECT 4.826 0.428 4.934 0.472 ;
      RECT 1.674 0.248 3.962 0.292 ;
      RECT 5.042 0.428 5.11 0.562 ;
      RECT 5.15 0.068 5.218 0.562 ;
      RECT 5.258 0.158 5.326 0.562 ;
      RECT 5.474 0.338 5.542 0.472 ;
      RECT 5.798 0.248 5.866 0.472 ;
    LAYER v1 ;
      RECT 5.802 0.428 5.862 0.472 ;
      RECT 5.478 0.428 5.538 0.472 ;
      RECT 5.262 0.428 5.322 0.472 ;
      RECT 5.046 0.428 5.106 0.472 ;
      RECT 4.83 0.428 4.89 0.472 ;
      RECT 3.966 0.428 4.026 0.472 ;
      RECT 3.75 0.428 3.81 0.472 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.726 0.428 0.786 0.472 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.078 0.428 0.138 0.472 ;
    LAYER v0 ;
      RECT 5.798 0.293 5.866 0.337 ;
      RECT 5.69 0.13 5.758 0.174 ;
      RECT 5.69 0.456 5.758 0.5 ;
      RECT 5.474 0.363 5.542 0.407 ;
      RECT 5.258 0.192 5.326 0.236 ;
      RECT 5.258 0.49 5.326 0.534 ;
      RECT 5.15 0.192 5.218 0.236 ;
      RECT 5.15 0.49 5.218 0.534 ;
      RECT 5.042 0.293 5.11 0.337 ;
      RECT 5.042 0.49 5.11 0.534 ;
      RECT 4.934 0.192 5.002 0.236 ;
      RECT 4.502 0.1715 4.57 0.2155 ;
      RECT 4.502 0.448 4.57 0.492 ;
      RECT 4.286 0.448 4.354 0.492 ;
      RECT 3.962 0.068 4.03 0.112 ;
      RECT 3.962 0.428 4.03 0.472 ;
      RECT 3.962 0.518 4.03 0.562 ;
      RECT 3.748 0.448 3.812 0.492 ;
      RECT 3.638 0.158 3.706 0.202 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.774 0.448 2.842 0.492 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.558 0.448 2.626 0.492 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.588 0.408 1.652 0.452 ;
      RECT 1.478 0.325 1.546 0.369 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.3685 1.114 0.4125 ;
      RECT 0.938 0.186 1.006 0.23 ;
      RECT 0.94 0.448 1.004 0.492 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.3155 0.79 0.3595 ;
      RECT 0.614 0.453 0.682 0.497 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.222 0.338 1.438 0.382 ;
      RECT 1.546 0.158 2.106 0.202 ;
      RECT 1.006 0.518 1.154 0.562 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.222 0.428 1.37 0.472 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.438 0.518 2.322 0.562 ;
      RECT 3.814 0.518 4.05 0.562 ;
      RECT 3.854 0.068 3.922 0.202 ;
      RECT 3.922 0.068 4.05 0.112 ;
      RECT 1.654 0.338 4.286 0.382 ;
      RECT 4.286 0.338 4.354 0.562 ;
      RECT 4.934 0.158 5.002 0.472 ;
      RECT 3.962 0.158 4.03 0.292 ;
      RECT 4.03 0.158 4.286 0.202 ;
      RECT 4.286 0.068 4.354 0.202 ;
      RECT 4.354 0.068 4.502 0.112 ;
      RECT 4.502 0.068 4.57 0.562 ;
      RECT 4.57 0.338 4.826 0.382 ;
      RECT 4.826 0.068 4.894 0.382 ;
      RECT 4.894 0.068 5.042 0.112 ;
      RECT 5.042 0.068 5.11 0.382 ;
      RECT 5.218 0.068 5.474 0.112 ;
      RECT 5.474 0.068 5.542 0.292 ;
      RECT 5.542 0.248 5.69 0.292 ;
      RECT 5.69 0.068 5.758 0.562 ;
  END
END b15fqn08fhn1n16x5

MACRO b15fqy003hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy003hn1n02x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.428 1.222 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
      LAYER m2 ;
        RECT 0.38 0.518 1.24 0.562 ;
      LAYER v1 ;
        RECT 0.402 0.518 0.462 0.562 ;
        RECT 1.158 0.518 1.218 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.498 0.466 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.498 2.086 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.382 ;
      LAYER v0 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.403 0.25 0.447 ;
        RECT 0.182 0.1915 0.25 0.2355 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.472 ;
      LAYER v0 ;
        RECT 2.666 0.293 2.734 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.76277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.5255555 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
        RECT 2.342 0.068 2.626 0.112 ;
      LAYER v0 ;
        RECT 2.45 0.068 2.518 0.112 ;
        RECT 2.558 0.498 2.626 0.542 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 1.046 0.338 1.114 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.506 0.403 0.574 0.447 ;
        RECT 1.046 0.402 1.114 0.446 ;
        RECT 1.37 0.403 1.438 0.447 ;
        RECT 1.802 0.47 1.87 0.514 ;
        RECT 2.234 0.393 2.302 0.437 ;
        RECT 2.774 0.403 2.842 0.447 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.234 -0.022 2.302 0.292 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.046 0.158 1.33 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.398 0.088 0.466 0.132 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.774 0.1945 2.842 0.2385 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 0.824 0.382 ;
      RECT 0.904 0.338 1.688 0.382 ;
      RECT 0.812 0.428 1.996 0.472 ;
      RECT 1.568 0.518 2.228 0.562 ;
      RECT 1.768 0.338 2.552 0.382 ;
      RECT 2.308 0.518 2.984 0.562 ;
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.382 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.83 0.248 1.262 0.292 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.37 0.158 1.586 0.202 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.91 0.068 1.978 0.472 ;
      RECT 1.478 0.518 1.762 0.562 ;
      RECT 1.694 0.068 1.762 0.472 ;
      RECT 1.802 0.248 1.87 0.382 ;
      RECT 2.126 0.428 2.194 0.562 ;
      RECT 2.342 0.428 2.41 0.562 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.882 0.158 2.95 0.562 ;
    LAYER v1 ;
      RECT 2.886 0.518 2.946 0.562 ;
      RECT 2.454 0.338 2.514 0.382 ;
      RECT 2.346 0.518 2.406 0.562 ;
      RECT 2.13 0.518 2.19 0.562 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.806 0.338 1.866 0.382 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 2.882 0.1945 2.95 0.2385 ;
      RECT 2.882 0.403 2.95 0.447 ;
      RECT 2.45 0.403 2.518 0.447 ;
      RECT 2.342 0.498 2.41 0.542 ;
      RECT 2.126 0.293 2.194 0.337 ;
      RECT 2.126 0.498 2.194 0.542 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.694 0.138 1.762 0.182 ;
      RECT 1.694 0.3835 1.762 0.4275 ;
      RECT 1.586 0.3835 1.654 0.4275 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.403 1.33 0.447 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.498 0.898 0.542 ;
      RECT 0.722 0.376 0.79 0.42 ;
      RECT 0.614 0.498 0.682 0.542 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.79 0.158 1.006 0.202 ;
      RECT 0.682 0.068 1.006 0.112 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.978 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.382 ;
  END
END b15fqy003hn1n02x5

MACRO b15fqy003hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy003hn1n03x5 0 0 ;
  SIZE 3.132 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 4.948889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 4.948889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.428 1.33 0.562 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.518 1.348 0.562 ;
      LAYER v1 ;
        RECT 0.51 0.518 0.57 0.562 ;
        RECT 1.266 0.518 1.326 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 1.262 0.498 1.33 0.542 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.158 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.498 2.194 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.158 2.518 0.382 ;
      LAYER v0 ;
        RECT 2.45 0.293 2.518 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.403 0.142 0.447 ;
        RECT 0.074 0.183 0.142 0.227 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.068 2.842 0.472 ;
      LAYER v0 ;
        RECT 2.774 0.293 2.842 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.76277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.5255555 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.562 ;
        RECT 2.45 0.068 2.734 0.112 ;
      LAYER v0 ;
        RECT 2.558 0.068 2.626 0.112 ;
        RECT 2.666 0.498 2.734 0.542 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.166 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.614 0.338 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.403 0.25 0.447 ;
        RECT 0.614 0.383 0.682 0.427 ;
        RECT 1.154 0.383 1.222 0.427 ;
        RECT 1.478 0.403 1.546 0.447 ;
        RECT 1.91 0.47 1.978 0.514 ;
        RECT 2.342 0.393 2.41 0.437 ;
        RECT 2.882 0.403 2.95 0.447 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.166 0.022 ;
        RECT 2.882 -0.022 2.95 0.292 ;
        RECT 2.342 -0.022 2.41 0.292 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.183 0.25 0.227 ;
        RECT 0.506 0.203 0.574 0.247 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.91 0.138 1.978 0.182 ;
        RECT 2.342 0.1695 2.41 0.2135 ;
        RECT 2.882 0.1955 2.95 0.2395 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 0.932 0.382 ;
      RECT 1.012 0.338 1.796 0.382 ;
      RECT 0.92 0.428 2.104 0.472 ;
      RECT 1.676 0.518 2.336 0.562 ;
      RECT 1.876 0.338 2.66 0.382 ;
      RECT 2.416 0.518 3.092 0.562 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 0.938 0.248 1.37 0.292 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.478 0.158 1.694 0.202 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 2.018 0.068 2.086 0.472 ;
      RECT 1.586 0.518 1.87 0.562 ;
      RECT 1.802 0.068 1.87 0.472 ;
      RECT 1.91 0.248 1.978 0.382 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.45 0.428 2.518 0.562 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 2.99 0.158 3.058 0.562 ;
    LAYER v1 ;
      RECT 2.994 0.518 3.054 0.562 ;
      RECT 2.562 0.338 2.622 0.382 ;
      RECT 2.454 0.518 2.514 0.562 ;
      RECT 2.238 0.518 2.298 0.562 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.698 0.518 1.758 0.562 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.402 0.338 0.462 0.382 ;
    LAYER v0 ;
      RECT 2.99 0.1955 3.058 0.2395 ;
      RECT 2.99 0.403 3.058 0.447 ;
      RECT 2.558 0.403 2.626 0.447 ;
      RECT 2.45 0.498 2.518 0.542 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.234 0.498 2.302 0.542 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.138 1.87 0.182 ;
      RECT 1.802 0.3835 1.87 0.4275 ;
      RECT 1.694 0.3835 1.762 0.4275 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.37 0.403 1.438 0.447 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.498 1.114 0.542 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.398 0.403 0.466 0.447 ;
      RECT 0.29 0.183 0.358 0.227 ;
      RECT 0.29 0.403 0.358 0.447 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.79 0.068 1.006 0.112 ;
      RECT 0.898 0.158 1.114 0.202 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 2.086 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.382 ;
  END
END b15fqy003hn1n03x5

MACRO b15fqy003hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy003hn1n04x5 0 0 ;
  SIZE 3.24 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 6.748611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 6.748611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.438 0.382 ;
        RECT 1.154 0.338 1.222 0.562 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.518 1.24 0.562 ;
      LAYER v1 ;
        RECT 0.51 0.518 0.57 0.562 ;
        RECT 1.158 0.518 1.218 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.158 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.498 2.302 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.158 2.626 0.382 ;
      LAYER v0 ;
        RECT 2.558 0.293 2.626 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.403 0.142 0.447 ;
        RECT 0.074 0.178 0.142 0.222 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.472 ;
      LAYER v0 ;
        RECT 2.882 0.293 2.95 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.76277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.5255555 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.068 2.842 0.562 ;
        RECT 2.558 0.068 2.842 0.112 ;
      LAYER v0 ;
        RECT 2.666 0.068 2.734 0.112 ;
        RECT 2.774 0.498 2.842 0.542 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.274 0.652 ;
        RECT 2.99 0.338 3.058 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.586 0.338 1.654 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.338 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.403 0.25 0.447 ;
        RECT 0.614 0.363 0.682 0.407 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.586 0.403 1.654 0.447 ;
        RECT 2.018 0.47 2.086 0.514 ;
        RECT 2.45 0.393 2.518 0.437 ;
        RECT 2.99 0.403 3.058 0.447 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.274 0.022 ;
        RECT 2.99 -0.022 3.058 0.292 ;
        RECT 2.45 -0.022 2.518 0.292 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.178 0.25 0.222 ;
        RECT 0.506 0.222 0.574 0.266 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.99 0.1955 3.058 0.2395 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 0.932 0.382 ;
      RECT 1.012 0.338 1.904 0.382 ;
      RECT 0.92 0.428 2.212 0.472 ;
      RECT 1.784 0.518 2.444 0.562 ;
      RECT 1.984 0.338 2.768 0.382 ;
      RECT 2.524 0.518 3.2 0.562 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.046 0.248 1.478 0.292 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.586 0.158 1.802 0.202 ;
      RECT 2.126 0.068 2.194 0.472 ;
      RECT 1.694 0.518 1.978 0.562 ;
      RECT 1.91 0.068 1.978 0.472 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 2.342 0.428 2.41 0.562 ;
      RECT 2.558 0.428 2.626 0.562 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 3.098 0.158 3.166 0.562 ;
    LAYER v1 ;
      RECT 3.102 0.518 3.162 0.562 ;
      RECT 2.67 0.338 2.73 0.382 ;
      RECT 2.562 0.518 2.622 0.562 ;
      RECT 2.346 0.518 2.406 0.562 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.806 0.338 1.866 0.382 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.402 0.338 0.462 0.382 ;
    LAYER v0 ;
      RECT 3.098 0.1955 3.166 0.2395 ;
      RECT 3.098 0.403 3.166 0.447 ;
      RECT 2.666 0.403 2.734 0.447 ;
      RECT 2.558 0.498 2.626 0.542 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.342 0.498 2.41 0.542 ;
      RECT 2.126 0.293 2.194 0.337 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.3835 1.978 0.4275 ;
      RECT 1.802 0.3835 1.87 0.4275 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.478 0.403 1.546 0.447 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.395 0.898 0.439 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.398 0.403 0.466 0.447 ;
      RECT 0.29 0.178 0.358 0.222 ;
      RECT 0.29 0.403 0.358 0.447 ;
    LAYER m1 ;
      RECT 0.83 0.518 1.046 0.562 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 0.898 0.158 1.114 0.202 ;
      RECT 1.222 0.338 1.438 0.382 ;
      RECT 1.478 0.248 1.546 0.562 ;
      RECT 0.79 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 1.546 0.068 1.762 0.112 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 2.194 0.068 2.342 0.112 ;
      RECT 2.342 0.068 2.41 0.382 ;
  END
END b15fqy003hn1n04x5

MACRO b15fqy003hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy003hn1n06x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    ANTENNADIFFAREA 0.03672 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.428 0.484 0.472 ;
      LAYER v1 ;
        RECT 0.078 0.428 0.138 0.472 ;
        RECT 0.294 0.428 0.354 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.074 0.179 0.142 0.223 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAGATEAREA 0.0117 LAYER m2 ;
      ANTENNAMAXAREACAR 0.3144445 LAYER m1 ;
      ANTENNAMAXAREACAR 4.950889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.2515555 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.3930555 LAYER m1 ;
      ANTENNAMAXAREACAR 6.188611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.338 1.654 0.562 ;
        RECT 1.458 0.338 1.654 0.382 ;
        RECT 0.398 0.428 0.466 0.562 ;
      LAYER m2 ;
        RECT 0.38 0.518 1.672 0.562 ;
      LAYER v1 ;
        RECT 0.402 0.518 0.462 0.562 ;
        RECT 1.59 0.518 1.65 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.498 0.466 0.542 ;
        RECT 1.478 0.338 1.546 0.382 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.248 2.41 0.382 ;
      LAYER v0 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.158 2.842 0.382 ;
      LAYER v0 ;
        RECT 2.774 0.293 2.842 0.337 ;
    END
  END d
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.068 3.166 0.472 ;
      LAYER v0 ;
        RECT 3.098 0.293 3.166 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.76277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.5255555 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.068 3.058 0.562 ;
        RECT 2.774 0.068 3.058 0.112 ;
      LAYER v0 ;
        RECT 2.882 0.068 2.95 0.112 ;
        RECT 2.99 0.498 3.058 0.542 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.206 0.338 3.274 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.498 0.25 0.542 ;
        RECT 0.614 0.467 0.682 0.511 ;
        RECT 1.262 0.503 1.33 0.547 ;
        RECT 1.802 0.403 1.87 0.447 ;
        RECT 2.234 0.4055 2.302 0.4495 ;
        RECT 2.666 0.393 2.734 0.437 ;
        RECT 3.206 0.403 3.274 0.447 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.206 -0.022 3.274 0.292 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.088 0.25 0.132 ;
        RECT 0.506 0.088 0.574 0.132 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 3.206 0.184 3.274 0.228 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.338 0.916 0.382 ;
      RECT 1.244 0.338 2.104 0.382 ;
      RECT 0.812 0.428 2.66 0.472 ;
      RECT 2.432 0.518 2.968 0.562 ;
      RECT 2.74 0.428 3.416 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.182 0.248 0.25 0.382 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.398 0.338 0.682 0.382 ;
      RECT 0.83 0.158 0.898 0.562 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.458 0.338 1.586 0.382 ;
      RECT 1.154 0.338 1.35 0.382 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.802 0.158 2.018 0.202 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 2.45 0.248 2.518 0.472 ;
      RECT 2.342 0.518 2.538 0.562 ;
      RECT 2.774 0.428 2.842 0.562 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 3.314 0.338 3.382 0.472 ;
    LAYER v1 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 2.886 0.518 2.946 0.562 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.454 0.428 2.514 0.472 ;
      RECT 2.454 0.518 2.514 0.562 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
      RECT 0.186 0.338 0.246 0.382 ;
    LAYER v0 ;
      RECT 3.314 0.403 3.382 0.447 ;
      RECT 2.882 0.403 2.95 0.447 ;
      RECT 2.774 0.498 2.842 0.542 ;
      RECT 2.558 0.293 2.626 0.337 ;
      RECT 2.45 0.293 2.518 0.337 ;
      RECT 2.45 0.518 2.518 0.562 ;
      RECT 2.018 0.3835 2.086 0.4275 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.694 0.403 1.762 0.447 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 1.046 0.467 1.114 0.511 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.467 0.898 0.511 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.088 0.682 0.132 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.182 0.293 0.25 0.337 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.898 0.158 1.114 0.202 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.114 0.248 1.694 0.292 ;
      RECT 1.694 0.248 1.762 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 0.79 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.438 0.158 1.694 0.202 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.91 0.518 2.126 0.562 ;
      RECT 1.762 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.562 ;
      RECT 2.194 0.158 2.558 0.202 ;
      RECT 2.558 0.158 2.626 0.382 ;
  END
END b15fqy003hn1n06x5

MACRO b15fqy003hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy003hn1n08x5 0 0 ;
  SIZE 3.888 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 7.788889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 7.788889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.338 1.762 0.382 ;
        RECT 1.37 0.518 1.546 0.562 ;
        RECT 1.478 0.338 1.546 0.562 ;
        RECT 0.506 0.248 0.574 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.518 1.472 0.562 ;
      LAYER v1 ;
        RECT 0.51 0.518 0.57 0.562 ;
        RECT 1.374 0.518 1.434 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.248 2.734 0.472 ;
      LAYER v0 ;
        RECT 2.666 0.338 2.734 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.248 3.274 0.292 ;
        RECT 3.206 0.158 3.274 0.292 ;
      LAYER v0 ;
        RECT 3.098 0.248 3.166 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.598 0.472 ;
      LAYER v0 ;
        RECT 3.53 0.293 3.598 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.76277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.5255555 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.068 3.49 0.562 ;
        RECT 3.206 0.068 3.49 0.112 ;
      LAYER v0 ;
        RECT 3.314 0.068 3.382 0.112 ;
        RECT 3.422 0.498 3.49 0.542 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.922 0.652 ;
        RECT 3.638 0.338 3.706 0.652 ;
        RECT 2.99 0.428 3.274 0.472 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.694 0.472 1.762 0.516 ;
        RECT 1.91 0.472 1.978 0.516 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 3.098 0.428 3.166 0.472 ;
        RECT 3.638 0.403 3.706 0.447 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.922 0.022 ;
        RECT 3.638 -0.022 3.706 0.292 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.614 0.1245 0.682 0.1685 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.91 0.048 1.978 0.092 ;
        RECT 2.666 0.138 2.734 0.182 ;
        RECT 3.098 0.048 3.166 0.092 ;
        RECT 3.638 0.183 3.706 0.227 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.596 0.248 1.04 0.292 ;
      RECT 1.552 0.518 2.32 0.562 ;
      RECT 1.12 0.248 2.876 0.292 ;
      RECT 1.46 0.068 3.076 0.112 ;
      RECT 3.172 0.518 3.848 0.562 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.37 0.518 1.478 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.242 0.158 1.978 0.202 ;
      RECT 2.018 0.158 2.234 0.202 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.882 0.068 2.95 0.382 ;
      RECT 2.342 0.068 2.41 0.472 ;
      RECT 2.774 0.068 2.842 0.562 ;
      RECT 2.99 0.068 3.058 0.202 ;
      RECT 3.098 0.518 3.382 0.562 ;
      RECT 3.746 0.338 3.814 0.562 ;
    LAYER v1 ;
      RECT 3.75 0.518 3.81 0.562 ;
      RECT 3.21 0.518 3.27 0.562 ;
      RECT 2.994 0.068 3.054 0.112 ;
      RECT 2.778 0.248 2.838 0.292 ;
      RECT 2.346 0.068 2.406 0.112 ;
      RECT 2.238 0.518 2.298 0.562 ;
      RECT 2.13 0.248 2.19 0.292 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.482 0.068 1.542 0.112 ;
      RECT 1.158 0.248 1.218 0.292 ;
      RECT 0.942 0.248 1.002 0.292 ;
      RECT 0.618 0.248 0.678 0.292 ;
    LAYER v0 ;
      RECT 3.746 0.403 3.814 0.447 ;
      RECT 3.314 0.248 3.382 0.292 ;
      RECT 3.206 0.518 3.274 0.562 ;
      RECT 2.99 0.138 3.058 0.182 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.774 0.138 2.842 0.182 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.344 0.088 2.408 0.132 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.472 1.87 0.516 ;
      RECT 1.586 0.472 1.654 0.516 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.154 0.473 1.222 0.517 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.006 0.158 1.134 0.202 ;
      RECT 1.114 0.248 1.33 0.292 ;
      RECT 0.898 0.068 1.654 0.112 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.546 0.338 1.762 0.382 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.248 1.438 0.382 ;
      RECT 1.438 0.248 1.802 0.292 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.87 0.248 2.018 0.292 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 2.234 0.158 2.302 0.562 ;
      RECT 2.95 0.338 3.314 0.382 ;
      RECT 3.314 0.158 3.382 0.382 ;
  END
END b15fqy003hn1n08x5

MACRO b15fqy003hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy003hn1n12x5 0 0 ;
  SIZE 4.536 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0207 LAYER m2 ;
      ANTENNAMAXAREACAR 0.61185175 LAYER m1 ;
      ANTENNAMAXAREACAR 5.1925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 0.61185175 LAYER m1 ;
      ANTENNAMAXAREACAR 5.1925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.338 1.978 0.382 ;
        RECT 1.694 0.338 1.762 0.562 ;
        RECT 0.614 0.248 0.682 0.562 ;
      LAYER m2 ;
        RECT 0.596 0.518 1.796 0.562 ;
      LAYER v1 ;
        RECT 0.618 0.518 0.678 0.562 ;
        RECT 1.698 0.518 1.758 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.248 4.246 0.562 ;
      LAYER v0 ;
        RECT 4.178 0.293 4.246 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.248 3.382 0.562 ;
      LAYER v0 ;
        RECT 3.314 0.293 3.382 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.338 3.922 0.382 ;
        RECT 3.854 0.158 3.922 0.382 ;
      LAYER v0 ;
        RECT 3.746 0.338 3.814 0.382 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 8.455 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.382 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.068 4.03 0.562 ;
      LAYER v0 ;
        RECT 3.962 0.472 4.03 0.516 ;
        RECT 3.962 0.099 4.03 0.143 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.57 0.652 ;
        RECT 4.286 0.428 4.354 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 2.126 0.338 2.194 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.83 0.4485 0.898 0.4925 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 1.802 0.473 1.87 0.517 ;
        RECT 2.126 0.473 2.194 0.517 ;
        RECT 2.342 0.473 2.41 0.517 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.746 0.472 3.814 0.516 ;
        RECT 4.286 0.473 4.354 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.57 0.022 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.746 -0.022 3.814 0.292 ;
        RECT 3.206 -0.022 3.274 0.112 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.722 0.1245 0.79 0.1685 ;
        RECT 2.126 0.048 2.194 0.092 ;
        RECT 2.99 0.138 3.058 0.182 ;
        RECT 3.208 0.048 3.272 0.092 ;
        RECT 3.746 0.183 3.814 0.227 ;
        RECT 4.178 0.099 4.246 0.143 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.704 0.338 1.148 0.382 ;
      RECT 1.876 0.518 2.768 0.562 ;
      RECT 3.62 0.518 3.94 0.562 ;
      RECT 1.228 0.338 4.372 0.382 ;
      RECT 1.568 0.068 4.496 0.112 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 1.154 0.338 1.438 0.382 ;
      RECT 0.938 0.068 1.006 0.472 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.91 0.428 1.978 0.562 ;
      RECT 1.154 0.248 1.478 0.292 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 1.566 0.158 2.41 0.202 ;
      RECT 2.45 0.248 2.518 0.472 ;
      RECT 2.666 0.158 2.734 0.382 ;
      RECT 2.342 0.068 2.774 0.112 ;
      RECT 3.098 0.158 3.166 0.472 ;
      RECT 2.882 0.068 2.95 0.562 ;
      RECT 3.422 0.248 3.49 0.562 ;
      RECT 3.854 0.428 3.922 0.562 ;
      RECT 4.07 0.068 4.138 0.562 ;
      RECT 4.286 0.248 4.354 0.382 ;
      RECT 4.394 0.068 4.462 0.562 ;
    LAYER v1 ;
      RECT 4.398 0.068 4.458 0.112 ;
      RECT 4.29 0.338 4.35 0.382 ;
      RECT 4.074 0.338 4.134 0.382 ;
      RECT 3.858 0.518 3.918 0.562 ;
      RECT 3.642 0.518 3.702 0.562 ;
      RECT 2.778 0.068 2.838 0.112 ;
      RECT 2.67 0.338 2.73 0.382 ;
      RECT 2.67 0.518 2.73 0.562 ;
      RECT 2.454 0.068 2.514 0.112 ;
      RECT 2.454 0.338 2.514 0.382 ;
      RECT 1.914 0.518 1.974 0.562 ;
      RECT 1.59 0.068 1.65 0.112 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
    LAYER v0 ;
      RECT 4.394 0.183 4.462 0.227 ;
      RECT 4.394 0.473 4.462 0.517 ;
      RECT 4.286 0.293 4.354 0.337 ;
      RECT 4.07 0.099 4.138 0.143 ;
      RECT 4.07 0.472 4.138 0.516 ;
      RECT 3.854 0.472 3.922 0.516 ;
      RECT 3.53 0.408 3.598 0.452 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.422 0.293 3.49 0.337 ;
      RECT 3.098 0.293 3.166 0.337 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.882 0.448 2.95 0.492 ;
      RECT 2.774 0.338 2.842 0.382 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.473 2.302 0.517 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 2.018 0.473 2.086 0.517 ;
      RECT 1.91 0.473 1.978 0.517 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.3485 1.546 0.3925 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.048 0.498 1.112 0.542 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.722 0.4485 0.79 0.4925 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.448 0.574 0.492 ;
    LAYER m1 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.428 1.35 0.472 ;
      RECT 1.114 0.158 1.458 0.202 ;
      RECT 1.006 0.068 1.654 0.112 ;
      RECT 1.762 0.338 1.978 0.382 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.546 0.248 2.018 0.292 ;
      RECT 2.018 0.248 2.086 0.562 ;
      RECT 2.086 0.248 2.234 0.292 ;
      RECT 2.234 0.248 2.302 0.562 ;
      RECT 2.626 0.518 2.842 0.562 ;
      RECT 2.774 0.068 2.842 0.472 ;
      RECT 3.166 0.158 3.53 0.202 ;
      RECT 3.53 0.158 3.598 0.472 ;
      RECT 3.49 0.518 3.706 0.562 ;
  END
END b15fqy003hn1n12x5

MACRO b15fqy003hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy003hn1n16x5 0 0 ;
  SIZE 5.4 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 5.1925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0342 LAYER m2 ;
      ANTENNAMAXAREACAR 5.1925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.338 2.518 0.382 ;
        RECT 2.018 0.338 2.086 0.562 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER m2 ;
        RECT 0.704 0.518 2.228 0.562 ;
      LAYER v1 ;
        RECT 0.726 0.518 0.786 0.562 ;
        RECT 2.022 0.518 2.082 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.3155 0.79 0.3595 ;
        RECT 2.342 0.338 2.41 0.382 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.042 0.248 5.11 0.562 ;
      LAYER v0 ;
        RECT 5.042 0.293 5.11 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.248 4.138 0.562 ;
      LAYER v0 ;
        RECT 4.07 0.293 4.138 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.502 0.338 4.786 0.382 ;
        RECT 4.718 0.158 4.786 0.382 ;
      LAYER v0 ;
        RECT 4.61 0.338 4.678 0.382 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 8.455 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.81833325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.826 0.068 4.894 0.562 ;
      LAYER v0 ;
        RECT 4.826 0.472 4.894 0.516 ;
        RECT 4.826 0.099 4.894 0.143 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.434 0.652 ;
        RECT 5.15 0.428 5.218 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.91 0.473 1.978 0.517 ;
        RECT 2.126 0.473 2.194 0.517 ;
        RECT 2.45 0.473 2.518 0.517 ;
        RECT 2.666 0.473 2.734 0.517 ;
        RECT 2.99 0.473 3.058 0.517 ;
        RECT 3.746 0.473 3.814 0.517 ;
        RECT 3.962 0.473 4.03 0.517 ;
        RECT 4.61 0.472 4.678 0.516 ;
        RECT 5.15 0.473 5.218 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.434 0.022 ;
        RECT 5.042 -0.022 5.11 0.202 ;
        RECT 4.61 -0.022 4.678 0.292 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 2.342 0.158 3.078 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.746 0.048 3.814 0.092 ;
        RECT 3.962 0.048 4.03 0.092 ;
        RECT 4.61 0.183 4.678 0.227 ;
        RECT 5.042 0.099 5.11 0.143 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.812 0.338 1.256 0.382 ;
      RECT 2.308 0.518 3.616 0.562 ;
      RECT 4.268 0.518 4.804 0.562 ;
      RECT 1.336 0.338 5.236 0.382 ;
      RECT 1.46 0.068 5.36 0.112 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.722 0.248 0.79 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 1.262 0.338 1.762 0.382 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 1.89 0.158 2.214 0.202 ;
      RECT 2.342 0.428 2.41 0.562 ;
      RECT 1.37 0.518 1.802 0.562 ;
      RECT 3.186 0.158 3.314 0.202 ;
      RECT 3.206 0.248 3.274 0.472 ;
      RECT 2.99 0.068 3.638 0.112 ;
      RECT 3.53 0.428 3.598 0.562 ;
      RECT 3.422 0.248 3.49 0.562 ;
      RECT 3.962 0.158 4.03 0.382 ;
      RECT 4.286 0.248 4.354 0.562 ;
      RECT 4.718 0.428 4.786 0.562 ;
      RECT 4.934 0.068 5.002 0.562 ;
      RECT 5.15 0.248 5.218 0.382 ;
      RECT 5.258 0.068 5.326 0.562 ;
    LAYER v1 ;
      RECT 5.262 0.068 5.322 0.112 ;
      RECT 5.154 0.338 5.214 0.382 ;
      RECT 4.938 0.338 4.998 0.382 ;
      RECT 4.722 0.518 4.782 0.562 ;
      RECT 4.29 0.518 4.35 0.562 ;
      RECT 3.642 0.068 3.702 0.112 ;
      RECT 3.534 0.518 3.594 0.562 ;
      RECT 3.318 0.518 3.378 0.562 ;
      RECT 3.21 0.338 3.27 0.382 ;
      RECT 3.102 0.068 3.162 0.112 ;
      RECT 2.346 0.518 2.406 0.562 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.482 0.068 1.542 0.112 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.834 0.338 0.894 0.382 ;
    LAYER v0 ;
      RECT 5.258 0.183 5.326 0.227 ;
      RECT 5.258 0.473 5.326 0.517 ;
      RECT 5.15 0.293 5.218 0.337 ;
      RECT 4.934 0.099 5.002 0.143 ;
      RECT 4.934 0.472 5.002 0.516 ;
      RECT 4.718 0.472 4.786 0.516 ;
      RECT 4.394 0.472 4.462 0.516 ;
      RECT 4.286 0.158 4.354 0.202 ;
      RECT 4.286 0.293 4.354 0.337 ;
      RECT 3.962 0.293 4.03 0.337 ;
      RECT 3.854 0.473 3.922 0.517 ;
      RECT 3.856 0.178 3.92 0.222 ;
      RECT 3.64 0.138 3.704 0.182 ;
      RECT 3.53 0.248 3.598 0.292 ;
      RECT 3.53 0.498 3.598 0.542 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.422 0.498 3.49 0.542 ;
      RECT 3.314 0.498 3.382 0.542 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.206 0.293 3.274 0.337 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 2.99 0.338 3.058 0.382 ;
      RECT 2.774 0.473 2.842 0.517 ;
      RECT 2.558 0.473 2.626 0.517 ;
      RECT 2.342 0.473 2.41 0.517 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.3455 1.87 0.3895 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.156 0.498 1.22 0.542 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.614 0.448 0.682 0.492 ;
    LAYER m1 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 1.222 0.428 1.674 0.472 ;
      RECT 1.222 0.158 1.782 0.202 ;
      RECT 1.114 0.068 1.782 0.112 ;
      RECT 2.086 0.338 2.518 0.382 ;
      RECT 1.478 0.248 1.802 0.292 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.87 0.248 2.558 0.292 ;
      RECT 2.558 0.248 2.626 0.562 ;
      RECT 2.626 0.248 2.774 0.292 ;
      RECT 2.774 0.248 2.842 0.562 ;
      RECT 2.842 0.338 3.166 0.382 ;
      RECT 3.314 0.158 3.382 0.562 ;
      RECT 3.382 0.158 3.51 0.202 ;
      RECT 3.638 0.068 3.706 0.202 ;
      RECT 3.49 0.248 3.854 0.292 ;
      RECT 3.854 0.158 3.922 0.562 ;
      RECT 4.03 0.158 4.394 0.202 ;
      RECT 4.394 0.158 4.462 0.562 ;
  END
END b15fqy003hn1n16x5

MACRO b15fqy00chn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00chn1n02x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.28277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.28277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.248 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.448 2.626 0.492 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.248 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.338 2.842 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 6.08 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.472 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.574 0.112 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.068 0.466 0.112 ;
    END
  END psb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.248 3.382 0.472 ;
        RECT 3.186 0.248 3.382 0.292 ;
      LAYER v0 ;
        RECT 3.206 0.248 3.274 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.338 3.274 0.382 ;
        RECT 2.99 0.068 3.058 0.382 ;
        RECT 2.774 0.068 3.058 0.112 ;
      LAYER v0 ;
        RECT 2.882 0.068 2.95 0.112 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 2.342 0.366 2.41 0.41 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 3.206 0.448 3.274 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.566 0.158 1.978 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 0.486 0.158 0.682 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 3.206 0.113 3.274 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 1.242 0.248 1.91 0.292 ;
      RECT 0.81 0.518 1.046 0.562 ;
      RECT 2.018 0.068 2.086 0.472 ;
    LAYER v0 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.882 0.2455 2.95 0.2895 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.168 2.086 0.212 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.2705 1.114 0.3145 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.83 0.2705 0.898 0.3145 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.398 0.363 0.466 0.407 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.702 0.292 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.428 0.938 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 0.898 0.068 1.782 0.112 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.33 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 2.234 0.562 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.086 0.248 2.45 0.292 ;
      RECT 2.45 0.158 2.518 0.292 ;
      RECT 2.518 0.158 2.882 0.202 ;
      RECT 2.882 0.158 2.95 0.472 ;
      RECT 2.95 0.428 3.078 0.472 ;
  END
END b15fqy00chn1n02x5

MACRO b15fqy00chn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00chn1n03x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.28277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.28277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.248 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.448 2.626 0.492 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.248 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.338 2.842 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 6.08 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.472 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.574 0.112 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.068 0.466 0.112 ;
    END
  END psb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.248 3.382 0.472 ;
        RECT 3.186 0.248 3.382 0.292 ;
      LAYER v0 ;
        RECT 3.206 0.248 3.274 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.338 3.274 0.382 ;
        RECT 2.99 0.068 3.058 0.382 ;
        RECT 2.774 0.068 3.058 0.112 ;
      LAYER v0 ;
        RECT 2.882 0.068 2.95 0.112 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 2.342 0.366 2.41 0.41 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 3.206 0.448 3.274 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.566 0.158 1.978 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 0.486 0.158 0.682 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 3.206 0.113 3.274 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 1.242 0.248 1.91 0.292 ;
      RECT 0.81 0.518 1.046 0.562 ;
      RECT 2.018 0.068 2.086 0.472 ;
    LAYER v0 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.882 0.2455 2.95 0.2895 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.168 2.086 0.212 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.2705 1.114 0.3145 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.83 0.2705 0.898 0.3145 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.398 0.363 0.466 0.407 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.702 0.292 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.428 0.938 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 0.898 0.068 1.782 0.112 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.33 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 2.234 0.562 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.086 0.248 2.45 0.292 ;
      RECT 2.45 0.158 2.518 0.292 ;
      RECT 2.518 0.158 2.882 0.202 ;
      RECT 2.882 0.158 2.95 0.472 ;
      RECT 2.95 0.428 3.078 0.472 ;
  END
END b15fqy00chn1n03x5

MACRO b15fqy00chn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00chn1n04x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.28277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.28277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.248 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.448 2.626 0.492 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.248 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.338 2.842 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 6.08 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.472 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.574 0.112 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.068 0.466 0.112 ;
    END
  END psb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.248 3.382 0.472 ;
        RECT 3.186 0.248 3.382 0.292 ;
      LAYER v0 ;
        RECT 3.206 0.248 3.274 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.338 3.274 0.382 ;
        RECT 2.99 0.068 3.058 0.382 ;
        RECT 2.774 0.068 3.058 0.112 ;
      LAYER v0 ;
        RECT 2.882 0.068 2.95 0.112 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 2.342 0.366 2.41 0.41 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 3.206 0.448 3.274 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.566 0.158 1.978 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 0.486 0.158 0.682 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 3.206 0.113 3.274 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 1.242 0.248 1.91 0.292 ;
      RECT 0.81 0.518 1.046 0.562 ;
      RECT 2.018 0.068 2.086 0.472 ;
    LAYER v0 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.882 0.2455 2.95 0.2895 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.018 0.1695 2.086 0.2135 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.2705 1.114 0.3145 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.83 0.2705 0.898 0.3145 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.398 0.363 0.466 0.407 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.702 0.292 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.428 0.938 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 0.898 0.068 1.782 0.112 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.33 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 2.234 0.562 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.086 0.248 2.45 0.292 ;
      RECT 2.45 0.158 2.518 0.292 ;
      RECT 2.518 0.158 2.882 0.202 ;
      RECT 2.882 0.158 2.95 0.472 ;
      RECT 2.95 0.428 3.078 0.472 ;
  END
END b15fqy00chn1n04x5

MACRO b15fqy00chn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00chn1n06x5 0 0 ;
  SIZE 3.672 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.248 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.481 2.842 0.525 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.248 3.058 0.562 ;
      LAYER v0 ;
        RECT 2.99 0.338 3.058 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.182 0.186 0.25 0.23 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.016 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END psb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.248 3.598 0.472 ;
        RECT 3.402 0.248 3.598 0.292 ;
      LAYER v0 ;
        RECT 3.422 0.248 3.49 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.116 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.338 3.49 0.382 ;
        RECT 3.206 0.068 3.274 0.382 ;
        RECT 2.99 0.068 3.274 0.112 ;
      LAYER v0 ;
        RECT 3.098 0.068 3.166 0.112 ;
        RECT 3.314 0.338 3.382 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.706 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.29 0.3905 0.358 0.4345 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.558 0.366 2.626 0.41 ;
        RECT 2.882 0.481 2.95 0.525 ;
        RECT 3.422 0.448 3.49 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.706 0.022 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 0.594 0.158 0.79 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.186 0.142 0.23 ;
        RECT 0.29 0.186 0.358 0.23 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.422 0.113 3.49 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.154 0.248 1.782 0.292 ;
      RECT 1.458 0.338 1.91 0.382 ;
      RECT 0.918 0.518 1.154 0.562 ;
      RECT 2.234 0.068 2.302 0.472 ;
    LAYER v0 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.2455 3.166 0.2895 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.234 0.1705 2.302 0.2145 ;
      RECT 2.234 0.408 2.302 0.452 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 2.018 0.3155 2.086 0.3595 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.358 1.222 0.402 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.938 0.2705 1.006 0.3145 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.363 0.574 0.407 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.248 0.81 0.292 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.006 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.158 1.802 0.202 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 1.87 0.068 1.998 0.112 ;
      RECT 1.91 0.158 1.978 0.382 ;
      RECT 1.978 0.158 2.126 0.202 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.518 1.37 0.562 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.438 0.428 2.018 0.472 ;
      RECT 2.018 0.248 2.086 0.562 ;
      RECT 2.086 0.518 2.45 0.562 ;
      RECT 2.45 0.428 2.518 0.562 ;
      RECT 2.302 0.248 2.666 0.292 ;
      RECT 2.666 0.158 2.734 0.292 ;
      RECT 2.734 0.158 3.098 0.202 ;
      RECT 3.098 0.158 3.166 0.472 ;
      RECT 3.166 0.428 3.294 0.472 ;
  END
END b15fqy00chn1n06x5

MACRO b15fqy00chn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00chn1n08x5 0 0 ;
  SIZE 4.104 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.43833325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.43833325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.158 2.842 0.472 ;
      LAYER v0 ;
        RECT 2.774 0.384 2.842 0.428 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.248 3.166 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.423 0.25 0.467 ;
        RECT 0.182 0.203 0.25 0.247 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.87666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END psb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.248 3.814 0.382 ;
      LAYER v0 ;
        RECT 3.746 0.2705 3.814 0.3145 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.158 3.922 0.382 ;
        RECT 3.53 0.158 3.922 0.202 ;
        RECT 3.53 0.068 3.598 0.382 ;
        RECT 3.206 0.068 3.598 0.112 ;
      LAYER v0 ;
        RECT 3.314 0.068 3.382 0.112 ;
        RECT 3.53 0.2705 3.598 0.3145 ;
        RECT 3.854 0.2705 3.922 0.3145 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.138 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.423 0.142 0.467 ;
        RECT 0.29 0.423 0.358 0.467 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.99 0.473 3.058 0.517 ;
        RECT 3.746 0.538 3.814 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.138 0.022 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 1.566 0.158 2.214 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 0.594 0.158 0.79 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
        RECT 0.29 0.113 0.358 0.157 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 3.098 0.048 3.166 0.092 ;
        RECT 3.746 0.048 3.814 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.458 0.338 2.018 0.382 ;
      RECT 0.918 0.518 1.154 0.562 ;
      RECT 2.666 0.068 2.734 0.472 ;
      RECT 2.882 0.158 2.95 0.562 ;
      RECT 3.314 0.248 3.382 0.472 ;
    LAYER v0 ;
      RECT 3.962 0.158 4.03 0.202 ;
      RECT 3.964 0.498 4.028 0.542 ;
      RECT 3.422 0.518 3.49 0.562 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 2.882 0.2025 2.95 0.2465 ;
      RECT 2.882 0.473 2.95 0.517 ;
      RECT 2.666 0.1775 2.734 0.2215 ;
      RECT 2.666 0.384 2.734 0.428 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.558 0.384 2.626 0.428 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.938 0.2705 1.006 0.3145 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.363 0.574 0.407 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.248 0.81 0.292 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.33 0.248 1.89 0.292 ;
      RECT 1.006 0.068 1.89 0.112 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 2.086 0.248 2.342 0.292 ;
      RECT 2.342 0.158 2.41 0.292 ;
      RECT 2.41 0.158 2.558 0.202 ;
      RECT 2.558 0.158 2.626 0.472 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.518 1.37 0.562 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.438 0.428 2.126 0.472 ;
      RECT 2.126 0.338 2.194 0.472 ;
      RECT 2.194 0.338 2.45 0.382 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.518 0.518 2.842 0.562 ;
      RECT 2.734 0.068 2.99 0.112 ;
      RECT 2.99 0.068 3.058 0.202 ;
      RECT 3.058 0.158 3.206 0.202 ;
      RECT 3.206 0.158 3.274 0.562 ;
      RECT 3.274 0.158 3.49 0.202 ;
      RECT 3.274 0.518 3.51 0.562 ;
      RECT 3.382 0.428 3.962 0.472 ;
      RECT 3.962 0.068 4.03 0.562 ;
  END
END b15fqy00chn1n08x5

MACRO b15fqy00chn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00chn1n12x5 0 0 ;
  SIZE 4.752 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.43833325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.43833325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.518 3.382 0.562 ;
        RECT 3.314 0.338 3.382 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.518 3.166 0.562 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.338 3.922 0.472 ;
        RECT 3.422 0.338 3.922 0.382 ;
      LAYER v0 ;
        RECT 3.53 0.338 3.598 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.408 0.142 0.452 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.408 0.358 0.452 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 3.9425 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 3.154 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END psb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.248 4.678 0.562 ;
        RECT 4.394 0.248 4.678 0.292 ;
      LAYER v0 ;
        RECT 4.502 0.248 4.57 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 10.735 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.68375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.338 4.57 0.382 ;
        RECT 4.286 0.068 4.354 0.382 ;
        RECT 3.726 0.068 4.354 0.112 ;
      LAYER v0 ;
        RECT 3.746 0.068 3.814 0.112 ;
        RECT 4.394 0.338 4.462 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.786 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 3.638 0.518 3.706 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.398 0.493 0.466 0.537 ;
        RECT 0.614 0.493 0.682 0.537 ;
        RECT 0.938 0.383 1.006 0.427 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.018 0.538 2.086 0.582 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 3.422 0.538 3.49 0.582 ;
        RECT 3.638 0.538 3.706 0.582 ;
        RECT 4.502 0.448 4.57 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.786 0.022 ;
        RECT 4.502 -0.022 4.57 0.202 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 1.89 0.158 2.626 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 3.422 0.048 3.49 0.092 ;
        RECT 4.502 0.113 4.57 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.782 0.338 2.882 0.382 ;
      RECT 1.134 0.518 1.478 0.562 ;
      RECT 3.422 0.428 3.746 0.472 ;
      RECT 3.422 0.158 4.05 0.202 ;
      RECT 2.99 0.338 3.058 0.472 ;
    LAYER v0 ;
      RECT 4.178 0.399 4.246 0.443 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 4.07 0.399 4.138 0.443 ;
      RECT 3.962 0.158 4.03 0.202 ;
      RECT 3.962 0.399 4.03 0.443 ;
      RECT 3.854 0.248 3.922 0.292 ;
      RECT 3.53 0.158 3.598 0.202 ;
      RECT 3.53 0.428 3.598 0.472 ;
      RECT 2.99 0.248 3.058 0.292 ;
      RECT 2.99 0.408 3.058 0.452 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.882 0.498 2.95 0.542 ;
      RECT 2.774 0.338 2.842 0.382 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.342 0.248 2.41 0.292 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.586 0.268 1.654 0.312 ;
      RECT 1.478 0.4055 1.546 0.4495 ;
      RECT 1.37 0.178 1.438 0.222 ;
      RECT 1.262 0.2705 1.33 0.3145 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.493 0.79 0.537 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.508 0.408 0.572 0.452 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.472 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.898 0.248 1.046 0.292 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.114 0.428 1.37 0.472 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 1.654 0.428 2.302 0.472 ;
      RECT 1.33 0.068 2.322 0.112 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.546 0.158 1.694 0.202 ;
      RECT 1.694 0.158 1.762 0.292 ;
      RECT 1.762 0.248 3.078 0.292 ;
      RECT 3.746 0.428 3.814 0.562 ;
      RECT 3.814 0.518 4.07 0.562 ;
      RECT 4.07 0.338 4.138 0.562 ;
      RECT 3.058 0.338 3.206 0.382 ;
      RECT 2.862 0.158 3.206 0.202 ;
      RECT 3.206 0.158 3.274 0.382 ;
      RECT 3.274 0.248 3.962 0.292 ;
      RECT 3.962 0.248 4.03 0.472 ;
      RECT 4.03 0.248 4.178 0.292 ;
      RECT 4.178 0.248 4.246 0.472 ;
  END
END b15fqy00chn1n12x5

MACRO b15fqy00chn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00chn1n16x5 0 0 ;
  SIZE 5.616 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0198 LAYER m2 ;
      ANTENNAMAXAREACAR 1.497037 LAYER m1 ;
      ANTENNAMAXAREACAR 5.734074 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 1.497037 LAYER m1 ;
      ANTENNAMAXAREACAR 5.734074 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.214 0.338 2.734 0.382 ;
        RECT 0.83 0.338 0.898 0.562 ;
      LAYER m2 ;
        RECT 0.812 0.338 2.32 0.382 ;
      LAYER v1 ;
        RECT 0.834 0.338 0.894 0.382 ;
        RECT 2.238 0.338 2.298 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 2.234 0.338 2.302 0.382 ;
        RECT 2.558 0.338 2.626 0.382 ;
    END
  END psb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.518 4.246 0.562 ;
        RECT 4.178 0.428 4.246 0.562 ;
      LAYER v0 ;
        RECT 4.18 0.448 4.244 0.492 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.338 4.482 0.382 ;
        RECT 4.07 0.158 4.138 0.382 ;
      LAYER v0 ;
        RECT 4.394 0.338 4.462 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.4495 0.25 0.4935 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.398 0.4495 0.466 0.4935 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.474 0.248 5.542 0.562 ;
        RECT 5.258 0.248 5.542 0.292 ;
      LAYER v0 ;
        RECT 5.366 0.248 5.434 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 10.735 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 2.147 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.15 0.338 5.434 0.382 ;
        RECT 5.15 0.068 5.218 0.382 ;
        RECT 4.59 0.068 5.218 0.112 ;
      LAYER v0 ;
        RECT 4.61 0.068 4.678 0.112 ;
        RECT 5.258 0.338 5.326 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.65 0.652 ;
        RECT 5.366 0.428 5.434 0.652 ;
        RECT 4.502 0.518 4.57 0.652 ;
        RECT 4.286 0.518 4.354 0.652 ;
        RECT 3.854 0.428 3.922 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.666 0.4505 2.734 0.4945 ;
        RECT 3.854 0.473 3.922 0.517 ;
        RECT 4.288 0.538 4.352 0.582 ;
        RECT 4.504 0.538 4.568 0.582 ;
        RECT 5.366 0.448 5.434 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.65 0.022 ;
        RECT 5.366 -0.022 5.434 0.202 ;
        RECT 4.286 -0.022 4.354 0.112 ;
        RECT 3.854 -0.022 3.922 0.202 ;
        RECT 2.214 0.158 3.166 0.202 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
        RECT 0.29 0.113 0.358 0.157 ;
        RECT 0.506 0.113 0.574 0.157 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.882 0.158 2.95 0.202 ;
        RECT 3.854 0.138 3.922 0.182 ;
        RECT 4.286 0.048 4.354 0.092 ;
        RECT 5.366 0.113 5.434 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 1.37 0.068 1.438 0.382 ;
      RECT 1.91 0.428 2.538 0.472 ;
      RECT 2.214 0.338 2.734 0.382 ;
      RECT 1.242 0.518 1.802 0.562 ;
      RECT 2.774 0.338 2.842 0.472 ;
      RECT 4.286 0.428 4.718 0.472 ;
      RECT 4.286 0.158 4.914 0.202 ;
      RECT 3.402 0.518 3.746 0.562 ;
    LAYER v0 ;
      RECT 5.042 0.399 5.11 0.443 ;
      RECT 4.934 0.248 5.002 0.292 ;
      RECT 4.934 0.399 5.002 0.443 ;
      RECT 4.826 0.158 4.894 0.202 ;
      RECT 4.826 0.399 4.894 0.443 ;
      RECT 4.718 0.248 4.786 0.292 ;
      RECT 4.394 0.158 4.462 0.202 ;
      RECT 4.394 0.428 4.462 0.472 ;
      RECT 3.53 0.428 3.598 0.472 ;
      RECT 3.422 0.248 3.49 0.292 ;
      RECT 3.422 0.338 3.49 0.382 ;
      RECT 3.422 0.518 3.49 0.562 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 2.99 0.338 3.058 0.382 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.776 0.358 2.84 0.402 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.293 1.438 0.337 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.614 0.223 0.682 0.267 ;
      RECT 0.614 0.4495 0.682 0.4935 ;
    LAYER m1 ;
      RECT 0.938 0.248 1.006 0.562 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.222 0.428 1.478 0.472 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.546 0.428 1.674 0.472 ;
      RECT 1.546 0.158 1.89 0.202 ;
      RECT 1.438 0.068 2.97 0.112 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.87 0.248 2.882 0.292 ;
      RECT 2.882 0.248 2.95 0.382 ;
      RECT 2.95 0.338 3.51 0.382 ;
      RECT 2.842 0.428 3.638 0.472 ;
      RECT 3.098 0.248 3.638 0.292 ;
      RECT 3.638 0.248 3.706 0.472 ;
      RECT 4.718 0.428 4.786 0.562 ;
      RECT 4.786 0.518 4.934 0.562 ;
      RECT 4.934 0.338 5.002 0.562 ;
      RECT 3.294 0.158 3.746 0.202 ;
      RECT 3.746 0.158 3.814 0.562 ;
      RECT 3.814 0.248 3.962 0.292 ;
      RECT 3.962 0.068 4.03 0.292 ;
      RECT 4.03 0.068 4.178 0.112 ;
      RECT 4.178 0.068 4.246 0.292 ;
      RECT 4.246 0.248 4.826 0.292 ;
      RECT 4.826 0.248 4.894 0.472 ;
      RECT 4.894 0.248 5.042 0.292 ;
      RECT 5.042 0.248 5.11 0.472 ;
  END
END b15fqy00chn1n16x5

MACRO b15fqy00fhn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00fhn1n02x5 0 0 ;
  SIZE 3.78 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 8.348889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 8.348889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.158 3.49 0.562 ;
        RECT 1.802 0.518 2.086 0.562 ;
      LAYER m2 ;
        RECT 1.892 0.518 3.616 0.562 ;
      LAYER v1 ;
        RECT 1.914 0.518 1.974 0.562 ;
        RECT 3.426 0.518 3.486 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.518 1.978 0.562 ;
        RECT 3.422 0.248 3.49 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.068 3.058 0.382 ;
        RECT 2.342 0.338 2.626 0.382 ;
      LAYER m2 ;
        RECT 2.432 0.338 3.076 0.382 ;
      LAYER v1 ;
        RECT 2.562 0.338 2.622 0.382 ;
        RECT 2.994 0.338 3.054 0.382 ;
      LAYER v0 ;
        RECT 2.45 0.338 2.518 0.382 ;
        RECT 2.99 0.088 3.058 0.132 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.498 1.006 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.068 3.706 0.562 ;
      LAYER v0 ;
        RECT 3.638 0.448 3.706 0.492 ;
        RECT 3.638 0.138 3.706 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.814 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 1.154 0.47 1.222 0.514 ;
        RECT 1.694 0.538 1.762 0.582 ;
        RECT 2.342 0.4575 2.41 0.5015 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.532 0.538 3.596 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.814 0.022 ;
        RECT 3.53 -0.022 3.598 0.202 ;
        RECT 3.098 -0.022 3.166 0.292 ;
        RECT 1.694 0.158 2.41 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.722 0.203 0.79 0.247 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 3.098 0.203 3.166 0.247 ;
        RECT 3.53 0.138 3.598 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 1.256 0.382 ;
      RECT 0.812 0.518 1.456 0.562 ;
      RECT 1.336 0.338 2.104 0.382 ;
      RECT 1.028 0.428 2.66 0.472 ;
      RECT 2.74 0.428 3.616 0.472 ;
    LAYER m1 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 0.83 0.068 0.898 0.562 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.262 0.068 1.33 0.472 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.262 0.518 1.566 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.802 0.518 2.086 0.562 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 2.342 0.338 2.626 0.382 ;
      RECT 2.45 0.428 2.666 0.472 ;
      RECT 2.558 0.158 2.774 0.202 ;
      RECT 1.91 0.068 2.882 0.112 ;
      RECT 3.206 0.248 3.274 0.562 ;
      RECT 2.99 0.068 3.058 0.382 ;
      RECT 3.098 0.428 3.166 0.562 ;
      RECT 3.422 0.158 3.49 0.562 ;
      RECT 3.53 0.248 3.598 0.472 ;
    LAYER v1 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 3.53 0.338 3.598 0.382 ;
      RECT 3.314 0.138 3.382 0.182 ;
      RECT 3.206 0.448 3.274 0.492 ;
      RECT 3.098 0.448 3.166 0.492 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.37 0.3835 1.438 0.4275 ;
      RECT 1.262 0.138 1.33 0.182 ;
      RECT 1.262 0.3835 1.33 0.4275 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.83 0.203 0.898 0.247 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.506 0.2075 0.574 0.2515 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 1.438 0.158 1.654 0.202 ;
      RECT 1.762 0.428 2.234 0.472 ;
      RECT 2.234 0.248 2.302 0.472 ;
      RECT 2.302 0.248 2.626 0.292 ;
      RECT 2.666 0.248 2.734 0.472 ;
      RECT 2.774 0.158 2.842 0.562 ;
      RECT 2.882 0.068 2.95 0.472 ;
      RECT 3.274 0.248 3.314 0.292 ;
      RECT 3.314 0.068 3.382 0.292 ;
  END
END b15fqy00fhn1n02x5

MACRO b15fqy00fhn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00fhn1n03x5 0 0 ;
  SIZE 3.996 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 6.679111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 6.679111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.158 3.706 0.562 ;
        RECT 1.802 0.518 2.086 0.562 ;
      LAYER m2 ;
        RECT 1.892 0.518 3.724 0.562 ;
      LAYER v1 ;
        RECT 1.914 0.518 1.974 0.562 ;
        RECT 3.642 0.518 3.702 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.518 1.978 0.562 ;
        RECT 3.638 0.248 3.706 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.068 3.274 0.382 ;
        RECT 2.646 0.338 2.842 0.382 ;
      LAYER m2 ;
        RECT 2.632 0.338 3.292 0.382 ;
      LAYER v1 ;
        RECT 2.778 0.338 2.838 0.382 ;
        RECT 3.21 0.338 3.27 0.382 ;
      LAYER v0 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 3.206 0.088 3.274 0.132 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.498 1.006 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.068 3.922 0.562 ;
      LAYER v0 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 3.854 0.138 3.922 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 1.154 0.47 1.222 0.514 ;
        RECT 1.694 0.538 1.762 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.558 0.538 2.626 0.582 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 3.748 0.538 3.812 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.03 0.022 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.314 -0.022 3.382 0.292 ;
        RECT 1.694 0.158 2.322 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.722 0.203 0.79 0.247 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 3.314 0.203 3.382 0.247 ;
        RECT 3.746 0.138 3.814 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 1.256 0.382 ;
      RECT 0.812 0.518 1.456 0.562 ;
      RECT 1.336 0.338 2.552 0.382 ;
      RECT 1.028 0.428 2.876 0.472 ;
      RECT 2.956 0.428 3.832 0.472 ;
    LAYER m1 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 0.83 0.068 0.898 0.562 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.262 0.068 1.33 0.472 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.262 0.518 1.566 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.802 0.518 2.086 0.562 ;
      RECT 2.342 0.338 2.538 0.382 ;
      RECT 2.646 0.338 2.842 0.382 ;
      RECT 2.666 0.428 2.882 0.472 ;
      RECT 2.774 0.158 2.99 0.202 ;
      RECT 1.91 0.068 3.098 0.112 ;
      RECT 3.422 0.248 3.49 0.562 ;
      RECT 3.206 0.068 3.274 0.382 ;
      RECT 3.314 0.428 3.382 0.562 ;
      RECT 3.638 0.158 3.706 0.562 ;
      RECT 3.746 0.248 3.814 0.472 ;
    LAYER v1 ;
      RECT 3.75 0.428 3.81 0.472 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 2.994 0.428 3.054 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.454 0.338 2.514 0.382 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 3.746 0.338 3.814 0.382 ;
      RECT 3.53 0.138 3.598 0.182 ;
      RECT 3.422 0.448 3.49 0.492 ;
      RECT 3.314 0.448 3.382 0.492 ;
      RECT 3.098 0.338 3.166 0.382 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.37 0.3835 1.438 0.4275 ;
      RECT 1.262 0.138 1.33 0.182 ;
      RECT 1.262 0.3835 1.33 0.4275 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.83 0.203 0.898 0.247 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.506 0.2075 0.574 0.2515 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 1.438 0.158 1.654 0.202 ;
      RECT 1.762 0.428 2.126 0.472 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.194 0.428 2.43 0.472 ;
      RECT 2.194 0.248 2.842 0.292 ;
      RECT 2.882 0.248 2.95 0.472 ;
      RECT 2.99 0.158 3.058 0.562 ;
      RECT 3.098 0.068 3.166 0.472 ;
      RECT 3.49 0.248 3.53 0.292 ;
      RECT 3.53 0.068 3.598 0.292 ;
  END
END b15fqy00fhn1n03x5

MACRO b15fqy00fhn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00fhn1n04x5 0 0 ;
  SIZE 3.996 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 5.751111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 5.751111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.158 3.706 0.562 ;
        RECT 1.802 0.518 2.086 0.562 ;
      LAYER m2 ;
        RECT 1.892 0.518 3.724 0.562 ;
      LAYER v1 ;
        RECT 1.914 0.518 1.974 0.562 ;
        RECT 3.642 0.518 3.702 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.518 1.978 0.562 ;
        RECT 3.638 0.248 3.706 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.068 3.274 0.382 ;
        RECT 2.646 0.338 2.842 0.382 ;
      LAYER m2 ;
        RECT 2.632 0.338 3.292 0.382 ;
      LAYER v1 ;
        RECT 2.778 0.338 2.838 0.382 ;
        RECT 3.21 0.338 3.27 0.382 ;
      LAYER v0 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 3.206 0.088 3.274 0.132 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.498 1.006 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.068 3.922 0.562 ;
      LAYER v0 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 3.854 0.138 3.922 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 1.154 0.47 1.222 0.514 ;
        RECT 1.694 0.538 1.762 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.558 0.538 2.626 0.582 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 3.748 0.538 3.812 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.03 0.022 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.314 -0.022 3.382 0.292 ;
        RECT 1.694 0.158 2.322 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.722 0.203 0.79 0.247 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 3.314 0.203 3.382 0.247 ;
        RECT 3.746 0.138 3.814 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 1.256 0.382 ;
      RECT 0.812 0.518 1.456 0.562 ;
      RECT 1.336 0.338 2.552 0.382 ;
      RECT 1.028 0.428 2.876 0.472 ;
      RECT 2.956 0.428 3.832 0.472 ;
    LAYER m1 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 0.83 0.068 0.898 0.562 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.262 0.068 1.33 0.472 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.262 0.518 1.566 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.802 0.518 2.086 0.562 ;
      RECT 2.342 0.338 2.538 0.382 ;
      RECT 2.646 0.338 2.842 0.382 ;
      RECT 2.666 0.428 2.882 0.472 ;
      RECT 2.774 0.158 2.99 0.202 ;
      RECT 1.91 0.068 3.098 0.112 ;
      RECT 3.422 0.248 3.49 0.562 ;
      RECT 3.206 0.068 3.274 0.382 ;
      RECT 3.314 0.428 3.382 0.562 ;
      RECT 3.638 0.158 3.706 0.562 ;
      RECT 3.746 0.248 3.814 0.472 ;
    LAYER v1 ;
      RECT 3.75 0.428 3.81 0.472 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 2.994 0.428 3.054 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.454 0.338 2.514 0.382 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 3.746 0.338 3.814 0.382 ;
      RECT 3.53 0.138 3.598 0.182 ;
      RECT 3.422 0.448 3.49 0.492 ;
      RECT 3.314 0.448 3.382 0.492 ;
      RECT 3.098 0.338 3.166 0.382 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.37 0.3835 1.438 0.4275 ;
      RECT 1.262 0.138 1.33 0.182 ;
      RECT 1.262 0.3835 1.33 0.4275 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.83 0.203 0.898 0.247 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.506 0.2075 0.574 0.2515 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 1.438 0.158 1.654 0.202 ;
      RECT 1.762 0.428 2.126 0.472 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 2.194 0.428 2.43 0.472 ;
      RECT 2.194 0.248 2.842 0.292 ;
      RECT 2.882 0.248 2.95 0.472 ;
      RECT 2.99 0.158 3.058 0.562 ;
      RECT 3.098 0.068 3.166 0.472 ;
      RECT 3.49 0.248 3.53 0.292 ;
      RECT 3.53 0.068 3.598 0.292 ;
  END
END b15fqy00fhn1n04x5

MACRO b15fqy00fhn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00fhn1n06x5 0 0 ;
  SIZE 4.32 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 6.679111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 6.679111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.158 3.922 0.562 ;
        RECT 1.802 0.518 2.086 0.562 ;
      LAYER m2 ;
        RECT 1.892 0.518 3.94 0.562 ;
      LAYER v1 ;
        RECT 1.914 0.518 1.974 0.562 ;
        RECT 3.858 0.518 3.918 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.518 1.978 0.562 ;
        RECT 3.854 0.248 3.922 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.068 3.49 0.382 ;
        RECT 2.862 0.338 3.058 0.382 ;
      LAYER m2 ;
        RECT 2.74 0.338 3.508 0.382 ;
      LAYER v1 ;
        RECT 2.994 0.338 3.054 0.382 ;
        RECT 3.426 0.338 3.486 0.382 ;
      LAYER v0 ;
        RECT 2.882 0.338 2.95 0.382 ;
        RECT 3.422 0.088 3.49 0.132 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.498 1.006 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.068 4.138 0.562 ;
      LAYER v0 ;
        RECT 4.07 0.448 4.138 0.492 ;
        RECT 4.07 0.138 4.138 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.354 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 1.154 0.47 1.222 0.514 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 2.236 0.428 2.3 0.472 ;
        RECT 2.776 0.538 2.84 0.582 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.746 0.448 3.814 0.492 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 4.178 0.448 4.246 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.354 0.022 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.53 -0.022 3.598 0.292 ;
        RECT 1.694 0.158 2.538 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.722 0.203 0.79 0.247 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 3.53 0.203 3.598 0.247 ;
        RECT 3.962 0.138 4.03 0.182 ;
        RECT 4.178 0.138 4.246 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 1.256 0.382 ;
      RECT 0.812 0.518 1.456 0.562 ;
      RECT 1.336 0.338 2.66 0.382 ;
      RECT 1.028 0.428 3.092 0.472 ;
      RECT 3.172 0.428 4.048 0.472 ;
    LAYER m1 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 0.83 0.068 0.898 0.562 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.262 0.068 1.33 0.472 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.262 0.518 1.566 0.562 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.802 0.518 2.086 0.562 ;
      RECT 2.45 0.338 2.754 0.382 ;
      RECT 2.862 0.338 3.058 0.382 ;
      RECT 2.99 0.428 3.098 0.472 ;
      RECT 2.99 0.158 3.206 0.202 ;
      RECT 1.91 0.068 3.314 0.112 ;
      RECT 3.638 0.248 3.706 0.562 ;
      RECT 3.422 0.068 3.49 0.382 ;
      RECT 3.53 0.428 3.598 0.562 ;
      RECT 3.854 0.158 3.922 0.562 ;
      RECT 3.962 0.248 4.03 0.472 ;
    LAYER v1 ;
      RECT 3.966 0.428 4.026 0.472 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 2.994 0.428 3.054 0.472 ;
      RECT 2.562 0.338 2.622 0.382 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 3.962 0.338 4.03 0.382 ;
      RECT 3.746 0.138 3.814 0.182 ;
      RECT 3.638 0.448 3.706 0.492 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 3.098 0.158 3.166 0.202 ;
      RECT 3.098 0.338 3.166 0.382 ;
      RECT 2.882 0.248 2.95 0.292 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.37 0.3835 1.438 0.4275 ;
      RECT 1.262 0.138 1.33 0.182 ;
      RECT 1.262 0.3835 1.33 0.4275 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.83 0.203 0.898 0.247 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.506 0.2075 0.574 0.2515 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 1.438 0.158 1.654 0.202 ;
      RECT 1.762 0.428 2.018 0.472 ;
      RECT 2.018 0.248 2.086 0.472 ;
      RECT 2.086 0.248 2.342 0.292 ;
      RECT 2.342 0.248 2.41 0.472 ;
      RECT 2.41 0.428 2.538 0.472 ;
      RECT 2.41 0.248 3.058 0.292 ;
      RECT 3.098 0.248 3.166 0.472 ;
      RECT 3.206 0.158 3.274 0.562 ;
      RECT 3.314 0.068 3.382 0.472 ;
      RECT 3.706 0.248 3.746 0.292 ;
      RECT 3.746 0.068 3.814 0.292 ;
  END
END b15fqy00fhn1n06x5

MACRO b15fqy00fhn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00fhn1n08x5 0 0 ;
  SIZE 4.86 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 5.751111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.009 LAYER m2 ;
      ANTENNAMAXAREACAR 5.751111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.158 4.462 0.562 ;
        RECT 2.018 0.518 2.302 0.562 ;
      LAYER m2 ;
        RECT 2.108 0.518 4.48 0.562 ;
      LAYER v1 ;
        RECT 2.13 0.518 2.19 0.562 ;
        RECT 4.398 0.518 4.458 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.518 2.194 0.562 ;
        RECT 4.394 0.248 4.462 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 6.648889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.068 4.03 0.382 ;
        RECT 3.294 0.338 3.598 0.382 ;
      LAYER m2 ;
        RECT 3.512 0.338 4.048 0.382 ;
      LAYER v1 ;
        RECT 3.534 0.338 3.594 0.382 ;
        RECT 3.966 0.338 4.026 0.382 ;
      LAYER v0 ;
        RECT 3.422 0.338 3.49 0.382 ;
        RECT 3.962 0.088 4.03 0.132 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.498 1.006 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.068 4.678 0.562 ;
      LAYER v0 ;
        RECT 4.61 0.448 4.678 0.492 ;
        RECT 4.61 0.138 4.678 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.894 0.652 ;
        RECT 4.718 0.428 4.786 0.652 ;
        RECT 4.502 0.518 4.57 0.652 ;
        RECT 4.286 0.428 4.354 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.342 0.3835 2.41 0.4275 ;
        RECT 2.56 0.428 2.624 0.472 ;
        RECT 3.314 0.538 3.382 0.582 ;
        RECT 3.962 0.448 4.03 0.492 ;
        RECT 4.286 0.448 4.354 0.492 ;
        RECT 4.504 0.538 4.568 0.582 ;
        RECT 4.718 0.448 4.786 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.894 0.022 ;
        RECT 4.718 -0.022 4.786 0.202 ;
        RECT 4.502 -0.022 4.57 0.202 ;
        RECT 4.07 -0.022 4.138 0.292 ;
        RECT 1.91 0.158 3.078 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.722 0.203 0.79 0.247 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 2.774 0.158 2.842 0.202 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 4.07 0.203 4.138 0.247 ;
        RECT 4.502 0.138 4.57 0.182 ;
        RECT 4.718 0.138 4.786 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 1.472 0.382 ;
      RECT 0.812 0.518 1.672 0.562 ;
      RECT 1.552 0.338 2.968 0.382 ;
      RECT 1.028 0.428 3.632 0.472 ;
      RECT 3.712 0.428 4.588 0.472 ;
    LAYER m1 ;
      RECT 0.83 0.068 0.898 0.562 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.262 0.248 1.33 0.382 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 1.586 0.518 1.782 0.562 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 2.018 0.518 2.302 0.562 ;
      RECT 2.774 0.338 3.186 0.382 ;
      RECT 3.294 0.338 3.598 0.382 ;
      RECT 3.422 0.428 3.638 0.472 ;
      RECT 3.53 0.158 3.746 0.202 ;
      RECT 2.126 0.068 3.854 0.112 ;
      RECT 4.178 0.248 4.246 0.562 ;
      RECT 3.962 0.068 4.03 0.382 ;
      RECT 4.07 0.428 4.138 0.562 ;
      RECT 4.394 0.158 4.462 0.562 ;
      RECT 4.502 0.248 4.57 0.472 ;
    LAYER v1 ;
      RECT 4.506 0.428 4.566 0.472 ;
      RECT 4.074 0.428 4.134 0.472 ;
      RECT 3.75 0.428 3.81 0.472 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 2.886 0.338 2.946 0.382 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 4.502 0.338 4.57 0.382 ;
      RECT 4.286 0.138 4.354 0.182 ;
      RECT 4.178 0.448 4.246 0.492 ;
      RECT 4.07 0.448 4.138 0.492 ;
      RECT 3.854 0.338 3.922 0.382 ;
      RECT 3.746 0.068 3.814 0.112 ;
      RECT 3.746 0.428 3.814 0.472 ;
      RECT 3.638 0.158 3.706 0.202 ;
      RECT 3.638 0.338 3.706 0.382 ;
      RECT 3.422 0.248 3.49 0.292 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.338 3.166 0.382 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.3835 1.654 0.4275 ;
      RECT 1.48 0.088 1.544 0.132 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.83 0.203 0.898 0.247 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.506 0.2075 0.574 0.2515 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.114 0.158 1.478 0.202 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 1.654 0.158 1.87 0.202 ;
      RECT 1.978 0.428 2.234 0.472 ;
      RECT 2.234 0.248 2.302 0.472 ;
      RECT 2.302 0.248 2.666 0.292 ;
      RECT 2.666 0.248 2.734 0.472 ;
      RECT 2.734 0.428 3.382 0.472 ;
      RECT 2.734 0.248 3.598 0.292 ;
      RECT 3.638 0.248 3.706 0.472 ;
      RECT 3.746 0.158 3.814 0.562 ;
      RECT 3.854 0.068 3.922 0.472 ;
      RECT 4.246 0.248 4.286 0.292 ;
      RECT 4.286 0.068 4.354 0.292 ;
  END
END b15fqy00fhn1n08x5

MACRO b15fqy00fhn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00fhn1n12x5 0 0 ;
  SIZE 5.94 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 5.565926 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 5.565926 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.366 0.158 5.434 0.562 ;
        RECT 2.666 0.428 2.734 0.562 ;
      LAYER m2 ;
        RECT 2.648 0.518 5.452 0.562 ;
      LAYER v1 ;
        RECT 2.67 0.518 2.73 0.562 ;
        RECT 5.37 0.518 5.43 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.49 2.734 0.534 ;
        RECT 5.366 0.248 5.434 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAGATEAREA 0.0207 LAYER m2 ;
      ANTENNAMAXAREACAR 2.49714275 LAYER m1 ;
      ANTENNAMAXAREACAR 6.640635 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.89396825 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
      ANTENNAMAXAREACAR 7.7474075 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.042 0.248 5.218 0.292 ;
        RECT 5.15 0.068 5.218 0.292 ;
        RECT 5.042 0.248 5.11 0.382 ;
        RECT 3.962 0.338 4.158 0.382 ;
      LAYER m2 ;
        RECT 4.036 0.338 5.128 0.382 ;
      LAYER v1 ;
        RECT 4.074 0.338 4.134 0.382 ;
        RECT 5.046 0.338 5.106 0.382 ;
      LAYER v0 ;
        RECT 4.07 0.338 4.138 0.382 ;
        RECT 5.15 0.138 5.218 0.182 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.798 0.068 5.866 0.562 ;
        RECT 5.582 0.338 5.866 0.382 ;
        RECT 5.582 0.068 5.65 0.562 ;
      LAYER v0 ;
        RECT 5.582 0.448 5.65 0.492 ;
        RECT 5.582 0.138 5.65 0.182 ;
        RECT 5.798 0.448 5.866 0.492 ;
        RECT 5.798 0.138 5.866 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.974 0.652 ;
        RECT 5.69 0.428 5.758 0.652 ;
        RECT 5.474 0.518 5.542 0.652 ;
        RECT 5.258 0.428 5.326 0.652 ;
        RECT 4.934 0.428 5.002 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.098 0.338 3.166 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.466 0.25 0.51 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 1.154 0.518 1.222 0.562 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.586 0.4575 1.654 0.5015 ;
        RECT 2.342 0.538 2.41 0.582 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 3.098 0.428 3.166 0.472 ;
        RECT 4.072 0.538 4.136 0.582 ;
        RECT 4.934 0.448 5.002 0.492 ;
        RECT 5.258 0.448 5.326 0.492 ;
        RECT 5.476 0.538 5.54 0.582 ;
        RECT 5.69 0.448 5.758 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.974 0.022 ;
        RECT 5.69 -0.022 5.758 0.292 ;
        RECT 5.474 -0.022 5.542 0.202 ;
        RECT 5.042 -0.022 5.11 0.202 ;
        RECT 2.342 0.158 3.618 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.2005 0.25 0.2445 ;
        RECT 0.722 0.203 0.79 0.247 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.586 0.2245 1.654 0.2685 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.882 0.158 2.95 0.202 ;
        RECT 3.098 0.158 3.166 0.202 ;
        RECT 3.314 0.158 3.382 0.202 ;
        RECT 3.53 0.158 3.598 0.202 ;
        RECT 5.042 0.138 5.11 0.182 ;
        RECT 5.474 0.138 5.542 0.182 ;
        RECT 5.69 0.138 5.758 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 1.456 0.382 ;
      RECT 0.812 0.518 1.888 0.562 ;
      RECT 2 0.338 3.956 0.382 ;
      RECT 1.028 0.428 4.604 0.472 ;
      RECT 4.684 0.428 5.56 0.472 ;
    LAYER m1 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 0.83 0.068 0.898 0.562 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 3.53 0.248 3.598 0.472 ;
      RECT 2.666 0.428 2.734 0.562 ;
      RECT 3.854 0.338 3.922 0.472 ;
      RECT 3.962 0.338 4.158 0.382 ;
      RECT 3.726 0.158 4.158 0.202 ;
      RECT 4.394 0.338 4.462 0.562 ;
      RECT 2.342 0.248 2.41 0.472 ;
      RECT 4.502 0.338 4.57 0.562 ;
      RECT 2.558 0.068 4.826 0.112 ;
      RECT 5.042 0.248 5.11 0.382 ;
      RECT 5.042 0.428 5.11 0.562 ;
      RECT 5.15 0.338 5.218 0.562 ;
      RECT 5.366 0.158 5.434 0.562 ;
      RECT 5.474 0.248 5.542 0.472 ;
    LAYER v1 ;
      RECT 5.478 0.428 5.538 0.472 ;
      RECT 5.046 0.428 5.106 0.472 ;
      RECT 4.722 0.428 4.782 0.472 ;
      RECT 4.398 0.428 4.458 0.472 ;
      RECT 3.858 0.338 3.918 0.382 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.374 0.338 1.434 0.382 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 5.474 0.338 5.542 0.382 ;
      RECT 5.258 0.138 5.326 0.182 ;
      RECT 5.15 0.448 5.218 0.492 ;
      RECT 5.042 0.448 5.11 0.492 ;
      RECT 4.826 0.338 4.894 0.382 ;
      RECT 4.72 0.448 4.784 0.492 ;
      RECT 4.61 0.158 4.678 0.202 ;
      RECT 4.61 0.3675 4.678 0.4115 ;
      RECT 4.502 0.068 4.57 0.112 ;
      RECT 4.502 0.248 4.57 0.292 ;
      RECT 4.504 0.448 4.568 0.492 ;
      RECT 4.394 0.158 4.462 0.202 ;
      RECT 4.394 0.3675 4.462 0.4115 ;
      RECT 4.178 0.248 4.246 0.292 ;
      RECT 4.178 0.428 4.246 0.472 ;
      RECT 4.07 0.158 4.138 0.202 ;
      RECT 3.962 0.248 4.03 0.292 ;
      RECT 3.854 0.3835 3.922 0.4275 ;
      RECT 3.854 0.518 3.922 0.562 ;
      RECT 3.746 0.158 3.814 0.202 ;
      RECT 3.53 0.383 3.598 0.427 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 1.91 0.203 1.978 0.247 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.694 0.4575 1.762 0.5015 ;
      RECT 1.478 0.2245 1.546 0.2685 ;
      RECT 1.478 0.4575 1.546 0.5015 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.203 0.898 0.247 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.506 0.2075 0.574 0.2515 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 1.546 0.338 1.694 0.382 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 1.762 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.292 ;
      RECT 1.978 0.338 2.018 0.382 ;
      RECT 2.018 0.158 2.086 0.382 ;
      RECT 2.086 0.158 2.302 0.202 ;
      RECT 3.53 0.518 3.962 0.562 ;
      RECT 3.962 0.428 4.03 0.562 ;
      RECT 4.03 0.428 4.286 0.472 ;
      RECT 3.598 0.248 4.286 0.292 ;
      RECT 4.286 0.248 4.354 0.472 ;
      RECT 4.354 0.248 4.61 0.292 ;
      RECT 4.61 0.248 4.678 0.472 ;
      RECT 2.41 0.428 2.558 0.472 ;
      RECT 2.558 0.248 2.626 0.472 ;
      RECT 2.626 0.248 3.314 0.292 ;
      RECT 3.314 0.248 3.382 0.562 ;
      RECT 3.382 0.518 3.53 0.562 ;
      RECT 3.382 0.248 3.53 0.292 ;
      RECT 4.57 0.518 4.718 0.562 ;
      RECT 4.374 0.158 4.718 0.202 ;
      RECT 4.718 0.158 4.786 0.562 ;
      RECT 4.826 0.068 4.894 0.472 ;
      RECT 5.11 0.248 5.15 0.292 ;
      RECT 5.15 0.068 5.218 0.292 ;
      RECT 5.218 0.338 5.258 0.382 ;
      RECT 5.258 0.068 5.326 0.382 ;
  END
END b15fqy00fhn1n12x5

MACRO b15fqy00fhn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy00fhn1n16x5 0 0 ;
  SIZE 7.02 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAGATEAREA 0.0135 LAYER m2 ;
      ANTENNAMAXAREACAR 0.711746 LAYER m1 ;
      ANTENNAMAXAREACAR 5.072381 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.89396825 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAGATEAREA 0.0135 LAYER m2 ;
      ANTENNAMAXAREACAR 0.711746 LAYER m1 ;
      ANTENNAMAXAREACAR 5.072381 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.89396825 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 6.338 0.158 6.406 0.562 ;
        RECT 3.098 0.428 3.166 0.562 ;
      LAYER m2 ;
        RECT 3.08 0.518 6.424 0.562 ;
      LAYER v1 ;
        RECT 3.102 0.518 3.162 0.562 ;
        RECT 6.342 0.518 6.402 0.562 ;
      LAYER v0 ;
        RECT 3.098 0.49 3.166 0.534 ;
        RECT 6.338 0.248 6.406 0.292 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAGATEAREA 0.0279 LAYER m2 ;
      ANTENNAMAXAREACAR 2.49714275 LAYER m1 ;
      ANTENNAMAXAREACAR 6.640635 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.89396825 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0351 LAYER m2 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
      ANTENNAMAXAREACAR 7.7474075 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.906 0.248 6.082 0.292 ;
        RECT 6.014 0.068 6.082 0.292 ;
        RECT 5.906 0.248 5.974 0.382 ;
        RECT 4.718 0.338 4.914 0.382 ;
      LAYER m2 ;
        RECT 4.792 0.338 5.992 0.382 ;
      LAYER v1 ;
        RECT 4.83 0.338 4.89 0.382 ;
        RECT 5.91 0.338 5.97 0.382 ;
      LAYER v0 ;
        RECT 4.826 0.338 4.894 0.382 ;
        RECT 6.014 0.138 6.082 0.182 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 6.77 0.068 6.838 0.562 ;
        RECT 6.554 0.338 6.838 0.382 ;
        RECT 6.554 0.068 6.622 0.562 ;
      LAYER v0 ;
        RECT 6.554 0.448 6.622 0.492 ;
        RECT 6.554 0.138 6.622 0.182 ;
        RECT 6.77 0.448 6.838 0.492 ;
        RECT 6.77 0.138 6.838 0.182 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 8.6925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.8975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 7.054 0.652 ;
        RECT 6.878 0.428 6.946 0.652 ;
        RECT 6.662 0.428 6.73 0.652 ;
        RECT 6.446 0.518 6.514 0.652 ;
        RECT 6.122 0.428 6.19 0.652 ;
        RECT 5.798 0.428 5.866 0.652 ;
        RECT 5.042 0.518 5.11 0.652 ;
        RECT 4.826 0.518 4.894 0.652 ;
        RECT 3.746 0.338 3.814 0.652 ;
        RECT 3.53 0.338 3.598 0.652 ;
        RECT 3.314 0.338 3.382 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.472 0.25 0.516 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.37 0.518 1.438 0.562 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.802 0.4575 1.87 0.5015 ;
        RECT 2.776 0.538 2.84 0.582 ;
        RECT 3.314 0.403 3.382 0.447 ;
        RECT 3.53 0.428 3.598 0.472 ;
        RECT 3.746 0.428 3.814 0.472 ;
        RECT 4.828 0.538 4.892 0.582 ;
        RECT 5.044 0.538 5.108 0.582 ;
        RECT 5.798 0.448 5.866 0.492 ;
        RECT 6.122 0.448 6.19 0.492 ;
        RECT 6.448 0.538 6.512 0.582 ;
        RECT 6.662 0.448 6.73 0.492 ;
        RECT 6.878 0.448 6.946 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 7.054 0.022 ;
        RECT 6.878 -0.022 6.946 0.292 ;
        RECT 6.662 -0.022 6.73 0.292 ;
        RECT 6.446 -0.022 6.514 0.202 ;
        RECT 5.906 -0.022 5.974 0.202 ;
        RECT 2.558 0.158 4.482 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.938 -0.022 1.006 0.292 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.802 0.203 1.87 0.247 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.882 0.158 2.95 0.202 ;
        RECT 3.314 0.158 3.382 0.202 ;
        RECT 3.53 0.158 3.598 0.202 ;
        RECT 3.746 0.158 3.814 0.202 ;
        RECT 3.962 0.158 4.03 0.202 ;
        RECT 4.178 0.158 4.246 0.202 ;
        RECT 4.394 0.158 4.462 0.202 ;
        RECT 5.906 0.138 5.974 0.182 ;
        RECT 6.446 0.138 6.514 0.182 ;
        RECT 6.662 0.138 6.73 0.182 ;
        RECT 6.878 0.138 6.946 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.704 0.338 1.672 0.382 ;
      RECT 1.028 0.518 1.996 0.562 ;
      RECT 2.432 0.338 4.712 0.382 ;
      RECT 1.244 0.428 5.36 0.472 ;
      RECT 5.44 0.428 6.532 0.472 ;
    LAYER m1 ;
      RECT 1.694 0.158 1.762 0.562 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.91 0.428 1.978 0.562 ;
      RECT 2.234 0.248 2.302 0.472 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 4.178 0.338 4.246 0.562 ;
      RECT 2.558 0.338 2.626 0.562 ;
      RECT 3.098 0.428 3.166 0.562 ;
      RECT 4.61 0.338 4.678 0.472 ;
      RECT 4.718 0.338 4.914 0.382 ;
      RECT 4.59 0.158 5.13 0.202 ;
      RECT 5.15 0.338 5.218 0.562 ;
      RECT 2.666 0.248 2.734 0.472 ;
      RECT 5.366 0.338 5.434 0.562 ;
      RECT 2.754 0.068 5.69 0.112 ;
      RECT 5.906 0.248 5.974 0.382 ;
      RECT 5.906 0.428 5.974 0.562 ;
      RECT 6.014 0.338 6.082 0.562 ;
      RECT 6.338 0.158 6.406 0.562 ;
      RECT 6.446 0.248 6.514 0.472 ;
    LAYER v1 ;
      RECT 6.45 0.428 6.51 0.472 ;
      RECT 5.91 0.428 5.97 0.472 ;
      RECT 5.586 0.428 5.646 0.472 ;
      RECT 5.154 0.428 5.214 0.472 ;
      RECT 4.614 0.338 4.674 0.382 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.454 0.338 2.514 0.382 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 1.914 0.518 1.974 0.562 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 1.05 0.518 1.11 0.562 ;
      RECT 0.726 0.338 0.786 0.382 ;
    LAYER v0 ;
      RECT 6.446 0.338 6.514 0.382 ;
      RECT 6.23 0.448 6.298 0.492 ;
      RECT 6.122 0.138 6.19 0.182 ;
      RECT 6.014 0.448 6.082 0.492 ;
      RECT 5.906 0.448 5.974 0.492 ;
      RECT 5.69 0.338 5.758 0.382 ;
      RECT 5.584 0.448 5.648 0.492 ;
      RECT 5.474 0.158 5.542 0.202 ;
      RECT 5.474 0.3675 5.542 0.4115 ;
      RECT 5.366 0.248 5.434 0.292 ;
      RECT 5.368 0.448 5.432 0.492 ;
      RECT 5.258 0.158 5.326 0.202 ;
      RECT 5.258 0.3675 5.326 0.4115 ;
      RECT 5.15 0.068 5.218 0.112 ;
      RECT 5.15 0.448 5.218 0.492 ;
      RECT 5.042 0.158 5.11 0.202 ;
      RECT 4.934 0.248 5.002 0.292 ;
      RECT 4.934 0.428 5.002 0.472 ;
      RECT 4.826 0.158 4.894 0.202 ;
      RECT 4.718 0.248 4.786 0.292 ;
      RECT 4.61 0.158 4.678 0.202 ;
      RECT 4.61 0.3835 4.678 0.4275 ;
      RECT 4.61 0.518 4.678 0.562 ;
      RECT 4.394 0.383 4.462 0.427 ;
      RECT 4.178 0.428 4.246 0.472 ;
      RECT 3.962 0.428 4.03 0.472 ;
      RECT 2.774 0.068 2.842 0.112 ;
      RECT 2.666 0.293 2.734 0.337 ;
      RECT 2.558 0.383 2.626 0.427 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.45 0.479 2.518 0.523 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.293 2.302 0.337 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.203 2.086 0.247 ;
      RECT 1.91 0.4575 1.978 0.5015 ;
      RECT 1.694 0.203 1.762 0.247 ;
      RECT 1.694 0.4575 1.762 0.5015 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 1.762 0.338 2.126 0.382 ;
      RECT 2.126 0.158 2.194 0.562 ;
      RECT 2.194 0.158 2.41 0.202 ;
      RECT 2.086 0.068 2.45 0.112 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 4.178 0.248 4.394 0.292 ;
      RECT 4.394 0.248 4.462 0.472 ;
      RECT 4.246 0.518 4.718 0.562 ;
      RECT 4.718 0.428 4.786 0.562 ;
      RECT 4.786 0.428 5.042 0.472 ;
      RECT 4.462 0.248 5.042 0.292 ;
      RECT 5.042 0.248 5.11 0.472 ;
      RECT 5.11 0.248 5.258 0.292 ;
      RECT 5.258 0.248 5.326 0.562 ;
      RECT 5.326 0.248 5.474 0.292 ;
      RECT 5.474 0.248 5.542 0.472 ;
      RECT 2.734 0.428 2.882 0.472 ;
      RECT 2.882 0.248 2.95 0.472 ;
      RECT 2.95 0.248 3.962 0.292 ;
      RECT 3.962 0.248 4.03 0.562 ;
      RECT 4.03 0.518 4.178 0.562 ;
      RECT 4.03 0.248 4.178 0.292 ;
      RECT 5.434 0.518 5.582 0.562 ;
      RECT 5.238 0.158 5.582 0.202 ;
      RECT 5.582 0.158 5.65 0.562 ;
      RECT 5.69 0.068 5.758 0.472 ;
      RECT 5.974 0.248 6.014 0.292 ;
      RECT 6.014 0.068 6.082 0.292 ;
      RECT 6.082 0.338 6.122 0.382 ;
      RECT 6.122 0.068 6.19 0.382 ;
      RECT 6.19 0.338 6.23 0.382 ;
      RECT 6.23 0.338 6.298 0.562 ;
  END
END b15fqy00fhn1n16x5

MACRO b15fqy043hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy043hn1n02x5 0 0 ;
  SIZE 4.32 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.338 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.498 2.518 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 6.4125 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 6.4125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.338 3.706 0.562 ;
      LAYER v0 ;
        RECT 3.638 0.498 3.706 0.542 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 3.058 0.382 ;
        RECT 2.99 0.068 3.058 0.382 ;
      LAYER v0 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 2.882 0.338 2.95 0.382 ;
        RECT 2.99 0.088 3.058 0.132 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.182 0.203 0.25 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.81875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 4.655 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.088 0.574 0.132 ;
    END
  END rb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.248 4.246 0.472 ;
        RECT 4.05 0.248 4.246 0.292 ;
      LAYER v0 ;
        RECT 4.07 0.248 4.138 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.338 4.138 0.382 ;
        RECT 3.854 0.068 3.922 0.382 ;
        RECT 3.726 0.068 3.922 0.112 ;
      LAYER v0 ;
        RECT 3.746 0.068 3.814 0.112 ;
        RECT 3.962 0.338 4.03 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.354 0.652 ;
        RECT 4.07 0.428 4.138 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.566 0.428 1.762 0.472 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.5235 0.142 0.5675 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 2.342 0.403 2.41 0.447 ;
        RECT 2.774 0.472 2.842 0.516 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 4.07 0.448 4.138 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.354 0.022 ;
        RECT 4.07 -0.022 4.138 0.202 ;
        RECT 3.314 -0.022 3.382 0.292 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.0915 0.142 0.1355 ;
        RECT 0.398 0.198 0.466 0.242 ;
        RECT 1.478 0.048 1.546 0.092 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 3.314 0.2 3.382 0.244 ;
        RECT 4.07 0.114 4.138 0.158 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.068 2.536 0.112 ;
      RECT 2.864 0.068 3.508 0.112 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.614 0.068 0.682 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.782 0.158 1.91 0.202 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 0.702 0.518 0.938 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 2.45 0.068 2.646 0.112 ;
      RECT 2.97 0.428 3.098 0.472 ;
      RECT 3.422 0.068 3.49 0.292 ;
      RECT 3.53 0.068 3.598 0.202 ;
    LAYER v1 ;
      RECT 3.426 0.068 3.486 0.112 ;
      RECT 2.886 0.068 2.946 0.112 ;
      RECT 2.454 0.068 2.514 0.112 ;
      RECT 0.618 0.068 0.678 0.112 ;
      RECT 0.294 0.068 0.354 0.112 ;
    LAYER v0 ;
      RECT 3.854 0.428 3.922 0.472 ;
      RECT 3.746 0.2405 3.814 0.2845 ;
      RECT 3.53 0.088 3.598 0.132 ;
      RECT 3.532 0.408 3.596 0.452 ;
      RECT 3.422 0.2 3.49 0.244 ;
      RECT 3.098 0.205 3.166 0.249 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.234 0.403 2.302 0.447 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.018 0.178 2.086 0.222 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 1.046 0.498 1.114 0.542 ;
      RECT 0.938 0.33 1.006 0.374 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.4 0.358 0.464 0.402 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
    LAYER m1 ;
      RECT 0.398 0.338 0.466 0.472 ;
      RECT 0.466 0.428 0.83 0.472 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.114 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.338 1.674 0.382 ;
      RECT 1.91 0.158 1.978 0.472 ;
      RECT 0.79 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.438 0.158 1.586 0.202 ;
      RECT 1.586 0.068 1.654 0.202 ;
      RECT 1.654 0.068 2.214 0.112 ;
      RECT 0.938 0.248 1.006 0.562 ;
      RECT 1.006 0.248 1.802 0.292 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.87 0.518 2.234 0.562 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 2.086 0.248 2.882 0.292 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 3.098 0.158 3.166 0.472 ;
      RECT 3.166 0.338 3.53 0.382 ;
      RECT 3.53 0.338 3.598 0.472 ;
      RECT 3.598 0.158 3.746 0.202 ;
      RECT 3.746 0.158 3.814 0.472 ;
      RECT 3.814 0.428 3.942 0.472 ;
  END
END b15fqy043hn1n02x5

MACRO b15fqy043hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy043hn1n03x5 0 0 ;
  SIZE 4.428 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.498 2.626 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 6.4125 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 6.4125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.338 3.814 0.562 ;
      LAYER v0 ;
        RECT 3.746 0.498 3.814 0.542 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.338 3.166 0.382 ;
        RECT 3.098 0.068 3.166 0.382 ;
      LAYER v0 ;
        RECT 2.774 0.338 2.842 0.382 ;
        RECT 2.99 0.338 3.058 0.382 ;
        RECT 3.098 0.088 3.166 0.132 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.38875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.111 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END rb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.248 4.354 0.472 ;
        RECT 4.158 0.248 4.354 0.292 ;
      LAYER v0 ;
        RECT 4.178 0.248 4.246 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.338 4.246 0.382 ;
        RECT 3.962 0.068 4.03 0.382 ;
        RECT 3.834 0.068 4.03 0.112 ;
      LAYER v0 ;
        RECT 3.854 0.068 3.922 0.112 ;
        RECT 4.07 0.338 4.138 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.462 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.674 0.428 1.87 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 2.45 0.403 2.518 0.447 ;
        RECT 2.882 0.472 2.95 0.516 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 4.178 0.448 4.246 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.462 0.022 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.422 -0.022 3.49 0.292 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.198 0.574 0.242 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.422 0.2 3.49 0.244 ;
        RECT 4.178 0.114 4.246 0.158 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.068 2.644 0.112 ;
      RECT 2.972 0.068 3.616 0.112 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.89 0.158 2.018 0.202 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 0.81 0.518 1.046 0.562 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 2.558 0.068 2.754 0.112 ;
      RECT 3.078 0.428 3.206 0.472 ;
      RECT 3.53 0.068 3.598 0.292 ;
      RECT 3.638 0.068 3.706 0.202 ;
    LAYER v1 ;
      RECT 3.534 0.068 3.594 0.112 ;
      RECT 2.994 0.068 3.054 0.112 ;
      RECT 2.562 0.068 2.622 0.112 ;
      RECT 0.726 0.068 0.786 0.112 ;
      RECT 0.294 0.068 0.354 0.112 ;
    LAYER v0 ;
      RECT 3.962 0.428 4.03 0.472 ;
      RECT 3.854 0.2405 3.922 0.2845 ;
      RECT 3.638 0.088 3.706 0.132 ;
      RECT 3.64 0.408 3.704 0.452 ;
      RECT 3.53 0.2 3.598 0.244 ;
      RECT 3.206 0.205 3.274 0.249 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.342 0.403 2.41 0.447 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.126 0.178 2.194 0.222 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 1.046 0.33 1.114 0.374 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.508 0.358 0.572 0.402 ;
      RECT 0.29 0.203 0.358 0.247 ;
      RECT 0.29 0.3905 0.358 0.4345 ;
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 0.574 0.428 0.938 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.222 0.338 1.478 0.382 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.546 0.338 1.782 0.382 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 0.898 0.068 1.478 0.112 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 1.546 0.158 1.694 0.202 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.762 0.068 2.322 0.112 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.248 1.91 0.292 ;
      RECT 1.91 0.248 1.978 0.562 ;
      RECT 1.978 0.518 2.342 0.562 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.194 0.248 2.99 0.292 ;
      RECT 2.99 0.068 3.058 0.292 ;
      RECT 3.206 0.158 3.274 0.472 ;
      RECT 3.274 0.338 3.638 0.382 ;
      RECT 3.638 0.338 3.706 0.472 ;
      RECT 3.706 0.158 3.854 0.202 ;
      RECT 3.854 0.158 3.922 0.472 ;
      RECT 3.922 0.428 4.05 0.472 ;
  END
END b15fqy043hn1n03x5

MACRO b15fqy043hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy043hn1n04x5 0 0 ;
  SIZE 4.428 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.498 2.626 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 6.4125 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 6.4125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.338 3.814 0.562 ;
      LAYER v0 ;
        RECT 3.746 0.498 3.814 0.542 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.068 3.294 0.112 ;
        RECT 2.666 0.338 3.166 0.382 ;
        RECT 3.098 0.068 3.166 0.382 ;
      LAYER v0 ;
        RECT 2.774 0.338 2.842 0.382 ;
        RECT 2.99 0.338 3.058 0.382 ;
        RECT 3.206 0.068 3.274 0.112 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.25916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END rb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.248 4.354 0.472 ;
        RECT 4.158 0.248 4.354 0.292 ;
      LAYER v0 ;
        RECT 4.178 0.248 4.246 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.338 4.246 0.382 ;
        RECT 3.962 0.068 4.03 0.382 ;
        RECT 3.834 0.068 4.03 0.112 ;
      LAYER v0 ;
        RECT 3.854 0.068 3.922 0.112 ;
        RECT 4.07 0.338 4.138 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.462 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.674 0.428 1.87 0.472 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 2.45 0.403 2.518 0.447 ;
        RECT 2.882 0.472 2.95 0.516 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 4.178 0.448 4.246 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.462 0.022 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.422 -0.022 3.49 0.292 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.198 0.574 0.242 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.422 0.2 3.49 0.244 ;
        RECT 4.178 0.114 4.246 0.158 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.068 2.644 0.112 ;
      RECT 2.972 0.068 3.616 0.112 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.89 0.158 2.018 0.202 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 0.81 0.518 1.046 0.562 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 2.558 0.068 2.754 0.112 ;
      RECT 3.078 0.428 3.206 0.472 ;
      RECT 3.53 0.068 3.598 0.292 ;
      RECT 3.638 0.068 3.706 0.202 ;
    LAYER v1 ;
      RECT 3.534 0.068 3.594 0.112 ;
      RECT 2.994 0.068 3.054 0.112 ;
      RECT 2.562 0.068 2.622 0.112 ;
      RECT 0.726 0.068 0.786 0.112 ;
      RECT 0.294 0.068 0.354 0.112 ;
    LAYER v0 ;
      RECT 3.962 0.428 4.03 0.472 ;
      RECT 3.854 0.2405 3.922 0.2845 ;
      RECT 3.638 0.088 3.706 0.132 ;
      RECT 3.64 0.408 3.704 0.452 ;
      RECT 3.53 0.2 3.598 0.244 ;
      RECT 3.206 0.205 3.274 0.249 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.342 0.403 2.41 0.447 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.126 0.178 2.194 0.222 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 1.046 0.33 1.114 0.374 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.508 0.358 0.572 0.402 ;
      RECT 0.29 0.203 0.358 0.247 ;
      RECT 0.29 0.3905 0.358 0.4345 ;
    LAYER m1 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 0.574 0.428 0.938 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.222 0.338 1.478 0.382 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.546 0.338 1.782 0.382 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 0.898 0.068 1.478 0.112 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 1.546 0.158 1.694 0.202 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.762 0.068 2.322 0.112 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.248 1.91 0.292 ;
      RECT 1.91 0.248 1.978 0.562 ;
      RECT 1.978 0.518 2.342 0.562 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.194 0.248 2.99 0.292 ;
      RECT 2.99 0.068 3.058 0.292 ;
      RECT 3.206 0.158 3.274 0.472 ;
      RECT 3.274 0.338 3.638 0.382 ;
      RECT 3.638 0.338 3.706 0.472 ;
      RECT 3.706 0.158 3.854 0.202 ;
      RECT 3.854 0.158 3.922 0.472 ;
      RECT 3.922 0.428 4.05 0.472 ;
  END
END b15fqy043hn1n04x5

MACRO b15fqy043hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy043hn1n06x5 0 0 ;
  SIZE 4.752 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.338 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.498 2.95 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 5.13 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 5.13 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.338 4.138 0.562 ;
      LAYER v0 ;
        RECT 4.07 0.498 4.138 0.542 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.068 3.618 0.112 ;
        RECT 2.99 0.338 3.49 0.382 ;
        RECT 3.422 0.068 3.49 0.382 ;
      LAYER v0 ;
        RECT 3.098 0.338 3.166 0.382 ;
        RECT 3.314 0.338 3.382 0.382 ;
        RECT 3.53 0.068 3.598 0.112 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.182 0.203 0.25 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.63916675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 3.274706 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.088 0.574 0.132 ;
    END
  END rb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.61 0.248 4.678 0.472 ;
        RECT 4.482 0.248 4.678 0.292 ;
      LAYER v0 ;
        RECT 4.502 0.248 4.57 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.338 4.57 0.382 ;
        RECT 4.286 0.068 4.354 0.382 ;
        RECT 4.158 0.068 4.354 0.112 ;
      LAYER v0 ;
        RECT 4.178 0.068 4.246 0.112 ;
        RECT 4.394 0.338 4.462 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.786 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.29 0.3905 0.358 0.4345 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.774 0.403 2.842 0.447 ;
        RECT 3.206 0.472 3.274 0.516 ;
        RECT 3.746 0.448 3.814 0.492 ;
        RECT 4.502 0.448 4.57 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.786 0.022 ;
        RECT 4.502 -0.022 4.57 0.202 ;
        RECT 3.746 -0.022 3.814 0.292 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 1.566 0.158 2.086 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.29 0.203 0.358 0.247 ;
        RECT 0.614 0.178 0.682 0.222 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 3.206 0.138 3.274 0.182 ;
        RECT 3.746 0.2055 3.814 0.2495 ;
        RECT 4.502 0.114 4.57 0.158 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.068 2.968 0.112 ;
      RECT 3.296 0.068 3.94 0.112 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.35 0.338 1.89 0.382 ;
      RECT 2.214 0.158 2.342 0.202 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 2.45 0.158 2.518 0.472 ;
      RECT 2.882 0.068 3.078 0.112 ;
      RECT 3.402 0.428 3.53 0.472 ;
      RECT 3.854 0.068 3.922 0.292 ;
      RECT 3.962 0.068 4.03 0.202 ;
    LAYER v1 ;
      RECT 3.858 0.068 3.918 0.112 ;
      RECT 3.318 0.068 3.378 0.112 ;
      RECT 2.886 0.068 2.946 0.112 ;
      RECT 0.834 0.068 0.894 0.112 ;
      RECT 0.402 0.068 0.462 0.112 ;
    LAYER v0 ;
      RECT 4.286 0.428 4.354 0.472 ;
      RECT 4.178 0.2405 4.246 0.2845 ;
      RECT 3.962 0.088 4.03 0.132 ;
      RECT 3.964 0.408 4.028 0.452 ;
      RECT 3.854 0.2055 3.922 0.2495 ;
      RECT 3.53 0.2075 3.598 0.2515 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 2.99 0.068 3.058 0.112 ;
      RECT 2.666 0.403 2.734 0.447 ;
      RECT 2.45 0.178 2.518 0.222 ;
      RECT 2.45 0.408 2.518 0.452 ;
      RECT 2.342 0.408 2.41 0.452 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 1.154 0.498 1.222 0.542 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.616 0.358 0.68 0.402 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.3905 0.466 0.4345 ;
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.472 ;
      RECT 0.682 0.428 1.046 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.006 0.068 1.89 0.112 ;
      RECT 2.342 0.158 2.41 0.472 ;
      RECT 1.222 0.158 1.37 0.202 ;
      RECT 1.37 0.158 1.438 0.292 ;
      RECT 1.438 0.248 2.234 0.292 ;
      RECT 2.234 0.248 2.302 0.562 ;
      RECT 2.302 0.518 2.666 0.562 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.518 0.248 3.314 0.292 ;
      RECT 3.314 0.068 3.382 0.292 ;
      RECT 3.53 0.158 3.598 0.472 ;
      RECT 3.598 0.338 3.962 0.382 ;
      RECT 3.962 0.338 4.03 0.472 ;
      RECT 4.03 0.158 4.178 0.202 ;
      RECT 4.178 0.158 4.246 0.472 ;
      RECT 4.246 0.428 4.374 0.472 ;
  END
END b15fqy043hn1n06x5

MACRO b15fqy043hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy043hn1n08x5 0 0 ;
  SIZE 4.968 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.862 0.518 3.058 0.562 ;
        RECT 2.99 0.338 3.058 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.518 2.95 0.562 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 1.06158725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 1.06158725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.248 3.814 0.472 ;
      LAYER v0 ;
        RECT 3.746 0.338 3.814 0.382 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.726 0.112 ;
        RECT 3.53 0.068 3.598 0.472 ;
        RECT 3.314 0.248 3.598 0.292 ;
        RECT 3.314 0.248 3.382 0.472 ;
      LAYER v0 ;
        RECT 3.314 0.338 3.382 0.382 ;
        RECT 3.53 0.338 3.598 0.382 ;
        RECT 3.638 0.068 3.706 0.112 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.1995 0.25 0.2435 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 4.001875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 3.2015 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.113 0.574 0.157 ;
    END
  END rb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.826 0.248 4.894 0.472 ;
        RECT 4.61 0.248 4.894 0.292 ;
      LAYER v0 ;
        RECT 4.718 0.248 4.786 0.292 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 7.79 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.116 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.502 0.338 4.786 0.382 ;
        RECT 4.502 0.068 4.57 0.382 ;
        RECT 4.374 0.068 4.57 0.112 ;
      LAYER v0 ;
        RECT 4.394 0.068 4.462 0.112 ;
        RECT 4.61 0.338 4.678 0.382 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.002 0.652 ;
        RECT 4.718 0.428 4.786 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.234 0.472 2.302 0.516 ;
        RECT 3.098 0.453 3.166 0.497 ;
        RECT 3.422 0.472 3.49 0.516 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 4.718 0.448 4.786 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.002 0.022 ;
        RECT 4.718 -0.022 4.786 0.202 ;
        RECT 3.962 -0.022 4.03 0.292 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 1.154 0.158 2.322 0.202 ;
        RECT 0.83 0.338 1.222 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
        RECT 0.83 -0.022 0.898 0.382 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.0975 0.142 0.1415 ;
        RECT 0.29 0.0975 0.358 0.1415 ;
        RECT 0.614 0.113 0.682 0.157 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.99 0.088 3.058 0.132 ;
        RECT 3.422 0.138 3.49 0.182 ;
        RECT 3.962 0.181 4.03 0.225 ;
        RECT 4.718 0.114 4.786 0.158 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.068 3.2 0.112 ;
      RECT 3.28 0.068 4.172 0.112 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 2.43 0.158 2.558 0.202 ;
      RECT 0.918 0.518 1.37 0.562 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 2.774 0.158 2.842 0.292 ;
      RECT 3.098 0.068 3.166 0.202 ;
      RECT 3.638 0.158 3.706 0.562 ;
      RECT 4.07 0.068 4.138 0.292 ;
      RECT 4.178 0.068 4.246 0.382 ;
    LAYER v1 ;
      RECT 4.074 0.068 4.134 0.112 ;
      RECT 3.318 0.068 3.378 0.112 ;
      RECT 3.102 0.068 3.162 0.112 ;
      RECT 0.726 0.068 0.786 0.112 ;
      RECT 0.402 0.068 0.462 0.112 ;
    LAYER v0 ;
      RECT 4.502 0.428 4.57 0.472 ;
      RECT 4.394 0.23 4.462 0.274 ;
      RECT 4.286 0.498 4.354 0.542 ;
      RECT 4.178 0.088 4.246 0.132 ;
      RECT 4.07 0.181 4.138 0.225 ;
      RECT 3.746 0.158 3.814 0.202 ;
      RECT 3.64 0.448 3.704 0.492 ;
      RECT 3.098 0.088 3.166 0.132 ;
      RECT 2.776 0.178 2.84 0.222 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.666 0.3155 2.734 0.3595 ;
      RECT 2.558 0.408 2.626 0.452 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.342 0.248 2.41 0.292 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.37 0.3605 1.438 0.4045 ;
      RECT 1.262 0.268 1.33 0.312 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.938 0.228 1.006 0.272 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.616 0.358 0.68 0.402 ;
      RECT 0.398 0.206 0.466 0.25 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.472 ;
      RECT 0.682 0.428 1.262 0.472 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.546 0.338 1.694 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.762 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.978 0.338 2.322 0.382 ;
      RECT 2.558 0.158 2.626 0.472 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.438 0.248 2.45 0.292 ;
      RECT 2.45 0.248 2.518 0.562 ;
      RECT 2.518 0.518 2.666 0.562 ;
      RECT 2.666 0.248 2.734 0.562 ;
      RECT 1.006 0.068 2.842 0.112 ;
      RECT 2.842 0.248 3.206 0.292 ;
      RECT 3.206 0.068 3.274 0.292 ;
      RECT 3.274 0.068 3.382 0.112 ;
      RECT 3.706 0.158 3.834 0.202 ;
      RECT 3.706 0.518 3.854 0.562 ;
      RECT 3.854 0.428 3.922 0.562 ;
      RECT 3.922 0.428 4.286 0.472 ;
      RECT 4.286 0.428 4.354 0.562 ;
      RECT 4.246 0.338 4.394 0.382 ;
      RECT 4.394 0.158 4.462 0.472 ;
      RECT 4.462 0.428 4.59 0.472 ;
  END
END b15fqy043hn1n08x5

MACRO b15fqy043hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy043hn1n12x5 0 0 ;
  SIZE 5.508 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0117 LAYER m2 ;
      ANTENNAMAXAREACAR 9.19365075 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0126 LAYER m2 ;
      ANTENNAMAXAREACAR 8.3505555 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.518 4.246 0.562 ;
        RECT 4.178 0.158 4.246 0.562 ;
        RECT 3.962 0.248 4.03 0.562 ;
        RECT 3.53 0.518 3.814 0.562 ;
        RECT 3.746 0.338 3.814 0.562 ;
      LAYER m2 ;
        RECT 3.728 0.428 4.172 0.472 ;
      LAYER v1 ;
        RECT 3.75 0.428 3.81 0.472 ;
        RECT 3.966 0.428 4.026 0.472 ;
      LAYER v0 ;
        RECT 3.638 0.518 3.706 0.562 ;
        RECT 3.962 0.293 4.03 0.337 ;
        RECT 4.178 0.248 4.246 0.292 ;
    END
  END den
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0207 LAYER m2 ;
      ANTENNAMAXAREACAR 2.82185175 LAYER m1 ;
      ANTENNAMAXAREACAR 4.418889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0279 LAYER m2 ;
      ANTENNAMAXAREACAR 2.82185175 LAYER m1 ;
      ANTENNAMAXAREACAR 4.418889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.428 2.43 0.472 ;
        RECT 0.594 0.428 0.79 0.472 ;
      LAYER m2 ;
        RECT 0.596 0.428 2.32 0.472 ;
      LAYER v1 ;
        RECT 0.618 0.428 0.678 0.472 ;
        RECT 2.238 0.428 2.298 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 2.342 0.428 2.41 0.472 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.158 3.49 0.382 ;
      LAYER v0 ;
        RECT 3.422 0.248 3.49 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.248 4.354 0.472 ;
      LAYER v0 ;
        RECT 4.286 0.338 4.354 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.562 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.1995 0.142 0.2435 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.29 0.1995 0.358 0.2435 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.15 0.248 5.218 0.472 ;
      LAYER v0 ;
        RECT 5.15 0.383 5.218 0.427 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.97916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.366 0.068 5.434 0.202 ;
      LAYER v0 ;
        RECT 5.366 0.088 5.434 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.542 0.652 ;
        RECT 5.258 0.518 5.326 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 4.394 0.518 4.462 0.652 ;
        RECT 3.854 0.338 3.922 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.83 0.338 0.898 0.472 ;
        RECT 0.398 0.338 0.898 0.382 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.832 0.408 0.896 0.452 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.666 0.538 2.734 0.582 ;
        RECT 3.422 0.538 3.49 0.582 ;
        RECT 3.854 0.4265 3.922 0.4705 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 4.612 0.538 4.676 0.582 ;
        RECT 5.26 0.538 5.324 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.542 0.022 ;
        RECT 5.258 -0.022 5.326 0.292 ;
        RECT 4.61 -0.022 4.678 0.202 ;
        RECT 4.394 -0.022 4.462 0.112 ;
        RECT 3.854 -0.022 3.922 0.112 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 1.782 0.158 2.842 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.0975 0.25 0.1415 ;
        RECT 0.398 0.0975 0.466 0.1415 ;
        RECT 0.722 0.113 0.79 0.157 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.856 0.048 3.92 0.092 ;
        RECT 4.396 0.048 4.46 0.092 ;
        RECT 4.61 0.133 4.678 0.177 ;
        RECT 5.258 0.183 5.326 0.227 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 2.864 0.428 3.292 0.472 ;
      RECT 0.488 0.068 3.848 0.112 ;
      RECT 3.928 0.068 4.588 0.112 ;
      RECT 4.252 0.428 4.928 0.472 ;
      RECT 5.008 0.428 5.468 0.472 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.594 0.428 0.79 0.472 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 2.234 0.428 2.43 0.472 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 2.322 0.518 2.558 0.562 ;
      RECT 3.53 0.518 3.746 0.562 ;
      RECT 3.206 0.428 3.274 0.562 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 3.746 0.068 3.814 0.202 ;
      RECT 3.962 0.248 4.03 0.562 ;
      RECT 4.07 0.068 4.138 0.472 ;
      RECT 4.718 0.338 4.786 0.562 ;
      RECT 4.502 0.068 4.57 0.562 ;
      RECT 4.826 0.338 4.894 0.472 ;
      RECT 4.718 0.158 4.786 0.292 ;
      RECT 5.366 0.248 5.434 0.562 ;
    LAYER v1 ;
      RECT 5.37 0.428 5.43 0.472 ;
      RECT 5.046 0.428 5.106 0.472 ;
      RECT 4.83 0.428 4.89 0.472 ;
      RECT 4.506 0.068 4.566 0.112 ;
      RECT 4.398 0.428 4.458 0.472 ;
      RECT 3.966 0.068 4.026 0.112 ;
      RECT 3.75 0.068 3.81 0.112 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 0.942 0.068 1.002 0.112 ;
      RECT 0.51 0.068 0.57 0.112 ;
    LAYER v0 ;
      RECT 5.366 0.293 5.434 0.337 ;
      RECT 5.042 0.158 5.11 0.202 ;
      RECT 5.042 0.293 5.11 0.337 ;
      RECT 4.934 0.408 5.002 0.452 ;
      RECT 4.826 0.408 4.894 0.452 ;
      RECT 4.718 0.408 4.786 0.452 ;
      RECT 4.72 0.228 4.784 0.272 ;
      RECT 4.502 0.133 4.57 0.177 ;
      RECT 4.502 0.453 4.57 0.497 ;
      RECT 4.178 0.068 4.246 0.112 ;
      RECT 4.07 0.3985 4.138 0.4425 ;
      RECT 3.746 0.138 3.814 0.182 ;
      RECT 3.206 0.473 3.274 0.517 ;
      RECT 3.098 0.473 3.166 0.517 ;
      RECT 2.99 0.338 3.058 0.382 ;
      RECT 2.882 0.338 2.95 0.382 ;
      RECT 2.884 0.138 2.948 0.182 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.342 0.518 2.41 0.562 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.408 1.438 0.452 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 1.048 0.138 1.112 0.182 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.206 0.574 0.25 ;
    LAYER m1 ;
      RECT 0.702 0.518 1.046 0.562 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.114 0.248 1.262 0.292 ;
      RECT 1.262 0.158 1.33 0.472 ;
      RECT 1.33 0.158 1.458 0.202 ;
      RECT 1.114 0.068 2.538 0.112 ;
      RECT 1.222 0.518 1.478 0.562 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.546 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.338 2.754 0.382 ;
      RECT 1.438 0.248 2.882 0.292 ;
      RECT 2.882 0.248 2.95 0.472 ;
      RECT 2.558 0.428 2.626 0.562 ;
      RECT 2.626 0.428 2.774 0.472 ;
      RECT 2.774 0.428 2.842 0.562 ;
      RECT 2.882 0.068 2.95 0.202 ;
      RECT 2.842 0.518 2.99 0.562 ;
      RECT 2.99 0.248 3.058 0.562 ;
      RECT 3.058 0.248 3.098 0.292 ;
      RECT 2.95 0.068 3.098 0.112 ;
      RECT 3.098 0.068 3.166 0.292 ;
      RECT 3.746 0.338 3.814 0.562 ;
      RECT 3.166 0.338 3.314 0.382 ;
      RECT 3.314 0.338 3.382 0.472 ;
      RECT 3.382 0.428 3.638 0.472 ;
      RECT 3.638 0.248 3.706 0.472 ;
      RECT 3.706 0.248 3.854 0.292 ;
      RECT 3.854 0.158 3.922 0.292 ;
      RECT 3.922 0.158 3.962 0.202 ;
      RECT 3.962 0.068 4.03 0.202 ;
      RECT 4.03 0.518 4.178 0.562 ;
      RECT 4.178 0.158 4.246 0.562 ;
      RECT 4.138 0.068 4.286 0.112 ;
      RECT 4.286 0.068 4.354 0.202 ;
      RECT 4.354 0.158 4.394 0.202 ;
      RECT 4.394 0.158 4.462 0.472 ;
      RECT 4.786 0.518 5.042 0.562 ;
      RECT 5.042 0.248 5.11 0.562 ;
      RECT 4.786 0.158 4.934 0.202 ;
      RECT 4.934 0.158 5.002 0.472 ;
      RECT 5.002 0.158 5.218 0.202 ;
  END
END b15fqy043hn1n12x5

MACRO b15fqy043hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy043hn1n16x5 0 0 ;
  SIZE 6.588 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.027 LAYER m2 ;
      ANTENNAMAXAREACAR 4.81333325 LAYER m1 ;
      ANTENNAMAXAREACAR 6.41037025 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0342 LAYER m2 ;
      ANTENNAMAXAREACAR 4.81333325 LAYER m1 ;
      ANTENNAMAXAREACAR 6.41037025 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.428 2.862 0.472 ;
        RECT 0.702 0.428 0.898 0.472 ;
      LAYER m2 ;
        RECT 0.704 0.428 2.752 0.472 ;
      LAYER v1 ;
        RECT 0.726 0.428 0.786 0.472 ;
        RECT 2.67 0.428 2.73 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 2.774 0.428 2.842 0.472 ;
    END
  END rb
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 1.83901225 LAYER m1 ;
      ANTENNAMAXAREACAR 4.55506175 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.69530875 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 1.655111 LAYER m1 ;
      ANTENNAMAXAREACAR 3.182889 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.7374075 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 6.446 0.068 6.514 0.382 ;
        RECT 5.798 0.068 6.298 0.112 ;
      LAYER m2 ;
        RECT 5.872 0.068 6.548 0.112 ;
      LAYER v1 ;
        RECT 5.91 0.068 5.97 0.112 ;
        RECT 6.45 0.068 6.51 0.112 ;
      LAYER v0 ;
        RECT 5.906 0.068 5.974 0.112 ;
        RECT 6.122 0.068 6.19 0.112 ;
    END
  END ssb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.158 4.03 0.382 ;
      LAYER v0 ;
        RECT 3.962 0.293 4.03 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.856508 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.856508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.258 0.248 5.454 0.292 ;
        RECT 5.258 0.068 5.326 0.292 ;
      LAYER v0 ;
        RECT 5.366 0.248 5.434 0.292 ;
    END
  END d
  PIN den
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 3.54666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 3.54666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.826 0.158 4.894 0.382 ;
        RECT 4.61 0.158 4.894 0.202 ;
        RECT 4.178 0.338 4.678 0.382 ;
        RECT 4.61 0.158 4.678 0.382 ;
      LAYER v0 ;
        RECT 4.286 0.338 4.354 0.382 ;
        RECT 4.502 0.338 4.57 0.382 ;
        RECT 4.826 0.248 4.894 0.292 ;
    END
  END den
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.1995 0.25 0.2435 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.1995 0.466 0.2435 ;
    END
  END o
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 6.23 0.248 6.298 0.472 ;
      LAYER v0 ;
        RECT 6.23 0.383 6.298 0.427 ;
    END
  END si
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.622 0.652 ;
        RECT 6.338 0.518 6.406 0.652 ;
        RECT 5.582 0.518 5.65 0.652 ;
        RECT 5.366 0.518 5.434 0.652 ;
        RECT 5.15 0.428 5.218 0.652 ;
        RECT 4.394 0.518 4.462 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 0.938 0.338 1.006 0.472 ;
        RECT 0.506 0.338 1.006 0.382 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.94 0.408 1.004 0.452 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.962 0.4795 4.03 0.5235 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 5.15 0.448 5.218 0.492 ;
        RECT 5.368 0.538 5.432 0.582 ;
        RECT 5.584 0.538 5.648 0.582 ;
        RECT 6.34 0.538 6.404 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.622 0.022 ;
        RECT 6.338 -0.022 6.406 0.292 ;
        RECT 5.582 -0.022 5.65 0.112 ;
        RECT 5.366 -0.022 5.434 0.112 ;
        RECT 5.15 -0.022 5.218 0.202 ;
        RECT 4.394 -0.022 4.462 0.202 ;
        RECT 4.07 -0.022 4.138 0.112 ;
        RECT 1.998 0.158 3.166 0.202 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.0975 0.142 0.1415 ;
        RECT 0.29 0.0975 0.358 0.1415 ;
        RECT 0.506 0.0975 0.574 0.1415 ;
        RECT 0.83 0.113 0.898 0.157 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 4.07 0.048 4.138 0.092 ;
        RECT 4.394 0.092 4.462 0.136 ;
        RECT 5.15 0.138 5.218 0.182 ;
        RECT 5.368 0.048 5.432 0.092 ;
        RECT 5.584 0.048 5.648 0.092 ;
        RECT 6.338 0.183 6.406 0.227 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.596 0.068 4.372 0.112 ;
      RECT 3.62 0.428 5.576 0.472 ;
      RECT 4.916 0.068 5.792 0.112 ;
      RECT 5.656 0.428 6.548 0.472 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.702 0.428 0.898 0.472 ;
      RECT 0.81 0.518 1.046 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 2.666 0.428 2.862 0.472 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.458 0.428 1.586 0.472 ;
      RECT 3.51 0.428 3.746 0.472 ;
      RECT 2.754 0.518 2.99 0.562 ;
      RECT 4.286 0.068 4.354 0.292 ;
      RECT 4.158 0.428 4.718 0.472 ;
      RECT 4.59 0.518 4.826 0.562 ;
      RECT 5.366 0.428 5.582 0.472 ;
      RECT 5.69 0.068 5.758 0.292 ;
      RECT 5.69 0.338 5.758 0.562 ;
      RECT 5.798 0.338 5.866 0.562 ;
      RECT 6.122 0.248 6.19 0.472 ;
      RECT 5.798 0.068 6.298 0.112 ;
      RECT 6.446 0.068 6.514 0.382 ;
      RECT 6.338 0.428 6.534 0.472 ;
    LAYER v1 ;
      RECT 6.342 0.428 6.402 0.472 ;
      RECT 6.126 0.428 6.186 0.472 ;
      RECT 5.694 0.068 5.754 0.112 ;
      RECT 5.694 0.428 5.754 0.472 ;
      RECT 5.478 0.428 5.538 0.472 ;
      RECT 4.938 0.068 4.998 0.112 ;
      RECT 4.29 0.068 4.35 0.112 ;
      RECT 3.642 0.428 3.702 0.472 ;
      RECT 1.05 0.068 1.11 0.112 ;
      RECT 0.618 0.068 0.678 0.112 ;
    LAYER v0 ;
      RECT 6.446 0.428 6.514 0.472 ;
      RECT 6.122 0.158 6.19 0.202 ;
      RECT 6.122 0.293 6.19 0.337 ;
      RECT 6.016 0.448 6.08 0.492 ;
      RECT 5.906 0.3375 5.974 0.3815 ;
      RECT 5.798 0.4285 5.866 0.4725 ;
      RECT 5.69 0.4285 5.758 0.4725 ;
      RECT 5.474 0.158 5.542 0.202 ;
      RECT 5.474 0.428 5.542 0.472 ;
      RECT 4.934 0.1525 5.002 0.1965 ;
      RECT 4.828 0.448 4.892 0.492 ;
      RECT 4.718 0.068 4.786 0.112 ;
      RECT 4.718 0.338 4.786 0.382 ;
      RECT 4.61 0.518 4.678 0.562 ;
      RECT 4.394 0.248 4.462 0.292 ;
      RECT 4.178 0.428 4.246 0.472 ;
      RECT 3.638 0.518 3.706 0.562 ;
      RECT 3.53 0.158 3.598 0.202 ;
      RECT 3.53 0.338 3.598 0.382 ;
      RECT 3.53 0.428 3.598 0.472 ;
      RECT 3.422 0.248 3.49 0.292 ;
      RECT 3.422 0.518 3.49 0.562 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.314 0.338 3.382 0.382 ;
      RECT 2.99 0.338 3.058 0.382 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.882 0.248 2.95 0.292 ;
      RECT 2.774 0.518 2.842 0.562 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.45 0.448 2.518 0.492 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.264 0.448 1.328 0.492 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.206 0.682 0.25 ;
    LAYER m1 ;
      RECT 0.83 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.114 0.338 1.478 0.382 ;
      RECT 1.262 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.546 0.158 1.782 0.202 ;
      RECT 1.222 0.248 1.35 0.292 ;
      RECT 1.222 0.068 2.97 0.112 ;
      RECT 1.33 0.518 1.694 0.562 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.762 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.086 0.338 2.45 0.382 ;
      RECT 2.45 0.338 2.518 0.562 ;
      RECT 2.518 0.338 3.078 0.382 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.654 0.248 3.206 0.292 ;
      RECT 3.206 0.248 3.274 0.382 ;
      RECT 3.274 0.338 3.618 0.382 ;
      RECT 3.402 0.248 3.746 0.292 ;
      RECT 3.746 0.248 3.814 0.472 ;
      RECT 2.99 0.428 3.058 0.562 ;
      RECT 3.058 0.428 3.314 0.472 ;
      RECT 3.314 0.428 3.382 0.562 ;
      RECT 3.382 0.518 3.854 0.562 ;
      RECT 3.206 0.158 3.854 0.202 ;
      RECT 3.854 0.158 3.922 0.562 ;
      RECT 4.354 0.248 4.482 0.292 ;
      RECT 4.718 0.248 4.786 0.472 ;
      RECT 4.826 0.428 4.894 0.562 ;
      RECT 4.698 0.068 4.934 0.112 ;
      RECT 4.934 0.068 5.002 0.292 ;
      RECT 4.894 0.518 5.042 0.562 ;
      RECT 5.002 0.248 5.042 0.292 ;
      RECT 5.042 0.248 5.11 0.562 ;
      RECT 5.366 0.158 5.582 0.202 ;
      RECT 5.582 0.158 5.65 0.472 ;
      RECT 5.758 0.248 5.906 0.292 ;
      RECT 5.906 0.248 5.974 0.472 ;
      RECT 5.866 0.518 6.014 0.562 ;
      RECT 6.014 0.158 6.082 0.562 ;
      RECT 6.082 0.158 6.298 0.202 ;
  END
END b15fqy043hn1n16x5

MACRO b15fqy08fhn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy08fhn1n02x5 0 0 ;
  SIZE 3.888 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 5.32 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 5.32 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.518 0.292 ;
      LAYER v0 ;
        RECT 2.45 0.228 2.518 0.272 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.248 3.274 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.338 3.274 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.4 0.142 0.444 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.15375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.15375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.398 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.496 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.654 0.202 ;
        RECT 1.046 0.068 1.114 0.202 ;
        RECT 0.83 0.068 1.114 0.112 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END rb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.598 0.292 ;
      LAYER v0 ;
        RECT 3.53 0.088 3.598 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.976 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.338 3.814 0.382 ;
        RECT 3.746 0.068 3.814 0.382 ;
        RECT 3.422 0.068 3.49 0.382 ;
      LAYER v0 ;
        RECT 3.422 0.088 3.49 0.132 ;
        RECT 3.53 0.338 3.598 0.382 ;
        RECT 3.746 0.088 3.814 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.922 0.652 ;
        RECT 3.638 0.428 3.706 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.383 0.466 0.427 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.234 0.358 2.302 0.402 ;
        RECT 2.558 0.473 2.626 0.517 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.638 0.448 3.706 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.922 0.022 ;
        RECT 3.638 -0.022 3.706 0.292 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.694 0.158 2.41 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 3.098 0.048 3.166 0.092 ;
        RECT 3.638 0.2025 3.706 0.2465 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.428 1.148 0.472 ;
      RECT 1.228 0.428 2.984 0.472 ;
      RECT 3.064 0.428 3.4 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 1.046 0.338 1.262 0.382 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.91 0.338 2.126 0.382 ;
      RECT 1.586 0.248 2.086 0.292 ;
      RECT 2.126 0.428 2.194 0.562 ;
      RECT 1.242 0.068 2.302 0.112 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 3.314 0.158 3.382 0.472 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.098 0.158 3.166 0.472 ;
    LAYER v1 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 2.67 0.428 2.73 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.186 0.428 0.246 0.472 ;
    LAYER v0 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 3.314 0.203 3.382 0.247 ;
      RECT 3.098 0.248 3.166 0.292 ;
      RECT 2.99 0.1575 3.058 0.2015 ;
      RECT 2.99 0.4575 3.058 0.5015 ;
      RECT 2.882 0.1575 2.95 0.2015 ;
      RECT 2.882 0.358 2.95 0.402 ;
      RECT 2.774 0.472 2.842 0.516 ;
      RECT 2.666 0.383 2.734 0.427 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.182 0.293 0.25 0.337 ;
    LAYER m1 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.358 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.574 0.338 0.938 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.114 0.518 1.37 0.562 ;
      RECT 1.154 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 2.086 0.562 ;
      RECT 2.126 0.248 2.194 0.382 ;
      RECT 2.194 0.248 2.342 0.292 ;
      RECT 2.342 0.248 2.41 0.382 ;
      RECT 2.41 0.338 2.558 0.382 ;
      RECT 2.558 0.248 2.626 0.382 ;
      RECT 2.626 0.248 2.774 0.292 ;
      RECT 2.774 0.248 2.842 0.562 ;
      RECT 2.842 0.248 2.882 0.292 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 3.382 0.428 3.51 0.472 ;
  END
END b15fqy08fhn1n02x5

MACRO b15fqy08fhn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy08fhn1n04x5 0 0 ;
  SIZE 3.888 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 5.32 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 5.32 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.518 0.292 ;
      LAYER v0 ;
        RECT 2.45 0.228 2.518 0.272 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.248 3.274 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.338 3.274 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.4 0.142 0.444 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 4.123 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 4.123 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.398 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 2.49714275 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.566 0.202 ;
        RECT 1.046 0.068 1.114 0.202 ;
        RECT 0.83 0.068 1.114 0.112 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END rb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.598 0.292 ;
      LAYER v0 ;
        RECT 3.53 0.088 3.598 0.132 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.976 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.338 3.814 0.382 ;
        RECT 3.746 0.068 3.814 0.382 ;
        RECT 3.422 0.068 3.49 0.382 ;
      LAYER v0 ;
        RECT 3.422 0.088 3.49 0.132 ;
        RECT 3.53 0.338 3.598 0.382 ;
        RECT 3.746 0.088 3.814 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.922 0.652 ;
        RECT 3.638 0.428 3.706 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.383 0.466 0.427 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 2.234 0.358 2.302 0.402 ;
        RECT 2.558 0.473 2.626 0.517 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.638 0.448 3.706 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.922 0.022 ;
        RECT 3.638 -0.022 3.706 0.292 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.782 0.158 2.41 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 3.098 0.048 3.166 0.092 ;
        RECT 3.638 0.2025 3.706 0.2465 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.428 1.148 0.472 ;
      RECT 1.228 0.428 2.984 0.472 ;
      RECT 3.064 0.428 3.4 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 1.046 0.338 1.262 0.382 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.91 0.338 2.126 0.382 ;
      RECT 1.674 0.248 1.998 0.292 ;
      RECT 2.126 0.428 2.194 0.562 ;
      RECT 1.242 0.068 2.214 0.112 ;
      RECT 2.666 0.338 2.734 0.562 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 3.314 0.158 3.382 0.472 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.098 0.158 3.166 0.472 ;
    LAYER v1 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 3.102 0.428 3.162 0.472 ;
      RECT 2.886 0.428 2.946 0.472 ;
      RECT 2.67 0.428 2.73 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.186 0.428 0.246 0.472 ;
    LAYER v0 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 3.314 0.203 3.382 0.247 ;
      RECT 3.098 0.248 3.166 0.292 ;
      RECT 2.99 0.1575 3.058 0.2015 ;
      RECT 2.99 0.4575 3.058 0.5015 ;
      RECT 2.882 0.1575 2.95 0.2015 ;
      RECT 2.882 0.358 2.95 0.402 ;
      RECT 2.774 0.472 2.842 0.516 ;
      RECT 2.666 0.383 2.734 0.427 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.506 0.498 0.574 0.542 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.182 0.293 0.25 0.337 ;
    LAYER m1 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.358 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.574 0.338 0.938 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.114 0.518 1.37 0.562 ;
      RECT 1.242 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 1.998 0.562 ;
      RECT 2.126 0.248 2.194 0.382 ;
      RECT 2.194 0.248 2.342 0.292 ;
      RECT 2.342 0.248 2.41 0.382 ;
      RECT 2.41 0.338 2.558 0.382 ;
      RECT 2.558 0.248 2.626 0.382 ;
      RECT 2.626 0.248 2.774 0.292 ;
      RECT 2.774 0.248 2.842 0.562 ;
      RECT 2.842 0.248 2.882 0.292 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 3.382 0.428 3.51 0.472 ;
  END
END b15fqy08fhn1n04x5

MACRO b15fqy08fhn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy08fhn1n08x5 0 0 ;
  SIZE 4.86 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.158 3.274 0.382 ;
        RECT 2.99 0.248 3.274 0.292 ;
      LAYER v0 ;
        RECT 3.098 0.248 3.166 0.292 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.248 4.246 0.562 ;
      LAYER v0 ;
        RECT 4.178 0.338 4.246 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.4 0.25 0.444 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 4.123 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 4.123 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.614 0.068 0.682 0.112 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.59916675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 1.199375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 2.214 0.112 ;
        RECT 0.938 0.068 1.006 0.292 ;
      LAYER v0 ;
        RECT 1.046 0.068 1.114 0.112 ;
        RECT 2.126 0.068 2.194 0.112 ;
    END
  END rb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.502 0.068 4.57 0.292 ;
      LAYER v0 ;
        RECT 4.502 0.113 4.57 0.157 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.338 4.786 0.382 ;
        RECT 4.718 0.068 4.786 0.382 ;
        RECT 4.394 0.068 4.462 0.382 ;
        RECT 4.266 0.068 4.462 0.112 ;
      LAYER v0 ;
        RECT 4.286 0.068 4.354 0.112 ;
        RECT 4.502 0.338 4.57 0.382 ;
        RECT 4.718 0.113 4.786 0.157 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.894 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.493 0.142 0.537 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.383 0.574 0.427 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 4.072 0.538 4.136 0.582 ;
        RECT 4.61 0.448 4.678 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.894 0.022 ;
        RECT 4.61 -0.022 4.678 0.292 ;
        RECT 4.07 -0.022 4.138 0.112 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.99 0.048 3.058 0.092 ;
        RECT 3.422 0.138 3.49 0.182 ;
        RECT 4.072 0.048 4.136 0.092 ;
        RECT 4.61 0.2025 4.678 0.2465 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.428 1.24 0.472 ;
      RECT 1.784 0.428 2.66 0.472 ;
      RECT 2.74 0.428 3.848 0.472 ;
      RECT 3.928 0.428 4.372 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 2.558 0.428 2.626 0.562 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 1.89 0.158 2.754 0.202 ;
      RECT 1.458 0.338 3.098 0.382 ;
      RECT 2.666 0.428 2.862 0.472 ;
      RECT 3.638 0.338 3.706 0.562 ;
      RECT 1.262 0.248 2.882 0.292 ;
      RECT 4.286 0.158 4.354 0.472 ;
      RECT 3.962 0.068 4.03 0.562 ;
      RECT 4.07 0.158 4.138 0.472 ;
    LAYER v1 ;
      RECT 4.29 0.428 4.35 0.472 ;
      RECT 4.074 0.428 4.134 0.472 ;
      RECT 3.642 0.428 3.702 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.158 0.428 1.218 0.472 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.294 0.428 0.354 0.472 ;
    LAYER v0 ;
      RECT 4.394 0.428 4.462 0.472 ;
      RECT 4.286 0.203 4.354 0.247 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 3.962 0.1575 4.03 0.2015 ;
      RECT 3.962 0.4575 4.03 0.5015 ;
      RECT 3.854 0.338 3.922 0.382 ;
      RECT 3.746 0.178 3.814 0.222 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.53 0.338 3.598 0.382 ;
      RECT 3.314 0.333 3.382 0.377 ;
      RECT 3.098 0.448 3.166 0.492 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.774 0.518 2.842 0.562 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.56 0.448 2.624 0.492 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.448 1.87 0.492 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.588 0.448 1.652 0.492 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.614 0.498 0.682 0.542 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.29 0.293 0.358 0.337 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.158 0.574 0.292 ;
      RECT 0.574 0.248 0.614 0.292 ;
      RECT 0.614 0.248 0.682 0.382 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.158 1.114 0.382 ;
      RECT 1.222 0.158 1.458 0.202 ;
      RECT 1.222 0.518 1.586 0.562 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 2.626 0.518 2.862 0.562 ;
      RECT 3.098 0.338 3.166 0.562 ;
      RECT 3.706 0.338 3.746 0.382 ;
      RECT 3.746 0.158 3.814 0.382 ;
      RECT 2.882 0.158 2.95 0.292 ;
      RECT 2.95 0.158 3.098 0.202 ;
      RECT 3.098 0.068 3.166 0.202 ;
      RECT 3.166 0.068 3.314 0.112 ;
      RECT 3.314 0.068 3.382 0.472 ;
      RECT 3.382 0.248 3.53 0.292 ;
      RECT 3.53 0.068 3.598 0.472 ;
      RECT 3.598 0.068 3.854 0.112 ;
      RECT 3.854 0.068 3.922 0.472 ;
      RECT 4.354 0.428 4.482 0.472 ;
  END
END b15fqy08fhn1n08x5

MACRO b15fqy08fhn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy08fhn1n16x5 0 0 ;
  SIZE 6.588 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.158 4.462 0.382 ;
        RECT 4.158 0.248 4.462 0.292 ;
      LAYER v0 ;
        RECT 4.178 0.248 4.246 0.292 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.798 0.158 5.866 0.382 ;
      LAYER v0 ;
        RECT 5.798 0.293 5.866 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.408 0.466 0.452 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0135 LAYER m1 ;
      ANTENNAMAXAREACAR 5.4014285 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0135 LAYER m1 ;
      ANTENNAMAXAREACAR 2.52066675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.3155 0.898 0.3595 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.027 LAYER m1 ;
      ANTENNAMAXAREACAR 3.04 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0342 LAYER m1 ;
      ANTENNAMAXAREACAR 3.04 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 2.322 0.112 ;
        RECT 1.37 0.068 1.438 0.292 ;
      LAYER v0 ;
        RECT 1.478 0.068 1.546 0.112 ;
        RECT 2.234 0.068 2.302 0.112 ;
    END
  END rb
  PIN si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 6.23 0.158 6.298 0.382 ;
      LAYER v0 ;
        RECT 6.23 0.293 6.298 0.337 ;
    END
  END si
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 8.2175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.73916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 6.122 0.068 6.19 0.382 ;
      LAYER v0 ;
        RECT 6.122 0.293 6.19 0.337 ;
        RECT 6.122 0.088 6.19 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.622 0.652 ;
        RECT 6.338 0.338 6.406 0.652 ;
        RECT 5.69 0.428 5.758 0.652 ;
        RECT 5.474 0.518 5.542 0.652 ;
        RECT 4.718 0.428 4.786 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.493 0.358 0.537 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 4.178 0.448 4.246 0.492 ;
        RECT 4.718 0.456 4.786 0.5 ;
        RECT 5.474 0.538 5.542 0.582 ;
        RECT 5.69 0.456 5.758 0.5 ;
        RECT 6.338 0.384 6.406 0.428 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.622 0.022 ;
        RECT 6.338 -0.022 6.406 0.292 ;
        RECT 5.69 -0.022 5.758 0.112 ;
        RECT 5.474 -0.022 5.542 0.112 ;
        RECT 4.61 -0.022 4.678 0.292 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.316 0.048 3.38 0.092 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.748 0.048 3.812 0.092 ;
        RECT 4.18 0.048 4.244 0.092 ;
        RECT 4.61 0.1715 4.678 0.2155 ;
        RECT 5.476 0.048 5.54 0.092 ;
        RECT 5.69 0.048 5.758 0.092 ;
        RECT 6.338 0.203 6.406 0.247 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.428 1.564 0.472 ;
      RECT 2.216 0.428 3.848 0.472 ;
      RECT 3.928 0.428 5.36 0.472 ;
      RECT 5.44 0.428 6.1 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.472 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 1.046 0.338 1.114 0.472 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 3.746 0.428 3.814 0.562 ;
      RECT 1.89 0.428 2.322 0.472 ;
      RECT 2.558 0.428 2.626 0.562 ;
      RECT 2.774 0.428 2.842 0.562 ;
      RECT 3.53 0.428 3.598 0.562 ;
      RECT 2.43 0.158 3.854 0.202 ;
      RECT 3.854 0.428 4.05 0.472 ;
      RECT 1.586 0.338 1.654 0.472 ;
      RECT 4.826 0.428 4.934 0.472 ;
      RECT 1.674 0.248 3.962 0.292 ;
      RECT 5.042 0.428 5.11 0.562 ;
      RECT 5.15 0.068 5.218 0.562 ;
      RECT 5.258 0.158 5.326 0.562 ;
      RECT 5.474 0.248 5.542 0.472 ;
      RECT 5.906 0.158 5.974 0.382 ;
    LAYER v1 ;
      RECT 6.018 0.428 6.078 0.472 ;
      RECT 5.478 0.428 5.538 0.472 ;
      RECT 5.262 0.428 5.322 0.472 ;
      RECT 5.046 0.428 5.106 0.472 ;
      RECT 4.83 0.428 4.89 0.472 ;
      RECT 3.966 0.428 4.026 0.472 ;
      RECT 3.75 0.428 3.81 0.472 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 2.778 0.428 2.838 0.472 ;
      RECT 2.562 0.428 2.622 0.472 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 0.726 0.428 0.786 0.472 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.078 0.428 0.138 0.472 ;
    LAYER v0 ;
      RECT 6.014 0.428 6.082 0.472 ;
      RECT 5.906 0.187 5.974 0.231 ;
      RECT 5.582 0.158 5.65 0.202 ;
      RECT 5.582 0.456 5.65 0.5 ;
      RECT 5.474 0.293 5.542 0.337 ;
      RECT 5.258 0.192 5.326 0.236 ;
      RECT 5.258 0.482 5.326 0.526 ;
      RECT 5.15 0.192 5.218 0.236 ;
      RECT 5.15 0.482 5.218 0.526 ;
      RECT 5.042 0.293 5.11 0.337 ;
      RECT 5.042 0.482 5.11 0.526 ;
      RECT 4.934 0.192 5.002 0.236 ;
      RECT 4.502 0.1715 4.57 0.2155 ;
      RECT 4.502 0.448 4.57 0.492 ;
      RECT 4.286 0.448 4.354 0.492 ;
      RECT 3.962 0.068 4.03 0.112 ;
      RECT 3.962 0.428 4.03 0.472 ;
      RECT 3.962 0.518 4.03 0.562 ;
      RECT 3.748 0.448 3.812 0.492 ;
      RECT 3.638 0.158 3.706 0.202 ;
      RECT 3.53 0.448 3.598 0.492 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.774 0.448 2.842 0.492 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.558 0.448 2.626 0.492 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.588 0.408 1.652 0.452 ;
      RECT 1.478 0.325 1.546 0.369 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.3685 1.114 0.4125 ;
      RECT 0.938 0.186 1.006 0.23 ;
      RECT 0.94 0.448 1.004 0.492 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.3155 0.79 0.3595 ;
      RECT 0.614 0.453 0.682 0.497 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.222 0.338 1.438 0.382 ;
      RECT 1.546 0.158 2.106 0.202 ;
      RECT 1.006 0.518 1.154 0.562 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.222 0.428 1.37 0.472 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.438 0.518 2.322 0.562 ;
      RECT 3.814 0.518 4.05 0.562 ;
      RECT 3.854 0.068 3.922 0.202 ;
      RECT 3.922 0.068 4.05 0.112 ;
      RECT 1.654 0.338 4.286 0.382 ;
      RECT 4.286 0.338 4.354 0.562 ;
      RECT 4.934 0.158 5.002 0.472 ;
      RECT 3.962 0.158 4.03 0.292 ;
      RECT 4.03 0.158 4.286 0.202 ;
      RECT 4.286 0.068 4.354 0.202 ;
      RECT 4.354 0.068 4.502 0.112 ;
      RECT 4.502 0.068 4.57 0.562 ;
      RECT 4.57 0.338 4.826 0.382 ;
      RECT 4.826 0.068 4.894 0.382 ;
      RECT 4.894 0.068 5.042 0.112 ;
      RECT 5.042 0.068 5.11 0.382 ;
      RECT 5.218 0.068 5.366 0.112 ;
      RECT 5.366 0.068 5.434 0.202 ;
      RECT 5.582 0.338 5.65 0.562 ;
      RECT 5.65 0.338 5.69 0.382 ;
      RECT 5.434 0.158 5.69 0.202 ;
      RECT 5.69 0.158 5.758 0.382 ;
      RECT 5.974 0.338 6.014 0.382 ;
      RECT 6.014 0.338 6.082 0.562 ;
  END
END b15fqy08fhn1n16x5

MACRO b15fqy203hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy203hn1n02x5 0 0 ;
  SIZE 5.616 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 4.948889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 3.29925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.15 0.428 5.218 0.562 ;
        RECT 4.394 0.338 4.462 0.562 ;
        RECT 1.154 0.338 1.222 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
      LAYER m2 ;
        RECT 0.38 0.518 5.236 0.562 ;
      LAYER v1 ;
        RECT 0.402 0.518 0.462 0.562 ;
        RECT 1.158 0.518 1.218 0.562 ;
        RECT 4.398 0.518 4.458 0.562 ;
        RECT 5.154 0.518 5.214 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.498 0.466 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
        RECT 4.394 0.498 4.462 0.542 ;
        RECT 5.15 0.498 5.218 0.542 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.068 3.49 0.382 ;
      LAYER v0 ;
        RECT 3.422 0.3155 3.49 0.3595 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.338 2.41 0.382 ;
        RECT 2.018 0.158 2.086 0.382 ;
      LAYER v0 ;
        RECT 2.234 0.338 2.302 0.382 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.068 3.274 0.382 ;
      LAYER v0 ;
        RECT 3.206 0.3155 3.274 0.3595 ;
    END
  END d2
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.3905 0.25 0.4345 ;
        RECT 0.182 0.1915 0.25 0.2355 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.366 0.158 5.434 0.562 ;
      LAYER v0 ;
        RECT 5.366 0.383 5.434 0.427 ;
        RECT 5.366 0.1915 5.434 0.2355 ;
    END
  END o2
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.292 ;
      LAYER v0 ;
        RECT 2.666 0.088 2.734 0.132 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.292 ;
      LAYER v0 ;
        RECT 2.882 0.088 2.95 0.132 ;
    END
  END si2
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 5.51 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 2.448889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 3.058 0.382 ;
        RECT 2.99 0.068 3.058 0.382 ;
        RECT 2.558 0.068 2.626 0.382 ;
        RECT 2.342 0.068 2.626 0.112 ;
      LAYER v0 ;
        RECT 2.45 0.068 2.518 0.112 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 2.882 0.338 2.95 0.382 ;
        RECT 2.99 0.088 3.058 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.65 0.652 ;
        RECT 5.474 0.518 5.542 0.652 ;
        RECT 5.042 0.338 5.11 0.652 ;
        RECT 4.502 0.338 4.57 0.652 ;
        RECT 4.178 0.338 4.246 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 1.046 0.338 1.114 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.506 0.403 0.574 0.447 ;
        RECT 1.046 0.402 1.114 0.446 ;
        RECT 1.37 0.377 1.438 0.421 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.234 0.473 2.302 0.517 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 3.422 0.471 3.49 0.515 ;
        RECT 3.746 0.471 3.814 0.515 ;
        RECT 4.178 0.408 4.246 0.452 ;
        RECT 4.502 0.402 4.57 0.446 ;
        RECT 5.042 0.403 5.11 0.447 ;
        RECT 5.476 0.538 5.54 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.65 0.022 ;
        RECT 5.474 -0.022 5.542 0.112 ;
        RECT 5.15 -0.022 5.218 0.202 ;
        RECT 4.394 -0.022 4.462 0.202 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.046 0.158 1.33 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.398 0.088 0.466 0.132 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.802 0.113 1.87 0.157 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.774 0.215 2.842 0.259 ;
        RECT 3.314 0.1135 3.382 0.1575 ;
        RECT 3.746 0.1135 3.814 0.1575 ;
        RECT 4.394 0.138 4.462 0.182 ;
        RECT 5.15 0.088 5.218 0.132 ;
        RECT 5.476 0.048 5.54 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 0.824 0.382 ;
      RECT 0.904 0.338 1.688 0.382 ;
      RECT 2.216 0.248 2.536 0.292 ;
      RECT 3.08 0.248 3.724 0.292 ;
      RECT 1.768 0.338 3.848 0.382 ;
      RECT 3.928 0.338 4.712 0.382 ;
      RECT 0.812 0.428 4.804 0.472 ;
      RECT 4.792 0.338 5.576 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.382 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 0.83 0.248 1.262 0.292 ;
      RECT 1.37 0.158 1.586 0.202 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.478 0.518 1.694 0.562 ;
      RECT 1.91 0.068 2.126 0.112 ;
      RECT 2.018 0.428 2.086 0.562 ;
      RECT 2.45 0.158 2.518 0.472 ;
      RECT 2.882 0.428 3.098 0.472 ;
      RECT 3.962 0.158 4.03 0.472 ;
      RECT 3.53 0.068 3.598 0.562 ;
      RECT 3.638 0.068 3.706 0.292 ;
      RECT 4.07 0.248 4.138 0.472 ;
      RECT 3.638 0.338 3.854 0.382 ;
      RECT 4.286 0.248 4.354 0.562 ;
      RECT 4.394 0.338 4.462 0.562 ;
      RECT 4.61 0.338 4.678 0.562 ;
      RECT 4.718 0.428 4.786 0.562 ;
      RECT 4.61 0.158 4.826 0.202 ;
      RECT 4.61 0.068 4.934 0.112 ;
      RECT 5.042 0.068 5.11 0.292 ;
      RECT 5.15 0.428 5.218 0.562 ;
      RECT 5.474 0.248 5.542 0.382 ;
    LAYER v1 ;
      RECT 5.478 0.338 5.538 0.382 ;
      RECT 4.83 0.338 4.89 0.382 ;
      RECT 4.722 0.428 4.782 0.472 ;
      RECT 4.614 0.338 4.674 0.382 ;
      RECT 4.074 0.428 4.134 0.472 ;
      RECT 3.966 0.338 4.026 0.382 ;
      RECT 3.75 0.338 3.81 0.382 ;
      RECT 3.642 0.248 3.702 0.292 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 3.102 0.248 3.162 0.292 ;
      RECT 2.454 0.248 2.514 0.292 ;
      RECT 2.238 0.248 2.298 0.292 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.59 0.338 1.65 0.382 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 5.474 0.293 5.542 0.337 ;
      RECT 5.258 0.088 5.326 0.132 ;
      RECT 5.258 0.498 5.326 0.542 ;
      RECT 5.042 0.088 5.11 0.132 ;
      RECT 4.934 0.498 5.002 0.542 ;
      RECT 4.826 0.363 4.894 0.407 ;
      RECT 4.718 0.068 4.786 0.112 ;
      RECT 4.718 0.158 4.786 0.202 ;
      RECT 4.718 0.498 4.786 0.542 ;
      RECT 4.61 0.248 4.678 0.292 ;
      RECT 4.61 0.498 4.678 0.542 ;
      RECT 4.286 0.408 4.354 0.452 ;
      RECT 4.178 0.068 4.246 0.112 ;
      RECT 4.07 0.158 4.138 0.202 ;
      RECT 4.07 0.293 4.138 0.337 ;
      RECT 3.962 0.383 4.03 0.427 ;
      RECT 3.962 0.518 4.03 0.562 ;
      RECT 3.638 0.1135 3.706 0.1575 ;
      RECT 3.53 0.1135 3.598 0.1575 ;
      RECT 3.53 0.471 3.598 0.515 ;
      RECT 3.098 0.208 3.166 0.252 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.45 0.203 2.518 0.247 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.91 0.1985 1.978 0.2425 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.586 0.3835 1.654 0.4275 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.377 1.33 0.421 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.498 0.898 0.542 ;
      RECT 0.722 0.363 0.79 0.407 ;
      RECT 0.614 0.498 0.682 0.542 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.79 0.158 1.006 0.202 ;
      RECT 0.682 0.068 1.222 0.112 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.37 0.068 1.694 0.112 ;
      RECT 1.694 0.068 1.762 0.562 ;
      RECT 1.762 0.338 1.91 0.382 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.194 0.248 2.41 0.292 ;
      RECT 2.518 0.428 2.734 0.472 ;
      RECT 3.098 0.158 3.166 0.472 ;
      RECT 4.03 0.158 4.246 0.202 ;
      RECT 3.854 0.068 3.922 0.562 ;
      RECT 3.922 0.518 4.138 0.562 ;
      RECT 3.922 0.068 4.354 0.112 ;
      RECT 4.354 0.248 4.786 0.292 ;
      RECT 4.826 0.158 4.894 0.472 ;
      RECT 4.934 0.068 5.002 0.562 ;
      RECT 5.11 0.248 5.258 0.292 ;
      RECT 5.258 0.068 5.326 0.562 ;
  END
END b15fqy203hn1n02x5

MACRO b15fqy203hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy203hn1n03x5 0 0 ;
  SIZE 5.832 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
      ANTENNAMAXAREACAR 8.401111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
      ANTENNAMAXAREACAR 8.401111 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.366 0.248 5.434 0.562 ;
        RECT 4.502 0.338 4.57 0.562 ;
        RECT 1.262 0.338 1.33 0.562 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER m2 ;
        RECT 0.38 0.518 5.452 0.562 ;
      LAYER v1 ;
        RECT 0.402 0.518 0.462 0.562 ;
        RECT 1.266 0.518 1.326 0.562 ;
        RECT 4.506 0.518 4.566 0.562 ;
        RECT 5.37 0.518 5.43 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
        RECT 1.262 0.498 1.33 0.542 ;
        RECT 4.502 0.498 4.57 0.542 ;
        RECT 5.366 0.293 5.434 0.337 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.598 0.382 ;
      LAYER v0 ;
        RECT 3.53 0.3155 3.598 0.3595 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.338 2.518 0.382 ;
        RECT 2.126 0.158 2.194 0.382 ;
      LAYER v0 ;
        RECT 2.342 0.338 2.41 0.382 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.068 3.382 0.382 ;
      LAYER v0 ;
        RECT 3.314 0.3155 3.382 0.3595 ;
    END
  END d2
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.383 0.142 0.427 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.69 0.158 5.758 0.562 ;
      LAYER v0 ;
        RECT 5.69 0.403 5.758 0.447 ;
        RECT 5.69 0.203 5.758 0.247 ;
    END
  END o2
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.068 2.842 0.292 ;
      LAYER v0 ;
        RECT 2.774 0.088 2.842 0.132 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.068 3.058 0.292 ;
      LAYER v0 ;
        RECT 2.99 0.088 3.058 0.132 ;
    END
  END si2
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 5.51 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 2.448889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.338 3.166 0.382 ;
        RECT 3.098 0.068 3.166 0.382 ;
        RECT 2.666 0.068 2.734 0.382 ;
        RECT 2.45 0.068 2.734 0.112 ;
      LAYER v0 ;
        RECT 2.558 0.068 2.626 0.112 ;
        RECT 2.774 0.338 2.842 0.382 ;
        RECT 2.99 0.338 3.058 0.382 ;
        RECT 3.098 0.088 3.166 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.866 0.652 ;
        RECT 5.582 0.338 5.65 0.652 ;
        RECT 5.15 0.338 5.218 0.652 ;
        RECT 4.61 0.338 4.678 0.652 ;
        RECT 4.286 0.338 4.354 0.652 ;
        RECT 3.854 0.428 3.922 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.614 0.338 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 0.614 0.403 0.682 0.447 ;
        RECT 1.154 0.402 1.222 0.446 ;
        RECT 1.478 0.377 1.546 0.421 ;
        RECT 1.91 0.538 1.978 0.582 ;
        RECT 2.342 0.473 2.41 0.517 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.53 0.471 3.598 0.515 ;
        RECT 3.854 0.471 3.922 0.515 ;
        RECT 4.286 0.408 4.354 0.452 ;
        RECT 4.61 0.402 4.678 0.446 ;
        RECT 5.15 0.403 5.218 0.447 ;
        RECT 5.582 0.403 5.65 0.447 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.866 0.022 ;
        RECT 5.582 -0.022 5.65 0.292 ;
        RECT 5.258 -0.022 5.326 0.202 ;
        RECT 4.502 -0.022 4.57 0.202 ;
        RECT 3.854 -0.022 3.922 0.202 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.882 -0.022 2.95 0.292 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.154 0.158 1.438 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.91 0.113 1.978 0.157 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.882 0.215 2.95 0.259 ;
        RECT 3.422 0.1135 3.49 0.1575 ;
        RECT 3.854 0.1135 3.922 0.1575 ;
        RECT 4.502 0.138 4.57 0.182 ;
        RECT 5.258 0.138 5.326 0.182 ;
        RECT 5.582 0.203 5.65 0.247 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 0.932 0.382 ;
      RECT 1.012 0.338 1.796 0.382 ;
      RECT 2.324 0.248 2.644 0.292 ;
      RECT 3.188 0.248 3.832 0.292 ;
      RECT 1.876 0.338 3.956 0.382 ;
      RECT 4.036 0.338 4.82 0.382 ;
      RECT 0.92 0.428 4.912 0.472 ;
      RECT 4.9 0.338 5.344 0.382 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.398 0.248 0.466 0.562 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 0.938 0.248 1.37 0.292 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.478 0.158 1.694 0.202 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.586 0.518 1.802 0.562 ;
      RECT 2.018 0.068 2.234 0.112 ;
      RECT 2.126 0.428 2.194 0.562 ;
      RECT 2.558 0.158 2.626 0.472 ;
      RECT 2.99 0.428 3.206 0.472 ;
      RECT 4.07 0.158 4.138 0.472 ;
      RECT 3.638 0.068 3.706 0.562 ;
      RECT 3.746 0.068 3.814 0.292 ;
      RECT 4.178 0.248 4.246 0.472 ;
      RECT 3.746 0.338 3.962 0.382 ;
      RECT 4.394 0.248 4.462 0.562 ;
      RECT 4.502 0.338 4.57 0.562 ;
      RECT 4.718 0.338 4.786 0.562 ;
      RECT 4.826 0.428 4.894 0.562 ;
      RECT 4.718 0.158 4.934 0.202 ;
      RECT 4.826 0.068 5.042 0.112 ;
      RECT 5.258 0.338 5.326 0.562 ;
      RECT 5.366 0.248 5.434 0.562 ;
      RECT 5.474 0.158 5.542 0.472 ;
    LAYER v1 ;
      RECT 5.262 0.338 5.322 0.382 ;
      RECT 4.938 0.338 4.998 0.382 ;
      RECT 4.83 0.428 4.89 0.472 ;
      RECT 4.722 0.338 4.782 0.382 ;
      RECT 4.182 0.428 4.242 0.472 ;
      RECT 4.074 0.338 4.134 0.382 ;
      RECT 3.858 0.338 3.918 0.382 ;
      RECT 3.75 0.248 3.81 0.292 ;
      RECT 3.642 0.428 3.702 0.472 ;
      RECT 3.21 0.248 3.27 0.292 ;
      RECT 2.562 0.248 2.622 0.292 ;
      RECT 2.346 0.248 2.406 0.292 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 5.474 0.203 5.542 0.247 ;
      RECT 5.474 0.403 5.542 0.447 ;
      RECT 5.258 0.403 5.326 0.447 ;
      RECT 5.042 0.498 5.11 0.542 ;
      RECT 4.934 0.068 5.002 0.112 ;
      RECT 4.934 0.363 5.002 0.407 ;
      RECT 4.826 0.158 4.894 0.202 ;
      RECT 4.826 0.498 4.894 0.542 ;
      RECT 4.718 0.248 4.786 0.292 ;
      RECT 4.718 0.498 4.786 0.542 ;
      RECT 4.394 0.408 4.462 0.452 ;
      RECT 4.286 0.068 4.354 0.112 ;
      RECT 4.178 0.158 4.246 0.202 ;
      RECT 4.178 0.293 4.246 0.337 ;
      RECT 4.07 0.383 4.138 0.427 ;
      RECT 4.07 0.518 4.138 0.562 ;
      RECT 3.746 0.1135 3.814 0.1575 ;
      RECT 3.638 0.1135 3.706 0.1575 ;
      RECT 3.638 0.471 3.706 0.515 ;
      RECT 3.206 0.208 3.274 0.252 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.558 0.203 2.626 0.247 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 2.018 0.1985 2.086 0.2425 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.694 0.3835 1.762 0.4275 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.37 0.377 1.438 0.421 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.498 1.114 0.542 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.83 0.363 0.898 0.407 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.506 0.403 0.574 0.447 ;
      RECT 0.29 0.203 0.358 0.247 ;
      RECT 0.29 0.383 0.358 0.427 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.79 0.068 1.006 0.112 ;
      RECT 0.898 0.158 1.114 0.202 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.478 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.87 0.338 2.018 0.382 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.302 0.248 2.518 0.292 ;
      RECT 2.626 0.428 2.842 0.472 ;
      RECT 3.206 0.158 3.274 0.472 ;
      RECT 4.138 0.158 4.354 0.202 ;
      RECT 3.962 0.068 4.03 0.562 ;
      RECT 4.03 0.518 4.246 0.562 ;
      RECT 4.03 0.068 4.462 0.112 ;
      RECT 4.462 0.248 4.894 0.292 ;
      RECT 4.934 0.158 5.002 0.472 ;
      RECT 5.042 0.068 5.11 0.562 ;
  END
END b15fqy203hn1n03x5

MACRO b15fqy203hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy203hn1n04x5 0 0 ;
  SIZE 6.048 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 5.05925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0216 LAYER m2 ;
      ANTENNAMAXAREACAR 5.048611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.474 0.428 5.542 0.562 ;
        RECT 4.826 0.338 4.894 0.562 ;
        RECT 4.61 0.338 4.894 0.382 ;
        RECT 1.154 0.338 1.438 0.382 ;
        RECT 1.154 0.338 1.222 0.562 ;
        RECT 0.506 0.428 0.574 0.562 ;
      LAYER m2 ;
        RECT 0.488 0.518 5.56 0.562 ;
      LAYER v1 ;
        RECT 0.51 0.518 0.57 0.562 ;
        RECT 1.158 0.518 1.218 0.562 ;
        RECT 4.83 0.518 4.89 0.562 ;
        RECT 5.478 0.518 5.538 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 4.718 0.338 4.786 0.382 ;
        RECT 5.474 0.498 5.542 0.542 ;
    END
  END rb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.068 3.706 0.382 ;
      LAYER v0 ;
        RECT 3.638 0.3155 3.706 0.3595 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.338 2.626 0.382 ;
        RECT 2.234 0.158 2.302 0.382 ;
      LAYER v0 ;
        RECT 2.45 0.338 2.518 0.382 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.068 3.49 0.382 ;
      LAYER v0 ;
        RECT 3.422 0.3155 3.49 0.3595 ;
    END
  END d2
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.158 0.142 0.202 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.906 0.068 5.974 0.562 ;
      LAYER v0 ;
        RECT 5.906 0.428 5.974 0.472 ;
        RECT 5.906 0.158 5.974 0.202 ;
    END
  END o2
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.292 ;
      LAYER v0 ;
        RECT 2.882 0.088 2.95 0.132 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.068 3.166 0.292 ;
      LAYER v0 ;
        RECT 3.098 0.088 3.166 0.132 ;
    END
  END si2
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 5.51 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 2.448889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.338 3.274 0.382 ;
        RECT 3.206 0.068 3.274 0.382 ;
        RECT 2.774 0.068 2.842 0.382 ;
        RECT 2.558 0.068 2.842 0.112 ;
      LAYER v0 ;
        RECT 2.666 0.068 2.734 0.112 ;
        RECT 2.882 0.338 2.95 0.382 ;
        RECT 3.098 0.338 3.166 0.382 ;
        RECT 3.206 0.088 3.274 0.132 ;
    END
  END ssb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.082 0.652 ;
        RECT 5.798 0.338 5.866 0.652 ;
        RECT 5.366 0.338 5.434 0.652 ;
        RECT 4.718 0.428 4.786 0.652 ;
        RECT 4.394 0.338 4.462 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.638 0.428 3.706 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.586 0.338 1.654 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.338 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.614 0.403 0.682 0.447 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.586 0.403 1.654 0.447 ;
        RECT 2.018 0.538 2.086 0.582 ;
        RECT 2.45 0.473 2.518 0.517 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.638 0.471 3.706 0.515 ;
        RECT 3.962 0.498 4.03 0.542 ;
        RECT 4.394 0.403 4.462 0.447 ;
        RECT 4.718 0.473 4.786 0.517 ;
        RECT 5.366 0.403 5.434 0.447 ;
        RECT 5.798 0.428 5.866 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.082 0.022 ;
        RECT 5.798 -0.022 5.866 0.292 ;
        RECT 5.474 -0.022 5.542 0.202 ;
        RECT 4.61 -0.022 4.678 0.112 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.53 -0.022 3.598 0.202 ;
        RECT 2.99 -0.022 3.058 0.292 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.018 -0.022 2.086 0.292 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.506 0.115 0.574 0.159 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 2.018 0.1985 2.086 0.2425 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 2.99 0.215 3.058 0.259 ;
        RECT 3.53 0.1135 3.598 0.1575 ;
        RECT 3.962 0.1135 4.03 0.1575 ;
        RECT 4.61 0.048 4.678 0.092 ;
        RECT 5.474 0.138 5.542 0.182 ;
        RECT 5.798 0.158 5.866 0.202 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.38 0.338 0.932 0.382 ;
      RECT 1.012 0.338 1.904 0.382 ;
      RECT 2.432 0.248 2.752 0.292 ;
      RECT 3.296 0.248 3.94 0.292 ;
      RECT 1.984 0.338 4.064 0.382 ;
      RECT 4.144 0.338 5.036 0.382 ;
      RECT 0.92 0.428 5.128 0.472 ;
      RECT 5.116 0.338 5.668 0.382 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.046 0.248 1.478 0.292 ;
      RECT 1.586 0.158 1.802 0.202 ;
      RECT 1.694 0.248 1.762 0.472 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 2.126 0.068 2.342 0.112 ;
      RECT 2.234 0.428 2.302 0.562 ;
      RECT 2.666 0.158 2.734 0.472 ;
      RECT 3.098 0.428 3.314 0.472 ;
      RECT 4.178 0.158 4.246 0.472 ;
      RECT 3.746 0.068 3.814 0.562 ;
      RECT 3.854 0.068 3.922 0.292 ;
      RECT 4.286 0.248 4.354 0.472 ;
      RECT 4.61 0.338 4.826 0.382 ;
      RECT 4.502 0.248 4.57 0.562 ;
      RECT 4.934 0.338 5.002 0.562 ;
      RECT 5.042 0.248 5.11 0.472 ;
      RECT 4.934 0.158 5.15 0.202 ;
      RECT 3.854 0.338 4.07 0.382 ;
      RECT 5.474 0.428 5.542 0.562 ;
      RECT 5.582 0.248 5.65 0.382 ;
      RECT 5.69 0.068 5.758 0.562 ;
    LAYER v1 ;
      RECT 5.586 0.338 5.646 0.382 ;
      RECT 5.154 0.338 5.214 0.382 ;
      RECT 5.046 0.428 5.106 0.472 ;
      RECT 4.938 0.338 4.998 0.382 ;
      RECT 4.29 0.428 4.35 0.472 ;
      RECT 4.182 0.338 4.242 0.382 ;
      RECT 3.966 0.338 4.026 0.382 ;
      RECT 3.858 0.248 3.918 0.292 ;
      RECT 3.75 0.428 3.81 0.472 ;
      RECT 3.318 0.248 3.378 0.292 ;
      RECT 2.67 0.248 2.73 0.292 ;
      RECT 2.454 0.248 2.514 0.292 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 2.13 0.338 2.19 0.382 ;
      RECT 1.806 0.338 1.866 0.382 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.402 0.338 0.462 0.382 ;
    LAYER v0 ;
      RECT 5.69 0.158 5.758 0.202 ;
      RECT 5.69 0.428 5.758 0.472 ;
      RECT 5.582 0.3085 5.65 0.3525 ;
      RECT 5.258 0.498 5.326 0.542 ;
      RECT 5.15 0.068 5.218 0.112 ;
      RECT 5.15 0.403 5.218 0.447 ;
      RECT 5.042 0.158 5.11 0.202 ;
      RECT 5.042 0.293 5.11 0.337 ;
      RECT 5.042 0.518 5.11 0.562 ;
      RECT 4.826 0.248 4.894 0.292 ;
      RECT 4.502 0.403 4.57 0.447 ;
      RECT 4.394 0.068 4.462 0.112 ;
      RECT 4.286 0.158 4.354 0.202 ;
      RECT 4.286 0.293 4.354 0.337 ;
      RECT 4.178 0.383 4.246 0.427 ;
      RECT 4.07 0.498 4.138 0.542 ;
      RECT 3.854 0.1135 3.922 0.1575 ;
      RECT 3.746 0.1135 3.814 0.1575 ;
      RECT 3.746 0.471 3.814 0.515 ;
      RECT 3.314 0.208 3.382 0.252 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.203 2.734 0.247 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.234 0.448 2.302 0.492 ;
      RECT 2.126 0.1985 2.194 0.2425 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 1.802 0.3835 1.87 0.4275 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.478 0.403 1.546 0.447 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.83 0.402 0.898 0.446 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.398 0.318 0.466 0.362 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
    LAYER m1 ;
      RECT 0.83 0.518 1.046 0.562 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 0.898 0.158 1.114 0.202 ;
      RECT 1.222 0.338 1.438 0.382 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 0.79 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 1.694 0.518 1.91 0.562 ;
      RECT 1.546 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 1.978 0.338 2.126 0.382 ;
      RECT 2.126 0.158 2.194 0.562 ;
      RECT 2.342 0.068 2.41 0.292 ;
      RECT 2.41 0.248 2.626 0.292 ;
      RECT 2.734 0.428 2.95 0.472 ;
      RECT 3.314 0.158 3.382 0.472 ;
      RECT 4.246 0.158 4.462 0.202 ;
      RECT 4.826 0.338 4.894 0.562 ;
      RECT 4.57 0.248 5.002 0.292 ;
      RECT 5.002 0.518 5.218 0.562 ;
      RECT 5.15 0.158 5.218 0.472 ;
      RECT 4.07 0.068 4.138 0.562 ;
      RECT 4.138 0.068 4.502 0.112 ;
      RECT 4.502 0.068 4.57 0.202 ;
      RECT 4.57 0.158 4.718 0.202 ;
      RECT 4.718 0.068 4.786 0.202 ;
      RECT 4.786 0.068 5.258 0.112 ;
      RECT 5.258 0.068 5.326 0.562 ;
  END
END b15fqy203hn1n04x5

MACRO b15fqy403hn1d02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy403hn1d02x5 0 0 ;
  SIZE 5.184 BY 1.26 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN d3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.878 2.842 1.012 ;
      LAYER m2 ;
        RECT 2.74 0.878 3.416 0.922 ;
      LAYER v1 ;
        RECT 2.778 0.878 2.838 0.922 ;
      LAYER v0 ;
        RECT 2.774 0.923 2.842 0.967 ;
    END
  END d3
  PIN d4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.878 2.626 1.012 ;
      LAYER m2 ;
        RECT 2.216 0.878 2.66 0.922 ;
      LAYER v1 ;
        RECT 2.562 0.878 2.622 0.922 ;
      LAYER v0 ;
        RECT 2.558 0.923 2.626 0.967 ;
    END
  END d4
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0288 LAYER m2 ;
      ANTENNAMAXAREACAR 3.56777775 LAYER m1 ;
      ANTENNAMAXAREACAR 4.83333325 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.036 LAYER m2 ;
      ANTENNAMAXAREACAR 3.56777775 LAYER m1 ;
      ANTENNAMAXAREACAR 4.83333325 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.718 0.698 4.786 0.832 ;
        RECT 3.962 0.698 4.03 0.832 ;
        RECT 1.154 0.698 1.222 0.832 ;
        RECT 0.398 0.698 0.466 0.832 ;
      LAYER m2 ;
        RECT 0.38 0.698 4.804 0.742 ;
      LAYER v1 ;
        RECT 0.402 0.698 0.462 0.742 ;
        RECT 1.158 0.698 1.218 0.742 ;
        RECT 3.966 0.698 4.026 0.742 ;
        RECT 4.722 0.698 4.782 0.742 ;
      LAYER v0 ;
        RECT 0.398 0.718 0.466 0.762 ;
        RECT 1.154 0.718 1.222 0.762 ;
        RECT 3.962 0.718 4.03 0.762 ;
        RECT 4.718 0.718 4.786 0.762 ;
    END
  END rb
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
      ANTENNAMAXAREACAR 2.7805555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 2.2244445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.158 2.95 0.382 ;
        RECT 2.45 0.158 2.518 0.382 ;
      LAYER m2 ;
        RECT 2.432 0.158 2.968 0.202 ;
      LAYER v1 ;
        RECT 2.454 0.158 2.514 0.202 ;
        RECT 2.886 0.158 2.946 0.202 ;
      LAYER v0 ;
        RECT 2.45 0.293 2.518 0.337 ;
        RECT 2.882 0.293 2.95 0.337 ;
    END
  END ssb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.788 1.978 1.012 ;
      LAYER v0 ;
        RECT 1.91 0.923 1.978 0.967 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.248 2.626 0.472 ;
      LAYER v0 ;
        RECT 2.558 0.293 2.626 0.337 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.248 2.842 0.382 ;
      LAYER v0 ;
        RECT 2.774 0.293 2.842 0.337 ;
    END
  END d2
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.403 0.25 0.447 ;
        RECT 0.182 0.1915 0.25 0.2355 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.934 0.158 5.002 0.562 ;
      LAYER v0 ;
        RECT 4.934 0.403 5.002 0.447 ;
        RECT 4.934 0.1915 5.002 0.2355 ;
    END
  END o2
  PIN o3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.934 0.698 5.002 1.102 ;
      LAYER v0 ;
        RECT 4.934 1.0245 5.002 1.0685 ;
        RECT 4.934 0.813 5.002 0.857 ;
    END
  END o3
  PIN o4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.698 0.25 1.102 ;
      LAYER v0 ;
        RECT 0.182 1.0245 0.25 1.0685 ;
        RECT 0.182 0.813 0.25 0.857 ;
    END
  END o4
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.158 2.302 0.382 ;
      LAYER v0 ;
        RECT 2.234 0.293 2.302 0.337 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.158 3.166 0.382 ;
      LAYER v0 ;
        RECT 3.098 0.293 3.166 0.337 ;
    END
  END si2
  PIN si3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.878 3.166 1.192 ;
      LAYER v0 ;
        RECT 3.098 0.923 3.166 0.967 ;
    END
  END si3
  PIN si4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.878 2.302 1.192 ;
      LAYER v0 ;
        RECT 2.234 0.923 2.302 0.967 ;
    END
  END si4
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.218 0.652 ;
        RECT 5.042 0.518 5.11 0.742 ;
        RECT 4.61 0.338 4.678 0.922 ;
        RECT 4.07 0.338 4.138 0.922 ;
        RECT 3.746 0.338 3.814 0.922 ;
        RECT 1.37 0.338 1.438 0.922 ;
        RECT 1.046 0.338 1.114 0.922 ;
        RECT 0.506 0.338 0.574 0.922 ;
        RECT 0.074 0.518 0.142 0.742 ;
      LAYER v0 ;
        RECT 0.076 0.678 0.14 0.722 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.506 0.813 0.574 0.857 ;
        RECT 0.506 0.403 0.574 0.447 ;
        RECT 1.046 0.814 1.114 0.858 ;
        RECT 1.046 0.402 1.114 0.446 ;
        RECT 1.37 0.839 1.438 0.883 ;
        RECT 1.37 0.377 1.438 0.421 ;
        RECT 1.802 0.608 1.87 0.652 ;
        RECT 2.126 0.608 2.194 0.652 ;
        RECT 2.666 0.608 2.734 0.652 ;
        RECT 2.99 0.608 3.058 0.652 ;
        RECT 3.206 0.608 3.274 0.652 ;
        RECT 3.746 0.813 3.814 0.857 ;
        RECT 3.746 0.403 3.814 0.447 ;
        RECT 4.07 0.814 4.138 0.858 ;
        RECT 4.07 0.402 4.138 0.446 ;
        RECT 4.61 0.813 4.678 0.857 ;
        RECT 4.61 0.403 4.678 0.447 ;
        RECT 5.044 0.678 5.108 0.722 ;
        RECT 5.044 0.538 5.108 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.218 0.022 ;
        RECT 5.042 -0.022 5.11 0.112 ;
        RECT 4.718 -0.022 4.786 0.202 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.126 -0.022 2.194 0.292 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.046 0.158 1.33 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
        RECT -0.034 1.238 5.218 1.282 ;
        RECT 5.042 1.148 5.11 1.282 ;
        RECT 4.718 1.058 4.786 1.282 ;
        RECT 3.962 1.058 4.03 1.282 ;
        RECT 3.314 0.968 3.382 1.282 ;
        RECT 2.666 1.148 2.734 1.282 ;
        RECT 2.126 0.968 2.194 1.282 ;
        RECT 1.91 1.058 1.978 1.282 ;
        RECT 1.262 1.058 1.33 1.282 ;
        RECT 1.046 1.058 1.33 1.102 ;
        RECT 0.398 1.058 0.466 1.282 ;
        RECT 0.074 1.148 0.142 1.282 ;
      LAYER v0 ;
        RECT 0.076 1.168 0.14 1.212 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.398 1.128 0.466 1.172 ;
        RECT 0.398 0.088 0.466 0.132 ;
        RECT 1.154 1.058 1.222 1.102 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.802 0.2025 1.87 0.2465 ;
        RECT 1.91 1.128 1.978 1.172 ;
        RECT 2.126 1.0135 2.194 1.0575 ;
        RECT 2.126 0.2025 2.194 0.2465 ;
        RECT 2.666 1.168 2.734 1.212 ;
        RECT 2.666 0.048 2.734 0.092 ;
        RECT 3.206 0.088 3.274 0.132 ;
        RECT 3.314 1.0375 3.382 1.0815 ;
        RECT 3.962 1.078 4.03 1.122 ;
        RECT 3.962 0.138 4.03 0.182 ;
        RECT 4.718 1.128 4.786 1.172 ;
        RECT 4.718 0.088 4.786 0.132 ;
        RECT 5.044 1.168 5.108 1.212 ;
        RECT 5.044 0.048 5.108 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.878 0.824 0.922 ;
      RECT 0.04 0.428 0.824 0.472 ;
      RECT 0.904 0.878 1.672 0.922 ;
      RECT 0.904 0.428 1.688 0.472 ;
      RECT 1.768 0.428 3.416 0.472 ;
      RECT 3.496 0.878 4.28 0.922 ;
      RECT 3.496 0.428 4.28 0.472 ;
      RECT 0.812 0.788 4.372 0.832 ;
      RECT 0.812 0.518 4.372 0.562 ;
      RECT 4.36 0.878 5.144 0.922 ;
      RECT 4.36 0.428 5.144 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.878 0.142 1.012 ;
      RECT 0.074 0.248 0.142 0.472 ;
      RECT 0.398 0.698 0.466 0.832 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.614 0.698 0.682 1.192 ;
      RECT 0.83 0.698 0.898 0.832 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.722 0.788 0.79 1.102 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.938 0.698 1.006 0.922 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.83 0.968 1.262 1.012 ;
      RECT 1.154 0.698 1.222 0.832 ;
      RECT 0.83 0.248 1.262 0.292 ;
      RECT 1.37 1.058 1.586 1.102 ;
      RECT 1.478 0.788 1.546 1.012 ;
      RECT 1.478 0.248 1.546 0.562 ;
      RECT 1.37 0.158 1.586 0.202 ;
      RECT 1.37 1.148 1.694 1.192 ;
      RECT 1.37 0.068 1.694 0.112 ;
      RECT 1.802 0.698 1.87 1.192 ;
      RECT 2.018 0.788 2.086 1.102 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 2.45 0.158 2.518 0.382 ;
      RECT 2.558 0.878 2.626 1.012 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.342 1.148 2.558 1.192 ;
      RECT 2.774 0.878 2.842 1.012 ;
      RECT 2.882 0.158 2.95 0.382 ;
      RECT 2.234 0.068 2.558 0.112 ;
      RECT 2.774 0.788 2.99 0.832 ;
      RECT 2.774 0.428 2.99 0.472 ;
      RECT 3.53 0.788 3.598 1.102 ;
      RECT 3.638 0.788 3.706 1.012 ;
      RECT 3.638 0.248 3.706 0.562 ;
      RECT 3.53 0.158 3.598 0.472 ;
      RECT 3.422 0.698 3.49 1.192 ;
      RECT 3.314 0.338 3.382 0.562 ;
      RECT 3.854 0.698 3.922 1.012 ;
      RECT 3.962 0.698 4.03 0.832 ;
      RECT 4.178 0.698 4.246 0.922 ;
      RECT 4.178 0.428 4.246 0.562 ;
      RECT 3.854 0.248 3.922 0.562 ;
      RECT 4.286 0.698 4.354 0.832 ;
      RECT 4.286 0.428 4.354 0.562 ;
      RECT 4.178 1.058 4.394 1.102 ;
      RECT 4.178 0.158 4.394 0.202 ;
      RECT 4.178 1.148 4.502 1.192 ;
      RECT 4.178 0.068 4.502 0.112 ;
      RECT 4.61 0.968 4.678 1.192 ;
      RECT 4.718 0.698 4.786 0.832 ;
      RECT 4.61 0.068 4.678 0.292 ;
      RECT 5.042 0.878 5.11 1.012 ;
      RECT 5.042 0.248 5.11 0.472 ;
    LAYER v1 ;
      RECT 5.046 0.428 5.106 0.472 ;
      RECT 5.046 0.878 5.106 0.922 ;
      RECT 4.398 0.428 4.458 0.472 ;
      RECT 4.398 0.878 4.458 0.922 ;
      RECT 4.29 0.518 4.35 0.562 ;
      RECT 4.29 0.788 4.35 0.832 ;
      RECT 4.182 0.428 4.242 0.472 ;
      RECT 4.182 0.878 4.242 0.922 ;
      RECT 3.642 0.518 3.702 0.562 ;
      RECT 3.642 0.788 3.702 0.832 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 3.534 0.878 3.594 0.922 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 2.022 0.788 2.082 0.832 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 1.59 0.878 1.65 0.922 ;
      RECT 1.482 0.518 1.542 0.562 ;
      RECT 1.482 0.788 1.542 0.832 ;
      RECT 0.942 0.428 1.002 0.472 ;
      RECT 0.942 0.878 1.002 0.922 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.834 0.788 0.894 0.832 ;
      RECT 0.726 0.428 0.786 0.472 ;
      RECT 0.726 0.878 0.786 0.922 ;
      RECT 0.078 0.428 0.138 0.472 ;
      RECT 0.078 0.878 0.138 0.922 ;
    LAYER v0 ;
      RECT 5.042 0.293 5.11 0.337 ;
      RECT 5.042 0.923 5.11 0.967 ;
      RECT 4.826 0.088 4.894 0.132 ;
      RECT 4.826 0.498 4.894 0.542 ;
      RECT 4.826 0.718 4.894 0.762 ;
      RECT 4.826 1.128 4.894 1.172 ;
      RECT 4.61 0.088 4.678 0.132 ;
      RECT 4.61 1.128 4.678 1.172 ;
      RECT 4.502 0.498 4.57 0.542 ;
      RECT 4.502 0.718 4.57 0.762 ;
      RECT 4.394 0.363 4.462 0.407 ;
      RECT 4.394 0.853 4.462 0.897 ;
      RECT 4.286 0.068 4.354 0.112 ;
      RECT 4.286 0.158 4.354 0.202 ;
      RECT 4.286 0.498 4.354 0.542 ;
      RECT 4.286 0.718 4.354 0.762 ;
      RECT 4.286 1.058 4.354 1.102 ;
      RECT 4.286 1.148 4.354 1.192 ;
      RECT 4.178 0.248 4.246 0.292 ;
      RECT 4.178 0.498 4.246 0.542 ;
      RECT 4.178 0.718 4.246 0.762 ;
      RECT 4.178 0.968 4.246 1.012 ;
      RECT 3.854 0.403 3.922 0.447 ;
      RECT 3.854 0.813 3.922 0.857 ;
      RECT 3.746 0.068 3.814 0.112 ;
      RECT 3.746 1.148 3.814 1.192 ;
      RECT 3.638 0.158 3.706 0.202 ;
      RECT 3.638 0.293 3.706 0.337 ;
      RECT 3.638 0.923 3.706 0.967 ;
      RECT 3.638 1.058 3.706 1.102 ;
      RECT 3.53 0.383 3.598 0.427 ;
      RECT 3.53 0.833 3.598 0.877 ;
      RECT 3.422 0.518 3.49 0.562 ;
      RECT 3.422 0.718 3.49 0.762 ;
      RECT 3.314 0.088 3.382 0.132 ;
      RECT 3.206 1.128 3.274 1.172 ;
      RECT 2.99 0.068 3.058 0.112 ;
      RECT 2.99 0.2025 3.058 0.2465 ;
      RECT 2.99 1.0135 3.058 1.0575 ;
      RECT 2.882 0.428 2.95 0.472 ;
      RECT 2.882 0.518 2.95 0.562 ;
      RECT 2.882 0.698 2.95 0.742 ;
      RECT 2.882 0.788 2.95 0.832 ;
      RECT 2.882 1.148 2.95 1.192 ;
      RECT 2.558 0.698 2.626 0.742 ;
      RECT 2.45 0.518 2.518 0.562 ;
      RECT 2.45 0.788 2.518 0.832 ;
      RECT 2.45 1.148 2.518 1.192 ;
      RECT 2.342 0.068 2.41 0.112 ;
      RECT 2.342 0.2025 2.41 0.2465 ;
      RECT 2.342 1.0135 2.41 1.0575 ;
      RECT 2.018 0.2025 2.086 0.2465 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 2.018 0.808 2.086 0.852 ;
      RECT 2.018 1.0135 2.086 1.0575 ;
      RECT 1.91 0.088 1.978 0.132 ;
      RECT 1.802 1.128 1.87 1.172 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.694 0.718 1.762 0.762 ;
      RECT 1.586 0.3835 1.654 0.4275 ;
      RECT 1.586 0.8325 1.654 0.8765 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.478 0.923 1.546 0.967 ;
      RECT 1.478 1.058 1.546 1.102 ;
      RECT 1.478 1.148 1.546 1.192 ;
      RECT 1.262 0.377 1.33 0.421 ;
      RECT 1.262 0.839 1.33 0.883 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.938 0.718 1.006 0.762 ;
      RECT 0.938 0.968 1.006 1.012 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.498 0.898 0.542 ;
      RECT 0.83 0.718 0.898 0.762 ;
      RECT 0.83 1.058 0.898 1.102 ;
      RECT 0.83 1.148 0.898 1.192 ;
      RECT 0.722 0.363 0.79 0.407 ;
      RECT 0.722 0.853 0.79 0.897 ;
      RECT 0.614 0.498 0.682 0.542 ;
      RECT 0.614 0.718 0.682 0.762 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.506 1.128 0.574 1.172 ;
      RECT 0.29 0.088 0.358 0.132 ;
      RECT 0.29 0.498 0.358 0.542 ;
      RECT 0.29 0.718 0.358 0.762 ;
      RECT 0.29 1.128 0.358 1.172 ;
      RECT 0.074 0.293 0.142 0.337 ;
      RECT 0.074 0.923 0.142 0.967 ;
    LAYER m1 ;
      RECT 0.29 0.698 0.358 1.192 ;
      RECT 0.358 0.968 0.506 1.012 ;
      RECT 0.506 0.968 0.574 1.192 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.682 1.148 1.006 1.192 ;
      RECT 0.79 1.058 1.006 1.102 ;
      RECT 0.79 0.158 1.006 0.202 ;
      RECT 0.682 0.068 1.006 0.112 ;
      RECT 1.262 0.788 1.33 1.012 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.586 0.788 1.654 1.102 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.694 0.698 1.762 1.192 ;
      RECT 1.694 0.068 1.762 0.382 ;
      RECT 1.586 0.518 1.802 0.562 ;
      RECT 1.762 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.698 2.342 0.742 ;
      RECT 2.342 0.698 2.41 1.102 ;
      RECT 2.41 0.788 2.626 0.832 ;
      RECT 1.978 0.518 2.342 0.562 ;
      RECT 2.342 0.158 2.41 0.562 ;
      RECT 2.41 0.518 2.626 0.562 ;
      RECT 2.558 1.058 2.626 1.192 ;
      RECT 2.626 1.058 2.666 1.102 ;
      RECT 2.45 0.698 2.666 0.742 ;
      RECT 2.666 0.698 2.734 1.102 ;
      RECT 2.734 1.058 2.774 1.102 ;
      RECT 2.774 1.058 2.842 1.192 ;
      RECT 2.842 1.148 3.058 1.192 ;
      RECT 2.734 0.698 3.058 0.742 ;
      RECT 2.558 0.068 2.626 0.202 ;
      RECT 2.626 0.158 2.666 0.202 ;
      RECT 2.666 0.158 2.734 0.562 ;
      RECT 2.734 0.158 2.774 0.202 ;
      RECT 2.774 0.068 2.842 0.202 ;
      RECT 2.734 0.518 3.058 0.562 ;
      RECT 2.842 0.068 3.166 0.112 ;
      RECT 2.99 0.788 3.058 1.102 ;
      RECT 3.058 0.788 3.206 0.832 ;
      RECT 3.206 0.788 3.274 1.192 ;
      RECT 2.99 0.158 3.058 0.472 ;
      RECT 3.058 0.428 3.206 0.472 ;
      RECT 3.206 0.248 3.274 0.472 ;
      RECT 3.274 0.248 3.314 0.292 ;
      RECT 3.314 0.068 3.382 0.292 ;
      RECT 3.598 1.058 3.726 1.102 ;
      RECT 3.598 0.158 3.726 0.202 ;
      RECT 3.49 1.148 3.922 1.192 ;
      RECT 3.382 0.338 3.422 0.382 ;
      RECT 3.422 0.068 3.49 0.382 ;
      RECT 3.382 0.518 3.598 0.562 ;
      RECT 3.49 0.068 3.922 0.112 ;
      RECT 3.922 0.968 4.354 1.012 ;
      RECT 3.922 0.248 4.354 0.292 ;
      RECT 4.394 0.788 4.462 1.102 ;
      RECT 4.394 0.158 4.462 0.472 ;
      RECT 4.502 0.698 4.57 1.192 ;
      RECT 4.502 0.068 4.57 0.562 ;
      RECT 4.678 0.968 4.826 1.012 ;
      RECT 4.826 0.698 4.894 1.192 ;
      RECT 4.678 0.248 4.826 0.292 ;
      RECT 4.826 0.068 4.894 0.562 ;
  END
END b15fqy403hn1d02x5

MACRO b15fqy403hn1d03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy403hn1d03x5 0 0 ;
  SIZE 5.4 BY 1.26 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN d3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.878 2.95 1.012 ;
      LAYER m2 ;
        RECT 2.848 0.878 3.524 0.922 ;
      LAYER v1 ;
        RECT 2.886 0.878 2.946 0.922 ;
      LAYER v0 ;
        RECT 2.882 0.923 2.95 0.967 ;
    END
  END d3
  PIN d4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.878 2.734 1.012 ;
      LAYER m2 ;
        RECT 2.324 0.878 2.768 0.922 ;
      LAYER v1 ;
        RECT 2.67 0.878 2.73 0.922 ;
      LAYER v0 ;
        RECT 2.666 0.923 2.734 0.967 ;
    END
  END d4
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0288 LAYER m2 ;
      ANTENNAMAXAREACAR 2.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 4.83333325 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.036 LAYER m2 ;
      ANTENNAMAXAREACAR 1.10666675 LAYER m1 ;
      ANTENNAMAXAREACAR 3.22222225 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.826 0.698 4.894 0.922 ;
        RECT 4.07 0.698 4.138 0.832 ;
        RECT 1.262 0.698 1.33 0.832 ;
        RECT 0.506 0.698 0.574 0.922 ;
      LAYER m2 ;
        RECT 0.38 0.698 4.912 0.742 ;
      LAYER v1 ;
        RECT 0.51 0.698 0.57 0.742 ;
        RECT 1.266 0.698 1.326 0.742 ;
        RECT 4.074 0.698 4.134 0.742 ;
        RECT 4.83 0.698 4.89 0.742 ;
      LAYER v0 ;
        RECT 0.506 0.718 0.574 0.762 ;
        RECT 1.262 0.718 1.33 0.762 ;
        RECT 4.07 0.718 4.138 0.762 ;
        RECT 4.826 0.718 4.894 0.762 ;
    END
  END rb
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
      ANTENNAMAXAREACAR 2.7805555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 2.2244445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.158 3.058 0.382 ;
        RECT 2.558 0.158 2.626 0.382 ;
      LAYER m2 ;
        RECT 2.54 0.158 3.076 0.202 ;
      LAYER v1 ;
        RECT 2.562 0.158 2.622 0.202 ;
        RECT 2.994 0.158 3.054 0.202 ;
      LAYER v0 ;
        RECT 2.558 0.293 2.626 0.337 ;
        RECT 2.99 0.293 3.058 0.337 ;
    END
  END ssb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.788 2.086 1.012 ;
      LAYER v0 ;
        RECT 2.018 0.923 2.086 0.967 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.248 2.734 0.472 ;
      LAYER v0 ;
        RECT 2.666 0.293 2.734 0.337 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.248 2.95 0.382 ;
      LAYER v0 ;
        RECT 2.882 0.293 2.95 0.337 ;
    END
  END d2
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.403 0.142 0.447 ;
        RECT 0.074 0.223 0.142 0.267 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.258 0.158 5.326 0.562 ;
      LAYER v0 ;
        RECT 5.258 0.403 5.326 0.447 ;
        RECT 5.258 0.223 5.326 0.267 ;
    END
  END o2
  PIN o3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.258 0.698 5.326 1.102 ;
      LAYER v0 ;
        RECT 5.258 0.993 5.326 1.037 ;
        RECT 5.258 0.813 5.326 0.857 ;
    END
  END o3
  PIN o4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.698 0.142 1.102 ;
      LAYER v0 ;
        RECT 0.074 0.993 0.142 1.037 ;
        RECT 0.074 0.813 0.142 0.857 ;
    END
  END o4
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.382 ;
      LAYER v0 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.158 3.274 0.382 ;
      LAYER v0 ;
        RECT 3.206 0.293 3.274 0.337 ;
    END
  END si2
  PIN si3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.878 3.274 1.192 ;
      LAYER v0 ;
        RECT 3.206 0.923 3.274 0.967 ;
    END
  END si3
  PIN si4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.878 2.41 1.192 ;
      LAYER v0 ;
        RECT 2.342 0.923 2.41 0.967 ;
    END
  END si4
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.434 0.652 ;
        RECT 5.15 0.338 5.218 0.922 ;
        RECT 4.718 0.338 4.786 0.922 ;
        RECT 4.178 0.338 4.246 0.922 ;
        RECT 3.854 0.338 3.922 0.922 ;
        RECT 1.478 0.338 1.546 0.922 ;
        RECT 1.154 0.338 1.222 0.922 ;
        RECT 0.614 0.338 0.682 0.922 ;
        RECT 0.182 0.338 0.25 0.922 ;
      LAYER v0 ;
        RECT 0.182 0.813 0.25 0.857 ;
        RECT 0.182 0.403 0.25 0.447 ;
        RECT 0.614 0.853 0.682 0.897 ;
        RECT 0.614 0.383 0.682 0.427 ;
        RECT 1.154 0.814 1.222 0.858 ;
        RECT 1.154 0.402 1.222 0.446 ;
        RECT 1.478 0.839 1.546 0.883 ;
        RECT 1.478 0.377 1.546 0.421 ;
        RECT 1.91 0.608 1.978 0.652 ;
        RECT 2.234 0.608 2.302 0.652 ;
        RECT 2.774 0.608 2.842 0.652 ;
        RECT 3.098 0.608 3.166 0.652 ;
        RECT 3.314 0.608 3.382 0.652 ;
        RECT 3.854 0.813 3.922 0.857 ;
        RECT 3.854 0.403 3.922 0.447 ;
        RECT 4.178 0.814 4.246 0.858 ;
        RECT 4.178 0.402 4.246 0.446 ;
        RECT 4.718 0.853 4.786 0.897 ;
        RECT 4.718 0.383 4.786 0.427 ;
        RECT 5.15 0.813 5.218 0.857 ;
        RECT 5.15 0.403 5.218 0.447 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.434 0.022 ;
        RECT 5.15 -0.022 5.218 0.292 ;
        RECT 4.826 -0.022 4.894 0.292 ;
        RECT 4.07 -0.022 4.138 0.202 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.234 -0.022 2.302 0.292 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.154 0.158 1.438 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
        RECT -0.034 1.238 5.434 1.282 ;
        RECT 5.15 0.968 5.218 1.282 ;
        RECT 4.826 0.968 4.894 1.282 ;
        RECT 4.07 1.058 4.138 1.282 ;
        RECT 3.422 0.968 3.49 1.282 ;
        RECT 2.774 1.148 2.842 1.282 ;
        RECT 2.234 0.968 2.302 1.282 ;
        RECT 2.018 1.058 2.086 1.282 ;
        RECT 1.37 1.058 1.438 1.282 ;
        RECT 1.154 1.058 1.438 1.102 ;
        RECT 0.506 0.968 0.574 1.282 ;
        RECT 0.182 0.968 0.25 1.282 ;
      LAYER v0 ;
        RECT 0.182 0.993 0.25 1.037 ;
        RECT 0.182 0.223 0.25 0.267 ;
        RECT 0.506 0.994 0.574 1.038 ;
        RECT 0.506 0.222 0.574 0.266 ;
        RECT 1.262 1.058 1.33 1.102 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.91 0.2025 1.978 0.2465 ;
        RECT 2.018 1.128 2.086 1.172 ;
        RECT 2.234 1.0135 2.302 1.0575 ;
        RECT 2.234 0.2025 2.302 0.2465 ;
        RECT 2.774 1.168 2.842 1.212 ;
        RECT 2.774 0.048 2.842 0.092 ;
        RECT 3.314 0.088 3.382 0.132 ;
        RECT 3.422 1.0375 3.49 1.0815 ;
        RECT 4.07 1.078 4.138 1.122 ;
        RECT 4.07 0.138 4.138 0.182 ;
        RECT 4.826 0.994 4.894 1.038 ;
        RECT 4.826 0.222 4.894 0.266 ;
        RECT 5.15 0.993 5.218 1.037 ;
        RECT 5.15 0.223 5.218 0.267 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.878 0.932 0.922 ;
      RECT 0.04 0.428 0.932 0.472 ;
      RECT 1.012 0.878 1.78 0.922 ;
      RECT 1.012 0.428 1.796 0.472 ;
      RECT 1.876 0.428 3.524 0.472 ;
      RECT 3.604 0.878 4.388 0.922 ;
      RECT 3.604 0.428 4.388 0.472 ;
      RECT 0.92 0.788 4.48 0.832 ;
      RECT 0.92 0.518 4.48 0.562 ;
      RECT 4.468 0.428 4.912 0.472 ;
      RECT 4.468 0.878 5.02 0.922 ;
    LAYER m1 ;
      RECT 0.29 0.788 0.358 1.102 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.398 0.698 0.466 0.922 ;
      RECT 0.506 0.698 0.574 0.922 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.938 0.698 1.006 0.832 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.83 0.788 0.898 1.102 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.046 0.698 1.114 0.922 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 0.938 0.968 1.37 1.012 ;
      RECT 1.262 0.698 1.33 0.832 ;
      RECT 0.938 0.248 1.37 0.292 ;
      RECT 1.478 1.058 1.694 1.102 ;
      RECT 1.586 0.788 1.654 1.012 ;
      RECT 1.586 0.248 1.654 0.562 ;
      RECT 1.478 0.158 1.694 0.202 ;
      RECT 1.478 1.148 1.802 1.192 ;
      RECT 1.478 0.068 1.802 0.112 ;
      RECT 1.91 0.698 1.978 1.192 ;
      RECT 2.126 0.788 2.194 1.102 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 2.558 0.158 2.626 0.382 ;
      RECT 2.666 0.878 2.734 1.012 ;
      RECT 2.018 0.068 2.086 0.562 ;
      RECT 2.45 1.148 2.666 1.192 ;
      RECT 2.882 0.878 2.95 1.012 ;
      RECT 2.99 0.158 3.058 0.382 ;
      RECT 2.342 0.068 2.666 0.112 ;
      RECT 2.882 0.788 3.098 0.832 ;
      RECT 2.882 0.428 3.098 0.472 ;
      RECT 3.638 0.788 3.706 1.102 ;
      RECT 3.746 0.788 3.814 1.012 ;
      RECT 3.746 0.248 3.814 0.562 ;
      RECT 3.638 0.158 3.706 0.472 ;
      RECT 3.53 0.698 3.598 1.192 ;
      RECT 3.422 0.338 3.49 0.562 ;
      RECT 3.962 0.698 4.03 1.012 ;
      RECT 4.07 0.698 4.138 0.832 ;
      RECT 4.286 0.698 4.354 0.922 ;
      RECT 4.286 0.428 4.354 0.562 ;
      RECT 3.962 0.248 4.03 0.562 ;
      RECT 4.394 0.698 4.462 0.832 ;
      RECT 4.394 0.428 4.462 0.562 ;
      RECT 4.286 1.058 4.502 1.102 ;
      RECT 4.286 0.158 4.502 0.202 ;
      RECT 4.394 1.148 4.61 1.192 ;
      RECT 4.394 0.068 4.61 0.112 ;
      RECT 4.826 0.698 4.894 0.922 ;
      RECT 4.826 0.338 4.894 0.472 ;
      RECT 4.934 0.788 5.002 0.922 ;
      RECT 5.042 0.788 5.11 1.102 ;
      RECT 5.042 0.158 5.11 0.472 ;
    LAYER v1 ;
      RECT 4.938 0.878 4.998 0.922 ;
      RECT 4.83 0.428 4.89 0.472 ;
      RECT 4.506 0.428 4.566 0.472 ;
      RECT 4.506 0.878 4.566 0.922 ;
      RECT 4.398 0.518 4.458 0.562 ;
      RECT 4.398 0.788 4.458 0.832 ;
      RECT 4.29 0.428 4.35 0.472 ;
      RECT 4.29 0.878 4.35 0.922 ;
      RECT 3.75 0.518 3.81 0.562 ;
      RECT 3.75 0.788 3.81 0.832 ;
      RECT 3.642 0.428 3.702 0.472 ;
      RECT 3.642 0.878 3.702 0.922 ;
      RECT 3.426 0.428 3.486 0.472 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 2.13 0.788 2.19 0.832 ;
      RECT 1.914 0.428 1.974 0.472 ;
      RECT 1.698 0.428 1.758 0.472 ;
      RECT 1.698 0.878 1.758 0.922 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.59 0.788 1.65 0.832 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 1.05 0.878 1.11 0.922 ;
      RECT 0.942 0.518 1.002 0.562 ;
      RECT 0.942 0.788 1.002 0.832 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.834 0.878 0.894 0.922 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.402 0.878 0.462 0.922 ;
    LAYER v0 ;
      RECT 5.042 0.223 5.11 0.267 ;
      RECT 5.042 0.403 5.11 0.447 ;
      RECT 5.042 0.813 5.11 0.857 ;
      RECT 5.042 0.993 5.11 1.037 ;
      RECT 4.934 0.813 5.002 0.857 ;
      RECT 4.826 0.383 4.894 0.427 ;
      RECT 4.61 0.498 4.678 0.542 ;
      RECT 4.61 0.718 4.678 0.762 ;
      RECT 4.502 0.068 4.57 0.112 ;
      RECT 4.502 0.363 4.57 0.407 ;
      RECT 4.502 0.853 4.57 0.897 ;
      RECT 4.502 1.148 4.57 1.192 ;
      RECT 4.394 0.158 4.462 0.202 ;
      RECT 4.394 0.498 4.462 0.542 ;
      RECT 4.394 0.718 4.462 0.762 ;
      RECT 4.394 1.058 4.462 1.102 ;
      RECT 4.286 0.248 4.354 0.292 ;
      RECT 4.286 0.498 4.354 0.542 ;
      RECT 4.286 0.718 4.354 0.762 ;
      RECT 4.286 0.968 4.354 1.012 ;
      RECT 3.962 0.403 4.03 0.447 ;
      RECT 3.962 0.813 4.03 0.857 ;
      RECT 3.854 0.068 3.922 0.112 ;
      RECT 3.854 1.148 3.922 1.192 ;
      RECT 3.746 0.158 3.814 0.202 ;
      RECT 3.746 0.293 3.814 0.337 ;
      RECT 3.746 0.923 3.814 0.967 ;
      RECT 3.746 1.058 3.814 1.102 ;
      RECT 3.638 0.383 3.706 0.427 ;
      RECT 3.638 0.833 3.706 0.877 ;
      RECT 3.53 0.518 3.598 0.562 ;
      RECT 3.53 0.718 3.598 0.762 ;
      RECT 3.422 0.088 3.49 0.132 ;
      RECT 3.314 1.128 3.382 1.172 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 3.098 0.2025 3.166 0.2465 ;
      RECT 3.098 1.0135 3.166 1.0575 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.99 0.518 3.058 0.562 ;
      RECT 2.99 0.698 3.058 0.742 ;
      RECT 2.99 0.788 3.058 0.832 ;
      RECT 2.99 1.148 3.058 1.192 ;
      RECT 2.666 0.698 2.734 0.742 ;
      RECT 2.558 0.518 2.626 0.562 ;
      RECT 2.558 0.788 2.626 0.832 ;
      RECT 2.558 1.148 2.626 1.192 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.45 0.2025 2.518 0.2465 ;
      RECT 2.45 1.0135 2.518 1.0575 ;
      RECT 2.126 0.2025 2.194 0.2465 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 2.126 0.808 2.194 0.852 ;
      RECT 2.126 1.0135 2.194 1.0575 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 1.91 1.128 1.978 1.172 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.802 0.718 1.87 0.762 ;
      RECT 1.694 0.3835 1.762 0.4275 ;
      RECT 1.694 0.8325 1.762 0.8765 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.586 0.923 1.654 0.967 ;
      RECT 1.586 1.058 1.654 1.102 ;
      RECT 1.586 1.148 1.654 1.192 ;
      RECT 1.37 0.377 1.438 0.421 ;
      RECT 1.37 0.839 1.438 0.883 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.498 1.114 0.542 ;
      RECT 1.046 0.718 1.114 0.762 ;
      RECT 1.046 0.968 1.114 1.012 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.938 0.718 1.006 0.762 ;
      RECT 0.938 1.058 1.006 1.102 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.83 0.363 0.898 0.407 ;
      RECT 0.83 0.853 0.898 0.897 ;
      RECT 0.83 1.148 0.898 1.192 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.722 0.718 0.79 0.762 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.398 0.813 0.466 0.857 ;
      RECT 0.29 0.223 0.358 0.267 ;
      RECT 0.29 0.403 0.358 0.447 ;
      RECT 0.29 0.813 0.358 0.857 ;
      RECT 0.29 0.993 0.358 1.037 ;
    LAYER m1 ;
      RECT 0.722 0.698 0.79 1.192 ;
      RECT 0.79 1.148 1.006 1.192 ;
      RECT 0.79 0.068 1.006 0.112 ;
      RECT 0.898 1.058 1.114 1.102 ;
      RECT 0.898 0.158 1.114 0.202 ;
      RECT 1.37 0.788 1.438 1.012 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.694 0.788 1.762 1.102 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.802 0.698 1.87 1.192 ;
      RECT 1.802 0.068 1.87 0.382 ;
      RECT 1.694 0.518 1.91 0.562 ;
      RECT 1.87 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.978 0.698 2.45 0.742 ;
      RECT 2.45 0.698 2.518 1.102 ;
      RECT 2.518 0.788 2.734 0.832 ;
      RECT 2.086 0.518 2.45 0.562 ;
      RECT 2.45 0.158 2.518 0.562 ;
      RECT 2.518 0.518 2.734 0.562 ;
      RECT 2.666 1.058 2.734 1.192 ;
      RECT 2.734 1.058 2.774 1.102 ;
      RECT 2.558 0.698 2.774 0.742 ;
      RECT 2.774 0.698 2.842 1.102 ;
      RECT 2.842 1.058 2.882 1.102 ;
      RECT 2.882 1.058 2.95 1.192 ;
      RECT 2.95 1.148 3.166 1.192 ;
      RECT 2.842 0.698 3.166 0.742 ;
      RECT 2.666 0.068 2.734 0.202 ;
      RECT 2.734 0.158 2.774 0.202 ;
      RECT 2.774 0.158 2.842 0.562 ;
      RECT 2.842 0.158 2.882 0.202 ;
      RECT 2.882 0.068 2.95 0.202 ;
      RECT 2.842 0.518 3.166 0.562 ;
      RECT 2.95 0.068 3.274 0.112 ;
      RECT 3.098 0.788 3.166 1.102 ;
      RECT 3.166 0.788 3.314 0.832 ;
      RECT 3.314 0.788 3.382 1.192 ;
      RECT 3.098 0.158 3.166 0.472 ;
      RECT 3.166 0.428 3.314 0.472 ;
      RECT 3.314 0.248 3.382 0.472 ;
      RECT 3.382 0.248 3.422 0.292 ;
      RECT 3.422 0.068 3.49 0.292 ;
      RECT 3.706 1.058 3.834 1.102 ;
      RECT 3.706 0.158 3.834 0.202 ;
      RECT 3.598 1.148 4.03 1.192 ;
      RECT 3.49 0.338 3.53 0.382 ;
      RECT 3.53 0.068 3.598 0.382 ;
      RECT 3.49 0.518 3.706 0.562 ;
      RECT 3.598 0.068 4.03 0.112 ;
      RECT 4.03 0.968 4.462 1.012 ;
      RECT 4.03 0.248 4.462 0.292 ;
      RECT 4.502 0.788 4.57 1.102 ;
      RECT 4.502 0.158 4.57 0.472 ;
      RECT 4.61 0.698 4.678 1.192 ;
      RECT 4.61 0.068 4.678 0.562 ;
  END
END b15fqy403hn1d03x5

MACRO b15fqy403hn1d04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15fqy403hn1d04x5 0 0 ;
  SIZE 5.616 BY 1.26 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN d3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.878 3.058 1.012 ;
      LAYER m2 ;
        RECT 2.956 0.878 3.632 0.922 ;
      LAYER v1 ;
        RECT 2.994 0.878 3.054 0.922 ;
      LAYER v0 ;
        RECT 2.99 0.923 3.058 0.967 ;
    END
  END d3
  PIN d4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0036 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 3.248889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.878 2.842 1.012 ;
      LAYER m2 ;
        RECT 2.432 0.878 2.876 0.922 ;
      LAYER v1 ;
        RECT 2.778 0.878 2.838 0.922 ;
      LAYER v0 ;
        RECT 2.774 0.923 2.842 0.967 ;
    END
  END d4
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.036 LAYER m2 ;
      ANTENNAMAXAREACAR 3.0681945 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAGATEAREA 0.0459 LAYER m2 ;
      ANTENNAMAXAREACAR 2.727284 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.69530875 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 5.042 0.698 5.11 0.922 ;
        RECT 4.178 0.878 4.462 0.922 ;
        RECT 4.394 0.698 4.462 0.922 ;
        RECT 1.154 0.878 1.438 0.922 ;
        RECT 1.154 0.698 1.222 0.922 ;
        RECT 0.506 0.698 0.574 0.922 ;
      LAYER m2 ;
        RECT 0.38 0.698 5.128 0.742 ;
      LAYER v1 ;
        RECT 0.51 0.698 0.57 0.742 ;
        RECT 1.158 0.698 1.218 0.742 ;
        RECT 4.398 0.698 4.458 0.742 ;
        RECT 5.046 0.698 5.106 0.742 ;
      LAYER v0 ;
        RECT 0.506 0.718 0.574 0.762 ;
        RECT 1.262 0.878 1.33 0.922 ;
        RECT 4.286 0.878 4.354 0.922 ;
        RECT 5.042 0.718 5.11 0.762 ;
    END
  END rb
  PIN ssb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
      ANTENNAMAXAREACAR 2.7805555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAGATEAREA 0.018 LAYER m2 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
      ANTENNAMAXAREACAR 2.2244445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.62577775 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.158 3.166 0.382 ;
        RECT 2.666 0.158 2.734 0.382 ;
      LAYER m2 ;
        RECT 2.648 0.158 3.184 0.202 ;
      LAYER v1 ;
        RECT 2.67 0.158 2.73 0.202 ;
        RECT 3.102 0.158 3.162 0.202 ;
      LAYER v0 ;
        RECT 2.666 0.293 2.734 0.337 ;
        RECT 3.098 0.293 3.166 0.337 ;
    END
  END ssb
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.788 2.194 1.012 ;
      LAYER v0 ;
        RECT 2.126 0.923 2.194 0.967 ;
    END
  END clk
  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.248 2.842 0.472 ;
      LAYER v0 ;
        RECT 2.774 0.293 2.842 0.337 ;
    END
  END d1
  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.99 0.248 3.058 0.382 ;
      LAYER v0 ;
        RECT 2.99 0.293 3.058 0.337 ;
    END
  END d2
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.158 0.142 0.202 ;
    END
  END o1
  PIN o2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.474 0.068 5.542 0.562 ;
      LAYER v0 ;
        RECT 5.474 0.4285 5.542 0.4725 ;
        RECT 5.474 0.158 5.542 0.202 ;
    END
  END o2
  PIN o3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.474 0.698 5.542 1.192 ;
      LAYER v0 ;
        RECT 5.474 1.058 5.542 1.102 ;
        RECT 5.474 0.813 5.542 0.857 ;
    END
  END o3
  PIN o4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.698 0.142 1.192 ;
      LAYER v0 ;
        RECT 0.074 1.058 0.142 1.102 ;
        RECT 0.074 0.788 0.142 0.832 ;
    END
  END o4
  PIN si1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.158 2.518 0.382 ;
      LAYER v0 ;
        RECT 2.45 0.293 2.518 0.337 ;
    END
  END si1
  PIN si2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.158 3.382 0.382 ;
      LAYER v0 ;
        RECT 3.314 0.293 3.382 0.337 ;
    END
  END si2
  PIN si3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.878 3.382 1.192 ;
      LAYER v0 ;
        RECT 3.314 0.923 3.382 0.967 ;
    END
  END si3
  PIN si4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.878 2.518 1.192 ;
      LAYER v0 ;
        RECT 2.45 0.923 2.518 0.967 ;
    END
  END si4
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.65 0.652 ;
        RECT 5.366 0.338 5.434 0.922 ;
        RECT 4.934 0.338 5.002 0.922 ;
        RECT 4.286 0.428 4.354 0.832 ;
        RECT 3.962 0.338 4.03 0.922 ;
        RECT 1.586 0.338 1.654 0.922 ;
        RECT 1.262 0.428 1.33 0.832 ;
        RECT 0.614 0.338 0.682 0.922 ;
        RECT 0.182 0.338 0.25 0.922 ;
      LAYER v0 ;
        RECT 0.182 0.788 0.25 0.832 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.614 0.853 0.682 0.897 ;
        RECT 0.614 0.383 0.682 0.427 ;
        RECT 1.262 0.743 1.33 0.787 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.586 0.813 1.654 0.857 ;
        RECT 1.586 0.403 1.654 0.447 ;
        RECT 2.018 0.608 2.086 0.652 ;
        RECT 2.342 0.608 2.41 0.652 ;
        RECT 2.882 0.608 2.95 0.652 ;
        RECT 3.206 0.608 3.274 0.652 ;
        RECT 3.422 0.608 3.49 0.652 ;
        RECT 3.962 0.813 4.03 0.857 ;
        RECT 3.962 0.403 4.03 0.447 ;
        RECT 4.286 0.743 4.354 0.787 ;
        RECT 4.286 0.448 4.354 0.492 ;
        RECT 4.934 0.853 5.002 0.897 ;
        RECT 4.934 0.383 5.002 0.427 ;
        RECT 5.366 0.813 5.434 0.857 ;
        RECT 5.366 0.4285 5.434 0.4725 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.65 0.022 ;
        RECT 5.366 -0.022 5.434 0.292 ;
        RECT 5.042 -0.022 5.11 0.292 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.342 -0.022 2.41 0.292 ;
        RECT 2.018 -0.022 2.086 0.292 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
        RECT -0.034 1.238 5.65 1.282 ;
        RECT 5.366 0.968 5.434 1.282 ;
        RECT 5.042 0.968 5.11 1.282 ;
        RECT 4.178 1.148 4.246 1.282 ;
        RECT 3.53 0.968 3.598 1.282 ;
        RECT 2.882 1.148 2.95 1.282 ;
        RECT 2.342 0.968 2.41 1.282 ;
        RECT 2.126 1.058 2.194 1.282 ;
        RECT 1.37 1.148 1.438 1.282 ;
        RECT 0.506 0.968 0.574 1.282 ;
        RECT 0.182 0.968 0.25 1.282 ;
      LAYER v0 ;
        RECT 0.182 1.058 0.25 1.102 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.506 0.994 0.574 1.038 ;
        RECT 0.506 0.222 0.574 0.266 ;
        RECT 1.37 1.168 1.438 1.212 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 2.018 0.2025 2.086 0.2465 ;
        RECT 2.126 1.128 2.194 1.172 ;
        RECT 2.342 1.0135 2.41 1.0575 ;
        RECT 2.342 0.2025 2.41 0.2465 ;
        RECT 2.882 1.168 2.95 1.212 ;
        RECT 2.882 0.048 2.95 0.092 ;
        RECT 3.422 0.088 3.49 0.132 ;
        RECT 3.53 1.0375 3.598 1.0815 ;
        RECT 4.178 1.168 4.246 1.212 ;
        RECT 4.178 0.048 4.246 0.092 ;
        RECT 5.042 0.994 5.11 1.038 ;
        RECT 5.042 0.203 5.11 0.247 ;
        RECT 5.366 1.058 5.434 1.102 ;
        RECT 5.366 0.158 5.434 0.202 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.878 0.932 0.922 ;
      RECT 0.04 0.428 0.932 0.472 ;
      RECT 1.012 0.878 1.888 0.922 ;
      RECT 1.012 0.428 1.904 0.472 ;
      RECT 1.984 0.428 3.632 0.472 ;
      RECT 3.712 0.878 4.604 0.922 ;
      RECT 3.712 0.428 4.604 0.472 ;
      RECT 0.92 0.788 4.696 0.832 ;
      RECT 0.92 0.518 4.696 0.562 ;
      RECT 4.684 0.428 5.128 0.472 ;
      RECT 4.684 0.878 5.236 0.922 ;
    LAYER m1 ;
      RECT 0.29 0.698 0.358 1.192 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.398 0.788 0.466 1.012 ;
      RECT 0.506 0.698 0.574 0.922 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 0.938 0.698 1.006 0.832 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.046 0.698 1.114 0.922 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.154 0.698 1.222 0.922 ;
      RECT 1.046 0.968 1.478 1.012 ;
      RECT 1.046 0.248 1.478 0.292 ;
      RECT 1.586 1.058 1.802 1.102 ;
      RECT 1.694 0.788 1.762 1.012 ;
      RECT 1.694 0.248 1.762 0.562 ;
      RECT 1.586 0.158 1.802 0.202 ;
      RECT 0.722 0.698 0.79 1.192 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 2.018 0.698 2.086 1.192 ;
      RECT 2.234 0.788 2.302 1.102 ;
      RECT 2.234 0.158 2.302 0.472 ;
      RECT 2.666 0.158 2.734 0.382 ;
      RECT 2.774 0.878 2.842 1.012 ;
      RECT 2.126 0.068 2.194 0.562 ;
      RECT 2.558 1.148 2.774 1.192 ;
      RECT 2.99 0.878 3.058 1.012 ;
      RECT 3.098 0.158 3.166 0.382 ;
      RECT 2.45 0.068 2.774 0.112 ;
      RECT 2.99 0.788 3.206 0.832 ;
      RECT 2.99 0.428 3.206 0.472 ;
      RECT 3.746 0.788 3.814 1.102 ;
      RECT 3.854 0.698 3.922 1.012 ;
      RECT 3.854 0.248 3.922 0.562 ;
      RECT 3.746 0.158 3.814 0.472 ;
      RECT 4.178 0.878 4.394 0.922 ;
      RECT 4.07 0.788 4.138 1.012 ;
      RECT 4.07 0.248 4.138 0.472 ;
      RECT 4.502 0.698 4.57 0.922 ;
      RECT 4.502 0.428 4.57 0.562 ;
      RECT 4.502 1.058 4.718 1.102 ;
      RECT 4.61 0.698 4.678 0.832 ;
      RECT 4.61 0.428 4.678 0.562 ;
      RECT 4.502 0.158 4.718 0.202 ;
      RECT 3.638 0.698 3.706 1.192 ;
      RECT 3.53 0.338 3.598 0.562 ;
      RECT 5.042 0.698 5.11 0.922 ;
      RECT 5.042 0.338 5.11 0.472 ;
      RECT 5.15 0.788 5.218 0.922 ;
      RECT 5.258 0.788 5.326 1.192 ;
      RECT 5.258 0.068 5.326 0.562 ;
    LAYER v1 ;
      RECT 5.154 0.878 5.214 0.922 ;
      RECT 5.046 0.428 5.106 0.472 ;
      RECT 4.722 0.428 4.782 0.472 ;
      RECT 4.722 0.878 4.782 0.922 ;
      RECT 4.614 0.518 4.674 0.562 ;
      RECT 4.614 0.788 4.674 0.832 ;
      RECT 4.506 0.428 4.566 0.472 ;
      RECT 4.506 0.878 4.566 0.922 ;
      RECT 3.858 0.518 3.918 0.562 ;
      RECT 3.858 0.788 3.918 0.832 ;
      RECT 3.75 0.428 3.81 0.472 ;
      RECT 3.75 0.878 3.81 0.922 ;
      RECT 3.534 0.428 3.594 0.472 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 2.238 0.788 2.298 0.832 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.806 0.878 1.866 0.922 ;
      RECT 1.698 0.518 1.758 0.562 ;
      RECT 1.698 0.788 1.758 0.832 ;
      RECT 1.05 0.428 1.11 0.472 ;
      RECT 1.05 0.878 1.11 0.922 ;
      RECT 0.942 0.518 1.002 0.562 ;
      RECT 0.942 0.788 1.002 0.832 ;
      RECT 0.834 0.428 0.894 0.472 ;
      RECT 0.834 0.878 0.894 0.922 ;
      RECT 0.51 0.428 0.57 0.472 ;
      RECT 0.402 0.878 0.462 0.922 ;
    LAYER v0 ;
      RECT 5.258 0.158 5.326 0.202 ;
      RECT 5.258 0.4285 5.326 0.4725 ;
      RECT 5.258 0.813 5.326 0.857 ;
      RECT 5.258 1.058 5.326 1.102 ;
      RECT 5.15 0.813 5.218 0.857 ;
      RECT 5.042 0.383 5.11 0.427 ;
      RECT 4.826 0.498 4.894 0.542 ;
      RECT 4.826 0.718 4.894 0.762 ;
      RECT 4.718 0.363 4.786 0.407 ;
      RECT 4.718 0.853 4.786 0.897 ;
      RECT 4.61 0.068 4.678 0.112 ;
      RECT 4.61 0.158 4.678 0.202 ;
      RECT 4.61 0.498 4.678 0.542 ;
      RECT 4.61 0.718 4.678 0.762 ;
      RECT 4.61 1.058 4.678 1.102 ;
      RECT 4.61 1.148 4.678 1.192 ;
      RECT 4.502 0.498 4.57 0.542 ;
      RECT 4.502 0.718 4.57 0.762 ;
      RECT 4.394 0.248 4.462 0.292 ;
      RECT 4.394 0.968 4.462 1.012 ;
      RECT 4.07 0.403 4.138 0.447 ;
      RECT 4.07 0.813 4.138 0.857 ;
      RECT 3.962 0.068 4.03 0.112 ;
      RECT 3.962 1.148 4.03 1.192 ;
      RECT 3.854 0.158 3.922 0.202 ;
      RECT 3.854 0.293 3.922 0.337 ;
      RECT 3.854 0.923 3.922 0.967 ;
      RECT 3.854 1.058 3.922 1.102 ;
      RECT 3.746 0.383 3.814 0.427 ;
      RECT 3.746 0.833 3.814 0.877 ;
      RECT 3.638 0.518 3.706 0.562 ;
      RECT 3.638 0.718 3.706 0.762 ;
      RECT 3.53 0.088 3.598 0.132 ;
      RECT 3.422 1.128 3.49 1.172 ;
      RECT 3.206 0.068 3.274 0.112 ;
      RECT 3.206 0.2025 3.274 0.2465 ;
      RECT 3.206 1.0135 3.274 1.0575 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 3.098 0.518 3.166 0.562 ;
      RECT 3.098 0.698 3.166 0.742 ;
      RECT 3.098 0.788 3.166 0.832 ;
      RECT 3.098 1.148 3.166 1.192 ;
      RECT 2.774 0.698 2.842 0.742 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.666 0.788 2.734 0.832 ;
      RECT 2.666 1.148 2.734 1.192 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.558 0.2025 2.626 0.2465 ;
      RECT 2.558 1.0135 2.626 1.0575 ;
      RECT 2.234 0.2025 2.302 0.2465 ;
      RECT 2.234 0.408 2.302 0.452 ;
      RECT 2.234 0.808 2.302 0.852 ;
      RECT 2.234 1.0135 2.302 1.0575 ;
      RECT 2.126 0.088 2.194 0.132 ;
      RECT 2.018 1.128 2.086 1.172 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.91 0.718 1.978 0.762 ;
      RECT 1.802 0.3835 1.87 0.4275 ;
      RECT 1.802 0.8325 1.87 0.8765 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.694 0.923 1.762 0.967 ;
      RECT 1.694 1.058 1.762 1.102 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.586 1.148 1.654 1.192 ;
      RECT 1.478 0.403 1.546 0.447 ;
      RECT 1.478 0.813 1.546 0.857 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 1.154 0.968 1.222 1.012 ;
      RECT 1.046 0.498 1.114 0.542 ;
      RECT 1.046 0.718 1.114 0.762 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.498 1.006 0.542 ;
      RECT 0.938 0.718 1.006 0.762 ;
      RECT 0.938 1.058 1.006 1.102 ;
      RECT 0.938 1.148 1.006 1.192 ;
      RECT 0.83 0.363 0.898 0.407 ;
      RECT 0.83 0.853 0.898 0.897 ;
      RECT 0.722 0.498 0.79 0.542 ;
      RECT 0.722 0.718 0.79 0.762 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.398 0.898 0.466 0.942 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.29 0.788 0.358 0.832 ;
      RECT 0.29 1.058 0.358 1.102 ;
    LAYER m1 ;
      RECT 0.83 0.788 0.898 1.102 ;
      RECT 0.898 1.058 1.114 1.102 ;
      RECT 0.898 0.158 1.114 0.202 ;
      RECT 1.222 0.878 1.438 0.922 ;
      RECT 1.478 0.788 1.546 1.012 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.802 0.788 1.87 1.102 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 0.79 1.148 1.262 1.192 ;
      RECT 1.262 1.058 1.33 1.192 ;
      RECT 1.33 1.058 1.478 1.102 ;
      RECT 1.478 1.058 1.546 1.192 ;
      RECT 1.546 1.148 1.91 1.192 ;
      RECT 1.91 0.698 1.978 1.192 ;
      RECT 0.79 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.158 1.478 0.202 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 1.546 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.382 ;
      RECT 1.802 0.518 2.018 0.562 ;
      RECT 1.978 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.086 0.698 2.558 0.742 ;
      RECT 2.558 0.698 2.626 1.102 ;
      RECT 2.626 0.788 2.842 0.832 ;
      RECT 2.194 0.518 2.558 0.562 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 2.626 0.518 2.842 0.562 ;
      RECT 2.774 1.058 2.842 1.192 ;
      RECT 2.842 1.058 2.882 1.102 ;
      RECT 2.666 0.698 2.882 0.742 ;
      RECT 2.882 0.698 2.95 1.102 ;
      RECT 2.95 1.058 2.99 1.102 ;
      RECT 2.99 1.058 3.058 1.192 ;
      RECT 3.058 1.148 3.274 1.192 ;
      RECT 2.95 0.698 3.274 0.742 ;
      RECT 2.774 0.068 2.842 0.202 ;
      RECT 2.842 0.158 2.882 0.202 ;
      RECT 2.882 0.158 2.95 0.562 ;
      RECT 2.95 0.158 2.99 0.202 ;
      RECT 2.99 0.068 3.058 0.202 ;
      RECT 2.95 0.518 3.274 0.562 ;
      RECT 3.058 0.068 3.382 0.112 ;
      RECT 3.206 0.788 3.274 1.102 ;
      RECT 3.274 0.788 3.422 0.832 ;
      RECT 3.422 0.788 3.49 1.192 ;
      RECT 3.206 0.158 3.274 0.472 ;
      RECT 3.274 0.428 3.422 0.472 ;
      RECT 3.422 0.248 3.49 0.472 ;
      RECT 3.49 0.248 3.53 0.292 ;
      RECT 3.53 0.068 3.598 0.292 ;
      RECT 3.814 1.058 4.03 1.102 ;
      RECT 3.814 0.158 4.03 0.202 ;
      RECT 4.394 0.698 4.462 0.922 ;
      RECT 4.138 0.968 4.57 1.012 ;
      RECT 4.138 0.248 4.57 0.292 ;
      RECT 4.718 0.788 4.786 1.102 ;
      RECT 4.718 0.158 4.786 0.472 ;
      RECT 3.706 1.148 4.07 1.192 ;
      RECT 4.07 1.058 4.138 1.192 ;
      RECT 4.138 1.058 4.286 1.102 ;
      RECT 4.286 1.058 4.354 1.192 ;
      RECT 4.354 1.148 4.826 1.192 ;
      RECT 4.826 0.698 4.894 1.192 ;
      RECT 3.598 0.338 3.638 0.382 ;
      RECT 3.638 0.068 3.706 0.382 ;
      RECT 3.598 0.518 3.814 0.562 ;
      RECT 3.706 0.068 4.07 0.112 ;
      RECT 4.07 0.068 4.138 0.202 ;
      RECT 4.138 0.158 4.286 0.202 ;
      RECT 4.286 0.068 4.354 0.202 ;
      RECT 4.354 0.068 4.826 0.112 ;
      RECT 4.826 0.068 4.894 0.562 ;
  END
END b15fqy403hn1d04x5

MACRO b15lsn000hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn000hn1n02x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.65 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.382 ;
        RECT 0.398 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.222 0.292 ;
        RECT 1.154 0.068 1.222 0.292 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.383 1.114 0.427 ;
        RECT 1.154 0.113 1.222 0.157 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.83 0.473 0.898 0.517 ;
        RECT 1.154 0.488 1.222 0.532 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.722 0.203 0.79 0.247 ;
        RECT 1.046 0.113 1.114 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.938 0.068 1.006 0.562 ;
    LAYER v0 ;
      RECT 0.938 0.113 1.006 0.157 ;
      RECT 0.938 0.473 1.006 0.517 ;
      RECT 0.83 0.203 0.898 0.247 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.203 0.574 0.247 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.3405 0.142 0.3845 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.518 0.594 0.562 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.338 0.83 0.382 ;
      RECT 0.83 0.158 0.898 0.382 ;
  END
END b15lsn000hn1n02x5

MACRO b15lsn000hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn000hn1n03x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.75 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.898 0.382 ;
        RECT 0.614 0.068 0.682 0.382 ;
        RECT 0.398 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.158 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.3935 1.33 0.4375 ;
        RECT 1.262 0.178 1.33 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.154 0.3935 1.222 0.4375 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.83 0.1905 0.898 0.2345 ;
        RECT 1.154 0.178 1.222 0.222 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 1.046 0.158 1.114 0.472 ;
    LAYER v0 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 1.046 0.3935 1.114 0.4375 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.203 0.574 0.247 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.428 0.938 0.472 ;
      RECT 0.938 0.248 1.006 0.472 ;
  END
END b15lsn000hn1n03x5

MACRO b15lsn000hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn000hn1n04x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 5.32 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.9555555 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.594 0.338 0.79 0.382 ;
        RECT 0.722 0.068 0.79 0.382 ;
        RECT 0.486 0.068 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.338 0.358 0.382 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.562 ;
      LAYER v0 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.262 0.088 1.33 0.132 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.154 0.448 1.222 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.154 0.088 1.222 0.132 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 1.046 0.068 1.114 0.562 ;
    LAYER v0 ;
      RECT 1.046 0.088 1.114 0.132 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.518 0.594 0.562 ;
      RECT 0.466 0.248 0.682 0.292 ;
      RECT 0.466 0.428 0.83 0.472 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.338 0.938 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
  END
END b15lsn000hn1n04x5

MACRO b15lsn000hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn000hn1n06x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.7 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.53333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.898 0.382 ;
        RECT 0.614 0.068 0.682 0.382 ;
        RECT 0.398 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.158 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.3935 1.33 0.4375 ;
        RECT 1.262 0.178 1.33 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.154 0.3935 1.222 0.4375 ;
        RECT 1.37 0.3935 1.438 0.4375 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.83 0.1905 0.898 0.2345 ;
        RECT 1.154 0.178 1.222 0.222 ;
        RECT 1.37 0.178 1.438 0.222 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
    LAYER v0 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 1.046 0.3935 1.114 0.4375 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.203 0.574 0.247 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.428 0.938 0.472 ;
      RECT 0.938 0.248 1.006 0.472 ;
  END
END b15lsn000hn1n06x5

MACRO b15lsn000hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn000hn1n08x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.04 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.736 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.518 1.114 0.562 ;
        RECT 1.046 0.338 1.114 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.518 1.006 0.562 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.562 ;
      LAYER v0 ;
        RECT 1.262 0.43 1.33 0.474 ;
        RECT 1.262 0.163 1.33 0.207 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.614 0.428 0.81 0.472 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 1.154 0.43 1.222 0.474 ;
        RECT 1.37 0.43 1.438 0.474 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.154 0.163 1.222 0.207 ;
        RECT 1.37 0.163 1.438 0.207 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.29 0.248 0.358 0.562 ;
      RECT 0.702 0.338 0.938 0.382 ;
    LAYER v0 ;
      RECT 0.938 0.256 1.006 0.3 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.29 0.3155 0.358 0.3595 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 0.466 0.068 0.594 0.112 ;
      RECT 0.358 0.518 0.506 0.562 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.574 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 0.938 0.158 1.006 0.382 ;
  END
END b15lsn000hn1n08x5

MACRO b15lsn000hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn000hn1n12x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.287 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.73916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.222 0.562 ;
      LAYER v0 ;
        RECT 1.154 0.498 1.222 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.37 0.338 1.654 0.382 ;
        RECT 1.37 0.158 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.372 0.408 1.436 0.452 ;
        RECT 1.37 0.2015 1.438 0.2455 ;
        RECT 1.588 0.408 1.652 0.452 ;
        RECT 1.586 0.2015 1.654 0.2455 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.722 0.428 0.918 0.472 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.262 0.498 1.33 0.542 ;
        RECT 1.478 0.493 1.546 0.537 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.178 0.25 0.222 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.262 0.113 1.33 0.157 ;
        RECT 1.478 0.113 1.546 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.81 0.338 1.046 0.382 ;
      RECT 0.506 0.068 0.574 0.472 ;
    LAYER v0 ;
      RECT 1.048 0.088 1.112 0.132 ;
      RECT 1.048 0.408 1.112 0.452 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.506 0.408 0.574 0.452 ;
      RECT 0.398 0.293 0.466 0.337 ;
      RECT 0.29 0.178 0.358 0.222 ;
      RECT 0.29 0.408 0.358 0.452 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 0.682 0.248 1.026 0.292 ;
      RECT 1.046 0.338 1.114 0.472 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.79 0.158 1.046 0.202 ;
      RECT 1.046 0.068 1.114 0.202 ;
  END
END b15lsn000hn1n12x5

MACRO b15lsn000hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn000hn1n16x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.287 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.73916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.222 0.562 ;
      LAYER v0 ;
        RECT 1.154 0.498 1.222 0.542 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.37 0.338 1.654 0.382 ;
        RECT 1.37 0.158 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.372 0.408 1.436 0.452 ;
        RECT 1.37 0.194 1.438 0.238 ;
        RECT 1.588 0.408 1.652 0.452 ;
        RECT 1.586 0.194 1.654 0.238 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.722 0.428 0.918 0.472 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.262 0.498 1.33 0.542 ;
        RECT 1.478 0.493 1.546 0.537 ;
        RECT 1.694 0.493 1.762 0.537 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.262 0.113 1.33 0.157 ;
        RECT 1.478 0.113 1.546 0.157 ;
        RECT 1.694 0.113 1.762 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.81 0.338 1.046 0.382 ;
      RECT 0.506 0.158 0.574 0.472 ;
    LAYER v0 ;
      RECT 1.048 0.088 1.112 0.132 ;
      RECT 1.048 0.408 1.112 0.452 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.408 0.574 0.452 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.292 0.358 0.356 0.402 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.076 0.358 0.14 0.402 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 0.682 0.248 1.026 0.292 ;
      RECT 1.046 0.338 1.114 0.472 ;
      RECT 0.574 0.158 1.046 0.202 ;
      RECT 1.046 0.068 1.114 0.202 ;
  END
END b15lsn000hn1n16x5

MACRO b15lsn080hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn080hn1n02x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.53333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.7 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 0.79 0.562 ;
        RECT 0.722 0.158 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.383 1.33 0.427 ;
        RECT 1.262 0.138 1.33 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.938 0.383 1.006 0.427 ;
        RECT 1.154 0.383 1.222 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 1.046 0.068 1.114 0.472 ;
    LAYER v0 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.383 1.114 0.427 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.408 0.142 0.452 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.382 ;
  END
END b15lsn080hn1n02x5

MACRO b15lsn080hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn080hn1n03x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.53333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.7 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 0.79 0.562 ;
        RECT 0.722 0.158 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.408 1.33 0.452 ;
        RECT 1.262 0.133 1.33 0.177 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.154 0.408 1.222 0.452 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.938 0.133 1.006 0.177 ;
        RECT 1.154 0.133 1.222 0.177 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 1.046 0.068 1.114 0.472 ;
    LAYER v0 ;
      RECT 1.046 0.133 1.114 0.177 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.408 0.142 0.452 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.382 ;
  END
END b15lsn080hn1n03x5

MACRO b15lsn080hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn080hn1n04x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.53333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.7 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.898 0.292 ;
        RECT 0.398 0.518 0.682 0.562 ;
        RECT 0.614 0.248 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.158 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.3935 1.33 0.4375 ;
        RECT 1.262 0.202 1.33 0.246 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.83 0.388 0.898 0.432 ;
        RECT 1.154 0.492 1.222 0.536 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.154 0.116 1.222 0.16 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 1.046 0.158 1.114 0.562 ;
    LAYER v0 ;
      RECT 1.046 0.202 1.114 0.246 ;
      RECT 1.046 0.492 1.114 0.536 ;
      RECT 0.938 0.293 1.006 0.337 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 0.938 0.202 ;
      RECT 0.938 0.158 1.006 0.382 ;
  END
END b15lsn080hn1n04x5

MACRO b15lsn080hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn080hn1n06x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.918 0.292 ;
        RECT 0.29 0.518 0.574 0.562 ;
        RECT 0.506 0.248 0.574 0.562 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.562 ;
      LAYER v0 ;
        RECT 1.262 0.4205 1.33 0.4645 ;
        RECT 1.262 0.193 1.33 0.237 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.702 0.428 0.898 0.472 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 1.154 0.4205 1.222 0.4645 ;
        RECT 1.37 0.4205 1.438 0.4645 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.154 0.193 1.222 0.237 ;
        RECT 1.37 0.193 1.438 0.237 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.702 0.338 1.046 0.382 ;
    LAYER v0 ;
      RECT 1.046 0.193 1.114 0.237 ;
      RECT 1.046 0.4205 1.114 0.4645 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.158 0.594 0.202 ;
      RECT 1.046 0.158 1.114 0.562 ;
  END
END b15lsn080hn1n06x5

MACRO b15lsn080hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn080hn1n08x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.918 0.292 ;
        RECT 0.29 0.518 0.574 0.562 ;
        RECT 0.506 0.248 0.574 0.562 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.562 ;
      LAYER v0 ;
        RECT 1.262 0.453 1.33 0.497 ;
        RECT 1.262 0.1645 1.33 0.2085 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.702 0.428 0.898 0.472 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 1.154 0.453 1.222 0.497 ;
        RECT 1.37 0.453 1.438 0.497 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.154 0.1645 1.222 0.2085 ;
        RECT 1.37 0.1645 1.438 0.2085 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.702 0.338 1.046 0.382 ;
    LAYER v0 ;
      RECT 1.046 0.1645 1.114 0.2085 ;
      RECT 1.046 0.453 1.114 0.497 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.158 0.594 0.202 ;
      RECT 1.046 0.068 1.114 0.562 ;
  END
END b15lsn080hn1n08x5

MACRO b15lsn080hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn080hn1n12x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 5.51 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.204 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.918 0.112 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
        RECT 0.83 0.068 0.898 0.112 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.562 ;
        RECT 1.37 0.338 1.654 0.382 ;
        RECT 1.37 0.158 1.438 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.45 1.438 0.494 ;
        RECT 1.37 0.2025 1.438 0.2465 ;
        RECT 1.586 0.45 1.654 0.494 ;
        RECT 1.586 0.2025 1.654 0.2465 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.722 0.428 0.918 0.472 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.262 0.45 1.33 0.494 ;
        RECT 1.478 0.45 1.546 0.494 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.81 0.158 1.114 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.184 0.25 0.228 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.262 0.113 1.33 0.157 ;
        RECT 1.478 0.113 1.546 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.81 0.338 1.33 0.382 ;
    LAYER v0 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.29 0.184 0.358 0.228 ;
      RECT 0.29 0.448 0.358 0.492 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.248 1.134 0.292 ;
  END
END b15lsn080hn1n12x5

MACRO b15lsn080hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lsn080hn1n16x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 5.51 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.204 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.918 0.112 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
        RECT 0.83 0.068 0.898 0.112 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.562 ;
        RECT 1.37 0.338 1.654 0.382 ;
        RECT 1.37 0.158 1.438 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.453 1.438 0.497 ;
        RECT 1.37 0.194 1.438 0.238 ;
        RECT 1.586 0.453 1.654 0.497 ;
        RECT 1.586 0.194 1.654 0.238 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.722 0.428 0.918 0.472 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.262 0.453 1.33 0.497 ;
        RECT 1.478 0.453 1.546 0.497 ;
        RECT 1.694 0.453 1.762 0.497 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.81 0.158 1.114 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.262 0.113 1.33 0.157 ;
        RECT 1.478 0.113 1.546 0.157 ;
        RECT 1.694 0.113 1.762 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.81 0.338 1.33 0.382 ;
    LAYER v0 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.4035 0.574 0.4475 ;
      RECT 0.4 0.498 0.464 0.542 ;
      RECT 0.29 0.143 0.358 0.187 ;
      RECT 0.074 0.143 0.142 0.187 ;
      RECT 0.076 0.3535 0.14 0.3975 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.358 0.428 0.398 0.472 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.574 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.248 1.134 0.292 ;
  END
END b15lsn080hn1n16x5

MACRO b15lyn003hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn003hn1n02x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.562 ;
      LAYER v0 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.586 0.203 1.654 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.61 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.61 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.242 0.382 ;
        RECT 1.046 0.068 1.114 0.382 ;
        RECT 0.398 0.068 1.114 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.478 0.448 1.546 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.223 0.358 0.267 ;
        RECT 1.154 0.203 1.222 0.247 ;
        RECT 1.478 0.203 1.546 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.248 0.79 0.562 ;
      RECT 1.37 0.158 1.438 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.158 0.466 0.382 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.158 0.81 0.202 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.006 0.428 1.242 0.472 ;
  END
END b15lyn003hn1n02x5

MACRO b15lyn003hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn003hn1n03x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.895 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.46222225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.562 ;
      LAYER v0 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.586 0.203 1.654 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.61 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.40666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.242 0.382 ;
        RECT 1.046 0.068 1.114 0.382 ;
        RECT 0.398 0.068 1.114 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.478 0.448 1.546 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.223 0.358 0.267 ;
        RECT 1.154 0.203 1.222 0.247 ;
        RECT 1.478 0.203 1.546 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.248 0.79 0.562 ;
      RECT 1.37 0.158 1.438 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.158 0.466 0.382 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.158 0.81 0.202 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.006 0.428 1.242 0.472 ;
  END
END b15lyn003hn1n03x5

MACRO b15lyn003hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn003hn1n04x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.56777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.211 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.562 ;
      LAYER v0 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.586 0.223 1.654 0.267 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.04 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.242 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.398 0.068 1.114 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 1.154 0.248 1.222 0.292 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.478 0.448 1.546 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.133 0.358 0.177 ;
        RECT 1.154 0.113 1.222 0.157 ;
        RECT 1.478 0.1125 1.546 0.1565 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.248 0.79 0.562 ;
      RECT 1.37 0.158 1.438 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.223 1.438 0.267 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.158 0.466 0.382 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.158 0.81 0.202 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.006 0.338 1.154 0.382 ;
      RECT 1.154 0.338 1.222 0.562 ;
  END
END b15lyn003hn1n04x5

MACRO b15lyn003hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn003hn1n06x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.56777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.211 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.562 ;
      LAYER v0 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.586 0.183 1.654 0.227 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.04 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.242 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.398 0.068 1.114 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 1.154 0.248 1.222 0.292 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.292 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.133 0.358 0.177 ;
        RECT 1.154 0.113 1.222 0.157 ;
        RECT 1.478 0.183 1.546 0.227 ;
        RECT 1.694 0.183 1.762 0.227 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.248 0.79 0.562 ;
      RECT 1.37 0.158 1.438 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.183 1.438 0.227 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.158 0.466 0.382 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.158 0.81 0.202 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.006 0.338 1.154 0.382 ;
      RECT 1.154 0.338 1.222 0.562 ;
  END
END b15lyn003hn1n06x5

MACRO b15lyn003hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn003hn1n08x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 4.0744445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 7.334 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 0.722 0.178 0.79 0.222 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.562 ;
      LAYER v0 ;
        RECT 1.802 0.4275 1.87 0.4715 ;
        RECT 1.802 0.1585 1.87 0.2025 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.42 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.382 ;
        RECT 0.506 0.068 1.33 0.112 ;
      LAYER v0 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.694 0.4275 1.762 0.4715 ;
        RECT 1.91 0.4275 1.978 0.4715 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.694 -0.022 1.762 0.292 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.398 0.158 0.594 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.167 0.142 0.211 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 1.37 0.113 1.438 0.157 ;
        RECT 1.694 0.1585 1.762 0.2025 ;
        RECT 1.91 0.1585 1.978 0.2025 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.586 0.068 1.654 0.562 ;
    LAYER v0 ;
      RECT 1.586 0.1585 1.654 0.2025 ;
      RECT 1.586 0.4275 1.654 0.4715 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.29 0.167 0.358 0.211 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.158 0.898 0.562 ;
      RECT 1.006 0.428 1.546 0.472 ;
  END
END b15lyn003hn1n08x5

MACRO b15lyn003hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn003hn1n12x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 6.8875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.29583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 1.242 0.292 ;
        RECT 0.83 0.158 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.832 0.178 0.896 0.222 ;
        RECT 1.154 0.248 1.222 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.378 0.382 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.158 2.194 0.562 ;
        RECT 1.91 0.338 2.194 0.382 ;
        RECT 1.91 0.158 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 1.91 0.183 1.978 0.227 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.126 0.183 2.194 0.227 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.64666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.292 ;
        RECT 0.614 0.068 1.546 0.112 ;
        RECT 0.614 0.068 0.682 0.382 ;
        RECT 0.398 0.158 0.682 0.202 ;
        RECT 0.398 0.068 0.466 0.202 ;
        RECT 0.182 0.068 0.466 0.112 ;
        RECT 0.074 0.158 0.25 0.202 ;
        RECT 0.182 0.068 0.25 0.202 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 1.478 0.203 1.546 0.247 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 1.802 0.093 1.87 0.137 ;
        RECT 2.018 0.093 2.086 0.137 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.694 0.158 1.762 0.562 ;
    LAYER v0 ;
      RECT 1.694 0.183 1.762 0.227 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.154 0.4405 1.222 0.4845 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.358 1.006 0.402 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.292 0.178 0.356 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.292 ;
      RECT 0.074 0.428 0.506 0.472 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.428 0.614 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 0.938 0.158 1.37 0.202 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.438 0.338 1.478 0.382 ;
      RECT 1.478 0.338 1.546 0.562 ;
  END
END b15lyn003hn1n12x5

MACRO b15lyn003hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn003hn1n16x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 7.125 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.458 0.292 ;
        RECT 1.046 0.158 1.114 0.292 ;
      LAYER v0 ;
        RECT 1.048 0.178 1.112 0.222 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.562 ;
        RECT 2.126 0.338 2.41 0.382 ;
        RECT 2.126 0.158 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.126 0.203 2.194 0.247 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.342 0.203 2.41 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0189 LAYER m1 ;
      ANTENNAMAXAREACAR 1.36477125 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0252 LAYER m1 ;
      ANTENNAMAXAREACAR 0.966713 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.068 1.762 0.292 ;
        RECT 0.83 0.068 1.762 0.112 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.228 0.898 0.272 ;
        RECT 1.694 0.203 1.762 0.247 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.1475 0.79 0.1915 ;
        RECT 1.802 0.093 1.87 0.137 ;
        RECT 2.018 0.093 2.086 0.137 ;
        RECT 2.234 0.093 2.302 0.137 ;
        RECT 2.45 0.093 2.518 0.137 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.91 0.158 1.978 0.562 ;
    LAYER v0 ;
      RECT 1.91 0.203 1.978 0.247 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.154 0.3895 1.222 0.4335 ;
      RECT 0.614 0.1475 0.682 0.1915 ;
      RECT 0.614 0.453 0.682 0.497 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.453 0.466 0.497 ;
      RECT 0.29 0.248 0.358 0.292 ;
      RECT 0.182 0.068 0.25 0.112 ;
      RECT 0.182 0.453 0.25 0.497 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.25 0.338 0.29 0.382 ;
      RECT 0.054 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.382 ;
      RECT 0.358 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.338 0.938 0.382 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.006 0.518 1.154 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.242 0.158 1.586 0.202 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 1.654 0.338 1.694 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
  END
END b15lyn003hn1n16x5

MACRO b15lyn00chn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn00chn1n02x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.382 ;
        RECT 0.27 0.068 1.114 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.83 0.068 0.898 0.112 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.802 0.391 1.87 0.435 ;
        RECT 1.802 0.138 1.87 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.694 0.391 1.762 0.435 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.398 0.248 0.682 0.292 ;
        RECT 0.614 0.158 0.682 0.292 ;
        RECT 0.398 0.158 0.466 0.292 ;
        RECT 0.074 0.158 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.616 0.178 0.68 0.222 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 1.694 0.138 1.762 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.562 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.586 0.068 1.654 0.472 ;
    LAYER v0 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.391 1.654 0.435 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.074 0.268 0.142 0.312 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 1.262 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.222 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
  END
END b15lyn00chn1n02x5

MACRO b15lyn00chn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn00chn1n03x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.382 ;
        RECT 0.27 0.068 1.114 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.83 0.068 0.898 0.112 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.802 0.391 1.87 0.435 ;
        RECT 1.802 0.138 1.87 0.182 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.694 0.391 1.762 0.435 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.398 0.248 0.682 0.292 ;
        RECT 0.614 0.158 0.682 0.292 ;
        RECT 0.398 0.158 0.466 0.292 ;
        RECT 0.074 0.158 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.616 0.178 0.68 0.222 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 1.694 0.138 1.762 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.562 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.586 0.068 1.654 0.472 ;
    LAYER v0 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.391 1.654 0.435 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.074 0.268 0.142 0.312 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 1.262 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.222 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
  END
END b15lyn00chn1n03x5

MACRO b15lyn00chn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn00chn1n04x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.29625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 10.5925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.273 0.898 0.317 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.434 1.978 0.478 ;
        RECT 1.91 0.113 1.978 0.157 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.6075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.6075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.574 0.202 ;
        RECT 0.506 0.068 0.574 0.202 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.158 0.466 0.202 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 1.478 0.478 1.546 0.522 ;
        RECT 1.802 0.434 1.87 0.478 ;
        RECT 2.018 0.434 2.086 0.478 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.802 0.113 1.87 0.157 ;
        RECT 2.018 0.113 2.086 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 1.694 0.068 1.762 0.562 ;
    LAYER v0 ;
      RECT 1.694 0.113 1.762 0.157 ;
      RECT 1.694 0.434 1.762 0.478 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.143 1.114 0.187 ;
      RECT 0.938 0.143 1.006 0.187 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.182 0.147 0.25 0.191 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.428 0.398 0.472 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.722 0.292 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.472 ;
      RECT 1.114 0.428 1.262 0.472 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.33 0.248 1.478 0.292 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.518 1.37 0.562 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.338 1.566 0.382 ;
  END
END b15lyn00chn1n04x5

MACRO b15lyn00chn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn00chn1n06x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.29625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 10.5925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.273 0.898 0.317 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.4025 1.978 0.4465 ;
        RECT 1.91 0.113 1.978 0.157 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.6075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.6075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.574 0.202 ;
        RECT 0.506 0.068 0.574 0.202 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.158 0.466 0.202 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 1.478 0.478 1.546 0.522 ;
        RECT 1.802 0.4025 1.87 0.4465 ;
        RECT 2.018 0.4025 2.086 0.4465 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.802 0.113 1.87 0.157 ;
        RECT 2.018 0.113 2.086 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.046 0.068 1.114 0.472 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 1.694 0.068 1.762 0.472 ;
    LAYER v0 ;
      RECT 1.694 0.113 1.762 0.157 ;
      RECT 1.694 0.4025 1.762 0.4465 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.143 1.114 0.187 ;
      RECT 0.938 0.143 1.006 0.187 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.182 0.147 0.25 0.191 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.428 0.398 0.472 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.722 0.292 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.472 ;
      RECT 1.114 0.428 1.262 0.472 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.33 0.248 1.478 0.292 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.518 1.37 0.562 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.338 1.566 0.382 ;
  END
END b15lyn00chn1n06x5

MACRO b15lyn00chn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn00chn1n08x5 0 0 ;
  SIZE 2.376 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.667 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 7.334 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.408 1.114 0.452 ;
        RECT 1.046 0.178 1.114 0.222 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.4305 2.194 0.4745 ;
        RECT 2.126 0.116 2.194 0.16 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.722 0.068 0.79 0.202 ;
        RECT 0.506 0.158 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.41 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.83 0.4725 0.898 0.5165 ;
        RECT 1.694 0.472 1.762 0.516 ;
        RECT 2.018 0.4305 2.086 0.4745 ;
        RECT 2.234 0.4305 2.302 0.4745 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.41 0.022 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.018 0.116 2.086 0.16 ;
        RECT 2.234 0.116 2.302 0.16 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 1.262 0.158 1.33 0.472 ;
      RECT 1.91 0.068 1.978 0.562 ;
    LAYER v0 ;
      RECT 1.91 0.116 1.978 0.16 ;
      RECT 1.91 0.4305 1.978 0.4745 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 0.722 0.4725 0.79 0.5165 ;
      RECT 0.398 0.157 0.466 0.201 ;
      RECT 0.182 0.157 0.25 0.201 ;
      RECT 0.184 0.408 0.248 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.248 0.682 0.382 ;
      RECT 0.682 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.006 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.472 ;
      RECT 0.79 0.338 0.938 0.382 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.006 0.518 1.586 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.654 0.338 1.782 0.382 ;
      RECT 1.33 0.428 1.478 0.472 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.546 0.248 1.782 0.292 ;
  END
END b15lyn00chn1n08x5

MACRO b15lyn00chn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn00chn1n12x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 6.175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.05833325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 1.438 0.382 ;
        RECT 1.026 0.068 1.438 0.112 ;
      LAYER v0 ;
        RECT 1.046 0.068 1.114 0.112 ;
        RECT 1.37 0.293 1.438 0.337 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.202 ;
        RECT 0.486 0.068 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.562 ;
        RECT 2.126 0.338 2.41 0.382 ;
        RECT 2.126 0.068 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.342 0.158 2.41 0.202 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.722 0.4775 0.79 0.5215 ;
        RECT 1.694 0.472 1.762 0.516 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.234 -0.022 2.302 0.292 ;
        RECT 2.018 -0.022 2.086 0.292 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 0.158 0.594 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.0705 0.358 0.1145 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 1.262 0.158 1.33 0.472 ;
      RECT 1.91 0.068 1.978 0.562 ;
    LAYER v0 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.1955 1.33 0.2395 ;
      RECT 1.154 0.308 1.222 0.352 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.408 0.574 0.452 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.182 0.338 0.25 0.382 ;
      RECT 0.074 0.068 0.142 0.112 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.378 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.006 0.428 1.154 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.428 0.398 0.472 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.518 1.586 0.562 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.654 0.338 1.782 0.382 ;
      RECT 1.33 0.428 1.478 0.472 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.546 0.248 1.782 0.292 ;
  END
END b15lyn00chn1n12x5

MACRO b15lyn00chn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn00chn1n16x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 7.8375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.6125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.338 1.654 0.382 ;
        RECT 1.586 0.158 1.654 0.382 ;
        RECT 1.262 0.158 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.586 0.248 1.654 0.292 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.382 ;
        RECT 0.054 0.248 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
        RECT 2.342 0.338 2.626 0.382 ;
        RECT 2.342 0.068 2.41 0.562 ;
      LAYER v0 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.558 0.158 2.626 0.202 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37071425 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.59916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.498 1.114 0.542 ;
    END
  END psb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.506 0.509 0.574 0.553 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.938 0.403 1.006 0.447 ;
        RECT 1.91 0.4385 1.978 0.4825 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.666 0.448 2.734 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.292 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.29 0.472 ;
      RECT 0.594 0.248 1.154 0.292 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 2.126 0.068 2.194 0.562 ;
    LAYER v0 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.163 1.546 0.207 ;
      RECT 1.37 0.163 1.438 0.207 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.518 0.25 0.562 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.398 0.562 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.054 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.358 0.158 1.154 0.202 ;
      RECT 1.154 0.068 1.222 0.202 ;
      RECT 1.222 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 1.222 0.518 1.802 0.562 ;
      RECT 1.802 0.248 1.87 0.562 ;
      RECT 1.566 0.428 1.694 0.472 ;
      RECT 1.546 0.068 1.694 0.112 ;
      RECT 1.694 0.068 1.762 0.472 ;
      RECT 1.762 0.158 2.086 0.202 ;
  END
END b15lyn00chn1n16x5

MACRO b15lyn00fhn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn00fhn1n02x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.95875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.95875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.574 0.562 ;
        RECT 0.182 0.068 0.574 0.112 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.518 0.466 0.562 ;
        RECT 0.398 0.068 0.466 0.112 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.3155 0.898 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.562 ;
      LAYER v0 ;
        RECT 1.802 0.473 1.87 0.517 ;
        RECT 1.802 0.14 1.87 0.184 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.158 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.3155 1.762 0.3595 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.3155 1.114 0.3595 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
        RECT 1.478 0.473 1.546 0.517 ;
        RECT 1.694 0.473 1.762 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.506 0.338 0.722 0.382 ;
      RECT 1.458 0.068 1.586 0.112 ;
    LAYER v0 ;
      RECT 1.586 0.473 1.654 0.517 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.3155 1.546 0.3595 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.292 0.178 0.356 0.222 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.466 0.428 1.37 0.472 ;
      RECT 1.154 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.006 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
  END
END b15lyn00fhn1n02x5

MACRO b15lyn00fhn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn00fhn1n04x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.95875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.95875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.574 0.562 ;
        RECT 0.182 0.068 0.574 0.112 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.518 0.466 0.562 ;
        RECT 0.398 0.068 0.466 0.112 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.3155 0.898 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.562 ;
      LAYER v0 ;
        RECT 1.802 0.473 1.87 0.517 ;
        RECT 1.802 0.14 1.87 0.184 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.158 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.3155 1.762 0.3595 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.3155 1.114 0.3595 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
        RECT 1.478 0.473 1.546 0.517 ;
        RECT 1.694 0.473 1.762 0.517 ;
        RECT 1.91 0.473 1.978 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 1.91 0.048 1.978 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.506 0.338 0.722 0.382 ;
      RECT 1.458 0.068 1.586 0.112 ;
    LAYER v0 ;
      RECT 1.586 0.473 1.654 0.517 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.3155 1.546 0.3595 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.292 0.178 0.356 0.222 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.466 0.428 1.37 0.472 ;
      RECT 1.154 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.006 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
      RECT 1.586 0.068 1.654 0.562 ;
  END
END b15lyn00fhn1n04x5

MACRO b15lyn00fhn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn00fhn1n08x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.95875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 6.1855555 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.574 0.562 ;
        RECT 0.182 0.068 0.574 0.112 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.518 0.466 0.562 ;
        RECT 0.398 0.068 0.466 0.112 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.3155 0.898 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.562 ;
        RECT 1.91 0.338 2.194 0.382 ;
        RECT 1.91 0.068 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.473 1.978 0.517 ;
        RECT 1.91 0.14 1.978 0.184 ;
        RECT 2.126 0.473 2.194 0.517 ;
        RECT 2.126 0.14 2.194 0.184 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.3155 1.87 0.3595 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.3155 1.222 0.3595 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.586 0.473 1.654 0.517 ;
        RECT 1.802 0.473 1.87 0.517 ;
        RECT 2.018 0.473 2.086 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.158 1.672 0.202 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.938 0.158 1.438 0.202 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.478 0.068 1.546 0.382 ;
    LAYER v1 ;
      RECT 1.482 0.158 1.542 0.202 ;
      RECT 0.726 0.158 0.786 0.202 ;
    LAYER v0 ;
      RECT 1.694 0.473 1.762 0.517 ;
      RECT 1.586 0.14 1.654 0.184 ;
      RECT 1.478 0.3155 1.546 0.3595 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.292 0.178 0.356 0.222 ;
    LAYER m1 ;
      RECT 0.506 0.338 0.722 0.382 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.466 0.428 1.546 0.472 ;
      RECT 1.654 0.338 1.694 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
  END
END b15lyn00fhn1n08x5

MACRO b15lyn00fhn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn00fhn1n16x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 6.1855555 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 5.060909 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.574 0.562 ;
        RECT 0.182 0.068 0.574 0.112 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.518 0.466 0.562 ;
        RECT 0.398 0.068 0.466 0.112 ;
    END
  END clk
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.3155 0.898 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.068 2.626 0.562 ;
        RECT 2.126 0.248 2.626 0.292 ;
        RECT 2.342 0.068 2.41 0.562 ;
        RECT 2.126 0.068 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.389 2.194 0.433 ;
        RECT 2.126 0.14 2.194 0.184 ;
        RECT 2.342 0.389 2.41 0.433 ;
        RECT 2.342 0.14 2.41 0.184 ;
        RECT 2.558 0.389 2.626 0.433 ;
        RECT 2.558 0.14 2.626 0.184 ;
    END
  END o
  PIN psb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.382 ;
      LAYER v0 ;
        RECT 2.018 0.293 2.086 0.337 ;
    END
  END psb
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.3155 1.222 0.3595 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.154 0.538 1.222 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.802 0.473 1.87 0.517 ;
        RECT 2.018 0.473 2.086 0.517 ;
        RECT 2.234 0.473 2.302 0.517 ;
        RECT 2.45 0.473 2.518 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.234 0.048 2.302 0.092 ;
        RECT 2.45 0.048 2.518 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.158 1.888 0.202 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.938 0.158 1.654 0.202 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.694 0.068 1.762 0.382 ;
    LAYER v1 ;
      RECT 1.698 0.158 1.758 0.202 ;
      RECT 0.726 0.158 0.786 0.202 ;
    LAYER v0 ;
      RECT 1.91 0.473 1.978 0.517 ;
      RECT 1.802 0.14 1.87 0.184 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.292 0.178 0.356 0.222 ;
    LAYER m1 ;
      RECT 0.506 0.338 0.722 0.382 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.466 0.428 1.762 0.472 ;
      RECT 1.87 0.248 1.91 0.292 ;
      RECT 1.91 0.248 1.978 0.562 ;
  END
END b15lyn00fhn1n16x5

MACRO b15lyn083hn1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn083hn1n02x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.1455555 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.53875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.562 ;
      LAYER v0 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.586 0.203 1.654 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 1.222 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 1.046 0.518 1.114 0.562 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.938 0.428 1.33 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.478 0.448 1.546 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.193 0.358 0.237 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.478 0.203 1.546 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 1.37 0.158 1.438 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.428 0.898 0.472 ;
      RECT 0.79 0.338 1.33 0.382 ;
  END
END b15lyn083hn1n02x5

MACRO b15lyn083hn1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn083hn1n03x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.46222225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.46222225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.562 ;
      LAYER v0 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.586 0.203 1.654 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 1.222 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 1.046 0.518 1.114 0.562 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.938 0.428 1.33 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.478 0.448 1.546 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.193 0.358 0.237 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.478 0.203 1.546 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 1.37 0.158 1.438 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.428 0.898 0.472 ;
      RECT 0.79 0.338 1.33 0.382 ;
  END
END b15lyn083hn1n03x5

MACRO b15lyn083hn1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn083hn1n04x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.088 0.574 0.132 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.562 ;
      LAYER v0 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.586 0.203 1.654 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 1.222 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 1.046 0.518 1.114 0.562 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.938 0.428 1.33 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.478 0.448 1.546 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.193 0.358 0.237 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.478 0.203 1.546 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 1.37 0.158 1.438 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.428 0.898 0.472 ;
      RECT 0.79 0.338 1.33 0.382 ;
  END
END b15lyn083hn1n04x5

MACRO b15lyn083hn1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn083hn1n06x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.088 0.574 0.132 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.562 ;
      LAYER v0 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.586 0.203 1.654 0.247 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 1.222 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 1.046 0.518 1.114 0.562 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.938 0.428 1.33 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.292 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.193 0.358 0.237 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.478 0.203 1.546 0.247 ;
        RECT 1.694 0.203 1.762 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 1.37 0.158 1.438 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.203 1.438 0.247 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.428 0.898 0.472 ;
      RECT 0.79 0.338 1.33 0.382 ;
  END
END b15lyn083hn1n06x5

MACRO b15lyn083hn1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn083hn1n08x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.755 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 5.51 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 0.722 0.178 0.79 0.222 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.562 ;
      LAYER v0 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 1.802 0.178 1.87 0.222 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.42 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 1.438 0.202 ;
        RECT 0.506 0.068 1.438 0.112 ;
      LAYER v0 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.262 0.068 1.33 0.112 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 1.694 -0.022 1.762 0.292 ;
        RECT 1.262 0.248 1.546 0.292 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 0.398 0.158 0.594 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.167 0.142 0.211 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.694 0.178 1.762 0.222 ;
        RECT 1.91 0.178 1.978 0.222 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.586 0.158 1.654 0.562 ;
    LAYER v0 ;
      RECT 1.586 0.178 1.654 0.222 ;
      RECT 1.586 0.448 1.654 0.492 ;
      RECT 1.37 0.448 1.438 0.492 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.29 0.167 0.358 0.211 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.158 0.898 0.562 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.006 0.518 1.154 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
  END
END b15lyn083hn1n08x5

MACRO b15lyn083hn1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn083hn1n12x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.4115385 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 6.27 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.472 ;
        RECT 0.83 0.248 1.222 0.292 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.358 0.898 0.402 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5811765 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.562 ;
        RECT 1.91 0.248 2.194 0.292 ;
        RECT 1.91 0.068 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 1.91 0.113 1.978 0.157 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.126 0.113 2.194 0.157 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 2.66 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0189 LAYER m1 ;
      ANTENNAMAXAREACAR 1.877647 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 1.438 0.292 ;
        RECT 0.614 0.068 1.438 0.112 ;
      LAYER v0 ;
        RECT 0.722 0.068 0.79 0.112 ;
        RECT 1.37 0.2255 1.438 0.2695 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.167 0.142 0.211 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 1.478 0.093 1.546 0.137 ;
        RECT 1.802 0.113 1.87 0.157 ;
        RECT 2.018 0.113 2.086 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.694 0.068 1.762 0.562 ;
    LAYER v0 ;
      RECT 1.694 0.113 1.762 0.157 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.048 0.448 1.112 0.492 ;
      RECT 0.938 0.358 1.006 0.402 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.074 0.428 0.506 0.472 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.562 ;
      RECT 0.79 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.046 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.338 1.478 0.382 ;
      RECT 1.478 0.338 1.546 0.562 ;
  END
END b15lyn083hn1n12x5

MACRO b15lyn083hn1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15lyn083hn1n16x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clkb
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.4115385 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 6.27 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.248 1.438 0.472 ;
        RECT 1.046 0.248 1.438 0.292 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.358 1.114 0.402 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END clkb
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.89818175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.682 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.562 ;
        RECT 2.126 0.248 2.41 0.292 ;
        RECT 2.126 0.068 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.126 0.113 2.194 0.157 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.342 0.113 2.41 0.157 ;
    END
  END o
  PIN rb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 2.14588225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0261 LAYER m1 ;
      ANTENNAMAXAREACAR 1.4592 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.068 1.654 0.292 ;
        RECT 0.83 0.068 1.654 0.112 ;
      LAYER v0 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 1.586 0.2255 1.654 0.2695 ;
    END
  END rb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 0.722 0.158 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.113 0.358 0.157 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.694 0.093 1.762 0.137 ;
        RECT 2.018 0.113 2.086 0.157 ;
        RECT 2.234 0.113 2.302 0.157 ;
        RECT 2.45 0.113 2.518 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.91 0.068 1.978 0.562 ;
    LAYER v0 ;
      RECT 1.91 0.113 1.978 0.157 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.264 0.448 1.328 0.492 ;
      RECT 1.154 0.358 1.222 0.402 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.074 0.428 0.722 0.472 ;
      RECT 0.25 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.562 ;
      RECT 1.006 0.518 1.154 0.562 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.33 0.518 1.478 0.562 ;
      RECT 1.262 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.546 0.338 1.694 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
  END
END b15lyn083hn1n16x5

END LIBRARY
