module test_io (
    inout port1,
    inout port2
);

    assign port2 = port1;

endmodule