module aes_cipher_top (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire net801;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire net800;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire net799;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire net798;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire net797;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire net796;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire net795;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire net794;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire net793;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire net792;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire net791;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire net790;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire net789;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire net788;
 wire _02242_;
 wire net787;
 wire net786;
 wire net785;
 wire net784;
 wire net783;
 wire net782;
 wire net781;
 wire net780;
 wire _02251_;
 wire net779;
 wire net778;
 wire net777;
 wire net776;
 wire net775;
 wire _02257_;
 wire net774;
 wire _02259_;
 wire net773;
 wire net772;
 wire _02262_;
 wire _02263_;
 wire net771;
 wire net770;
 wire net769;
 wire net768;
 wire net767;
 wire net766;
 wire net765;
 wire net764;
 wire net763;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire net762;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire net761;
 wire net760;
 wire net759;
 wire net758;
 wire _02286_;
 wire net757;
 wire net756;
 wire net755;
 wire _02290_;
 wire _02291_;
 wire net754;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire net753;
 wire net752;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire net751;
 wire net750;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire net749;
 wire net748;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire net747;
 wire _02313_;
 wire net746;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire net745;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire net744;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire net743;
 wire net742;
 wire net741;
 wire _02337_;
 wire _02338_;
 wire net740;
 wire _02340_;
 wire _02341_;
 wire net739;
 wire _02343_;
 wire net738;
 wire net737;
 wire _02346_;
 wire net736;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire net735;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire net734;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire net733;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire net732;
 wire net731;
 wire net730;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire net729;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire net728;
 wire net727;
 wire net726;
 wire _02385_;
 wire net725;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire net724;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire net723;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire net722;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire net721;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire net720;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire net719;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02422_;
 wire _02423_;
 wire net718;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire net717;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02433_;
 wire net716;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire net715;
 wire _02440_;
 wire _02441_;
 wire net714;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02455_;
 wire net713;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire net712;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire net711;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire net710;
 wire _02475_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire net709;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire net708;
 wire _02496_;
 wire net707;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire net706;
 wire _02504_;
 wire _02505_;
 wire net705;
 wire _02507_;
 wire net704;
 wire net703;
 wire net702;
 wire net701;
 wire net700;
 wire net699;
 wire _02515_;
 wire net698;
 wire _02517_;
 wire net697;
 wire net696;
 wire net695;
 wire net694;
 wire net693;
 wire _02524_;
 wire net692;
 wire _02526_;
 wire _02527_;
 wire net691;
 wire _02529_;
 wire net690;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire net689;
 wire net688;
 wire net687;
 wire net686;
 wire net685;
 wire net684;
 wire _02541_;
 wire _02543_;
 wire net683;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire net682;
 wire _02550_;
 wire net681;
 wire net680;
 wire _02554_;
 wire _02555_;
 wire net679;
 wire _02557_;
 wire net678;
 wire _02559_;
 wire net677;
 wire net676;
 wire _02562_;
 wire _02563_;
 wire net675;
 wire _02566_;
 wire _02567_;
 wire net674;
 wire _02569_;
 wire net673;
 wire net672;
 wire net671;
 wire _02573_;
 wire net670;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire net669;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire net668;
 wire _02583_;
 wire net667;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire net666;
 wire net665;
 wire net664;
 wire net663;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire net662;
 wire _02600_;
 wire net661;
 wire _02602_;
 wire net660;
 wire _02604_;
 wire _02605_;
 wire net659;
 wire net658;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire net657;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire net656;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire net655;
 wire _02622_;
 wire _02623_;
 wire net654;
 wire _02625_;
 wire net653;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire net652;
 wire net651;
 wire _02634_;
 wire _02635_;
 wire net650;
 wire _02637_;
 wire net649;
 wire _02639_;
 wire _02640_;
 wire _02642_;
 wire _02643_;
 wire net648;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02653_;
 wire _02654_;
 wire net647;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire net646;
 wire _02661_;
 wire _02662_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire net645;
 wire _02674_;
 wire net644;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire net643;
 wire _02683_;
 wire _02684_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire net642;
 wire _02692_;
 wire net641;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire net640;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire net639;
 wire net638;
 wire _02705_;
 wire net637;
 wire net636;
 wire _02709_;
 wire net635;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire net634;
 wire _02716_;
 wire net633;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire net632;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire net631;
 wire _02731_;
 wire _02732_;
 wire net630;
 wire _02734_;
 wire net629;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire net628;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire net627;
 wire net626;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire net625;
 wire net624;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire net623;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire net622;
 wire net621;
 wire net620;
 wire net619;
 wire net618;
 wire _02779_;
 wire net617;
 wire _02781_;
 wire _02782_;
 wire net616;
 wire _02784_;
 wire net615;
 wire net614;
 wire _02787_;
 wire _02788_;
 wire net613;
 wire net612;
 wire _02791_;
 wire net611;
 wire net610;
 wire _02794_;
 wire net609;
 wire net608;
 wire _02798_;
 wire _02799_;
 wire net607;
 wire net606;
 wire net605;
 wire net604;
 wire net603;
 wire net602;
 wire _02807_;
 wire _02808_;
 wire net601;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire net600;
 wire net599;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire net598;
 wire _02822_;
 wire net597;
 wire _02824_;
 wire _02825_;
 wire net596;
 wire _02827_;
 wire _02829_;
 wire net595;
 wire _02831_;
 wire net594;
 wire _02833_;
 wire _02834_;
 wire net593;
 wire net592;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire net591;
 wire net590;
 wire _02843_;
 wire _02844_;
 wire net589;
 wire net588;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire net587;
 wire _02853_;
 wire _02854_;
 wire net586;
 wire _02856_;
 wire net585;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02862_;
 wire net584;
 wire _02864_;
 wire net583;
 wire net582;
 wire _02867_;
 wire _02868_;
 wire net581;
 wire _02870_;
 wire _02871_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire net580;
 wire _02885_;
 wire _02886_;
 wire net579;
 wire net578;
 wire net577;
 wire net576;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire net575;
 wire _02904_;
 wire net574;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire net573;
 wire _02911_;
 wire net572;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire net571;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire net570;
 wire _02923_;
 wire _02924_;
 wire net569;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire net568;
 wire net567;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire net566;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire net565;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire net564;
 wire _02953_;
 wire _02954_;
 wire net563;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire net562;
 wire _02960_;
 wire _02961_;
 wire net561;
 wire net560;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire net559;
 wire _02970_;
 wire net558;
 wire _02973_;
 wire _02974_;
 wire net557;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire net556;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire net555;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire net554;
 wire _02992_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire net553;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire net552;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire net551;
 wire _03023_;
 wire _03024_;
 wire net550;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire net549;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire net548;
 wire _03036_;
 wire net547;
 wire net546;
 wire net545;
 wire net544;
 wire net543;
 wire net542;
 wire _03044_;
 wire net541;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire net540;
 wire _03050_;
 wire net539;
 wire net538;
 wire _03053_;
 wire net537;
 wire net536;
 wire net535;
 wire _03057_;
 wire net534;
 wire _03059_;
 wire net533;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire net532;
 wire net531;
 wire net530;
 wire _03067_;
 wire _03068_;
 wire net529;
 wire _03071_;
 wire net528;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire net527;
 wire _03077_;
 wire net526;
 wire _03079_;
 wire net525;
 wire _03082_;
 wire _03083_;
 wire net524;
 wire net523;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire net522;
 wire _03092_;
 wire net521;
 wire net520;
 wire _03095_;
 wire net519;
 wire _03097_;
 wire net518;
 wire _03099_;
 wire _03100_;
 wire net517;
 wire _03102_;
 wire net516;
 wire net515;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire net514;
 wire net513;
 wire net512;
 wire _03116_;
 wire net511;
 wire net510;
 wire net509;
 wire net508;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire net507;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire net506;
 wire _03132_;
 wire net505;
 wire _03134_;
 wire _03135_;
 wire _03137_;
 wire _03138_;
 wire net504;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire net503;
 wire _03152_;
 wire net502;
 wire net501;
 wire _03155_;
 wire net500;
 wire _03157_;
 wire _03159_;
 wire _03160_;
 wire net499;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire net498;
 wire _03175_;
 wire net497;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire net496;
 wire net495;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire net494;
 wire _03189_;
 wire net493;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire net492;
 wire net491;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire net490;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire net489;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire net488;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire net487;
 wire net486;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire net485;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire net484;
 wire _03261_;
 wire net483;
 wire _03263_;
 wire net482;
 wire net481;
 wire net480;
 wire _03267_;
 wire _03268_;
 wire net479;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire net478;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03324_;
 wire _03325_;
 wire net477;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire net476;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire net475;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire net474;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire net473;
 wire net472;
 wire _03421_;
 wire _03422_;
 wire net471;
 wire _03424_;
 wire _03425_;
 wire net470;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire net469;
 wire net468;
 wire net467;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire net466;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire net465;
 wire _03485_;
 wire _03486_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire net464;
 wire _03493_;
 wire _03494_;
 wire net463;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire net462;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire net461;
 wire net460;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire net459;
 wire _03519_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire net458;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire net457;
 wire _03556_;
 wire _03557_;
 wire net456;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire net455;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire net454;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire net453;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire net452;
 wire _03640_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire net451;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire net450;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire net449;
 wire _03683_;
 wire net448;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire net447;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire net446;
 wire net445;
 wire net444;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire net443;
 wire _03750_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire net442;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire net441;
 wire _03773_;
 wire net440;
 wire _03775_;
 wire net439;
 wire _03777_;
 wire net438;
 wire _03779_;
 wire net437;
 wire net436;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire net435;
 wire _03786_;
 wire _03787_;
 wire net434;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire net433;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire net432;
 wire net431;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire net430;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire net429;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire net428;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire net427;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire net426;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire net425;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire net424;
 wire net423;
 wire net422;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire net421;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire net420;
 wire _03898_;
 wire _03899_;
 wire net419;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03906_;
 wire net418;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire net417;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire net416;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire net415;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire net414;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire net413;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04509_;
 wire net412;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire net411;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05793_;
 wire net410;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire net409;
 wire net408;
 wire net407;
 wire net406;
 wire net405;
 wire _05820_;
 wire _05821_;
 wire net404;
 wire net403;
 wire net402;
 wire net401;
 wire net400;
 wire _05827_;
 wire net399;
 wire _05829_;
 wire net398;
 wire _05831_;
 wire _05832_;
 wire net397;
 wire net396;
 wire _05835_;
 wire net395;
 wire net394;
 wire net393;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire net392;
 wire _05846_;
 wire net391;
 wire _05848_;
 wire net390;
 wire net389;
 wire _05851_;
 wire net388;
 wire _05853_;
 wire _05854_;
 wire net387;
 wire _05856_;
 wire net386;
 wire net385;
 wire net384;
 wire _05860_;
 wire _05861_;
 wire net383;
 wire net382;
 wire _05864_;
 wire net381;
 wire net380;
 wire _05867_;
 wire net379;
 wire net378;
 wire _05870_;
 wire net377;
 wire net376;
 wire net375;
 wire net374;
 wire _05875_;
 wire net373;
 wire net372;
 wire net371;
 wire net370;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire net369;
 wire net368;
 wire net367;
 wire _05891_;
 wire net366;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire net365;
 wire net364;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire net363;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire net362;
 wire net361;
 wire net360;
 wire _05915_;
 wire net359;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire net358;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire net357;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire net356;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire net355;
 wire _05937_;
 wire net354;
 wire _05939_;
 wire net353;
 wire _05941_;
 wire _05942_;
 wire net352;
 wire net351;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire net350;
 wire _05949_;
 wire net349;
 wire net348;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire net347;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire net346;
 wire net345;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire net344;
 wire _05971_;
 wire _05972_;
 wire net343;
 wire _05974_;
 wire _05975_;
 wire net342;
 wire _05977_;
 wire _05978_;
 wire net341;
 wire _05980_;
 wire net340;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire net339;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire net338;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire net337;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire net336;
 wire _06009_;
 wire net335;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire net334;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire net333;
 wire net332;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire net331;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire net330;
 wire _06056_;
 wire net329;
 wire _06058_;
 wire net328;
 wire _06060_;
 wire net327;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire net326;
 wire _06070_;
 wire net325;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire net324;
 wire _06081_;
 wire _06082_;
 wire net323;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire net322;
 wire _06091_;
 wire net321;
 wire net320;
 wire net319;
 wire _06095_;
 wire _06096_;
 wire net318;
 wire net317;
 wire net316;
 wire _06100_;
 wire _06101_;
 wire net315;
 wire _06103_;
 wire net314;
 wire _06105_;
 wire net313;
 wire _06108_;
 wire _06109_;
 wire net312;
 wire _06111_;
 wire net311;
 wire net310;
 wire _06114_;
 wire net309;
 wire net308;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire net307;
 wire _06121_;
 wire net306;
 wire net305;
 wire net304;
 wire _06125_;
 wire net303;
 wire _06127_;
 wire _06128_;
 wire net302;
 wire net301;
 wire net300;
 wire net299;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire net298;
 wire net297;
 wire net296;
 wire _06139_;
 wire _06140_;
 wire net295;
 wire net294;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire net293;
 wire net292;
 wire _06150_;
 wire net291;
 wire net290;
 wire net289;
 wire net288;
 wire _06155_;
 wire _06156_;
 wire net287;
 wire _06158_;
 wire net286;
 wire net285;
 wire _06161_;
 wire net284;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire net283;
 wire _06169_;
 wire net282;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire net281;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire net280;
 wire net279;
 wire net278;
 wire _06183_;
 wire net277;
 wire net276;
 wire net275;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire net274;
 wire net273;
 wire net272;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire net271;
 wire _06197_;
 wire net270;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire net269;
 wire _06203_;
 wire net268;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire net267;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire net266;
 wire _06223_;
 wire _06224_;
 wire net265;
 wire net264;
 wire _06227_;
 wire _06228_;
 wire net263;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire net262;
 wire _06235_;
 wire _06236_;
 wire net261;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire net260;
 wire net259;
 wire _06248_;
 wire _06249_;
 wire net258;
 wire net257;
 wire net256;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire net255;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire net254;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire net253;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire net252;
 wire net251;
 wire _06282_;
 wire net250;
 wire _06284_;
 wire net249;
 wire _06286_;
 wire _06287_;
 wire net248;
 wire _06289_;
 wire net247;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire net246;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire net245;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire net244;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire net243;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire net242;
 wire net241;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire net240;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire net239;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire net238;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire net237;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire net236;
 wire _06375_;
 wire net235;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire net234;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire net233;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire net232;
 wire _06401_;
 wire _06402_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire net231;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire net230;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire net229;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire net228;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire net227;
 wire _06476_;
 wire net226;
 wire net225;
 wire net224;
 wire _06480_;
 wire net223;
 wire net222;
 wire net221;
 wire net220;
 wire net219;
 wire net218;
 wire net217;
 wire _06488_;
 wire net216;
 wire net215;
 wire _06491_;
 wire net214;
 wire net213;
 wire net212;
 wire _06495_;
 wire _06496_;
 wire net211;
 wire net210;
 wire _06499_;
 wire net209;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire net208;
 wire net207;
 wire net206;
 wire net205;
 wire net204;
 wire _06509_;
 wire net203;
 wire net202;
 wire net201;
 wire _06513_;
 wire _06514_;
 wire net200;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire net199;
 wire _06522_;
 wire net198;
 wire _06524_;
 wire _06525_;
 wire net197;
 wire _06527_;
 wire net196;
 wire _06529_;
 wire _06530_;
 wire net195;
 wire net194;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire net193;
 wire _06538_;
 wire _06539_;
 wire net192;
 wire _06541_;
 wire _06542_;
 wire net191;
 wire net190;
 wire _06545_;
 wire _06546_;
 wire net189;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire net188;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire net187;
 wire _06560_;
 wire net186;
 wire net185;
 wire net184;
 wire net183;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire net182;
 wire net181;
 wire net180;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire net179;
 wire net178;
 wire _06577_;
 wire net177;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire net176;
 wire net175;
 wire _06584_;
 wire net174;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire net173;
 wire net172;
 wire _06593_;
 wire _06594_;
 wire net171;
 wire _06596_;
 wire _06597_;
 wire net170;
 wire net169;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire net168;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire net167;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire net166;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire net165;
 wire net164;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire net163;
 wire _06623_;
 wire _06624_;
 wire net162;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire net161;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire net160;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06645_;
 wire net159;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire net158;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire net157;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire net156;
 wire _06661_;
 wire net155;
 wire _06663_;
 wire net154;
 wire net153;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire net152;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06678_;
 wire net151;
 wire net150;
 wire _06681_;
 wire _06682_;
 wire net149;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire net148;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire net147;
 wire net146;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire net145;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire net144;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire net143;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire net142;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire net141;
 wire _06743_;
 wire net140;
 wire net139;
 wire net138;
 wire net137;
 wire _06748_;
 wire net136;
 wire net135;
 wire net134;
 wire net133;
 wire net132;
 wire _06754_;
 wire net131;
 wire _06756_;
 wire net130;
 wire _06758_;
 wire net129;
 wire _06760_;
 wire _06761_;
 wire net128;
 wire net127;
 wire net126;
 wire _06765_;
 wire net125;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire net124;
 wire _06771_;
 wire net123;
 wire net122;
 wire net121;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire net120;
 wire _06781_;
 wire net119;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire net118;
 wire net117;
 wire _06790_;
 wire net116;
 wire _06792_;
 wire net115;
 wire net114;
 wire _06795_;
 wire net113;
 wire net112;
 wire _06798_;
 wire net111;
 wire _06800_;
 wire net110;
 wire net109;
 wire net108;
 wire _06804_;
 wire _06805_;
 wire net107;
 wire _06807_;
 wire net106;
 wire _06809_;
 wire net105;
 wire net104;
 wire net103;
 wire _06813_;
 wire net102;
 wire net101;
 wire net100;
 wire _06817_;
 wire net99;
 wire net98;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire net97;
 wire _06826_;
 wire net96;
 wire _06828_;
 wire net95;
 wire net94;
 wire _06831_;
 wire _06832_;
 wire net93;
 wire net92;
 wire net91;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire net90;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire net89;
 wire _06846_;
 wire _06847_;
 wire net88;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire net87;
 wire net86;
 wire net85;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire net84;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire net83;
 wire net82;
 wire _06872_;
 wire net81;
 wire net80;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire net79;
 wire net78;
 wire _06881_;
 wire _06882_;
 wire net77;
 wire net76;
 wire net75;
 wire _06886_;
 wire net74;
 wire _06888_;
 wire _06889_;
 wire net73;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire net72;
 wire _06896_;
 wire _06897_;
 wire net71;
 wire _06899_;
 wire net70;
 wire _06901_;
 wire net69;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire net68;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire net67;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire net66;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire net65;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire net64;
 wire net63;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire net62;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire net61;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire net60;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire net59;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire net58;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire net57;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire net56;
 wire _06988_;
 wire net55;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire net54;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire net53;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire net52;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire net51;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire net50;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire net49;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire net48;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire net47;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire net46;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire net45;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire net44;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire net43;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire net42;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire net41;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire net40;
 wire _07269_;
 wire _07270_;
 wire net39;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire net38;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire net37;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire net36;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire net35;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire net34;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire net33;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire net32;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire net31;
 wire _07497_;
 wire _07498_;
 wire net30;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire net29;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire net28;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire net27;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire net26;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire net25;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire net24;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire net23;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09456_;
 wire net22;
 wire net21;
 wire net20;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire net19;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire net18;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire net17;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire net16;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire net15;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire net14;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire net13;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire net12;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire net11;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire net10;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire net9;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire net8;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire net7;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire net6;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire net5;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire net4;
 wire _09581_;
 wire net3;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire net2;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire net1;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09627_;
 wire _09628_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09778_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09856_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09863_;
 wire _09867_;
 wire _09868_;
 wire _09870_;
 wire _09871_;
 wire _09873_;
 wire _09876_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09887_;
 wire _09888_;
 wire _09891_;
 wire _09892_;
 wire _09894_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09905_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09928_;
 wire _09931_;
 wire _09932_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09956_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09974_;
 wire _09975_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10020_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10084_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10096_;
 wire _10097_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10553_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10709_;
 wire _10710_;
 wire _10718_;
 wire _10720_;
 wire _10721_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10738_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10745_;
 wire _10748_;
 wire _10750_;
 wire _10751_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10773_;
 wire _10774_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10781_;
 wire _10783_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10802_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10854_;
 wire _10855_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10907_;
 wire _10909_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10929_;
 wire _10930_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10952_;
 wire _10953_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10974_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11391_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11556_;
 wire _11559_;
 wire _11561_;
 wire _11564_;
 wire _11565_;
 wire _11567_;
 wire _11569_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11579_;
 wire _11581_;
 wire _11584_;
 wire _11586_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11597_;
 wire _11599_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11613_;
 wire _11614_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11626_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11633_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11641_;
 wire _11643_;
 wire _11644_;
 wire _11646_;
 wire _11648_;
 wire _11649_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11660_;
 wire _11661_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11681_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11715_;
 wire _11716_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11760_;
 wire _11762_;
 wire _11763_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11808_;
 wire _11809_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11972_;
 wire _11973_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12400_;
 wire _12401_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12441_;
 wire _12442_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12511_;
 wire _12515_;
 wire _12519_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12531_;
 wire _12538_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12547_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12560_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12576_;
 wire _12577_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12584_;
 wire _12586_;
 wire _12587_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12629_;
 wire _12632_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12654_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12673_;
 wire _12675_;
 wire _12677_;
 wire _12679_;
 wire _12680_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12692_;
 wire _12693_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12782_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12796_;
 wire _12798_;
 wire _12800_;
 wire _12803_;
 wire _12811_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12822_;
 wire _12825_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12832_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12844_;
 wire _12848_;
 wire _12850_;
 wire _12851_;
 wire _12853_;
 wire _12857_;
 wire _12858_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12867_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12877_;
 wire _12879_;
 wire _12881_;
 wire _12883_;
 wire _12885_;
 wire _12886_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12896_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12904_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12919_;
 wire _12922_;
 wire _12924_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12931_;
 wire _12932_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12942_;
 wire _12945_;
 wire _12946_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12970_;
 wire _12971_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13022_;
 wire _13030_;
 wire _13033_;
 wire _13037_;
 wire _13038_;
 wire _13040_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13050_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13057_;
 wire _13062_;
 wire _13063_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13072_;
 wire _13075_;
 wire _13076_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13086_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13100_;
 wire _13101_;
 wire _13104_;
 wire _13106_;
 wire _13108_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13120_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13134_;
 wire _13135_;
 wire _13137_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13146_;
 wire _13147_;
 wire _13149_;
 wire _13150_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13165_;
 wire _13166_;
 wire _13171_;
 wire _13173_;
 wire _13174_;
 wire _13176_;
 wire _13178_;
 wire _13179_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13189_;
 wire _13191_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13277_;
 wire _13279_;
 wire _13280_;
 wire _13282_;
 wire _13283_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13302_;
 wire _13306_;
 wire _13310_;
 wire _13311_;
 wire _13313_;
 wire _13315_;
 wire _13318_;
 wire _13320_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13330_;
 wire _13336_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13343_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13349_;
 wire _13350_;
 wire _13352_;
 wire _13353_;
 wire _13355_;
 wire _13358_;
 wire _13361_;
 wire _13362_;
 wire _13364_;
 wire _13367_;
 wire _13368_;
 wire _13371_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13377_;
 wire _13378_;
 wire _13380_;
 wire _13382_;
 wire _13383_;
 wire _13385_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13392_;
 wire _13393_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13420_;
 wire _13421_;
 wire _13423_;
 wire _13425_;
 wire _13427_;
 wire _13428_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13441_;
 wire _13442_;
 wire _13444_;
 wire _13445_;
 wire _13447_;
 wire _13448_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13454_;
 wire _13455_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13466_;
 wire _13467_;
 wire _13469_;
 wire _13472_;
 wire _13473_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13582_;
 wire _13583_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13670_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13862_;
 wire _13863_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire _15891_;
 wire _15892_;
 wire _15893_;
 wire _15894_;
 wire _15895_;
 wire _15896_;
 wire _15897_;
 wire _15898_;
 wire _15899_;
 wire _15900_;
 wire _15901_;
 wire _15902_;
 wire _15903_;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire _15908_;
 wire _15909_;
 wire _15910_;
 wire _15911_;
 wire _15912_;
 wire _15913_;
 wire _15914_;
 wire _15915_;
 wire _15916_;
 wire _15917_;
 wire _15918_;
 wire _15919_;
 wire _15920_;
 wire _15921_;
 wire _15923_;
 wire _15924_;
 wire _15925_;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15939_;
 wire _15943_;
 wire _15947_;
 wire _15948_;
 wire _15952_;
 wire _15955_;
 wire _15956_;
 wire _15959_;
 wire _15963_;
 wire _15964_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15980_;
 wire _15985_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15993_;
 wire _15995_;
 wire _15997_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16004_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16013_;
 wire _16014_;
 wire _16018_;
 wire _16021_;
 wire _16023_;
 wire _16025_;
 wire _16026_;
 wire _16027_;
 wire _16028_;
 wire _16031_;
 wire _16032_;
 wire _16033_;
 wire _16034_;
 wire _16035_;
 wire _16037_;
 wire _16040_;
 wire _16042_;
 wire _16044_;
 wire _16045_;
 wire _16047_;
 wire _16049_;
 wire _16052_;
 wire _16053_;
 wire _16058_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16064_;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16071_;
 wire _16072_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16080_;
 wire _16082_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16106_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire _16139_;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16152_;
 wire _16153_;
 wire _16155_;
 wire _16156_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire _16164_;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16181_;
 wire _16185_;
 wire _16186_;
 wire _16189_;
 wire _16191_;
 wire _16193_;
 wire _16194_;
 wire _16195_;
 wire _16199_;
 wire _16202_;
 wire _16203_;
 wire _16206_;
 wire _16209_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16219_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire _16225_;
 wire _16226_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16237_;
 wire _16239_;
 wire _16240_;
 wire _16244_;
 wire _16247_;
 wire _16248_;
 wire _16250_;
 wire _16251_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16263_;
 wire _16266_;
 wire _16269_;
 wire _16270_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16282_;
 wire _16283_;
 wire _16285_;
 wire _16287_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16295_;
 wire _16296_;
 wire _16299_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16305_;
 wire _16307_;
 wire _16308_;
 wire _16310_;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16325_;
 wire _16326_;
 wire _16327_;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16332_;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire _16365_;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire _16406_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire _16412_;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16429_;
 wire _16432_;
 wire _16435_;
 wire _16438_;
 wire _16439_;
 wire _16441_;
 wire _16442_;
 wire _16446_;
 wire _16453_;
 wire _16454_;
 wire _16456_;
 wire _16458_;
 wire _16460_;
 wire _16461_;
 wire _16464_;
 wire _16466_;
 wire _16468_;
 wire _16473_;
 wire _16475_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16494_;
 wire _16495_;
 wire _16497_;
 wire _16498_;
 wire _16500_;
 wire clknet_opt_1_1_clk;
 wire _16503_;
 wire _16504_;
 wire clknet_opt_1_0_clk;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire clknet_1_1__leaf_clk;
 wire _16510_;
 wire _16511_;
 wire clknet_1_0__leaf_clk;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire clknet_0_clk;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_16_clk;
 wire _16535_;
 wire _16536_;
 wire clknet_leaf_15_clk;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire clknet_leaf_14_clk;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire clknet_leaf_13_clk;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_9_clk;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_7_clk;
 wire _16561_;
 wire clknet_leaf_6_clk;
 wire _16563_;
 wire _16564_;
 wire clknet_leaf_5_clk;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_3_clk;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire clknet_leaf_2_clk;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire clknet_leaf_1_clk;
 wire _16579_;
 wire clknet_leaf_0_clk;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire net948;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire net947;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire net946;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire net945;
 wire _16637_;
 wire _16638_;
 wire net944;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire net943;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire net942;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire net941;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire net940;
 wire net939;
 wire _16693_;
 wire net938;
 wire net937;
 wire net936;
 wire net935;
 wire net934;
 wire net933;
 wire net932;
 wire net931;
 wire _16702_;
 wire net930;
 wire net929;
 wire net928;
 wire net927;
 wire net926;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire net925;
 wire _16713_;
 wire net924;
 wire _16715_;
 wire net923;
 wire net922;
 wire net921;
 wire _16719_;
 wire net920;
 wire _16721_;
 wire net919;
 wire net918;
 wire net917;
 wire _16725_;
 wire _16726_;
 wire net916;
 wire _16728_;
 wire _16729_;
 wire net915;
 wire _16731_;
 wire net914;
 wire net913;
 wire net912;
 wire _16735_;
 wire net911;
 wire net910;
 wire net909;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire net908;
 wire _16746_;
 wire net907;
 wire _16748_;
 wire net906;
 wire _16750_;
 wire _16751_;
 wire net905;
 wire net904;
 wire net903;
 wire _16755_;
 wire net902;
 wire net901;
 wire _16758_;
 wire net900;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire net899;
 wire net898;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire net897;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire net896;
 wire net895;
 wire _16778_;
 wire net894;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire net893;
 wire net892;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire net891;
 wire _16798_;
 wire net890;
 wire _16800_;
 wire net889;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire net888;
 wire _16806_;
 wire _16807_;
 wire net887;
 wire net886;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire net885;
 wire net884;
 wire net883;
 wire net882;
 wire _16820_;
 wire net881;
 wire net880;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire net879;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire net878;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire net877;
 wire _16838_;
 wire _16839_;
 wire net876;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire net875;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire net874;
 wire net873;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire net872;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire net871;
 wire _16877_;
 wire net870;
 wire net869;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire net868;
 wire net867;
 wire net866;
 wire _16887_;
 wire _16888_;
 wire net865;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire net864;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire net863;
 wire _16912_;
 wire net862;
 wire _16914_;
 wire _16915_;
 wire net861;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire net860;
 wire _16921_;
 wire _16922_;
 wire net859;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire net858;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire net857;
 wire _16944_;
 wire net856;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire net855;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire net854;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire net853;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire net852;
 wire _16993_;
 wire net851;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire net850;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire net849;
 wire net848;
 wire _17076_;
 wire _17077_;
 wire net847;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire net846;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire net845;
 wire net844;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire net843;
 wire net842;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire _17121_;
 wire _17122_;
 wire net841;
 wire _17124_;
 wire _17125_;
 wire net840;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire net839;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire net838;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire net837;
 wire net836;
 wire _17143_;
 wire net835;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire net834;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire net833;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire net832;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire net831;
 wire net830;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire net829;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire net828;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire net827;
 wire net826;
 wire _17292_;
 wire net825;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire net824;
 wire net823;
 wire _17307_;
 wire net822;
 wire _17309_;
 wire net821;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire net820;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire net819;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire net818;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire net817;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire net816;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire net815;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire net814;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire net813;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire net812;
 wire net811;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire net810;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire net809;
 wire net808;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire net807;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire net806;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire net805;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire net804;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire net803;
 wire _17589_;
 wire _17590_;
 wire net802;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire \dcnt[0] ;
 wire \dcnt[1] ;
 wire \dcnt[2] ;
 wire \dcnt[3] ;
 wire ld_r;
 wire \text_in_r[0] ;
 wire \text_in_r[100] ;
 wire \text_in_r[101] ;
 wire \text_in_r[102] ;
 wire \text_in_r[103] ;
 wire \text_in_r[104] ;
 wire \text_in_r[105] ;
 wire \text_in_r[106] ;
 wire \text_in_r[107] ;
 wire \text_in_r[108] ;
 wire \text_in_r[109] ;
 wire \text_in_r[10] ;
 wire \text_in_r[110] ;
 wire \text_in_r[111] ;
 wire \text_in_r[112] ;
 wire \text_in_r[113] ;
 wire \text_in_r[114] ;
 wire \text_in_r[115] ;
 wire \text_in_r[116] ;
 wire \text_in_r[117] ;
 wire \text_in_r[118] ;
 wire \text_in_r[119] ;
 wire \text_in_r[11] ;
 wire \text_in_r[120] ;
 wire \text_in_r[121] ;
 wire \text_in_r[122] ;
 wire \text_in_r[123] ;
 wire \text_in_r[124] ;
 wire \text_in_r[125] ;
 wire \text_in_r[126] ;
 wire \text_in_r[127] ;
 wire \text_in_r[12] ;
 wire \text_in_r[13] ;
 wire \text_in_r[14] ;
 wire \text_in_r[15] ;
 wire \text_in_r[16] ;
 wire \text_in_r[17] ;
 wire \text_in_r[18] ;
 wire \text_in_r[19] ;
 wire \text_in_r[1] ;
 wire \text_in_r[20] ;
 wire \text_in_r[21] ;
 wire \text_in_r[22] ;
 wire \text_in_r[23] ;
 wire \text_in_r[24] ;
 wire \text_in_r[25] ;
 wire \text_in_r[26] ;
 wire \text_in_r[27] ;
 wire \text_in_r[28] ;
 wire \text_in_r[29] ;
 wire \text_in_r[2] ;
 wire \text_in_r[30] ;
 wire \text_in_r[31] ;
 wire \text_in_r[32] ;
 wire \text_in_r[33] ;
 wire \text_in_r[34] ;
 wire \text_in_r[35] ;
 wire \text_in_r[36] ;
 wire \text_in_r[37] ;
 wire \text_in_r[38] ;
 wire \text_in_r[39] ;
 wire \text_in_r[3] ;
 wire \text_in_r[40] ;
 wire \text_in_r[41] ;
 wire \text_in_r[42] ;
 wire \text_in_r[43] ;
 wire \text_in_r[44] ;
 wire \text_in_r[45] ;
 wire \text_in_r[46] ;
 wire \text_in_r[47] ;
 wire \text_in_r[48] ;
 wire \text_in_r[49] ;
 wire \text_in_r[4] ;
 wire \text_in_r[50] ;
 wire \text_in_r[51] ;
 wire \text_in_r[52] ;
 wire \text_in_r[53] ;
 wire \text_in_r[54] ;
 wire \text_in_r[55] ;
 wire \text_in_r[56] ;
 wire \text_in_r[57] ;
 wire \text_in_r[58] ;
 wire \text_in_r[59] ;
 wire \text_in_r[5] ;
 wire \text_in_r[60] ;
 wire \text_in_r[61] ;
 wire \text_in_r[62] ;
 wire \text_in_r[63] ;
 wire \text_in_r[64] ;
 wire \text_in_r[65] ;
 wire \text_in_r[66] ;
 wire \text_in_r[67] ;
 wire \text_in_r[68] ;
 wire \text_in_r[69] ;
 wire \text_in_r[6] ;
 wire \text_in_r[70] ;
 wire \text_in_r[71] ;
 wire \text_in_r[72] ;
 wire \text_in_r[73] ;
 wire \text_in_r[74] ;
 wire \text_in_r[75] ;
 wire \text_in_r[76] ;
 wire \text_in_r[77] ;
 wire \text_in_r[78] ;
 wire \text_in_r[79] ;
 wire \text_in_r[7] ;
 wire \text_in_r[80] ;
 wire \text_in_r[81] ;
 wire \text_in_r[82] ;
 wire \text_in_r[83] ;
 wire \text_in_r[84] ;
 wire \text_in_r[85] ;
 wire \text_in_r[86] ;
 wire \text_in_r[87] ;
 wire \text_in_r[88] ;
 wire \text_in_r[89] ;
 wire \text_in_r[8] ;
 wire \text_in_r[90] ;
 wire \text_in_r[91] ;
 wire \text_in_r[92] ;
 wire \text_in_r[93] ;
 wire \text_in_r[94] ;
 wire \text_in_r[95] ;
 wire \text_in_r[96] ;
 wire \text_in_r[97] ;
 wire \text_in_r[98] ;
 wire \text_in_r[99] ;
 wire \text_in_r[9] ;
 wire \u0.r0.out[24] ;
 wire \u0.r0.out[25] ;
 wire \u0.r0.out[26] ;
 wire \u0.r0.out[27] ;
 wire \u0.r0.out[28] ;
 wire \u0.r0.out[29] ;
 wire \u0.r0.out[30] ;
 wire \u0.r0.out[31] ;
 wire \u0.r0.rcnt[0] ;
 wire \u0.r0.rcnt[1] ;
 wire \u0.r0.rcnt[2] ;
 wire \u0.r0.rcnt[3] ;
 wire \u0.tmp_w[0] ;
 wire \u0.tmp_w[10] ;
 wire \u0.tmp_w[11] ;
 wire \u0.tmp_w[12] ;
 wire \u0.tmp_w[13] ;
 wire \u0.tmp_w[14] ;
 wire \u0.tmp_w[15] ;
 wire \u0.tmp_w[16] ;
 wire \u0.tmp_w[17] ;
 wire \u0.tmp_w[18] ;
 wire \u0.tmp_w[19] ;
 wire \u0.tmp_w[1] ;
 wire \u0.tmp_w[20] ;
 wire \u0.tmp_w[21] ;
 wire \u0.tmp_w[22] ;
 wire \u0.tmp_w[23] ;
 wire \u0.tmp_w[24] ;
 wire \u0.tmp_w[25] ;
 wire \u0.tmp_w[26] ;
 wire \u0.tmp_w[27] ;
 wire \u0.tmp_w[28] ;
 wire \u0.tmp_w[29] ;
 wire \u0.tmp_w[2] ;
 wire \u0.tmp_w[30] ;
 wire \u0.tmp_w[31] ;
 wire \u0.tmp_w[3] ;
 wire \u0.tmp_w[4] ;
 wire \u0.tmp_w[5] ;
 wire \u0.tmp_w[6] ;
 wire \u0.tmp_w[7] ;
 wire \u0.tmp_w[8] ;
 wire \u0.tmp_w[9] ;
 wire \u0.w[0][0] ;
 wire \u0.w[0][10] ;
 wire \u0.w[0][11] ;
 wire \u0.w[0][12] ;
 wire \u0.w[0][13] ;
 wire \u0.w[0][14] ;
 wire \u0.w[0][15] ;
 wire \u0.w[0][16] ;
 wire \u0.w[0][17] ;
 wire \u0.w[0][18] ;
 wire \u0.w[0][19] ;
 wire \u0.w[0][1] ;
 wire \u0.w[0][20] ;
 wire \u0.w[0][21] ;
 wire \u0.w[0][22] ;
 wire \u0.w[0][23] ;
 wire \u0.w[0][24] ;
 wire \u0.w[0][25] ;
 wire \u0.w[0][26] ;
 wire \u0.w[0][27] ;
 wire \u0.w[0][28] ;
 wire \u0.w[0][29] ;
 wire \u0.w[0][2] ;
 wire \u0.w[0][30] ;
 wire \u0.w[0][31] ;
 wire \u0.w[0][3] ;
 wire \u0.w[0][4] ;
 wire \u0.w[0][5] ;
 wire \u0.w[0][6] ;
 wire \u0.w[0][7] ;
 wire \u0.w[0][8] ;
 wire \u0.w[0][9] ;
 wire \u0.w[1][0] ;
 wire \u0.w[1][10] ;
 wire \u0.w[1][11] ;
 wire \u0.w[1][12] ;
 wire \u0.w[1][13] ;
 wire \u0.w[1][14] ;
 wire \u0.w[1][15] ;
 wire \u0.w[1][16] ;
 wire \u0.w[1][17] ;
 wire \u0.w[1][18] ;
 wire \u0.w[1][19] ;
 wire \u0.w[1][1] ;
 wire \u0.w[1][20] ;
 wire \u0.w[1][21] ;
 wire \u0.w[1][22] ;
 wire \u0.w[1][23] ;
 wire \u0.w[1][24] ;
 wire \u0.w[1][25] ;
 wire \u0.w[1][26] ;
 wire \u0.w[1][27] ;
 wire \u0.w[1][28] ;
 wire \u0.w[1][29] ;
 wire \u0.w[1][2] ;
 wire \u0.w[1][30] ;
 wire \u0.w[1][31] ;
 wire \u0.w[1][3] ;
 wire \u0.w[1][4] ;
 wire \u0.w[1][5] ;
 wire \u0.w[1][6] ;
 wire \u0.w[1][7] ;
 wire \u0.w[1][8] ;
 wire \u0.w[1][9] ;
 wire \u0.w[2][0] ;
 wire \u0.w[2][10] ;
 wire \u0.w[2][11] ;
 wire \u0.w[2][12] ;
 wire \u0.w[2][13] ;
 wire \u0.w[2][14] ;
 wire \u0.w[2][15] ;
 wire \u0.w[2][16] ;
 wire \u0.w[2][17] ;
 wire \u0.w[2][18] ;
 wire \u0.w[2][19] ;
 wire \u0.w[2][1] ;
 wire \u0.w[2][20] ;
 wire \u0.w[2][21] ;
 wire \u0.w[2][22] ;
 wire \u0.w[2][23] ;
 wire \u0.w[2][24] ;
 wire \u0.w[2][25] ;
 wire \u0.w[2][26] ;
 wire \u0.w[2][27] ;
 wire \u0.w[2][28] ;
 wire \u0.w[2][29] ;
 wire \u0.w[2][2] ;
 wire \u0.w[2][30] ;
 wire \u0.w[2][31] ;
 wire \u0.w[2][3] ;
 wire \u0.w[2][4] ;
 wire \u0.w[2][5] ;
 wire \u0.w[2][6] ;
 wire \u0.w[2][7] ;
 wire \u0.w[2][8] ;
 wire \u0.w[2][9] ;
 wire \us00.a[0] ;
 wire \us00.a[1] ;
 wire \us00.a[2] ;
 wire \us00.a[3] ;
 wire \us00.a[4] ;
 wire \us00.a[5] ;
 wire \us00.a[6] ;
 wire \us00.a[7] ;
 wire \us01.a[0] ;
 wire \us01.a[1] ;
 wire \us01.a[2] ;
 wire \us01.a[3] ;
 wire \us01.a[4] ;
 wire \us01.a[5] ;
 wire \us01.a[6] ;
 wire \us01.a[7] ;
 wire \us02.a[0] ;
 wire \us02.a[1] ;
 wire \us02.a[2] ;
 wire \us02.a[3] ;
 wire \us02.a[4] ;
 wire \us02.a[5] ;
 wire \us02.a[6] ;
 wire \us02.a[7] ;
 wire \us03.a[0] ;
 wire \us03.a[1] ;
 wire \us03.a[2] ;
 wire \us03.a[3] ;
 wire \us03.a[4] ;
 wire \us03.a[5] ;
 wire \us03.a[6] ;
 wire \us03.a[7] ;
 wire \us10.a[0] ;
 wire \us10.a[1] ;
 wire \us10.a[2] ;
 wire \us10.a[3] ;
 wire \us10.a[4] ;
 wire \us10.a[5] ;
 wire \us10.a[6] ;
 wire \us10.a[7] ;
 wire \us11.a[0] ;
 wire \us11.a[1] ;
 wire \us11.a[2] ;
 wire \us11.a[3] ;
 wire \us11.a[4] ;
 wire \us11.a[5] ;
 wire \us11.a[6] ;
 wire \us11.a[7] ;
 wire \us12.a[0] ;
 wire \us12.a[1] ;
 wire \us12.a[2] ;
 wire \us12.a[3] ;
 wire \us12.a[4] ;
 wire \us12.a[5] ;
 wire \us12.a[6] ;
 wire \us12.a[7] ;
 wire \us13.a[0] ;
 wire \us13.a[1] ;
 wire \us13.a[2] ;
 wire \us13.a[3] ;
 wire \us13.a[4] ;
 wire \us13.a[5] ;
 wire \us13.a[6] ;
 wire \us13.a[7] ;
 wire \us20.a[0] ;
 wire \us20.a[1] ;
 wire \us20.a[2] ;
 wire \us20.a[3] ;
 wire \us20.a[4] ;
 wire \us20.a[5] ;
 wire \us20.a[6] ;
 wire \us20.a[7] ;
 wire \us21.a[0] ;
 wire \us21.a[1] ;
 wire \us21.a[2] ;
 wire \us21.a[3] ;
 wire \us21.a[4] ;
 wire \us21.a[5] ;
 wire \us21.a[6] ;
 wire \us21.a[7] ;
 wire \us22.a[0] ;
 wire \us22.a[1] ;
 wire \us22.a[2] ;
 wire \us22.a[3] ;
 wire \us22.a[4] ;
 wire \us22.a[5] ;
 wire \us22.a[6] ;
 wire \us22.a[7] ;
 wire \us23.a[0] ;
 wire \us23.a[1] ;
 wire \us23.a[2] ;
 wire \us23.a[3] ;
 wire \us23.a[4] ;
 wire \us23.a[5] ;
 wire \us23.a[6] ;
 wire \us23.a[7] ;
 wire \us30.a[0] ;
 wire \us30.a[1] ;
 wire \us30.a[2] ;
 wire \us30.a[3] ;
 wire \us30.a[4] ;
 wire \us30.a[5] ;
 wire \us30.a[6] ;
 wire \us30.a[7] ;
 wire \us31.a[0] ;
 wire \us31.a[1] ;
 wire \us31.a[2] ;
 wire \us31.a[3] ;
 wire \us31.a[4] ;
 wire \us31.a[5] ;
 wire \us31.a[6] ;
 wire \us31.a[7] ;
 wire \us32.a[0] ;
 wire \us32.a[1] ;
 wire \us32.a[2] ;
 wire \us32.a[3] ;
 wire \us32.a[4] ;
 wire \us32.a[5] ;
 wire \us32.a[6] ;
 wire \us32.a[7] ;
 wire \us33.a[0] ;
 wire \us33.a[1] ;
 wire \us33.a[2] ;
 wire \us33.a[3] ;
 wire \us33.a[4] ;
 wire \us33.a[5] ;
 wire \us33.a[6] ;
 wire \us33.a[7] ;

 b15inv040ah1n02x5 _17617_ (.a(net1),
    .o1(_02399_));
 b15zdnd11an1n64x5 FILLER_1_1624 ();
 b15zdnd00an1n01x5 FILLER_1_1603 ();
 b15zdnd00an1n02x5 FILLER_1_1601 ();
 b15zdnd11an1n08x5 FILLER_1_1593 ();
 b15zdnd11an1n04x5 FILLER_1_1569 ();
 b15zdnd11an1n04x5 FILLER_1_1560 ();
 b15zdnd00an1n01x5 FILLER_1_1539 ();
 b15zdnd11an1n16x5 FILLER_1_1523 ();
 b15zdnd11an1n32x5 FILLER_1_1491 ();
 b15zdnd00an1n01x5 FILLER_1_1486 ();
 b15zdnd11an1n16x5 FILLER_1_1470 ();
 b15zdnd11an1n32x5 FILLER_1_1438 ();
 b15zdnd00an1n02x5 FILLER_1_1432 ();
 b15zdnd11an1n08x5 FILLER_1_1424 ();
 b15zdnd11an1n32x5 FILLER_1_1392 ();
 b15nona23aq1n24x5 _17633_ (.a(net415),
    .b(net412),
    .c(net405),
    .d(net409),
    .out0(_02575_));
 b15norp02ar1n02x5 _17634_ (.a(net427),
    .b(_02575_),
    .o1(_02586_));
 b15nonb02as1n16x5 _17635_ (.a(net405),
    .b(net410),
    .out0(_02597_));
 b15zdnd11an1n04x5 FILLER_1_1384 ();
 b15norp02as1n48x5 _17637_ (.a(net416),
    .b(\u0.tmp_w[29] ),
    .o1(_02619_));
 b15and002ah1n16x5 _17638_ (.a(_02597_),
    .b(_02619_),
    .o(_02630_));
 b15zdnd00an1n02x5 FILLER_1_1362 ();
 b15zdnd11an1n08x5 FILLER_1_1354 ();
 b15zdnd00an1n01x5 FILLER_1_1348 ();
 b15aoai13ar1n02x5 _17642_ (.a(\u0.tmp_w[26] ),
    .b(_02586_),
    .c(_02630_),
    .d(net427),
    .o1(_02674_));
 b15zdnd11an1n04x5 FILLER_1_1344 ();
 b15inv020ah1n64x5 _17644_ (.a(net419),
    .o1(_02696_));
 b15zdnd00an1n01x5 FILLER_1_1338 ();
 b15zdnd11an1n04x5 FILLER_1_1334 ();
 b15zdnd00an1n01x5 FILLER_1_1327 ();
 b15zdnd11an1n08x5 FILLER_1_1319 ();
 b15zdnd11an1n04x5 FILLER_1_1311 ();
 b15aoi012ar1n02x5 _17650_ (.a(_02696_),
    .b(_02630_),
    .c(net432),
    .o1(_02762_));
 b15and002ar1n02x5 _17651_ (.a(_02674_),
    .b(_02762_),
    .o(_02773_));
 b15inv000al1n48x5 _17652_ (.a(net431),
    .o1(_02784_));
 b15zdnd00an1n01x5 FILLER_1_1304 ();
 b15zdnd00an1n02x5 FILLER_1_1302 ();
 b15zdnd11an1n04x5 FILLER_1_1298 ();
 b15zdnd00an1n01x5 FILLER_1_1293 ();
 b15nona23ah1n16x5 _17657_ (.a(net412),
    .b(net409),
    .c(net405),
    .d(net415),
    .out0(_02839_));
 b15nanb02as1n24x5 _17658_ (.a(net423),
    .b(net425),
    .out0(_02850_));
 b15zdnd11an1n04x5 FILLER_1_1289 ();
 b15zdnd11an1n04x5 FILLER_1_1281 ();
 b15zdnd00an1n01x5 FILLER_1_1276 ();
 b15nona23al1n32x5 _17662_ (.a(net415),
    .b(net409),
    .c(net405),
    .d(net412),
    .out0(_02894_));
 b15zdnd11an1n04x5 FILLER_1_1272 ();
 b15nanb02as1n24x5 _17664_ (.a(net428),
    .b(net424),
    .out0(_02916_));
 b15oai022ar1n02x5 _17665_ (.a(_02839_),
    .b(_02850_),
    .c(_02894_),
    .d(_02916_),
    .o1(_02927_));
 b15nand02ar1n02x5 _17666_ (.a(_02784_),
    .b(_02927_),
    .o1(_02938_));
 b15nonb02as1n16x5 _17667_ (.a(net428),
    .b(net424),
    .out0(_02949_));
 b15nor004as1n12x5 _17668_ (.a(\u0.tmp_w[28] ),
    .b(\u0.tmp_w[29] ),
    .c(\u0.tmp_w[31] ),
    .d(net408),
    .o1(_02960_));
 b15zdnd11an1n04x5 FILLER_1_1263 ();
 b15nand02ah1n04x5 _17670_ (.a(_02949_),
    .b(_02960_),
    .o1(_02982_));
 b15zdnd11an1n04x5 FILLER_1_1255 ();
 b15nano23as1n24x5 _17672_ (.a(net412),
    .b(net409),
    .c(net405),
    .d(net415),
    .out0(_03004_));
 b15zdnd00an1n01x5 FILLER_1_1248 ();
 b15inv040an1n36x5 _17674_ (.a(net427),
    .o1(_03026_));
 b15zdnd00an1n02x5 FILLER_1_1246 ();
 b15aoai13ar1n02x5 _17676_ (.a(net424),
    .b(_03004_),
    .c(_02630_),
    .d(_03026_),
    .o1(_03048_));
 b15nand04al1n02x5 _17677_ (.a(_02696_),
    .b(_02938_),
    .c(_02982_),
    .d(_03048_),
    .o1(_03059_));
 b15zdnd11an1n04x5 FILLER_1_1242 ();
 b15zdnd11an1n04x5 FILLER_1_1234 ();
 b15nona23as1n32x5 _17680_ (.a(net415),
    .b(net405),
    .c(net409),
    .d(net412),
    .out0(_03092_));
 b15zdnd11an1n04x5 FILLER_1_1226 ();
 b15zdnd11an1n08x5 FILLER_1_1218 ();
 b15xnr002ar1n16x5 _17683_ (.a(net408),
    .b(net422),
    .out0(_03125_));
 b15zdnd11an1n04x5 FILLER_1_1207 ();
 b15nanb02al1n24x5 _17685_ (.a(net425),
    .b(\u0.tmp_w[28] ),
    .out0(_03147_));
 b15zdnd00an1n01x5 FILLER_1_1201 ();
 b15zdnd00an1n02x5 FILLER_1_1199 ();
 b15nanb02as1n12x5 _17688_ (.a(net407),
    .b(net422),
    .out0(_03180_));
 b15obai22aq1n12x5 _17689_ (.a(_03125_),
    .b(_03147_),
    .c(\u0.tmp_w[28] ),
    .d(_03180_),
    .out0(_03191_));
 b15nonb02as1n16x5 _17690_ (.a(net423),
    .b(net425),
    .out0(_03202_));
 b15nor002an1n24x5 _17691_ (.a(net416),
    .b(net408),
    .o1(_03213_));
 b15aoi022as1n08x5 _17692_ (.a(\u0.tmp_w[31] ),
    .b(_03191_),
    .c(_03202_),
    .d(_03213_),
    .o1(_03224_));
 b15zdnd11an1n04x5 FILLER_1_1195 ();
 b15zdnd11an1n04x5 FILLER_1_1186 ();
 b15oaoi13al1n08x5 _17695_ (.a(_02784_),
    .b(_03092_),
    .c(_03224_),
    .d(\u0.tmp_w[29] ),
    .o1(_03257_));
 b15oab012aq1n04x5 _17696_ (.a(_02773_),
    .b(_03059_),
    .c(_03257_),
    .out0(_03268_));
 b15zdnd11an1n04x5 FILLER_1_1178 ();
 b15zdnd11an1n08x5 FILLER_1_1164 ();
 b15nandp2ar1n32x5 _17699_ (.a(net428),
    .b(net420),
    .o1(_03301_));
 b15oai012ar1n02x5 _17700_ (.a(\u0.tmp_w[26] ),
    .b(_02839_),
    .c(_03301_),
    .o1(_03312_));
 b15zdnd00an1n01x5 FILLER_1_1159 ();
 b15norp02ar1n48x5 _17702_ (.a(net428),
    .b(net420),
    .o1(_03334_));
 b15oai012ar1n02x5 _17703_ (.a(_03301_),
    .b(_03334_),
    .c(net432),
    .o1(_03345_));
 b15nanb02ah1n24x5 _17704_ (.a(net414),
    .b(net412),
    .out0(_03356_));
 b15orn002al1n16x5 _17705_ (.a(net404),
    .b(net410),
    .o(_03367_));
 b15norp02an1n24x5 _17706_ (.a(_03356_),
    .b(_03367_),
    .o1(_03378_));
 b15aoi012ah1n02x5 _17707_ (.a(_03312_),
    .b(_03345_),
    .c(_03378_),
    .o1(_03389_));
 b15zdnd00an1n02x5 FILLER_1_1157 ();
 b15zdnd11an1n04x5 FILLER_1_1153 ();
 b15norp03aq1n16x5 _17710_ (.a(net405),
    .b(net409),
    .c(net418),
    .o1(_03421_));
 b15nonb02as1n16x5 _17711_ (.a(net431),
    .b(net428),
    .out0(_03432_));
 b15nonb02as1n16x5 _17712_ (.a(\u0.tmp_w[29] ),
    .b(\u0.tmp_w[28] ),
    .out0(_03443_));
 b15nonb02as1n16x5 _17713_ (.a(net416),
    .b(\u0.tmp_w[29] ),
    .out0(_03454_));
 b15zdnd00an1n01x5 FILLER_1_1148 ();
 b15oai112ah1n16x5 _17715_ (.a(_03421_),
    .b(_03432_),
    .c(_03443_),
    .d(_03454_),
    .o1(_03476_));
 b15zdnd00an1n02x5 FILLER_1_1146 ();
 b15orn002ah1n08x5 _17717_ (.a(net430),
    .b(net419),
    .o(_03498_));
 b15zdnd11an1n08x5 FILLER_1_1138 ();
 b15zdnd11an1n04x5 FILLER_1_1127 ();
 b15nano23as1n24x5 _17720_ (.a(net405),
    .b(net409),
    .c(net415),
    .d(net412),
    .out0(_03531_));
 b15nand02ar1n02x5 _17721_ (.a(net427),
    .b(_03531_),
    .o1(_03542_));
 b15and002aq1n32x5 _17722_ (.a(\u0.tmp_w[31] ),
    .b(net409),
    .o(_03553_));
 b15nand02ar1n32x5 _17723_ (.a(_03443_),
    .b(_03553_),
    .o1(_03564_));
 b15oaoi13an1n02x5 _17724_ (.a(_03498_),
    .b(_03542_),
    .c(net427),
    .d(_03564_),
    .o1(_03575_));
 b15nanb02as1n24x5 _17725_ (.a(net420),
    .b(net428),
    .out0(_03586_));
 b15oai022ar1n02x5 _17726_ (.a(_02696_),
    .b(_02575_),
    .c(_03564_),
    .d(_03586_),
    .o1(_03597_));
 b15zdnd11an1n04x5 FILLER_1_1119 ();
 b15zdnd11an1n04x5 FILLER_1_1111 ();
 b15aoi012ah1n02x5 _17729_ (.a(_03575_),
    .b(_03597_),
    .c(net432),
    .o1(_03630_));
 b15zdnd11an1n04x5 FILLER_1_1103 ();
 b15zdnd11an1n08x5 FILLER_1_1095 ();
 b15zdnd11an1n04x5 FILLER_1_1086 ();
 b15and003ah1n12x5 _17733_ (.a(\u0.tmp_w[28] ),
    .b(\u0.tmp_w[29] ),
    .c(net419),
    .o(_03674_));
 b15aoi012aq1n02x5 _17734_ (.a(\u0.tmp_w[26] ),
    .b(_03553_),
    .c(_03674_),
    .o1(_03685_));
 b15aoi022aq1n08x5 _17735_ (.a(_03389_),
    .b(_03476_),
    .c(_03630_),
    .d(_03685_),
    .o1(_03696_));
 b15zdnd11an1n04x5 FILLER_1_1078 ();
 b15and002ah1n16x5 _17737_ (.a(net416),
    .b(net406),
    .o(_03718_));
 b15nor002ah1n16x5 _17738_ (.a(net410),
    .b(net428),
    .o1(_03729_));
 b15nonb03ah1n08x5 _17739_ (.a(net410),
    .b(net404),
    .c(net415),
    .out0(_03740_));
 b15zdnd11an1n04x5 FILLER_1_1070 ();
 b15and002as1n08x5 _17741_ (.a(net426),
    .b(net417),
    .o(_03762_));
 b15aoi022ar1n02x5 _17742_ (.a(_03718_),
    .b(_03729_),
    .c(_03740_),
    .d(_03762_),
    .o1(_03773_));
 b15nand02al1n12x5 _17743_ (.a(net413),
    .b(net422),
    .o1(_03784_));
 b15norp03ah1n02x5 _17744_ (.a(net432),
    .b(_03773_),
    .c(_03784_),
    .o1(_03795_));
 b15nanb02as1n24x5 _17745_ (.a(net411),
    .b(net415),
    .out0(_03806_));
 b15nandp2ah1n16x5 _17746_ (.a(net404),
    .b(net407),
    .o1(_03817_));
 b15nor002an1n08x5 _17747_ (.a(_03806_),
    .b(_03817_),
    .o1(_03828_));
 b15andc04aq1n12x5 _17748_ (.a(net415),
    .b(net412),
    .c(net405),
    .d(net409),
    .o(_03839_));
 b15nonb03aq1n12x5 _17749_ (.a(net421),
    .b(net417),
    .c(net426),
    .out0(_03850_));
 b15aoi022ar1n02x5 _17750_ (.a(_03762_),
    .b(_03828_),
    .c(_03839_),
    .d(_03850_),
    .o1(_03861_));
 b15oab012aq1n06x5 _17751_ (.a(_03795_),
    .b(_03861_),
    .c(net432),
    .out0(_03872_));
 b15zdnd11an1n08x5 FILLER_1_1062 ();
 b15norp03ar1n02x5 _17753_ (.a(\u0.tmp_w[29] ),
    .b(net423),
    .c(net419),
    .o1(_03894_));
 b15zdnd11an1n08x5 FILLER_1_1050 ();
 b15zdnd11an1n04x5 FILLER_1_1042 ();
 b15zdnd11an1n16x5 FILLER_1_1026 ();
 b15aoi012an1n02x5 _17757_ (.a(_03894_),
    .b(net419),
    .c(\u0.tmp_w[29] ),
    .o1(_03937_));
 b15zdnd00an1n02x5 FILLER_1_1019 ();
 b15nonb02aq1n12x5 _17759_ (.a(net407),
    .b(net432),
    .out0(_03959_));
 b15nand03al1n12x5 _17760_ (.a(net427),
    .b(_03718_),
    .c(_03959_),
    .o1(_03970_));
 b15zdnd11an1n08x5 FILLER_1_1011 ();
 b15zdnd00an1n01x5 FILLER_1_1006 ();
 b15zdnd11an1n04x5 FILLER_1_1002 ();
 b15nonb02as1n04x5 _17764_ (.a(net409),
    .b(net416),
    .out0(_04014_));
 b15and002aq1n16x5 _17765_ (.a(\u0.tmp_w[29] ),
    .b(\u0.tmp_w[31] ),
    .o(_04025_));
 b15nandp3ar1n03x5 _17766_ (.a(net419),
    .b(_04014_),
    .c(_04025_),
    .o1(_04036_));
 b15nona22al1n32x5 _17767_ (.a(net427),
    .b(net423),
    .c(net430),
    .out0(_04047_));
 b15nanb02aq1n12x5 _17768_ (.a(net430),
    .b(net423),
    .out0(_04058_));
 b15nand02al1n02x5 _17769_ (.a(_04047_),
    .b(_04058_),
    .o1(_04069_));
 b15oai022an1n06x5 _17770_ (.a(_03937_),
    .b(_03970_),
    .c(_04036_),
    .d(_04069_),
    .o1(_04080_));
 b15nanb02as1n24x5 _17771_ (.a(net406),
    .b(net409),
    .out0(_04091_));
 b15nand02al1n48x5 _17772_ (.a(\u0.tmp_w[28] ),
    .b(net413),
    .o1(_04102_));
 b15nor002an1n24x5 _17773_ (.a(_04091_),
    .b(_04102_),
    .o1(_04113_));
 b15zdnd00an1n01x5 FILLER_1_997 ();
 b15oai012ar1n02x5 _17775_ (.a(net430),
    .b(_02696_),
    .c(_03202_),
    .o1(_04135_));
 b15orn002as1n16x5 _17776_ (.a(net425),
    .b(net423),
    .o(_04146_));
 b15oai012an1n04x5 _17777_ (.a(_04135_),
    .b(_04146_),
    .c(net418),
    .o1(_04157_));
 b15inv000aq1n48x5 _17778_ (.a(net422),
    .o1(_04168_));
 b15nandp2ah1n08x5 _17779_ (.a(net430),
    .b(_04168_),
    .o1(_04179_));
 b15zdnd11an1n04x5 FILLER_1_993 ();
 b15nand02al1n16x5 _17781_ (.a(net423),
    .b(net419),
    .o1(_04201_));
 b15zdnd11an1n08x5 FILLER_1_985 ();
 b15oaoi13aq1n03x5 _17783_ (.a(_03026_),
    .b(_04179_),
    .c(_04201_),
    .d(net430),
    .o1(_04223_));
 b15oaoi13as1n04x5 _17784_ (.a(_04080_),
    .b(_04113_),
    .c(_04157_),
    .d(_04223_),
    .o1(_04234_));
 b15zdnd11an1n04x5 FILLER_1_977 ();
 b15zdnd00an1n02x5 FILLER_1_971 ();
 b15nano23as1n24x5 _17787_ (.a(net415),
    .b(net412),
    .c(net405),
    .d(net409),
    .out0(_04267_));
 b15nandp2al1n08x5 _17788_ (.a(\u0.tmp_w[26] ),
    .b(_04267_),
    .o1(_04278_));
 b15oai012al1n06x5 _17789_ (.a(_02982_),
    .b(_04278_),
    .c(net427),
    .o1(_04289_));
 b15zdnd11an1n04x5 FILLER_1_967 ();
 b15nona23as1n32x5 _17791_ (.a(\u0.tmp_w[29] ),
    .b(\u0.tmp_w[31] ),
    .c(net408),
    .d(\u0.tmp_w[28] ),
    .out0(_04311_));
 b15aoai13ah1n03x5 _17792_ (.a(net432),
    .b(_02696_),
    .c(_04311_),
    .d(net427),
    .o1(_04322_));
 b15zdnd00an1n01x5 FILLER_1_962 ();
 b15nonb03aq1n04x5 _17794_ (.a(net409),
    .b(net405),
    .c(net412),
    .out0(_04343_));
 b15aboi22ah1n06x5 _17795_ (.a(\u0.tmp_w[26] ),
    .b(net420),
    .c(net415),
    .d(\u0.tmp_w[25] ),
    .out0(_04354_));
 b15oai122as1n16x5 _17796_ (.a(_04343_),
    .b(_04354_),
    .c(\u0.tmp_w[24] ),
    .d(_03586_),
    .e(net415),
    .o1(_04365_));
 b15nonb02ah1n16x5 _17797_ (.a(net410),
    .b(net405),
    .out0(_04376_));
 b15nandp2al1n12x5 _17798_ (.a(_04376_),
    .b(_02619_),
    .o1(_04387_));
 b15aoi012ar1n04x5 _17799_ (.a(_04365_),
    .b(_04387_),
    .c(_03026_),
    .o1(_04398_));
 b15nanb02ar1n04x5 _17800_ (.a(net426),
    .b(net404),
    .out0(_04409_));
 b15orn002ah1n03x5 _17801_ (.a(net404),
    .b(net421),
    .o(_04420_));
 b15oai022ar1n02x5 _17802_ (.a(_03806_),
    .b(_04409_),
    .c(_04420_),
    .d(_03356_),
    .o1(_04431_));
 b15and002as1n04x5 _17803_ (.a(net407),
    .b(net417),
    .o(_04442_));
 b15nonb02aq1n12x5 _17804_ (.a(net405),
    .b(net419),
    .out0(_04453_));
 b15norp02ar1n08x5 _17805_ (.a(_03125_),
    .b(_04102_),
    .o1(_04464_));
 b15ao0022an1n06x5 _17806_ (.a(_04431_),
    .b(_04442_),
    .c(_04453_),
    .d(_04464_),
    .o(_04475_));
 b15aoi222ah1n08x5 _17807_ (.a(net419),
    .b(_04289_),
    .c(_04322_),
    .d(_04398_),
    .e(_04475_),
    .f(net432),
    .o1(_04486_));
 b15nanb03as1n16x5 _17808_ (.a(net419),
    .b(net423),
    .c(net427),
    .out0(_04497_));
 b15zdnd00an1n02x5 FILLER_1_960 ();
 b15oai112ah1n08x5 _17810_ (.a(_02597_),
    .b(_02850_),
    .c(net430),
    .d(_03202_),
    .o1(_04519_));
 b15zdnd11an1n64x5 FILLER_1_896 ();
 b15nand02ah1n04x5 _17812_ (.a(net418),
    .b(_03443_),
    .o1(_04541_));
 b15oai022al1n16x5 _17813_ (.a(_04311_),
    .b(_04497_),
    .c(_04519_),
    .d(_04541_),
    .o1(_04552_));
 b15zdnd11an1n64x5 FILLER_1_832 ();
 b15nanb02aq1n24x5 _17815_ (.a(net428),
    .b(net417),
    .out0(_04574_));
 b15nandp2ar1n24x5 _17816_ (.a(_02597_),
    .b(_02619_),
    .o1(_04585_));
 b15oai122an1n16x5 _17817_ (.a(_04365_),
    .b(_04574_),
    .c(_03092_),
    .d(_04585_),
    .e(_03498_),
    .o1(_04596_));
 b15nandp3ah1n04x5 _17818_ (.a(net419),
    .b(_03454_),
    .c(_03553_),
    .o1(_04607_));
 b15and002al1n04x5 _17819_ (.a(net430),
    .b(net418),
    .o(_04618_));
 b15norp02aq1n48x5 _17820_ (.a(\u0.tmp_w[31] ),
    .b(net408),
    .o1(_04629_));
 b15zdnd11an1n04x5 FILLER_1_824 ();
 b15aoi012al1n04x5 _17822_ (.a(_04618_),
    .b(_04629_),
    .c(_03443_),
    .o1(_04650_));
 b15nor003as1n04x5 _17823_ (.a(net416),
    .b(net405),
    .c(net409),
    .o1(_04661_));
 b15nanb02ah1n08x5 _17824_ (.a(net430),
    .b(net419),
    .out0(_04672_));
 b15oai122as1n04x5 _17825_ (.a(_04661_),
    .b(_04672_),
    .c(net425),
    .d(_03586_),
    .e(_02784_),
    .o1(_04683_));
 b15and002aq1n24x5 _17826_ (.a(net414),
    .b(net411),
    .o(_04694_));
 b15nandp2as1n04x5 _17827_ (.a(_03553_),
    .b(_04694_),
    .o1(_04705_));
 b15oai122as1n08x5 _17828_ (.a(_04607_),
    .b(_04650_),
    .c(_04683_),
    .d(_04705_),
    .e(_03586_),
    .o1(_04716_));
 b15oaoi13an1n08x5 _17829_ (.a(_04552_),
    .b(_04168_),
    .c(_04596_),
    .d(_04716_),
    .o1(_04727_));
 b15nand04ah1n12x5 _17830_ (.a(_03872_),
    .b(_04234_),
    .c(_04486_),
    .d(_04727_),
    .o1(_04738_));
 b15nand02ah1n32x5 _17831_ (.a(net431),
    .b(net428),
    .o1(_04749_));
 b15norp02al1n24x5 _17832_ (.a(net427),
    .b(\u0.tmp_w[26] ),
    .o1(_04760_));
 b15aoi022ar1n02x5 _17833_ (.a(net423),
    .b(_03531_),
    .c(_04760_),
    .d(_04267_),
    .o1(_04771_));
 b15zdnd11an1n08x5 FILLER_1_816 ();
 b15oai022al1n02x5 _17835_ (.a(_04278_),
    .b(_04749_),
    .c(_04771_),
    .d(net430),
    .o1(_04793_));
 b15xor002as1n16x5 _17836_ (.a(net429),
    .b(net426),
    .out0(_04804_));
 b15nandp3ar1n02x5 _17837_ (.a(net423),
    .b(_02960_),
    .c(_04804_),
    .o1(_04815_));
 b15nandp2an1n16x5 _17838_ (.a(_03454_),
    .b(_04629_),
    .o1(_04826_));
 b15oai013ar1n02x5 _17839_ (.a(_04815_),
    .b(_04804_),
    .c(_04826_),
    .d(net423),
    .o1(_04837_));
 b15zdnd11an1n64x5 FILLER_1_752 ();
 b15nand02aq1n32x5 _17841_ (.a(net430),
    .b(net423),
    .o1(_04859_));
 b15nand04al1n02x5 _17842_ (.a(net427),
    .b(_03454_),
    .c(_04629_),
    .d(_04859_),
    .o1(_04870_));
 b15oai012aq1n04x5 _17843_ (.a(_04870_),
    .b(_03564_),
    .c(_02916_),
    .o1(_04881_));
 b15nor002ah1n16x5 _17844_ (.a(net431),
    .b(net424),
    .o1(_04892_));
 b15aoi013an1n03x5 _17845_ (.a(net418),
    .b(_02597_),
    .c(_04694_),
    .d(_04892_),
    .o1(_04903_));
 b15nanb02al1n08x5 _17846_ (.a(net409),
    .b(net427),
    .out0(_04914_));
 b15nandp3an1n03x5 _17847_ (.a(net416),
    .b(net413),
    .c(net406),
    .o1(_04925_));
 b15nanb02an1n08x5 _17848_ (.a(_04925_),
    .b(_04168_),
    .out0(_04936_));
 b15nonb02ar1n08x5 _17849_ (.a(net421),
    .b(net404),
    .out0(_04947_));
 b15nand02al1n08x5 _17850_ (.a(_02619_),
    .b(_04947_),
    .o1(_04958_));
 b15aoai13as1n08x5 _17851_ (.a(_04903_),
    .b(_04914_),
    .c(_04936_),
    .d(_04958_),
    .o1(_04968_));
 b15oaoi13ah1n03x5 _17852_ (.a(_04793_),
    .b(_04837_),
    .c(_04881_),
    .d(_04968_),
    .o1(_04979_));
 b15nand02ar1n24x5 _17853_ (.a(_04629_),
    .b(_04694_),
    .o1(_04990_));
 b15aoi022ar1n02x5 _17854_ (.a(_02960_),
    .b(_04760_),
    .c(_04267_),
    .d(net427),
    .o1(_05001_));
 b15oa0022as1n02x5 _17855_ (.a(_04179_),
    .b(_04990_),
    .c(_05001_),
    .d(net430),
    .o(_05012_));
 b15nor002ah1n02x5 _17856_ (.a(_04968_),
    .b(_04881_),
    .o1(_05023_));
 b15aoi022an1n12x5 _17857_ (.a(net419),
    .b(_04979_),
    .c(_05012_),
    .d(_05023_),
    .o1(_05034_));
 b15nor004as1n12x5 _17858_ (.a(_03268_),
    .b(_03696_),
    .c(_04738_),
    .d(_05034_),
    .o1(_05045_));
 b15xor002ah1n03x5 _17859_ (.a(\u0.w[0][0] ),
    .b(_05045_),
    .out0(_05056_));
 b15xor002as1n03x5 _17860_ (.a(\u0.w[1][0] ),
    .b(_05056_),
    .out0(_05067_));
 b15xor002al1n03x5 _17861_ (.a(\u0.w[2][0] ),
    .b(_05067_),
    .out0(_05078_));
 b15xor002ar1n02x5 _17862_ (.a(\u0.tmp_w[0] ),
    .b(_05078_),
    .out0(_05089_));
 b15zdnd11an1n64x5 FILLER_1_688 ();
 b15zdnd11an1n64x5 FILLER_1_624 ();
 b15zdnd11an1n64x5 FILLER_1_560 ();
 b15mdn022ar1n02x5 _17866_ (.a(_02399_),
    .b(_05089_),
    .o1(_00353_),
    .sa(net948));
 b15zdnd11an1n64x5 FILLER_1_496 ();
 b15zdnd11an1n64x5 FILLER_1_432 ();
 b15nand02ar1n02x5 _17869_ (.a(net944),
    .b(net40),
    .o1(_05165_));
 b15zdnd11an1n32x5 FILLER_1_384 ();
 b15zdnd11an1n64x5 FILLER_1_320 ();
 b15zdnd11an1n64x5 FILLER_1_256 ();
 b15zdnd11an1n64x5 FILLER_1_192 ();
 b15zdnd11an1n64x5 FILLER_1_128 ();
 b15inv040al1n03x5 _17875_ (.a(\u0.tmp_w[31] ),
    .o1(_05231_));
 b15zdnd11an1n64x5 FILLER_1_64 ();
 b15nandp2ah1n16x5 _17877_ (.a(net409),
    .b(net430),
    .o1(_05252_));
 b15nand04al1n02x5 _17878_ (.a(_05231_),
    .b(net419),
    .c(_02619_),
    .d(_05252_),
    .o1(_05263_));
 b15norp02aq1n48x5 _17879_ (.a(net423),
    .b(net419),
    .o1(_05274_));
 b15zdnd11an1n64x5 FILLER_1_0 ();
 b15norp02ar1n48x5 _17881_ (.a(net413),
    .b(net406),
    .o1(_05296_));
 b15oai112ar1n02x5 _17882_ (.a(_03213_),
    .b(_05274_),
    .c(_05296_),
    .d(_04025_),
    .o1(_05307_));
 b15nandp3ah1n02x5 _17883_ (.a(net425),
    .b(_05263_),
    .c(_05307_),
    .o1(_05318_));
 b15nandp3ar1n02x5 _17884_ (.a(_02619_),
    .b(_03421_),
    .c(_04892_),
    .o1(_05329_));
 b15oai012aq1n03x5 _17885_ (.a(_05329_),
    .b(_04990_),
    .c(_04201_),
    .o1(_05340_));
 b15nano23as1n24x5 _17886_ (.a(net414),
    .b(net404),
    .c(net410),
    .d(net411),
    .out0(_05351_));
 b15norp02ar1n02x5 _17887_ (.a(_05351_),
    .b(_05274_),
    .o1(_05362_));
 b15aoi012al1n04x5 _17888_ (.a(_05362_),
    .b(_04826_),
    .c(_05274_),
    .o1(_05373_));
 b15oai013ah1n04x5 _17889_ (.a(_05318_),
    .b(_05340_),
    .c(_05373_),
    .d(net425),
    .o1(_05384_));
 b15nanb02as1n24x5 _17890_ (.a(net414),
    .b(net410),
    .out0(_05395_));
 b15nand02aq1n04x5 _17891_ (.a(net421),
    .b(_02696_),
    .o1(_05406_));
 b15zdnd00an1n02x5 FILLER_0_2274 ();
 b15nonb02as1n16x5 _17893_ (.a(net406),
    .b(net413),
    .out0(_05428_));
 b15nonb02ar1n02x5 _17894_ (.a(net413),
    .b(net429),
    .out0(_05439_));
 b15aoi022ar1n04x5 _17895_ (.a(net429),
    .b(_05428_),
    .c(_05439_),
    .d(_04409_),
    .o1(_05450_));
 b15norp03aq1n08x5 _17896_ (.a(_05395_),
    .b(_05406_),
    .c(_05450_),
    .o1(_05461_));
 b15orn002aq1n12x5 _17897_ (.a(net429),
    .b(net426),
    .o(_05472_));
 b15oai112aq1n02x5 _17898_ (.a(_05274_),
    .b(_05472_),
    .c(_04267_),
    .d(_03004_),
    .o1(_05483_));
 b15nonb02as1n16x5 _17899_ (.a(net421),
    .b(net418),
    .out0(_05493_));
 b15nanb02as1n24x5 _17900_ (.a(net424),
    .b(net420),
    .out0(_05504_));
 b15zdnd11an1n16x5 FILLER_0_2258 ();
 b15nor002ah1n16x5 _17902_ (.a(net429),
    .b(net426),
    .o1(_05526_));
 b15nona23ar1n04x5 _17903_ (.a(_05493_),
    .b(_04311_),
    .c(_05504_),
    .d(_05526_),
    .out0(_05537_));
 b15and002aq1n03x5 _17904_ (.a(net408),
    .b(net430),
    .o(_05548_));
 b15and002aq1n03x5 _17905_ (.a(net406),
    .b(net425),
    .o(_05559_));
 b15nor003ar1n02x5 _17906_ (.a(net406),
    .b(net425),
    .c(net423),
    .o1(_05570_));
 b15oai112as1n04x5 _17907_ (.a(_03674_),
    .b(_05548_),
    .c(_05559_),
    .d(_05570_),
    .o1(_05581_));
 b15orn002an1n03x5 _17908_ (.a(\u0.tmp_w[28] ),
    .b(net425),
    .o(_05592_));
 b15nand04an1n03x5 _17909_ (.a(_05274_),
    .b(_05428_),
    .c(_05548_),
    .d(_05592_),
    .o1(_05603_));
 b15nand04aq1n03x5 _17910_ (.a(_05483_),
    .b(_05537_),
    .c(_05581_),
    .d(_05603_),
    .o1(_05614_));
 b15and002an1n16x5 _17911_ (.a(net427),
    .b(net423),
    .o(_05625_));
 b15aoi013an1n02x5 _17912_ (.a(net430),
    .b(net418),
    .c(_04267_),
    .d(_05625_),
    .o1(_05636_));
 b15nona22ar1n04x5 _17913_ (.a(\u0.tmp_w[28] ),
    .b(\u0.tmp_w[29] ),
    .c(net408),
    .out0(_05647_));
 b15nanb03ar1n02x5 _17914_ (.a(net408),
    .b(\u0.tmp_w[29] ),
    .c(\u0.tmp_w[28] ),
    .out0(_05658_));
 b15oai022an1n02x5 _17915_ (.a(_04146_),
    .b(_05647_),
    .c(_05658_),
    .d(_03202_),
    .o1(_05669_));
 b15aob012ar1n03x5 _17916_ (.a(_05636_),
    .b(_05669_),
    .c(_04453_),
    .out0(_05680_));
 b15zdnd11an1n32x5 FILLER_0_2226 ();
 b15nand02an1n32x5 _17918_ (.a(net425),
    .b(net423),
    .o1(_05699_));
 b15oab012ar1n02x5 _17919_ (.a(_02784_),
    .b(_04311_),
    .c(_05699_),
    .out0(_05708_));
 b15nanb02as1n16x5 _17920_ (.a(net407),
    .b(net418),
    .out0(_05718_));
 b15nanb02al1n08x5 _17921_ (.a(net418),
    .b(net409),
    .out0(_05727_));
 b15cmbn22ar1n02x5 _17922_ (.clk1(_05718_),
    .clk2(_05727_),
    .clkout(_05736_),
    .s(net406));
 b15oai013as1n02x5 _17923_ (.a(_05708_),
    .b(_05736_),
    .c(_04102_),
    .d(net422),
    .o1(_05746_));
 b15aoi112ar1n04x5 _17924_ (.a(_05461_),
    .b(_05614_),
    .c(_05680_),
    .d(_05746_),
    .o1(_05755_));
 b15zdnd11an1n64x5 FILLER_0_2162 ();
 b15nand02ar1n02x5 _17926_ (.a(net407),
    .b(_04694_),
    .o1(_05774_));
 b15nonb02as1n16x5 _17927_ (.a(net428),
    .b(net431),
    .out0(_05783_));
 b15zdnd00an1n01x5 FILLER_0_2153 ();
 b15oai012ah1n02x5 _17929_ (.a(net404),
    .b(_03334_),
    .c(_05783_),
    .o1(_05801_));
 b15nand02al1n02x5 _17930_ (.a(_02696_),
    .b(_05526_),
    .o1(_05810_));
 b15aoai13al1n04x5 _17931_ (.a(net421),
    .b(_05774_),
    .c(_05801_),
    .d(_05810_),
    .o1(_05820_));
 b15orn002ar1n24x5 _17932_ (.a(net411),
    .b(net404),
    .o(_05831_));
 b15norp02ar1n32x5 _17933_ (.a(_05395_),
    .b(_05831_),
    .o1(_05842_));
 b15nanb02as1n24x5 _17934_ (.a(net429),
    .b(net426),
    .out0(_05853_));
 b15norp02ar1n02x5 _17935_ (.a(net417),
    .b(_05853_),
    .o1(_05864_));
 b15aoi022an1n04x5 _17936_ (.a(net417),
    .b(_05842_),
    .c(_05864_),
    .d(_02630_),
    .o1(_05875_));
 b15aob012ar1n12x5 _17937_ (.a(_05820_),
    .b(_05875_),
    .c(_04168_),
    .out0(_05886_));
 b15nonb02as1n16x5 _17938_ (.a(net413),
    .b(net406),
    .out0(_05897_));
 b15mdn022ar1n03x5 _17939_ (.a(_05897_),
    .b(_05428_),
    .o1(_05908_),
    .sa(net416));
 b15qgbno2an1n05x5 _17940_ (.o1(_05919_),
    .a(net409),
    .b(net418));
 b15nand02ar1n02x5 _17941_ (.a(net430),
    .b(_05919_),
    .o1(_05930_));
 b15aoi022al1n06x5 _17942_ (.a(_02619_),
    .b(_03334_),
    .c(_03674_),
    .d(_04804_),
    .o1(_05941_));
 b15nanb02as1n24x5 _17943_ (.a(net410),
    .b(net404),
    .out0(_05952_));
 b15oai022ar1n04x5 _17944_ (.a(_05908_),
    .b(_05930_),
    .c(_05941_),
    .d(_05952_),
    .o1(_05963_));
 b15aoi012ar1n02x5 _17945_ (.a(_04629_),
    .b(_03959_),
    .c(net406),
    .o1(_05974_));
 b15zdnd11an1n04x5 FILLER_0_2149 ();
 b15oai022ar1n02x5 _17947_ (.a(_03817_),
    .b(_05472_),
    .c(_05974_),
    .d(net416),
    .o1(_05996_));
 b15norp02aq1n03x5 _17948_ (.a(net413),
    .b(_02696_),
    .o1(_06007_));
 b15aoai13as1n02x5 _17949_ (.a(net422),
    .b(_05963_),
    .c(_05996_),
    .d(_06007_),
    .o1(_06018_));
 b15nand04an1n08x5 _17950_ (.a(_05384_),
    .b(_05755_),
    .c(_05886_),
    .d(_06018_),
    .o1(_06029_));
 b15zdnd11an1n08x5 FILLER_0_2141 ();
 b15zdnd11an1n16x5 FILLER_0_2125 ();
 b15nor002al1n04x5 _17953_ (.a(net408),
    .b(net430),
    .o1(_06062_));
 b15aoi013al1n03x5 _17954_ (.a(net419),
    .b(_05296_),
    .c(_06062_),
    .d(net423),
    .o1(_06073_));
 b15nano23al1n24x5 _17955_ (.a(\u0.tmp_w[29] ),
    .b(\u0.tmp_w[31] ),
    .c(net408),
    .d(\u0.tmp_w[28] ),
    .out0(_06084_));
 b15aoi022al1n06x5 _17956_ (.a(net430),
    .b(_06084_),
    .c(_02960_),
    .d(net423),
    .o1(_06095_));
 b15zdnd11an1n32x5 FILLER_0_2093 ();
 b15oai012ah1n08x5 _17958_ (.a(_06073_),
    .b(_06095_),
    .c(net425),
    .o1(_06117_));
 b15nor002an1n06x5 _17959_ (.a(_03806_),
    .b(_03367_),
    .o1(_06128_));
 b15nand02an1n04x5 _17960_ (.a(_06128_),
    .b(_05783_),
    .o1(_06139_));
 b15orn002ar1n24x5 _17961_ (.a(net407),
    .b(net421),
    .o(_06150_));
 b15nanb02as1n08x5 _17962_ (.a(net414),
    .b(net404),
    .out0(_06161_));
 b15nand02ah1n06x5 _17963_ (.a(net410),
    .b(net424),
    .o1(_06172_));
 b15nanb02as1n24x5 _17964_ (.a(net404),
    .b(net414),
    .out0(_06183_));
 b15oai022al1n16x5 _17965_ (.a(_06150_),
    .b(_06161_),
    .c(_06172_),
    .d(_06183_),
    .o1(_06194_));
 b15norp02al1n12x5 _17966_ (.a(_03202_),
    .b(_02949_),
    .o1(_06205_));
 b15oai112al1n08x5 _17967_ (.a(net412),
    .b(_06194_),
    .c(_06205_),
    .d(net431),
    .o1(_06216_));
 b15aoi022ah1n04x5 _17968_ (.a(net424),
    .b(_05351_),
    .c(_03432_),
    .d(_05842_),
    .o1(_06227_));
 b15nand04as1n12x5 _17969_ (.a(net420),
    .b(_06139_),
    .c(_06216_),
    .d(_06227_),
    .o1(_06238_));
 b15nandp2ar1n03x5 _17970_ (.a(net432),
    .b(_06205_),
    .o1(_06249_));
 b15nor002as1n08x5 _17971_ (.a(_03356_),
    .b(_03817_),
    .o1(_06260_));
 b15oai112as1n06x5 _17972_ (.a(_02784_),
    .b(_05699_),
    .c(_06260_),
    .d(net426),
    .o1(_06271_));
 b15aoi022ah1n08x5 _17973_ (.a(_04585_),
    .b(_03564_),
    .c(_06249_),
    .d(_06271_),
    .o1(_06282_));
 b15norp03an1n08x5 _17974_ (.a(net411),
    .b(net407),
    .c(net426),
    .o1(_06293_));
 b15zdnd11an1n64x5 FILLER_0_2029 ();
 b15oai012aq1n03x5 _17976_ (.a(net407),
    .b(net426),
    .c(net411),
    .o1(_06315_));
 b15nona23as1n08x5 _17977_ (.a(_06293_),
    .b(_06183_),
    .c(_06315_),
    .d(_05853_),
    .out0(_06326_));
 b15oaoi13an1n04x5 _17978_ (.a(net422),
    .b(_06326_),
    .c(_05853_),
    .d(_04311_),
    .o1(_06337_));
 b15oai013ar1n12x5 _17979_ (.a(_06117_),
    .b(_06238_),
    .c(_06282_),
    .d(_06337_),
    .o1(_06348_));
 b15nand02ar1n02x5 _17980_ (.a(_04859_),
    .b(_05897_),
    .o1(_06359_));
 b15nor003aq1n03x5 _17981_ (.a(\u0.tmp_w[28] ),
    .b(net430),
    .c(net423),
    .o1(_06370_));
 b15nanb02an1n12x5 _17982_ (.a(net413),
    .b(net406),
    .out0(_06381_));
 b15oai012ar1n02x5 _17983_ (.a(_06359_),
    .b(_06370_),
    .c(_06381_),
    .o1(_06392_));
 b15zdnd11an1n64x5 FILLER_0_1965 ();
 b15xor002ah1n03x5 _17985_ (.a(net430),
    .b(net423),
    .out0(_06414_));
 b15nand02ar1n02x5 _17986_ (.a(\u0.tmp_w[28] ),
    .b(_06414_),
    .o1(_06425_));
 b15and002aq1n12x5 _17987_ (.a(net407),
    .b(net427),
    .o(_06436_));
 b15aoi013ar1n02x5 _17988_ (.a(_02696_),
    .b(_06392_),
    .c(_06425_),
    .d(_06436_),
    .o1(_06447_));
 b15nor002ah1n02x5 _17989_ (.a(net422),
    .b(_02839_),
    .o1(_06458_));
 b15oai012ar1n02x5 _17990_ (.a(_04058_),
    .b(_05625_),
    .c(_02784_),
    .o1(_06469_));
 b15aoi022an1n02x5 _17991_ (.a(_06458_),
    .b(_05783_),
    .c(_06469_),
    .d(_05842_),
    .o1(_06480_));
 b15nand02an1n24x5 _17992_ (.a(_03454_),
    .b(_03553_),
    .o1(_06491_));
 b15nandp2an1n03x5 _17993_ (.a(net422),
    .b(_05472_),
    .o1(_06502_));
 b15oab012ar1n03x5 _17994_ (.a(_03378_),
    .b(_06491_),
    .c(_06502_),
    .out0(_06513_));
 b15oaoi13aq1n03x5 _17995_ (.a(_02784_),
    .b(_04146_),
    .c(_05699_),
    .d(_03828_),
    .o1(_06524_));
 b15oai012ah1n06x5 _17996_ (.a(_06480_),
    .b(_06513_),
    .c(_06524_),
    .o1(_06535_));
 b15oabi12an1n03x5 _17997_ (.a(_06447_),
    .b(_06535_),
    .c(net419),
    .out0(_06546_));
 b15nanb03al1n08x5 _17998_ (.a(_06029_),
    .b(_06348_),
    .c(_06546_),
    .out0(_06557_));
 b15xnr002ah1n03x5 _17999_ (.a(\u0.w[0][1] ),
    .b(_06557_),
    .out0(_06568_));
 b15xor002an1n04x5 _18000_ (.a(\u0.w[1][1] ),
    .b(_06568_),
    .out0(_06579_));
 b15xor002as1n02x5 _18001_ (.a(\u0.w[2][1] ),
    .b(_06579_),
    .out0(_06590_));
 b15xor002ar1n02x5 _18002_ (.a(\u0.tmp_w[1] ),
    .b(_06590_),
    .out0(_06601_));
 b15zdnd11an1n64x5 FILLER_0_1901 ();
 b15oai012ar1n02x5 _18004_ (.a(_05165_),
    .b(_06601_),
    .c(net944),
    .o1(_00364_));
 b15nand02ar1n02x5 _18005_ (.a(net944),
    .b(net51),
    .o1(_06633_));
 b15zdnd11an1n64x5 FILLER_0_1837 ();
 b15zdnd11an1n64x5 FILLER_0_1773 ();
 b15zdnd11an1n64x5 FILLER_0_1709 ();
 b15zdnd11an1n64x5 FILLER_0_1645 ();
 b15nano22ar1n02x5 _18010_ (.a(net432),
    .b(net419),
    .c(net405),
    .out0(_06688_));
 b15oai112ar1n02x5 _18011_ (.a(net412),
    .b(_03213_),
    .c(_04453_),
    .d(_06688_),
    .o1(_06699_));
 b15oaoi13an1n03x5 _18012_ (.a(_03026_),
    .b(_06699_),
    .c(_06491_),
    .d(net419),
    .o1(_06710_));
 b15aoi013al1n03x5 _18013_ (.a(_04168_),
    .b(_06084_),
    .c(net430),
    .d(_03026_),
    .o1(_06721_));
 b15aoi022an1n06x5 _18014_ (.a(_02696_),
    .b(_02619_),
    .c(_03674_),
    .d(_06062_),
    .o1(_06732_));
 b15oai012ar1n12x5 _18015_ (.a(_06721_),
    .b(_06732_),
    .c(_05231_),
    .o1(_06743_));
 b15nano23an1n03x5 _18016_ (.a(net407),
    .b(net426),
    .c(net429),
    .d(net411),
    .out0(_06754_));
 b15nor003aq1n06x5 _18017_ (.a(net414),
    .b(net404),
    .c(net417),
    .o1(_06765_));
 b15aoai13al1n08x5 _18018_ (.a(_06754_),
    .b(_06765_),
    .c(net417),
    .d(_03718_),
    .o1(_06776_));
 b15nandp2as1n12x5 _18019_ (.a(net416),
    .b(net404),
    .o1(_06787_));
 b15nand03aq1n06x5 _18020_ (.a(net413),
    .b(_03498_),
    .c(_06436_),
    .o1(_06798_));
 b15orn003ar1n04x5 _18021_ (.a(net413),
    .b(_05783_),
    .c(_05718_),
    .o(_06809_));
 b15aoai13ah1n08x5 _18022_ (.a(_06776_),
    .b(_06787_),
    .c(_06798_),
    .d(_06809_),
    .o1(_06820_));
 b15oai022ah1n06x5 _18023_ (.a(_06710_),
    .b(_06743_),
    .c(_06820_),
    .d(net422),
    .o1(_06831_));
 b15oaoi13al1n03x5 _18024_ (.a(_02784_),
    .b(_04278_),
    .c(_04826_),
    .d(\u0.tmp_w[26] ),
    .o1(_06842_));
 b15oaoi13ah1n02x5 _18025_ (.a(_04146_),
    .b(_04826_),
    .c(_04990_),
    .d(net432),
    .o1(_06853_));
 b15norp03ar1n08x5 _18026_ (.a(_02696_),
    .b(_06842_),
    .c(_06853_),
    .o1(_06864_));
 b15nanb03ar1n02x5 _18027_ (.a(net404),
    .b(net410),
    .c(net414),
    .out0(_06875_));
 b15oai022an1n02x5 _18028_ (.a(_06150_),
    .b(_06161_),
    .c(_06875_),
    .d(_02916_),
    .o1(_06886_));
 b15nano22aq1n08x5 _18029_ (.a(net429),
    .b(_06886_),
    .c(net411),
    .out0(_06897_));
 b15aoi112ar1n06x5 _18030_ (.a(_04968_),
    .b(_06897_),
    .c(_02630_),
    .d(_04760_),
    .o1(_06908_));
 b15nonb02ah1n16x5 _18031_ (.a(net424),
    .b(net431),
    .out0(_06919_));
 b15oai012ar1n02x5 _18032_ (.a(_05952_),
    .b(_05252_),
    .c(net405),
    .o1(_06930_));
 b15norp02ar1n02x5 _18033_ (.a(net424),
    .b(_03806_),
    .o1(_06941_));
 b15aoi022al1n04x5 _18034_ (.a(_06260_),
    .b(_06919_),
    .c(_06930_),
    .d(_06941_),
    .o1(_06952_));
 b15nanb02an1n04x5 _18035_ (.a(_06952_),
    .b(net426),
    .out0(_06963_));
 b15aoai13al1n08x5 _18036_ (.a(_06831_),
    .b(_06864_),
    .c(_06908_),
    .d(_06963_),
    .o1(_06974_));
 b15norp03ar1n04x5 _18037_ (.a(net428),
    .b(_02696_),
    .c(_02575_),
    .o1(_06985_));
 b15nand02al1n12x5 _18038_ (.a(net412),
    .b(net405),
    .o1(_06996_));
 b15nor003ah1n02x5 _18039_ (.a(_05395_),
    .b(_06996_),
    .c(_04497_),
    .o1(_07007_));
 b15oai012ah1n06x5 _18040_ (.a(net431),
    .b(_06985_),
    .c(_07007_),
    .o1(_07017_));
 b15nandp3ar1n08x5 _18041_ (.a(net420),
    .b(_02949_),
    .c(_03531_),
    .o1(_07028_));
 b15nonb02as1n16x5 _18042_ (.a(net418),
    .b(net421),
    .out0(_07039_));
 b15nand03ah1n03x5 _18043_ (.a(_03959_),
    .b(_07039_),
    .c(_05897_),
    .o1(_07050_));
 b15oaoi13as1n08x5 _18044_ (.a(_05592_),
    .b(_07050_),
    .c(_03180_),
    .d(_06381_),
    .o1(_07061_));
 b15nor002ah1n02x5 _18045_ (.a(net415),
    .b(_05504_),
    .o1(_07072_));
 b15and002ah1n16x5 _18046_ (.a(net431),
    .b(net428),
    .o(_07083_));
 b15nandp3ar1n02x5 _18047_ (.a(net412),
    .b(_04376_),
    .c(_07083_),
    .o1(_07094_));
 b15oai012aq1n04x5 _18048_ (.a(_07094_),
    .b(_05952_),
    .c(net412),
    .o1(_07105_));
 b15nandp3as1n04x5 _18049_ (.a(net432),
    .b(_03301_),
    .c(_04146_),
    .o1(_07116_));
 b15oai012an1n04x5 _18050_ (.a(_07116_),
    .b(_05504_),
    .c(net426),
    .o1(_07127_));
 b15aoi122ah1n04x5 _18051_ (.a(_07061_),
    .b(_07072_),
    .c(_07105_),
    .d(_07127_),
    .e(_04113_),
    .o1(_07138_));
 b15nand04al1n04x5 _18052_ (.a(net430),
    .b(_03454_),
    .c(_04629_),
    .d(_05274_),
    .o1(_07149_));
 b15zdnd11an1n04x5 FILLER_0_1637 ();
 b15nandp3al1n04x5 _18054_ (.a(_03454_),
    .b(_04629_),
    .c(_05493_),
    .o1(_07171_));
 b15nanb02al1n04x5 _18055_ (.a(_04311_),
    .b(_07039_),
    .out0(_07182_));
 b15aoai13aq1n08x5 _18056_ (.a(_07149_),
    .b(net430),
    .c(_07171_),
    .d(_07182_),
    .o1(_07193_));
 b15nonb03ah1n03x5 _18057_ (.a(net407),
    .b(net427),
    .c(net413),
    .out0(_07204_));
 b15nor002as1n08x5 _18058_ (.a(net416),
    .b(net406),
    .o1(_07215_));
 b15aoi022ah1n04x5 _18059_ (.a(_05493_),
    .b(_07215_),
    .c(_07039_),
    .d(_03718_),
    .o1(_07226_));
 b15and002ah1n12x5 _18060_ (.a(net421),
    .b(net418),
    .o(_07237_));
 b15nonb03al1n04x5 _18061_ (.a(net411),
    .b(net418),
    .c(net416),
    .out0(_07248_));
 b15aoi022aq1n08x5 _18062_ (.a(_03454_),
    .b(_07237_),
    .c(_07248_),
    .d(_02850_),
    .o1(_07259_));
 b15obai22as1n12x5 _18063_ (.a(_07204_),
    .b(_07226_),
    .c(_07259_),
    .d(_04091_),
    .out0(_07270_));
 b15aoi022al1n24x5 _18064_ (.a(net425),
    .b(_07193_),
    .c(_07270_),
    .d(net430),
    .o1(_07281_));
 b15nand04ah1n12x5 _18065_ (.a(_07017_),
    .b(_07028_),
    .c(_07138_),
    .d(_07281_),
    .o1(_07292_));
 b15nand02ar1n16x5 _18066_ (.a(_02597_),
    .b(_04694_),
    .o1(_07303_));
 b15aoi012ar1n02x5 _18067_ (.a(_07083_),
    .b(_07303_),
    .c(_02696_),
    .o1(_07314_));
 b15oai012as1n03x5 _18068_ (.a(_07237_),
    .b(_05526_),
    .c(_03092_),
    .o1(_07325_));
 b15and002an1n04x5 _18069_ (.a(_02597_),
    .b(_03674_),
    .o(_07336_));
 b15oai112ah1n06x5 _18070_ (.a(_07314_),
    .b(_07325_),
    .c(net424),
    .d(_07336_),
    .o1(_07347_));
 b15aoi012al1n02x5 _18071_ (.a(net432),
    .b(_02894_),
    .c(_04387_),
    .o1(_07358_));
 b15aoai13ar1n06x5 _18072_ (.a(_03762_),
    .b(_07358_),
    .c(_05842_),
    .d(net424),
    .o1(_07369_));
 b15nand04al1n12x5 _18073_ (.a(_03586_),
    .b(_03839_),
    .c(_04047_),
    .d(_04672_),
    .o1(_07380_));
 b15nandp3ar1n03x5 _18074_ (.a(_03454_),
    .b(_03729_),
    .c(_07237_),
    .o1(_07391_));
 b15oai112al1n06x5 _18075_ (.a(_07380_),
    .b(_07391_),
    .c(_02575_),
    .d(_03586_),
    .o1(_07402_));
 b15nandp2al1n03x5 _18076_ (.a(net415),
    .b(_02696_),
    .o1(_07413_));
 b15oai022ah1n04x5 _18077_ (.a(net415),
    .b(_05504_),
    .c(_07413_),
    .d(_06919_),
    .o1(_07424_));
 b15aoi013al1n06x5 _18078_ (.a(_07402_),
    .b(_07424_),
    .c(_05897_),
    .d(_03729_),
    .o1(_07435_));
 b15aoi012ar1n02x5 _18079_ (.a(net422),
    .b(_02696_),
    .c(_05853_),
    .o1(_07446_));
 b15nand03an1n04x5 _18080_ (.a(_02696_),
    .b(_03443_),
    .c(_04629_),
    .o1(_07457_));
 b15oaoi13aq1n03x5 _18081_ (.a(_07446_),
    .b(_07457_),
    .c(_03432_),
    .d(_04607_),
    .o1(_07468_));
 b15nandp2ah1n05x5 _18082_ (.a(_03443_),
    .b(_04629_),
    .o1(_07479_));
 b15oai022an1n04x5 _18083_ (.a(_07479_),
    .b(_05504_),
    .c(_04497_),
    .d(_04990_),
    .o1(_07490_));
 b15aoi012ah1n06x5 _18084_ (.a(_07468_),
    .b(_07490_),
    .c(_02784_),
    .o1(_07500_));
 b15nand04ah1n12x5 _18085_ (.a(_07347_),
    .b(_07369_),
    .c(_07435_),
    .d(_07500_),
    .o1(_07511_));
 b15oai012ar1n02x5 _18086_ (.a(_02960_),
    .b(_03334_),
    .c(_02784_),
    .o1(_07522_));
 b15oaoi13ar1n02x5 _18087_ (.a(net424),
    .b(_07522_),
    .c(_06491_),
    .d(net420),
    .o1(_07533_));
 b15aoi012al1n06x5 _18088_ (.a(_02960_),
    .b(_04014_),
    .c(_04025_),
    .o1(_07544_));
 b15oai022an1n04x5 _18089_ (.a(_03564_),
    .b(_07083_),
    .c(_07544_),
    .d(_04168_),
    .o1(_07555_));
 b15aoi012ar1n02x5 _18090_ (.a(_07533_),
    .b(_07555_),
    .c(net420),
    .o1(_07566_));
 b15aoi012al1n04x5 _18091_ (.a(_07566_),
    .b(_06205_),
    .c(_02784_),
    .o1(_07577_));
 b15nor004as1n12x5 _18092_ (.a(_06974_),
    .b(_07292_),
    .c(_07511_),
    .d(_07577_),
    .o1(_07588_));
 b15xor002an1n16x5 _18093_ (.a(\u0.w[0][2] ),
    .b(_07588_),
    .out0(_07599_));
 b15xor002as1n16x5 _18094_ (.a(\u0.w[1][2] ),
    .b(_07599_),
    .out0(_07610_));
 b15xor002as1n16x5 _18095_ (.a(\u0.w[2][2] ),
    .b(_07610_),
    .out0(_07621_));
 b15xor002an1n16x5 _18096_ (.a(net512),
    .b(_07621_),
    .out0(_07632_));
 b15oai012ar1n02x5 _18097_ (.a(_06633_),
    .b(_07632_),
    .c(net944),
    .o1(_00375_));
 b15nand02ar1n02x5 _18098_ (.a(net947),
    .b(net62),
    .o1(_07653_));
 b15zdnd11an1n04x5 FILLER_0_1629 ();
 b15zdnd11an1n16x5 FILLER_0_1608 ();
 b15zdnd11an1n04x5 FILLER_0_1600 ();
 b15nandp2ah1n03x5 _18102_ (.a(_07039_),
    .b(_05428_),
    .o1(_07697_));
 b15nonb03aq1n02x5 _18103_ (.a(net407),
    .b(net426),
    .c(net416),
    .out0(_07708_));
 b15inv020ar1n32x5 _18104_ (.a(net407),
    .o1(_07719_));
 b15aoi013al1n06x5 _18105_ (.a(_07708_),
    .b(_04804_),
    .c(_07719_),
    .d(net416),
    .o1(_07730_));
 b15aoi012ar1n06x5 _18106_ (.a(_06436_),
    .b(_03432_),
    .c(_07719_),
    .o1(_07741_));
 b15nandp3al1n08x5 _18107_ (.a(net418),
    .b(_03443_),
    .c(_04947_),
    .o1(_07752_));
 b15oai022an1n16x5 _18108_ (.a(_07697_),
    .b(_07730_),
    .c(_07741_),
    .d(_07752_),
    .o1(_07763_));
 b15nand03ar1n06x5 _18109_ (.a(_02597_),
    .b(_02619_),
    .c(_03850_),
    .o1(_07774_));
 b15nor002an1n06x5 _18110_ (.a(net406),
    .b(net418),
    .o1(_07785_));
 b15and003ar1n02x5 _18111_ (.a(net411),
    .b(net404),
    .c(net417),
    .o(_07796_));
 b15aoi022al1n02x5 _18112_ (.a(_07785_),
    .b(_06293_),
    .c(_06436_),
    .d(_07796_),
    .o1(_07807_));
 b15inv000ar1n24x5 _18113_ (.a(net416),
    .o1(_07818_));
 b15oaoi13al1n03x5 _18114_ (.a(net429),
    .b(_07774_),
    .c(_07807_),
    .d(_07818_),
    .o1(_07829_));
 b15nand02ar1n02x5 _18115_ (.a(net427),
    .b(_05351_),
    .o1(_07840_));
 b15nand02aq1n06x5 _18116_ (.a(net411),
    .b(net407),
    .o1(_07851_));
 b15nanb02aq1n24x5 _18117_ (.a(net426),
    .b(net429),
    .out0(_07862_));
 b15aoi022ar1n02x5 _18118_ (.a(_07862_),
    .b(_03718_),
    .c(_07215_),
    .d(_05472_),
    .o1(_07873_));
 b15oai012as1n04x5 _18119_ (.a(_07840_),
    .b(_07851_),
    .c(_07873_),
    .o1(_07884_));
 b15aoi112as1n04x5 _18120_ (.a(_07763_),
    .b(_07829_),
    .c(_07884_),
    .d(_05274_),
    .o1(_07894_));
 b15aoi022ar1n04x5 _18121_ (.a(_04168_),
    .b(_06084_),
    .c(_02960_),
    .d(_06919_),
    .o1(_07905_));
 b15norp02al1n04x5 _18122_ (.a(net418),
    .b(_07905_),
    .o1(_07916_));
 b15nand02ar1n02x5 _18123_ (.a(net411),
    .b(_05493_),
    .o1(_07927_));
 b15nanb02al1n04x5 _18124_ (.a(net411),
    .b(net418),
    .out0(_07938_));
 b15aoi112an1n03x5 _18125_ (.a(_06787_),
    .b(_05252_),
    .c(_07927_),
    .d(_07938_),
    .o1(_07949_));
 b15nandp3ah1n08x5 _18126_ (.a(_03454_),
    .b(_03553_),
    .c(_07237_),
    .o1(_07960_));
 b15and002as1n04x5 _18127_ (.a(\u0.tmp_w[29] ),
    .b(net423),
    .o(_07971_));
 b15aoi022ar1n04x5 _18128_ (.a(net406),
    .b(_07971_),
    .c(_05296_),
    .d(_07039_),
    .o1(_07982_));
 b15nand02an1n02x5 _18129_ (.a(net432),
    .b(_03213_),
    .o1(_07993_));
 b15oai112al1n08x5 _18130_ (.a(net427),
    .b(_07960_),
    .c(_07982_),
    .d(_07993_),
    .o1(_08004_));
 b15norp03aq1n12x5 _18131_ (.a(_07916_),
    .b(_07949_),
    .c(_08004_),
    .o1(_08015_));
 b15norp02as1n08x5 _18132_ (.a(net430),
    .b(_04278_),
    .o1(_08026_));
 b15and002as1n04x5 _18133_ (.a(net414),
    .b(net410),
    .o(_08037_));
 b15nand03aq1n02x5 _18134_ (.a(_05274_),
    .b(_05428_),
    .c(_08037_),
    .o1(_08048_));
 b15aoi022ar1n06x5 _18135_ (.a(_07237_),
    .b(_05428_),
    .c(_07785_),
    .d(net411),
    .o1(_08059_));
 b15oai013al1n06x5 _18136_ (.a(_08048_),
    .b(_08059_),
    .c(net407),
    .d(net414),
    .o1(_08070_));
 b15aoi112al1n06x5 _18137_ (.a(net426),
    .b(_08026_),
    .c(_08070_),
    .d(net429),
    .o1(_08081_));
 b15oai012ar1n16x5 _18138_ (.a(_07894_),
    .b(_08015_),
    .c(_08081_),
    .o1(_08092_));
 b15orn002al1n04x5 _18139_ (.a(net428),
    .b(net420),
    .o(_08103_));
 b15nor003aq1n02x5 _18140_ (.a(net410),
    .b(_08103_),
    .c(_06996_),
    .o1(_08114_));
 b15aoi012an1n04x5 _18141_ (.a(_08114_),
    .b(_05296_),
    .c(net420),
    .o1(_08125_));
 b15oai022ar1n02x5 _18142_ (.a(_04574_),
    .b(_04826_),
    .c(_08125_),
    .d(net415),
    .o1(_08136_));
 b15and002ar1n04x5 _18143_ (.a(_06919_),
    .b(_08136_),
    .o(_08147_));
 b15aoi112ah1n02x5 _18144_ (.a(net417),
    .b(_04387_),
    .c(_06205_),
    .d(net432),
    .o1(_08158_));
 b15nand02al1n02x5 _18145_ (.a(net432),
    .b(_03004_),
    .o1(_08169_));
 b15oai022ar1n02x5 _18146_ (.a(_05699_),
    .b(_07303_),
    .c(_08169_),
    .d(_05504_),
    .o1(_08180_));
 b15nanb02ah1n08x5 _18147_ (.a(net429),
    .b(net407),
    .out0(_08191_));
 b15oai022ar1n02x5 _18148_ (.a(net412),
    .b(_03367_),
    .c(_06996_),
    .d(_08191_),
    .o1(_08202_));
 b15aob012ar1n02x5 _18149_ (.a(_08169_),
    .b(_08202_),
    .c(net415),
    .out0(_08213_));
 b15aoi112an1n03x5 _18150_ (.a(_08158_),
    .b(_08180_),
    .c(_08213_),
    .d(_03850_),
    .o1(_08224_));
 b15nand04ar1n02x5 _18151_ (.a(net432),
    .b(_03454_),
    .c(_03553_),
    .d(_05493_),
    .o1(_08235_));
 b15oaoi13al1n02x5 _18152_ (.a(_03026_),
    .b(_08235_),
    .c(_05504_),
    .d(_04585_),
    .o1(_08246_));
 b15nanb02al1n04x5 _18153_ (.a(net407),
    .b(net414),
    .out0(_08256_));
 b15oai022aq1n08x5 _18154_ (.a(_07862_),
    .b(_05395_),
    .c(_08256_),
    .d(_04804_),
    .o1(_08267_));
 b15aoi013ah1n02x5 _18155_ (.a(_08246_),
    .b(_08267_),
    .c(_07039_),
    .d(_05296_),
    .o1(_08278_));
 b15nandp3ar1n02x5 _18156_ (.a(net422),
    .b(_02597_),
    .c(_03498_),
    .o1(_08289_));
 b15oaoi13an1n02x5 _18157_ (.a(_03806_),
    .b(_08289_),
    .c(_02696_),
    .d(_04091_),
    .o1(_08300_));
 b15aoai13an1n02x5 _18158_ (.a(_02784_),
    .b(_03334_),
    .c(_07039_),
    .d(net426),
    .o1(_08311_));
 b15norp02ar1n02x5 _18159_ (.a(_03564_),
    .b(_05493_),
    .o1(_08322_));
 b15aoi013an1n03x5 _18160_ (.a(_08300_),
    .b(_08311_),
    .c(_08322_),
    .d(_07116_),
    .o1(_08333_));
 b15nonb03aq1n04x5 _18161_ (.a(net404),
    .b(net426),
    .c(net416),
    .out0(_08344_));
 b15and003aq1n04x5 _18162_ (.a(net411),
    .b(net407),
    .c(net421),
    .o(_08355_));
 b15nor003ar1n08x5 _18163_ (.a(net411),
    .b(net407),
    .c(net421),
    .o1(_08366_));
 b15oai012as1n08x5 _18164_ (.a(_08344_),
    .b(_08355_),
    .c(_08366_),
    .o1(_08377_));
 b15oaoi13aq1n02x5 _18165_ (.a(net418),
    .b(_08377_),
    .c(_04058_),
    .d(_03564_),
    .o1(_08388_));
 b15nand04ar1n02x5 _18166_ (.a(net427),
    .b(_02696_),
    .c(_03454_),
    .d(_04629_),
    .o1(_08399_));
 b15nandp2al1n08x5 _18167_ (.a(net432),
    .b(net418),
    .o1(_08410_));
 b15oaoi13as1n02x5 _18168_ (.a(net421),
    .b(_08399_),
    .c(_08410_),
    .d(_04705_),
    .o1(_08421_));
 b15aoi013an1n02x5 _18169_ (.a(_02784_),
    .b(_04168_),
    .c(_02619_),
    .d(_04453_),
    .o1(_08432_));
 b15aoi012an1n02x5 _18170_ (.a(_03740_),
    .b(_02597_),
    .c(net414),
    .o1(_08443_));
 b15oai013al1n06x5 _18171_ (.a(_08432_),
    .b(_08443_),
    .c(_03784_),
    .d(_02696_),
    .o1(_08454_));
 b15nandp3ar1n02x5 _18172_ (.a(_03454_),
    .b(_03553_),
    .c(_03850_),
    .o1(_08465_));
 b15oai112as1n02x5 _18173_ (.a(_02784_),
    .b(_08465_),
    .c(_03301_),
    .d(_04585_),
    .o1(_08476_));
 b15aoi112an1n04x5 _18174_ (.a(_08388_),
    .b(_08421_),
    .c(_08454_),
    .d(_08476_),
    .o1(_08487_));
 b15nand04al1n08x5 _18175_ (.a(_08224_),
    .b(_08278_),
    .c(_08333_),
    .d(_08487_),
    .o1(_08498_));
 b15oai022ar1n02x5 _18176_ (.a(_03180_),
    .b(_04102_),
    .c(_05647_),
    .d(net425),
    .o1(_08509_));
 b15and003an1n02x5 _18177_ (.a(net406),
    .b(_02784_),
    .c(_08509_),
    .o(_08520_));
 b15aoi022al1n02x5 _18178_ (.a(_03147_),
    .b(_07971_),
    .c(_05699_),
    .d(_02619_),
    .o1(_08531_));
 b15oai012al1n06x5 _18179_ (.a(_04936_),
    .b(_08531_),
    .c(net406),
    .o1(_08542_));
 b15nonb02an1n06x5 _18180_ (.a(net432),
    .b(net407),
    .out0(_08553_));
 b15aoai13al1n08x5 _18181_ (.a(_02696_),
    .b(_08520_),
    .c(_08542_),
    .d(_08553_),
    .o1(_08563_));
 b15nor004as1n02x5 _18182_ (.a(_04168_),
    .b(_04091_),
    .c(_04102_),
    .d(_05853_),
    .o1(_08574_));
 b15aoi112ah1n02x5 _18183_ (.a(_05252_),
    .b(_06183_),
    .c(net412),
    .d(_05625_),
    .o1(_08585_));
 b15aoi112al1n04x5 _18184_ (.a(net418),
    .b(_08574_),
    .c(_08585_),
    .d(_04146_),
    .o1(_08596_));
 b15nor003al1n03x5 _18185_ (.a(net406),
    .b(_02916_),
    .c(_04102_),
    .o1(_08607_));
 b15aoai13aq1n06x5 _18186_ (.a(_05548_),
    .b(_08607_),
    .c(_05559_),
    .d(_02619_),
    .o1(_08618_));
 b15aoi012ar1n02x5 _18187_ (.a(_02696_),
    .b(_03531_),
    .c(net421),
    .o1(_08629_));
 b15and002al1n04x5 _18188_ (.a(_08618_),
    .b(_08629_),
    .o(_08640_));
 b15nor002aq1n03x5 _18189_ (.a(_08191_),
    .b(_06183_),
    .o1(_08651_));
 b15orn002ar1n02x5 _18190_ (.a(_07818_),
    .b(_04804_),
    .o(_08662_));
 b15oaoi13al1n04x5 _18191_ (.a(_05952_),
    .b(_08662_),
    .c(_05853_),
    .d(net414),
    .o1(_08673_));
 b15oai112ah1n12x5 _18192_ (.a(net413),
    .b(_04168_),
    .c(_08651_),
    .d(_08673_),
    .o1(_08684_));
 b15aoai13al1n08x5 _18193_ (.a(_08563_),
    .b(_08596_),
    .c(_08640_),
    .d(_08684_),
    .o1(_08695_));
 b15nor004an1n12x5 _18194_ (.a(_08092_),
    .b(_08147_),
    .c(_08498_),
    .d(_08695_),
    .o1(_08706_));
 b15xor002an1n08x5 _18195_ (.a(\u0.w[0][3] ),
    .b(net403),
    .out0(_08717_));
 b15xor002ah1n06x5 _18196_ (.a(\u0.w[1][3] ),
    .b(_08717_),
    .out0(_08728_));
 b15xor002ah1n08x5 _18197_ (.a(\u0.w[2][3] ),
    .b(_08728_),
    .out0(_08739_));
 b15xor002ar1n02x5 _18198_ (.a(\u0.tmp_w[3] ),
    .b(_08739_),
    .out0(_08750_));
 b15oai012ar1n02x5 _18199_ (.a(_07653_),
    .b(_08750_),
    .c(net947),
    .o1(_00378_));
 b15nand02ar1n02x5 _18200_ (.a(net943),
    .b(net73),
    .o1(_08771_));
 b15zdnd11an1n04x5 FILLER_0_1591 ();
 b15zdnd11an1n08x5 FILLER_0_1583 ();
 b15zdnd11an1n16x5 FILLER_0_1567 ();
 b15aoi022ah1n08x5 _18204_ (.a(_07818_),
    .b(_04025_),
    .c(_04947_),
    .d(_03454_),
    .o1(_08815_));
 b15nona23as1n02x5 _18205_ (.a(_07719_),
    .b(_08815_),
    .c(net430),
    .d(_05699_),
    .out0(_08826_));
 b15oaoi13as1n08x5 _18206_ (.a(net419),
    .b(_08826_),
    .c(_07479_),
    .d(net430),
    .o1(_08836_));
 b15oai112aq1n06x5 _18207_ (.a(net415),
    .b(_07719_),
    .c(_03202_),
    .d(_07083_),
    .o1(_08847_));
 b15aoai13as1n06x5 _18208_ (.a(net410),
    .b(_06919_),
    .c(_02949_),
    .d(net431),
    .o1(_08858_));
 b15oai012an1n02x5 _18209_ (.a(_08847_),
    .b(_08858_),
    .c(net415),
    .o1(_08869_));
 b15aoi013as1n03x5 _18210_ (.a(_08836_),
    .b(_08869_),
    .c(_02696_),
    .d(_05296_),
    .o1(_08880_));
 b15oai122ar1n12x5 _18211_ (.a(net417),
    .b(_03564_),
    .c(_04146_),
    .d(_04990_),
    .e(_05699_),
    .o1(_08891_));
 b15aoai13ah1n02x5 _18212_ (.a(_07971_),
    .b(_04661_),
    .c(net416),
    .d(_03553_),
    .o1(_08902_));
 b15nanb03ar1n02x5 _18213_ (.a(net409),
    .b(net425),
    .c(net405),
    .out0(_08913_));
 b15oai013ar1n02x5 _18214_ (.a(_08913_),
    .b(net423),
    .c(_07719_),
    .d(net405),
    .o1(_08924_));
 b15aob012as1n06x5 _18215_ (.a(_08902_),
    .b(_08924_),
    .c(_02619_),
    .out0(_08935_));
 b15nand03al1n06x5 _18216_ (.a(net412),
    .b(net404),
    .c(net407),
    .o1(_08946_));
 b15oaoi13aq1n04x5 _18217_ (.a(_03147_),
    .b(_08946_),
    .c(_06150_),
    .d(_05831_),
    .o1(_08957_));
 b15aoai13ar1n02x5 _18218_ (.a(net431),
    .b(_08957_),
    .c(_02630_),
    .d(net424),
    .o1(_08968_));
 b15oai012al1n02x5 _18219_ (.a(_02784_),
    .b(net428),
    .c(_02839_),
    .o1(_08979_));
 b15oai112ar1n04x5 _18220_ (.a(net424),
    .b(_08979_),
    .c(_06260_),
    .d(_05351_),
    .o1(_08990_));
 b15nona23aq1n04x5 _18221_ (.a(_08891_),
    .b(_08935_),
    .c(_08968_),
    .d(_08990_),
    .out0(_09001_));
 b15and002ar1n02x5 _18222_ (.a(_02949_),
    .b(_03740_),
    .o(_09012_));
 b15norp03ar1n04x5 _18223_ (.a(net410),
    .b(_02916_),
    .c(_06787_),
    .o1(_09023_));
 b15oai112ar1n08x5 _18224_ (.a(net412),
    .b(net431),
    .c(_09012_),
    .d(_09023_),
    .o1(_09034_));
 b15xor002an1n12x5 _18225_ (.a(net428),
    .b(net424),
    .out0(_09045_));
 b15oai013ah1n06x5 _18226_ (.a(_09034_),
    .b(_09045_),
    .c(_03092_),
    .d(net431),
    .o1(_09056_));
 b15oai012ar1n08x5 _18227_ (.a(_09001_),
    .b(_09056_),
    .c(net420),
    .o1(_09067_));
 b15nor004ah1n02x5 _18228_ (.a(_03026_),
    .b(_02696_),
    .c(_03356_),
    .d(_03367_),
    .o1(_09078_));
 b15oai013as1n02x5 _18229_ (.a(net431),
    .b(net420),
    .c(_02894_),
    .d(_09045_),
    .o1(_09089_));
 b15nona23an1n12x5 _18230_ (.a(net421),
    .b(net418),
    .c(net411),
    .d(net404),
    .out0(_09099_));
 b15oai022an1n12x5 _18231_ (.a(_03092_),
    .b(_04201_),
    .c(_09099_),
    .d(_04914_),
    .o1(_09110_));
 b15oai013an1n02x5 _18232_ (.a(_02784_),
    .b(_03356_),
    .c(_03367_),
    .d(_04574_),
    .o1(_09121_));
 b15oai022an1n06x5 _18233_ (.a(_09078_),
    .b(_09089_),
    .c(_09110_),
    .d(_09121_),
    .o1(_09132_));
 b15norp02ar1n02x5 _18234_ (.a(net420),
    .b(_02575_),
    .o1(_09143_));
 b15aoai13ah1n02x5 _18235_ (.a(net424),
    .b(_09143_),
    .c(_06128_),
    .d(net420),
    .o1(_09154_));
 b15aoi022an1n04x5 _18236_ (.a(_03334_),
    .b(_04113_),
    .c(_07336_),
    .d(_02949_),
    .o1(_09165_));
 b15aoai13ah1n03x5 _18237_ (.a(_09132_),
    .b(net431),
    .c(_09154_),
    .d(_09165_),
    .o1(_09176_));
 b15nona23ah1n02x5 _18238_ (.a(net415),
    .b(net412),
    .c(net431),
    .d(net420),
    .out0(_09187_));
 b15oai013ar1n02x5 _18239_ (.a(_09187_),
    .b(_05783_),
    .c(_04102_),
    .d(net420),
    .o1(_09198_));
 b15aoi012al1n02x5 _18240_ (.a(_04168_),
    .b(_04629_),
    .c(_09198_),
    .o1(_09209_));
 b15nor003an1n02x5 _18241_ (.a(_05395_),
    .b(_06996_),
    .c(_03586_),
    .o1(_09220_));
 b15nanb02al1n24x5 _18242_ (.a(net407),
    .b(net411),
    .out0(_09231_));
 b15oai022ah1n08x5 _18243_ (.a(_08410_),
    .b(_09231_),
    .c(_05727_),
    .d(net412),
    .o1(_09242_));
 b15norp02ar1n03x5 _18244_ (.a(net426),
    .b(_06183_),
    .o1(_09253_));
 b15aoi112an1n04x5 _18245_ (.a(net424),
    .b(_09220_),
    .c(_09242_),
    .d(_09253_),
    .o1(_09264_));
 b15oai112ah1n06x5 _18246_ (.a(_07017_),
    .b(_07028_),
    .c(_09209_),
    .d(_09264_),
    .o1(_09275_));
 b15and002aq1n04x5 _18247_ (.a(net429),
    .b(net421),
    .o(_09286_));
 b15norp02ar1n02x5 _18248_ (.a(_04311_),
    .b(_09286_),
    .o1(_09297_));
 b15oai012ar1n03x5 _18249_ (.a(_03762_),
    .b(_09297_),
    .c(_06458_),
    .o1(_09308_));
 b15aoai13an1n02x5 _18250_ (.a(net422),
    .b(_04113_),
    .c(_03334_),
    .d(_02630_),
    .o1(_09319_));
 b15oai012al1n02x5 _18251_ (.a(_02784_),
    .b(net426),
    .c(_05274_),
    .o1(_09328_));
 b15aoi013an1n03x5 _18252_ (.a(_06491_),
    .b(_04047_),
    .c(_09328_),
    .d(_03301_),
    .o1(_09337_));
 b15nonb02al1n02x5 _18253_ (.a(net418),
    .b(net426),
    .out0(_09346_));
 b15nor003al1n03x5 _18254_ (.a(net411),
    .b(net407),
    .c(net429),
    .o1(_09355_));
 b15oai112as1n08x5 _18255_ (.a(_07215_),
    .b(_09346_),
    .c(_08355_),
    .d(_09355_),
    .o1(_09365_));
 b15oai112ah1n08x5 _18256_ (.a(net407),
    .b(_05897_),
    .c(_04749_),
    .d(_07818_),
    .o1(_09374_));
 b15oai012ar1n08x5 _18257_ (.a(_07039_),
    .b(net429),
    .c(net416),
    .o1(_09383_));
 b15nandp2ah1n05x5 _18258_ (.a(_02619_),
    .b(_03421_),
    .o1(_09392_));
 b15xor002ah1n03x5 _18259_ (.a(net421),
    .b(_05526_),
    .out0(_09401_));
 b15oai122as1n16x5 _18260_ (.a(_09365_),
    .b(_09374_),
    .c(_09383_),
    .d(_09392_),
    .e(_09401_),
    .o1(_09410_));
 b15nano23aq1n08x5 _18261_ (.a(_09308_),
    .b(_09319_),
    .c(_09337_),
    .d(_09410_),
    .out0(_09419_));
 b15aoai13aq1n03x5 _18262_ (.a(net425),
    .b(_06370_),
    .c(_06414_),
    .d(\u0.tmp_w[28] ),
    .o1(_09428_));
 b15oai012ar1n12x5 _18263_ (.a(_09428_),
    .b(_04859_),
    .c(\u0.tmp_w[28] ),
    .o1(_09434_));
 b15aoi013as1n08x5 _18264_ (.a(_04552_),
    .b(_05428_),
    .c(_05919_),
    .d(_09434_),
    .o1(_09435_));
 b15nona23ar1n24x5 _18265_ (.a(_09176_),
    .b(_09275_),
    .c(_09419_),
    .d(_09435_),
    .out0(_09436_));
 b15aoi022al1n04x5 _18266_ (.a(_03531_),
    .b(_05274_),
    .c(_06919_),
    .d(_03839_),
    .o1(_09437_));
 b15aoi013an1n08x5 _18267_ (.a(_06765_),
    .b(_03718_),
    .c(net417),
    .d(net429),
    .o1(_09438_));
 b15oaoi13as1n08x5 _18268_ (.a(net426),
    .b(_09437_),
    .c(_09438_),
    .d(_09231_),
    .o1(_09439_));
 b15nano23as1n24x5 _18269_ (.a(_08880_),
    .b(_09067_),
    .c(_09436_),
    .d(_09439_),
    .out0(_09440_));
 b15xor002as1n16x5 _18270_ (.a(\u0.w[0][4] ),
    .b(_09440_),
    .out0(_09441_));
 b15xor002an1n16x5 _18271_ (.a(\u0.w[1][4] ),
    .b(_09441_),
    .out0(_09442_));
 b15xor002as1n16x5 _18272_ (.a(\u0.w[2][4] ),
    .b(_09442_),
    .out0(_09443_));
 b15xor002ar1n02x5 _18273_ (.a(\u0.tmp_w[4] ),
    .b(_09443_),
    .out0(_09444_));
 b15oai012ar1n02x5 _18274_ (.a(_08771_),
    .b(_09444_),
    .c(net943),
    .o1(_00379_));
 b15inv040ah1n02x5 _18275_ (.a(net84),
    .o1(_09445_));
 b15zdnd00an1n01x5 FILLER_0_1562 ();
 b15zdnd00an1n02x5 FILLER_0_1560 ();
 b15zdnd11an1n04x5 FILLER_0_1556 ();
 b15nand04ar1n02x5 _18279_ (.a(net428),
    .b(net424),
    .c(_04376_),
    .d(_04694_),
    .o1(_09469_));
 b15nonb03al1n04x5 _18280_ (.a(net404),
    .b(net410),
    .c(net431),
    .out0(_09475_));
 b15oaoi13ar1n02x5 _18281_ (.a(_09475_),
    .b(net424),
    .c(_04376_),
    .d(_02597_),
    .o1(_09482_));
 b15oai013al1n02x5 _18282_ (.a(_09469_),
    .b(_09482_),
    .c(_03806_),
    .d(net428),
    .o1(_09489_));
 b15oai112ar1n02x5 _18283_ (.a(net412),
    .b(_02597_),
    .c(_07083_),
    .d(_04892_),
    .o1(_09495_));
 b15oai012ar1n02x5 _18284_ (.a(_09495_),
    .b(_08858_),
    .c(_05831_),
    .o1(_09502_));
 b15nand02ah1n04x5 _18285_ (.a(_03443_),
    .b(_04859_),
    .o1(_09508_));
 b15nor002an1n03x5 _18286_ (.a(_04168_),
    .b(_05783_),
    .o1(_09515_));
 b15oai022ar1n08x5 _18287_ (.a(net426),
    .b(_09508_),
    .c(_09515_),
    .d(_03806_),
    .o1(_09521_));
 b15aoi122an1n02x5 _18288_ (.a(_09489_),
    .b(_09502_),
    .c(net415),
    .d(_03553_),
    .e(_09521_),
    .o1(_09527_));
 b15orn002aq1n03x5 _18289_ (.a(net420),
    .b(_09527_),
    .o(_09534_));
 b15nonb02al1n12x5 _18290_ (.a(net431),
    .b(net417),
    .out0(_09540_));
 b15norp02ah1n02x5 _18291_ (.a(net411),
    .b(_05718_),
    .o1(_09547_));
 b15mdn022as1n03x5 _18292_ (.a(_06183_),
    .b(_06161_),
    .o1(_09553_),
    .sa(_04804_));
 b15aoi022ah1n06x5 _18293_ (.a(_05842_),
    .b(_09540_),
    .c(_09547_),
    .d(_09553_),
    .o1(_09559_));
 b15norp03ar1n02x5 _18294_ (.a(net407),
    .b(net429),
    .c(net417),
    .o1(_09566_));
 b15aoi022ar1n02x5 _18295_ (.a(_04694_),
    .b(_04442_),
    .c(_09566_),
    .d(_02619_),
    .o1(_09573_));
 b15orn003ah1n02x5 _18296_ (.a(net404),
    .b(_05783_),
    .c(_09573_),
    .o(_09579_));
 b15oai013al1n04x5 _18297_ (.a(_04168_),
    .b(_03806_),
    .c(_03817_),
    .d(_04574_),
    .o1(_09586_));
 b15nanb03ar1n02x5 _18298_ (.a(net411),
    .b(net404),
    .c(net417),
    .out0(_09592_));
 b15aob012ar1n02x5 _18299_ (.a(_09592_),
    .b(_05897_),
    .c(_03334_),
    .out0(_09598_));
 b15qgbao4an1n05x5 _18300_ (.o1(_09605_),
    .a(_09586_),
    .b(_09598_),
    .c(_08037_),
    .d(net429));
 b15aoi022ah1n12x5 _18301_ (.a(net421),
    .b(_09559_),
    .c(_09579_),
    .d(_09605_),
    .o1(_09611_));
 b15nand02al1n06x5 _18302_ (.a(net417),
    .b(_03378_),
    .o1(_09617_));
 b15ao0022ar1n02x5 _18303_ (.a(_04629_),
    .b(_05274_),
    .c(_04442_),
    .d(net404),
    .o(_09623_));
 b15aoi022an1n06x5 _18304_ (.a(_05274_),
    .b(_05842_),
    .c(_09623_),
    .d(_04694_),
    .o1(_09630_));
 b15oaoi13as1n04x5 _18305_ (.a(net432),
    .b(_09617_),
    .c(_09630_),
    .d(_04760_),
    .o1(_09637_));
 b15nand03al1n12x5 _18306_ (.a(net411),
    .b(net404),
    .c(net428),
    .o1(_09644_));
 b15aoi012an1n06x5 _18307_ (.a(_05395_),
    .b(_05831_),
    .c(_09644_),
    .o1(_09650_));
 b15aoi012ar1n02x5 _18308_ (.a(_03531_),
    .b(_09650_),
    .c(net420),
    .o1(_09655_));
 b15oai012ar1n02x5 _18309_ (.a(_05699_),
    .b(_09650_),
    .c(_05504_),
    .o1(_09656_));
 b15aoi012an1n02x5 _18310_ (.a(_09655_),
    .b(_09656_),
    .c(net431),
    .o1(_09657_));
 b15oai112al1n02x5 _18311_ (.a(net424),
    .b(_08103_),
    .c(_09650_),
    .d(_02696_),
    .o1(_09658_));
 b15oai112as1n04x5 _18312_ (.a(_02784_),
    .b(_09658_),
    .c(_02575_),
    .d(net424),
    .o1(_09659_));
 b15aoi112ah1n04x5 _18313_ (.a(_09611_),
    .b(_09637_),
    .c(_09657_),
    .d(_09659_),
    .o1(_09660_));
 b15norp02ar1n02x5 _18314_ (.a(_03092_),
    .b(_05493_),
    .o1(_09661_));
 b15oai022ar1n02x5 _18315_ (.a(_04091_),
    .b(_03784_),
    .c(_06381_),
    .d(_06150_),
    .o1(_09662_));
 b15and003as1n04x5 _18316_ (.a(\u0.tmp_w[28] ),
    .b(net418),
    .c(_09662_),
    .o(_09663_));
 b15aoai13ar1n03x5 _18317_ (.a(net432),
    .b(_09661_),
    .c(_09663_),
    .d(_03026_),
    .o1(_09664_));
 b15nand02an1n03x5 _18318_ (.a(net418),
    .b(_06084_),
    .o1(_09665_));
 b15oai013an1n04x5 _18319_ (.a(_09665_),
    .b(_04179_),
    .c(_04585_),
    .d(net418),
    .o1(_09666_));
 b15oai012ar1n02x5 _18320_ (.a(_04267_),
    .b(_07083_),
    .c(net422),
    .o1(_09667_));
 b15oai012as1n03x5 _18321_ (.a(_09667_),
    .b(_07479_),
    .c(net422),
    .o1(_09668_));
 b15aoi222ah1n06x5 _18322_ (.a(net427),
    .b(_09666_),
    .c(_09668_),
    .d(net418),
    .e(_09663_),
    .f(_05783_),
    .o1(_09669_));
 b15oai022ar1n02x5 _18323_ (.a(net432),
    .b(_03202_),
    .c(_07862_),
    .d(_03839_),
    .o1(_09670_));
 b15oai022ar1n02x5 _18324_ (.a(net412),
    .b(_03367_),
    .c(_08946_),
    .d(_02949_),
    .o1(_09671_));
 b15nona22an1n02x5 _18325_ (.a(_07413_),
    .b(_09670_),
    .c(_09671_),
    .out0(_09672_));
 b15nor003ar1n02x5 _18326_ (.a(net414),
    .b(_05952_),
    .c(_05526_),
    .o1(_09673_));
 b15nand02al1n02x5 _18327_ (.a(net407),
    .b(_07862_),
    .o1(_09674_));
 b15oab012as1n03x5 _18328_ (.a(_09673_),
    .b(_09674_),
    .c(_06183_),
    .out0(_09675_));
 b15oai013aq1n08x5 _18329_ (.a(_09672_),
    .b(_09675_),
    .c(_05504_),
    .d(net412),
    .o1(_09676_));
 b15and002as1n04x5 _18330_ (.a(_05831_),
    .b(_09644_),
    .o(_09677_));
 b15nandp3ar1n03x5 _18331_ (.a(_03213_),
    .b(_05493_),
    .c(_04749_),
    .o1(_09678_));
 b15aoi012ah1n02x5 _18332_ (.a(_08366_),
    .b(_03959_),
    .c(net411),
    .o1(_09679_));
 b15oab012al1n02x5 _18333_ (.a(net418),
    .b(net427),
    .c(net429),
    .out0(_09680_));
 b15nandp2an1n02x5 _18334_ (.a(_07215_),
    .b(_09680_),
    .o1(_09681_));
 b15oai022ah1n06x5 _18335_ (.a(_09677_),
    .b(_09678_),
    .c(_09679_),
    .d(_09681_),
    .o1(_09682_));
 b15nor002aq1n03x5 _18336_ (.a(_03026_),
    .b(_06414_),
    .o1(_09683_));
 b15oaoi13an1n03x5 _18337_ (.a(_09683_),
    .b(_07457_),
    .c(_07303_),
    .d(_04201_),
    .o1(_09684_));
 b15nor004ar1n02x5 _18338_ (.a(_05952_),
    .b(_03432_),
    .c(_04102_),
    .d(_05504_),
    .o1(_09685_));
 b15aoi012ar1n02x5 _18339_ (.a(_05718_),
    .b(net421),
    .c(net414),
    .o1(_09686_));
 b15aoi013al1n02x5 _18340_ (.a(_09685_),
    .b(_09686_),
    .c(_07862_),
    .d(_05296_),
    .o1(_09687_));
 b15nand03ar1n03x5 _18341_ (.a(_06084_),
    .b(_05274_),
    .c(_04749_),
    .o1(_09688_));
 b15nona23ah1n04x5 _18342_ (.a(_09682_),
    .b(_09684_),
    .c(_09687_),
    .d(_09688_),
    .out0(_09689_));
 b15nano23as1n08x5 _18343_ (.a(_09664_),
    .b(_09669_),
    .c(_09676_),
    .d(_09689_),
    .out0(_09690_));
 b15and003aq1n24x5 _18344_ (.a(_09534_),
    .b(_09660_),
    .c(_09690_),
    .o(_09691_));
 b15xor002as1n16x5 _18345_ (.a(\u0.w[0][5] ),
    .b(_09691_),
    .out0(_09692_));
 b15xor002aq1n12x5 _18346_ (.a(\u0.w[1][5] ),
    .b(_09692_),
    .out0(_09693_));
 b15xor002ah1n02x5 _18347_ (.a(\u0.w[2][5] ),
    .b(_09693_),
    .out0(_09694_));
 b15xor002ar1n02x5 _18348_ (.a(\u0.tmp_w[5] ),
    .b(_09694_),
    .out0(_09695_));
 b15mdn022ar1n02x5 _18349_ (.a(_09445_),
    .b(_09695_),
    .o1(_00380_),
    .sa(net937));
 b15nand02ar1n02x5 _18350_ (.a(net937),
    .b(net95),
    .o1(_09696_));
 b15zdnd11an1n04x5 FILLER_0_1548 ();
 b15zdnd00an1n01x5 FILLER_0_1541 ();
 b15zdnd00an1n02x5 FILLER_0_1539 ();
 b15zdnd11an1n04x5 FILLER_0_1535 ();
 b15aoi022ar1n02x5 _18355_ (.a(_03828_),
    .b(_04892_),
    .c(_09286_),
    .d(_02630_),
    .o1(_09701_));
 b15nand04an1n03x5 _18356_ (.a(net404),
    .b(_03454_),
    .c(_09674_),
    .d(_09515_),
    .o1(_09702_));
 b15xor002ar1n02x5 _18357_ (.a(net414),
    .b(net421),
    .out0(_09703_));
 b15aoi013an1n02x5 _18358_ (.a(_02696_),
    .b(_03729_),
    .c(_05428_),
    .d(_09703_),
    .o1(_09704_));
 b15nand03aq1n03x5 _18359_ (.a(_09701_),
    .b(_09702_),
    .c(_09704_),
    .o1(_09705_));
 b15aoi022ar1n02x5 _18360_ (.a(net421),
    .b(_03004_),
    .c(_03828_),
    .d(_04892_),
    .o1(_09706_));
 b15oai012ah1n02x5 _18361_ (.a(_02696_),
    .b(_09706_),
    .c(net426),
    .o1(_09707_));
 b15nor003ar1n02x5 _18362_ (.a(net407),
    .b(_05472_),
    .c(_06161_),
    .o1(_09708_));
 b15aoi013ar1n02x5 _18363_ (.a(net421),
    .b(_05395_),
    .c(_08256_),
    .d(_05428_),
    .o1(_09709_));
 b15oab012al1n02x5 _18364_ (.a(_09708_),
    .b(_09709_),
    .c(_04749_),
    .out0(_09710_));
 b15aoi012an1n02x5 _18365_ (.a(_09710_),
    .b(_02894_),
    .c(net421),
    .o1(_09711_));
 b15oai012aq1n08x5 _18366_ (.a(_09705_),
    .b(_09707_),
    .c(_09711_),
    .o1(_09712_));
 b15nandp3ar1n02x5 _18367_ (.a(_04376_),
    .b(_04694_),
    .c(_05493_),
    .o1(_09713_));
 b15aoi012al1n02x5 _18368_ (.a(_02784_),
    .b(_09665_),
    .c(_09713_),
    .o1(_09714_));
 b15aoi022al1n06x5 _18369_ (.a(_03378_),
    .b(_07039_),
    .c(_04618_),
    .d(_04267_),
    .o1(_09715_));
 b15nandp3an1n03x5 _18370_ (.a(net422),
    .b(net418),
    .c(_06084_),
    .o1(_09716_));
 b15nona23ar1n12x5 _18371_ (.a(_03026_),
    .b(_09714_),
    .c(_09715_),
    .d(_09716_),
    .out0(_09717_));
 b15nona23ar1n04x5 _18372_ (.a(net406),
    .b(_03125_),
    .c(_03443_),
    .d(net418),
    .out0(_09718_));
 b15nor002aq1n08x5 _18373_ (.a(_07719_),
    .b(_04168_),
    .o1(_09719_));
 b15nanb03ar1n02x5 _18374_ (.a(net422),
    .b(net407),
    .c(net406),
    .out0(_09720_));
 b15oai012al1n02x5 _18375_ (.a(_09720_),
    .b(_03180_),
    .c(net406),
    .o1(_09721_));
 b15aoi022ah1n04x5 _18376_ (.a(_07215_),
    .b(_09719_),
    .c(_09721_),
    .d(\u0.tmp_w[28] ),
    .o1(_09722_));
 b15nandp2ah1n02x5 _18377_ (.a(net413),
    .b(net418),
    .o1(_09723_));
 b15oai013al1n08x5 _18378_ (.a(_09718_),
    .b(_09722_),
    .c(_09723_),
    .d(net432),
    .o1(_09724_));
 b15oai012al1n06x5 _18379_ (.a(_03817_),
    .b(_04179_),
    .c(_03367_),
    .o1(_09725_));
 b15oai022ar1n02x5 _18380_ (.a(_04091_),
    .b(_07938_),
    .c(_09099_),
    .d(net407),
    .o1(_09726_));
 b15ao0022an1n02x5 _18381_ (.a(_07248_),
    .b(_09725_),
    .c(_09726_),
    .d(net416),
    .o(_09727_));
 b15oai013an1n08x5 _18382_ (.a(_09717_),
    .b(_09724_),
    .c(_09727_),
    .d(net427),
    .o1(_09728_));
 b15aoi012ar1n02x5 _18383_ (.a(_02784_),
    .b(_04146_),
    .c(_04497_),
    .o1(_09729_));
 b15norp02ar1n02x5 _18384_ (.a(_05625_),
    .b(_04672_),
    .o1(_09730_));
 b15oai012as1n04x5 _18385_ (.a(_03531_),
    .b(_09729_),
    .c(_09730_),
    .o1(_09731_));
 b15nor002an1n03x5 _18386_ (.a(net427),
    .b(_03092_),
    .o1(_09732_));
 b15aoi112ar1n08x5 _18387_ (.a(net430),
    .b(_09732_),
    .c(_02960_),
    .d(net427),
    .o1(_09733_));
 b15oai012ar1n08x5 _18388_ (.a(_05274_),
    .b(_02960_),
    .c(_03004_),
    .o1(_09734_));
 b15oai012ar1n16x5 _18389_ (.a(_09731_),
    .b(_09733_),
    .c(_09734_),
    .o1(_09735_));
 b15nandp3ar1n02x5 _18390_ (.a(net416),
    .b(_04047_),
    .c(_05699_),
    .o1(_09736_));
 b15oai112ah1n02x5 _18391_ (.a(_07818_),
    .b(_04859_),
    .c(_02850_),
    .d(net432),
    .o1(_09737_));
 b15nand04as1n04x5 _18392_ (.a(_04629_),
    .b(_06007_),
    .c(_09736_),
    .d(_09737_),
    .o1(_09738_));
 b15norp02ar1n02x5 _18393_ (.a(net413),
    .b(_08191_),
    .o1(_09739_));
 b15aoi013an1n02x5 _18394_ (.a(_09739_),
    .b(_04804_),
    .c(_07719_),
    .d(net413),
    .o1(_09740_));
 b15oai013an1n03x5 _18395_ (.a(_09738_),
    .b(_09740_),
    .c(_06787_),
    .d(_05406_),
    .o1(_09741_));
 b15oai022as1n02x5 _18396_ (.a(_02839_),
    .b(_02850_),
    .c(_04585_),
    .d(_04058_),
    .o1(_09742_));
 b15aoai13as1n03x5 _18397_ (.a(net432),
    .b(_04760_),
    .c(_04826_),
    .d(net427),
    .o1(_09743_));
 b15oai012ar1n08x5 _18398_ (.a(_04826_),
    .b(_06502_),
    .c(_04387_),
    .o1(_09744_));
 b15aoai13as1n08x5 _18399_ (.a(_02696_),
    .b(_09742_),
    .c(_09743_),
    .d(_09744_),
    .o1(_09745_));
 b15nand04ah1n12x5 _18400_ (.a(net418),
    .b(_03202_),
    .c(_04014_),
    .d(_04025_),
    .o1(_09746_));
 b15oa0022ar1n02x5 _18401_ (.a(_02916_),
    .b(_06787_),
    .c(_04420_),
    .d(net416),
    .o(_09747_));
 b15oai013an1n03x5 _18402_ (.a(_09746_),
    .b(_09747_),
    .c(_07851_),
    .d(_08410_),
    .o1(_09748_));
 b15aoi112as1n02x5 _18403_ (.a(_05625_),
    .b(_05718_),
    .c(_04958_),
    .d(_04925_),
    .o1(_09749_));
 b15nanb02as1n04x5 _18404_ (.a(\u0.tmp_w[28] ),
    .b(net418),
    .out0(_09750_));
 b15aoi112ar1n02x5 _18405_ (.a(_06381_),
    .b(_06150_),
    .c(_09750_),
    .d(_03147_),
    .o1(_09751_));
 b15and003ar1n02x5 _18406_ (.a(_03026_),
    .b(_02960_),
    .c(_05274_),
    .o(_09752_));
 b15oab012al1n04x5 _18407_ (.a(net432),
    .b(_09751_),
    .c(_09752_),
    .out0(_09753_));
 b15nor003aq1n06x5 _18408_ (.a(_09748_),
    .b(_09749_),
    .c(_09753_),
    .o1(_09754_));
 b15nona23al1n16x5 _18409_ (.a(_09735_),
    .b(_09741_),
    .c(_09745_),
    .d(_09754_),
    .out0(_09755_));
 b15nandp2ar1n05x5 _18410_ (.a(net418),
    .b(_04113_),
    .o1(_09756_));
 b15nor004ar1n04x5 _18411_ (.a(net432),
    .b(_02696_),
    .c(_04091_),
    .d(_04102_),
    .o1(_09757_));
 b15aoi012ar1n06x5 _18412_ (.a(_09757_),
    .b(_05493_),
    .c(_03378_),
    .o1(_09758_));
 b15oai022an1n16x5 _18413_ (.a(_04859_),
    .b(_09756_),
    .c(_09758_),
    .d(_03026_),
    .o1(_09759_));
 b15nand02ar1n02x5 _18414_ (.a(net416),
    .b(net407),
    .o1(_09760_));
 b15aoi022ar1n02x5 _18415_ (.a(net418),
    .b(_05296_),
    .c(_09680_),
    .d(_04025_),
    .o1(_09761_));
 b15oai112ah1n02x5 _18416_ (.a(net421),
    .b(_09392_),
    .c(_09760_),
    .d(_09761_),
    .o1(_09762_));
 b15oaoi13an1n02x5 _18417_ (.a(_07204_),
    .b(net413),
    .c(_03959_),
    .d(_08553_),
    .o1(_09763_));
 b15nand02an1n02x5 _18418_ (.a(net416),
    .b(_07785_),
    .o1(_09764_));
 b15aoi022ar1n02x5 _18419_ (.a(_04025_),
    .b(_03729_),
    .c(_03959_),
    .d(_05296_),
    .o1(_09765_));
 b15oai022al1n04x5 _18420_ (.a(_09763_),
    .b(_09764_),
    .c(_09750_),
    .d(_09765_),
    .o1(_09766_));
 b15oai012aq1n06x5 _18421_ (.a(_09762_),
    .b(_09766_),
    .c(net421),
    .o1(_09767_));
 b15oai112aq1n12x5 _18422_ (.a(_02696_),
    .b(_04311_),
    .c(_07303_),
    .d(net421),
    .o1(_09768_));
 b15oaoi13aq1n08x5 _18423_ (.a(_05395_),
    .b(_09644_),
    .c(_05831_),
    .d(_02916_),
    .o1(_09769_));
 b15oai112al1n08x5 _18424_ (.a(net429),
    .b(_09768_),
    .c(_09769_),
    .d(_02696_),
    .o1(_09770_));
 b15nanb03aq1n12x5 _18425_ (.a(_09759_),
    .b(_09767_),
    .c(_09770_),
    .out0(_09771_));
 b15nano23as1n24x5 _18426_ (.a(_09712_),
    .b(_09728_),
    .c(_09755_),
    .d(_09771_),
    .out0(_09772_));
 b15xor002aq1n08x5 _18427_ (.a(\u0.w[0][6] ),
    .b(_09772_),
    .out0(_09773_));
 b15xor002as1n08x5 _18428_ (.a(\u0.w[1][6] ),
    .b(_09773_),
    .out0(_09774_));
 b15xor002an1n03x5 _18429_ (.a(\u0.w[2][6] ),
    .b(_09774_),
    .out0(_09775_));
 b15xor002ar1n02x5 _18430_ (.a(\u0.tmp_w[6] ),
    .b(_09775_),
    .out0(_09776_));
 b15oai012ar1n02x5 _18431_ (.a(_09696_),
    .b(_09776_),
    .c(net937),
    .o1(_00381_));
 b15zdnd00an1n01x5 FILLER_0_1530 ();
 b15nand02ar1n02x5 _18433_ (.a(net938),
    .b(net106),
    .o1(_09778_));
 b15zdnd00an1n02x5 FILLER_0_1528 ();
 b15zdnd11an1n04x5 FILLER_0_1524 ();
 b15zdnd11an1n08x5 FILLER_0_1516 ();
 b15aoai13al1n02x5 _18437_ (.a(_08037_),
    .b(_03432_),
    .c(net411),
    .d(_05853_),
    .o1(_09782_));
 b15norp03ar1n02x5 _18438_ (.a(net414),
    .b(net410),
    .c(_04804_),
    .o1(_09783_));
 b15aoi012aq1n02x5 _18439_ (.a(_09783_),
    .b(_08037_),
    .c(_05783_),
    .o1(_09784_));
 b15oaoi13an1n04x5 _18440_ (.a(net404),
    .b(_09782_),
    .c(_09784_),
    .d(net411),
    .o1(_09785_));
 b15aoai13aq1n08x5 _18441_ (.a(_05493_),
    .b(_09785_),
    .c(net426),
    .d(_05351_),
    .o1(_09786_));
 b15nonb02ah1n04x5 _18442_ (.a(net404),
    .b(net414),
    .out0(_09787_));
 b15oab012ar1n02x5 _18443_ (.a(_06172_),
    .b(net428),
    .c(net411),
    .out0(_09788_));
 b15aoi013an1n03x5 _18444_ (.a(net431),
    .b(net417),
    .c(_09787_),
    .d(_09788_),
    .o1(_09789_));
 b15nanb02al1n02x5 _18445_ (.a(net417),
    .b(net411),
    .out0(_09790_));
 b15nand03al1n03x5 _18446_ (.a(_09787_),
    .b(_09719_),
    .c(_09790_),
    .o1(_09791_));
 b15oaoi13an1n04x5 _18447_ (.a(_09789_),
    .b(_09791_),
    .c(_06491_),
    .d(_03301_),
    .o1(_09792_));
 b15oai012al1n06x5 _18448_ (.a(net411),
    .b(_03432_),
    .c(_05783_),
    .o1(_09793_));
 b15oai012aq1n04x5 _18449_ (.a(_03586_),
    .b(_05504_),
    .c(net426),
    .o1(_09794_));
 b15nandp2ar1n02x5 _18450_ (.a(_03004_),
    .b(_09794_),
    .o1(_09795_));
 b15norp02ar1n08x5 _18451_ (.a(_05952_),
    .b(_04102_),
    .o1(_09796_));
 b15mdn022an1n02x5 _18452_ (.a(_05842_),
    .b(_09796_),
    .o1(_09797_),
    .sa(net417));
 b15oai012aq1n06x5 _18453_ (.a(_09795_),
    .b(_09797_),
    .c(_04168_),
    .o1(_09798_));
 b15aoi122an1n08x5 _18454_ (.a(_07763_),
    .b(_09792_),
    .c(_09793_),
    .d(_09798_),
    .e(net429),
    .o1(_09799_));
 b15aoai13as1n02x5 _18455_ (.a(net431),
    .b(_04267_),
    .c(_02630_),
    .d(_02949_),
    .o1(_09800_));
 b15nano22ar1n02x5 _18456_ (.a(net431),
    .b(net424),
    .c(net411),
    .out0(_09801_));
 b15oai112ar1n02x5 _18457_ (.a(_03729_),
    .b(_09787_),
    .c(_09801_),
    .d(_04892_),
    .o1(_09802_));
 b15and002an1n03x5 _18458_ (.a(_02696_),
    .b(_09802_),
    .o(_09803_));
 b15oab012ar1n02x5 _18459_ (.a(net431),
    .b(_02960_),
    .c(_04267_),
    .out0(_09804_));
 b15aoai13ah1n02x5 _18460_ (.a(net424),
    .b(_09804_),
    .c(_02960_),
    .d(_03026_),
    .o1(_09805_));
 b15nano23ar1n02x5 _18461_ (.a(net416),
    .b(net426),
    .c(net421),
    .d(net404),
    .out0(_09806_));
 b15oab012aq1n06x5 _18462_ (.a(_09231_),
    .b(_08344_),
    .c(_09806_),
    .out0(_09807_));
 b15oai013aq1n08x5 _18463_ (.a(net420),
    .b(_02839_),
    .c(_04749_),
    .d(_04168_),
    .o1(_09808_));
 b15oai012ar1n02x5 _18464_ (.a(_03356_),
    .b(_02916_),
    .c(_03806_),
    .o1(_09809_));
 b15aoi112aq1n03x5 _18465_ (.a(_09807_),
    .b(_09808_),
    .c(_09809_),
    .d(_09475_),
    .o1(_09810_));
 b15aoi022ar1n08x5 _18466_ (.a(_09800_),
    .b(_09803_),
    .c(_09805_),
    .d(_09810_),
    .o1(_09811_));
 b15nandp3ah1n02x5 _18467_ (.a(_02784_),
    .b(_03531_),
    .c(_05274_),
    .o1(_09812_));
 b15aoi012as1n02x5 _18468_ (.a(net426),
    .b(_07960_),
    .c(_09812_),
    .o1(_09813_));
 b15oai012an1n04x5 _18469_ (.a(_09790_),
    .b(_03301_),
    .c(net411),
    .o1(_09814_));
 b15aoi022ar1n02x5 _18470_ (.a(_03762_),
    .b(_09796_),
    .c(_09814_),
    .d(_03740_),
    .o1(_09815_));
 b15aoi012al1n04x5 _18471_ (.a(_04168_),
    .b(_05783_),
    .c(_07336_),
    .o1(_09816_));
 b15nor002al1n02x5 _18472_ (.a(_09815_),
    .b(_09816_),
    .o1(_09817_));
 b15mdn022ar1n02x5 _18473_ (.a(_02916_),
    .b(_05853_),
    .o1(_09818_),
    .sa(net413));
 b15aoi022al1n02x5 _18474_ (.a(_02619_),
    .b(_05625_),
    .c(_09818_),
    .d(net414),
    .o1(_09819_));
 b15nor003an1n03x5 _18475_ (.a(net417),
    .b(_03817_),
    .c(_09819_),
    .o1(_09820_));
 b15nor004an1n06x5 _18476_ (.a(_09811_),
    .b(_09813_),
    .c(_09817_),
    .d(_09820_),
    .o1(_09821_));
 b15oai112ah1n06x5 _18477_ (.a(_03454_),
    .b(_09540_),
    .c(_04376_),
    .d(_02597_),
    .o1(_09822_));
 b15aoi013aq1n03x5 _18478_ (.a(_06293_),
    .b(_07862_),
    .c(net407),
    .d(net411),
    .o1(_09823_));
 b15nandp2al1n03x5 _18479_ (.a(net417),
    .b(_09787_),
    .o1(_09824_));
 b15oaoi13aq1n04x5 _18480_ (.a(net424),
    .b(_09822_),
    .c(_09823_),
    .d(_09824_),
    .o1(_09825_));
 b15norp02ar1n02x5 _18481_ (.a(_05831_),
    .b(_05252_),
    .o1(_09826_));
 b15nand04aq1n03x5 _18482_ (.a(net415),
    .b(net428),
    .c(net424),
    .d(net420),
    .o1(_09827_));
 b15oai013ar1n08x5 _18483_ (.a(_09827_),
    .b(_09045_),
    .c(net420),
    .d(net415),
    .o1(_09828_));
 b15oai013aq1n02x5 _18484_ (.a(_04047_),
    .b(_07039_),
    .c(net432),
    .d(_05493_),
    .o1(_09829_));
 b15aoi022ar1n02x5 _18485_ (.a(_09826_),
    .b(_09828_),
    .c(_09829_),
    .d(_03839_),
    .o1(_09830_));
 b15norp02ar1n02x5 _18486_ (.a(net429),
    .b(_04574_),
    .o1(_09831_));
 b15aoi022ar1n02x5 _18487_ (.a(net413),
    .b(_03213_),
    .c(_03454_),
    .d(_04442_),
    .o1(_09832_));
 b15orn003al1n02x5 _18488_ (.a(_04420_),
    .b(_09831_),
    .c(_09832_),
    .o(_09833_));
 b15aoai13an1n03x5 _18489_ (.a(_09830_),
    .b(_09833_),
    .c(_07083_),
    .d(_09617_),
    .o1(_09834_));
 b15aoi022an1n04x5 _18490_ (.a(_08103_),
    .b(_06919_),
    .c(_09540_),
    .d(_09045_),
    .o1(_09835_));
 b15nor002ar1n02x5 _18491_ (.a(_04574_),
    .b(_06183_),
    .o1(_09836_));
 b15nanb03al1n02x5 _18492_ (.a(net424),
    .b(net410),
    .c(net412),
    .out0(_09837_));
 b15oai012ar1n06x5 _18493_ (.a(_09837_),
    .b(net410),
    .c(net412),
    .o1(_09838_));
 b15aoi222aq1n06x5 _18494_ (.a(_03334_),
    .b(_09796_),
    .c(_06128_),
    .d(_09835_),
    .e(_09836_),
    .f(_09838_),
    .o1(_09839_));
 b15oaoi13ah1n02x5 _18495_ (.a(_04113_),
    .b(_06260_),
    .c(_02850_),
    .d(_02784_),
    .o1(_09840_));
 b15oai012aq1n02x5 _18496_ (.a(_02696_),
    .b(_06260_),
    .c(_04168_),
    .o1(_09841_));
 b15aoi012ar1n02x5 _18497_ (.a(net432),
    .b(_02916_),
    .c(_06260_),
    .o1(_09842_));
 b15oai013ar1n06x5 _18498_ (.a(_09839_),
    .b(_09840_),
    .c(_09841_),
    .d(_09842_),
    .o1(_09843_));
 b15nor004aq1n06x5 _18499_ (.a(_09759_),
    .b(_09825_),
    .c(_09834_),
    .d(_09843_),
    .o1(_09844_));
 b15nand04as1n16x5 _18500_ (.a(_09786_),
    .b(_09799_),
    .c(_09821_),
    .d(_09844_),
    .o1(_09845_));
 b15xnr002aq1n12x5 _18501_ (.a(\u0.w[0][7] ),
    .b(_09845_),
    .out0(_09846_));
 b15xor002as1n12x5 _18502_ (.a(\u0.w[1][7] ),
    .b(_09846_),
    .out0(_09847_));
 b15xor002as1n03x5 _18503_ (.a(\u0.w[2][7] ),
    .b(_09847_),
    .out0(_09848_));
 b15xor002ar1n02x5 _18504_ (.a(\u0.tmp_w[7] ),
    .b(_09848_),
    .out0(_09849_));
 b15oai012ar1n02x5 _18505_ (.a(_09778_),
    .b(_09849_),
    .c(net938),
    .o1(_00382_));
 b15nand02ar1n02x5 _18506_ (.a(net947),
    .b(net117),
    .o1(_09850_));
 b15zdnd11an1n04x5 FILLER_0_1508 ();
 b15zdnd00an1n02x5 FILLER_0_1502 ();
 b15zdnd11an1n04x5 FILLER_0_1498 ();
 b15zdnd00an1n02x5 FILLER_0_1490 ();
 b15zdnd11an1n04x5 FILLER_0_1486 ();
 b15nandp2an1n32x5 _18512_ (.a(net510),
    .b(\u0.tmp_w[3] ),
    .o1(_09856_));
 b15zdnd00an1n01x5 FILLER_0_1481 ();
 b15nonb02as1n16x5 _18514_ (.a(net500),
    .b(net504),
    .out0(_09858_));
 b15norp02as1n48x5 _18515_ (.a(net496),
    .b(net492),
    .o1(_09859_));
 b15nandp2ah1n24x5 _18516_ (.a(_09858_),
    .b(_09859_),
    .o1(_09860_));
 b15oai012ar1n02x5 _18517_ (.a(net516),
    .b(_09856_),
    .c(_09860_),
    .o1(_09861_));
 b15zdnd11an1n04x5 FILLER_0_1477 ();
 b15nonb02an1n16x5 _18519_ (.a(net518),
    .b(net512),
    .out0(_09863_));
 b15zdnd11an1n04x5 FILLER_0_1469 ();
 b15zdnd11an1n08x5 FILLER_0_1461 ();
 b15zdnd11an1n04x5 FILLER_0_1453 ();
 b15and003ah1n08x5 _18523_ (.a(net500),
    .b(net496),
    .c(net492),
    .o(_09867_));
 b15nor002ah1n32x5 _18524_ (.a(net507),
    .b(net506),
    .o1(_09868_));
 b15zdnd00an1n02x5 FILLER_0_1444 ();
 b15nand02ar1n02x5 _18526_ (.a(_09867_),
    .b(_09868_),
    .o1(_09870_));
 b15nonb02an1n16x5 _18527_ (.a(net504),
    .b(net500),
    .out0(_09871_));
 b15zdnd00an1n02x5 FILLER_0_1434 ();
 b15norp02ar1n02x5 _18529_ (.a(_09871_),
    .b(_09858_),
    .o1(_09873_));
 b15zdnd00an1n01x5 FILLER_0_1429 ();
 b15zdnd11an1n08x5 FILLER_0_1421 ();
 b15nonb02as1n16x5 _18532_ (.a(net510),
    .b(net509),
    .out0(_09876_));
 b15zdnd11an1n04x5 FILLER_0_1413 ();
 b15zdnd11an1n04x5 FILLER_0_1405 ();
 b15zdnd11an1n04x5 FILLER_0_1397 ();
 b15orn002aq1n24x5 _18536_ (.a(net520),
    .b(net515),
    .o(_09880_));
 b15nand03ar1n02x5 _18537_ (.a(_09859_),
    .b(_09876_),
    .c(_09880_),
    .o1(_09881_));
 b15oai022ar1n04x5 _18538_ (.a(_09863_),
    .b(_09870_),
    .c(_09873_),
    .d(_09881_),
    .o1(_09882_));
 b15oai012as1n02x5 _18539_ (.a(_09861_),
    .b(_09882_),
    .c(net516),
    .o1(_09883_));
 b15zdnd11an1n04x5 FILLER_0_1389 ();
 b15zdnd00an1n01x5 FILLER_0_1384 ();
 b15zdnd00an1n02x5 FILLER_0_1382 ();
 b15orn002aq1n16x5 _18543_ (.a(net520),
    .b(net513),
    .o(_09887_));
 b15inv040an1n60x5 _18544_ (.a(net519),
    .o1(_09888_));
 b15zdnd11an1n04x5 FILLER_0_1378 ();
 b15zdnd11an1n04x5 FILLER_0_1370 ();
 b15oai112ar1n02x5 _18547_ (.a(net516),
    .b(_09887_),
    .c(_09856_),
    .d(_09888_),
    .o1(_09891_));
 b15inv000as1n56x5 _18548_ (.a(net513),
    .o1(_09892_));
 b15zdnd00an1n01x5 FILLER_0_1365 ();
 b15nanb02as1n24x5 _18550_ (.a(net492),
    .b(net496),
    .out0(_09894_));
 b15zdnd11an1n04x5 FILLER_0_1361 ();
 b15nand02an1n24x5 _18552_ (.a(net504),
    .b(net499),
    .o1(_09896_));
 b15norp02an1n12x5 _18553_ (.a(_09894_),
    .b(_09896_),
    .o1(_09897_));
 b15nor002as1n03x5 _18554_ (.a(_09892_),
    .b(_09897_),
    .o1(_09898_));
 b15nonb02as1n16x5 _18555_ (.a(net509),
    .b(net510),
    .out0(_09899_));
 b15oai013ar1n02x5 _18556_ (.a(_09891_),
    .b(_09898_),
    .c(_09899_),
    .d(net516),
    .o1(_09900_));
 b15inv000ah1n32x5 _18557_ (.a(\u0.tmp_w[4] ),
    .o1(_09901_));
 b15zdnd11an1n08x5 FILLER_0_1353 ();
 b15zdnd11an1n04x5 FILLER_0_1345 ();
 b15zdnd11an1n04x5 FILLER_0_1337 ();
 b15nanb02as1n24x5 _18561_ (.a(net517),
    .b(net513),
    .out0(_09905_));
 b15zdnd11an1n04x5 FILLER_0_1329 ();
 b15nano23as1n24x5 _18563_ (.a(net506),
    .b(net495),
    .c(net491),
    .d(net499),
    .out0(_09907_));
 b15nanb02as1n24x5 _18564_ (.a(net508),
    .b(net516),
    .out0(_09908_));
 b15oaoi13aq1n03x5 _18565_ (.a(net519),
    .b(_09905_),
    .c(_09907_),
    .d(_09908_),
    .o1(_09909_));
 b15nonb02as1n16x5 _18566_ (.a(net507),
    .b(net499),
    .out0(_09910_));
 b15nor004ar1n08x5 _18567_ (.a(_09901_),
    .b(_09894_),
    .c(_09909_),
    .d(_09910_),
    .o1(_09911_));
 b15aob012ar1n08x5 _18568_ (.a(_09883_),
    .b(_09900_),
    .c(_09911_),
    .out0(_09912_));
 b15zdnd00an1n02x5 FILLER_0_1323 ();
 b15nona22ah1n32x5 _18570_ (.a(net502),
    .b(net491),
    .c(net495),
    .out0(_09914_));
 b15nor002ah1n12x5 _18571_ (.a(net504),
    .b(_09914_),
    .o1(_09915_));
 b15norp02al1n24x5 _18572_ (.a(net516),
    .b(net508),
    .o1(_09916_));
 b15nand02ar1n02x5 _18573_ (.a(_09915_),
    .b(_09916_),
    .o1(_09917_));
 b15nanb02as1n24x5 _18574_ (.a(net515),
    .b(net508),
    .out0(_09918_));
 b15mdn022ar1n02x5 _18575_ (.a(_09908_),
    .b(_09918_),
    .o1(_09919_),
    .sa(net520));
 b15oaoi13as1n02x5 _18576_ (.a(net513),
    .b(_09917_),
    .c(_09919_),
    .d(_09860_),
    .o1(_09920_));
 b15norp02an1n16x5 _18577_ (.a(net518),
    .b(net512),
    .o1(_09921_));
 b15nanb02as1n24x5 _18578_ (.a(net506),
    .b(net509),
    .out0(_09922_));
 b15and003ar1n02x5 _18579_ (.a(net519),
    .b(net515),
    .c(net511),
    .o(_09923_));
 b15nor004al1n04x5 _18580_ (.a(_09921_),
    .b(_09914_),
    .c(_09922_),
    .d(_09923_),
    .o1(_09924_));
 b15nanb02as1n24x5 _18581_ (.a(net495),
    .b(net491),
    .out0(_09925_));
 b15ornc04as1n24x5 _18582_ (.a(net504),
    .b(net500),
    .c(net496),
    .d(net492),
    .o(_09926_));
 b15zdnd11an1n08x5 FILLER_0_1315 ();
 b15oai022al1n12x5 _18584_ (.a(_09896_),
    .b(_09925_),
    .c(_09926_),
    .d(net517),
    .o1(_09928_));
 b15zdnd11an1n04x5 FILLER_0_1307 ();
 b15zdnd11an1n04x5 FILLER_0_1299 ();
 b15qbfno2bn1n16x5 _18587_ (.a(net511),
    .b(net508),
    .o1(_09931_));
 b15inv000al1n80x5 _18588_ (.a(net516),
    .o1(_09932_));
 b15zdnd00an1n01x5 FILLER_0_1291 ();
 b15nandp2al1n08x5 _18590_ (.a(net519),
    .b(_09932_),
    .o1(_09934_));
 b15aoi013an1n06x5 _18591_ (.a(_09924_),
    .b(_09928_),
    .c(_09931_),
    .d(_09934_),
    .o1(_09935_));
 b15nonb02as1n16x5 _18592_ (.a(net510),
    .b(net515),
    .out0(_09936_));
 b15zdnd11an1n04x5 FILLER_0_1287 ();
 b15and002ar1n24x5 _18594_ (.a(net496),
    .b(net492),
    .o(_09938_));
 b15nanb02as1n24x5 _18595_ (.a(net518),
    .b(net514),
    .out0(_09939_));
 b15and002as1n16x5 _18596_ (.a(net514),
    .b(net512),
    .o(_09940_));
 b15oai012ar1n02x5 _18597_ (.a(_09939_),
    .b(_09940_),
    .c(_09888_),
    .o1(_09941_));
 b15aoi022al1n02x5 _18598_ (.a(_09936_),
    .b(_09938_),
    .c(_09941_),
    .d(_09859_),
    .o1(_09942_));
 b15oai013ah1n04x5 _18599_ (.a(_09935_),
    .b(_09922_),
    .c(_09942_),
    .d(net500),
    .o1(_09943_));
 b15zdnd00an1n02x5 FILLER_0_1281 ();
 b15nano23as1n24x5 _18601_ (.a(net504),
    .b(net492),
    .c(net496),
    .d(net500),
    .out0(_09945_));
 b15nanb02al1n06x5 _18602_ (.a(_09856_),
    .b(_09945_),
    .out0(_09946_));
 b15nandp3ar1n02x5 _18603_ (.a(_09863_),
    .b(_09867_),
    .c(_09868_),
    .o1(_09947_));
 b15aoi012ar1n02x5 _18604_ (.a(_09932_),
    .b(_09946_),
    .c(_09947_),
    .o1(_09948_));
 b15nonb02as1n16x5 _18605_ (.a(net507),
    .b(\u0.tmp_w[4] ),
    .out0(_09949_));
 b15zdnd11an1n04x5 FILLER_0_1277 ();
 b15nano22ah1n24x5 _18607_ (.a(net495),
    .b(net491),
    .c(net499),
    .out0(_09951_));
 b15nand03an1n06x5 _18608_ (.a(net519),
    .b(_09949_),
    .c(_09951_),
    .o1(_09952_));
 b15nandp2ah1n16x5 _18609_ (.a(_09871_),
    .b(_09859_),
    .o1(_09953_));
 b15oai012ar1n04x5 _18610_ (.a(_09952_),
    .b(_09953_),
    .c(_09908_),
    .o1(_09954_));
 b15zdnd00an1n01x5 FILLER_0_1271 ();
 b15aoi012ah1n02x5 _18612_ (.a(_09948_),
    .b(_09954_),
    .c(_09892_),
    .o1(_09956_));
 b15zdnd00an1n02x5 FILLER_0_1269 ();
 b15zdnd11an1n04x5 FILLER_0_1265 ();
 b15zdnd11an1n04x5 FILLER_0_1257 ();
 b15zdnd11an1n04x5 FILLER_0_1249 ();
 b15zdnd00an1n01x5 FILLER_0_1242 ();
 b15nano23as1n24x5 _18618_ (.a(net501),
    .b(net497),
    .c(net494),
    .d(net505),
    .out0(_09962_));
 b15oaoi13aq1n03x5 _18619_ (.a(net520),
    .b(net511),
    .c(_09962_),
    .d(_09932_),
    .o1(_09963_));
 b15nonb02as1n16x5 _18620_ (.a(net494),
    .b(net497),
    .out0(_09964_));
 b15zdnd11an1n04x5 FILLER_0_1238 ();
 b15zdnd00an1n01x5 FILLER_0_1232 ();
 b15norp02ar1n32x5 _18623_ (.a(net505),
    .b(net501),
    .o1(_09967_));
 b15aoi013an1n03x5 _18624_ (.a(_09962_),
    .b(_09964_),
    .c(_09967_),
    .d(net511),
    .o1(_09968_));
 b15nor003al1n08x5 _18625_ (.a(net508),
    .b(_09963_),
    .c(_09968_),
    .o1(_09969_));
 b15nonb03ah1n08x5 _18626_ (.a(net493),
    .b(net495),
    .c(net506),
    .out0(_09970_));
 b15zdnd00an1n02x5 FILLER_0_1230 ();
 b15zdnd11an1n08x5 FILLER_0_1222 ();
 b15zdnd11an1n04x5 FILLER_0_1214 ();
 b15nano22al1n06x5 _18630_ (.a(net506),
    .b(net498),
    .c(net493),
    .out0(_09974_));
 b15oai112aq1n08x5 _18631_ (.a(_09910_),
    .b(_09863_),
    .c(_09970_),
    .d(_09974_),
    .o1(_09975_));
 b15zdnd11an1n04x5 FILLER_0_1206 ();
 b15nonb03as1n12x5 _18633_ (.a(net498),
    .b(net493),
    .c(net502),
    .out0(_09977_));
 b15nano22ah1n24x5 _18634_ (.a(net502),
    .b(net493),
    .c(net495),
    .out0(_09978_));
 b15aoi012al1n06x5 _18635_ (.a(_09977_),
    .b(_09978_),
    .c(net512),
    .o1(_09979_));
 b15orn002al1n16x5 _18636_ (.a(net509),
    .b(net506),
    .o(_09980_));
 b15oai013as1n12x5 _18637_ (.a(_09975_),
    .b(_09979_),
    .c(_09980_),
    .d(_09880_),
    .o1(_09981_));
 b15nanb02as1n24x5 _18638_ (.a(net500),
    .b(net504),
    .out0(_09982_));
 b15nanb02as1n24x5 _18639_ (.a(net504),
    .b(net500),
    .out0(_09983_));
 b15nand04aq1n16x5 _18640_ (.a(net516),
    .b(_09982_),
    .c(_09983_),
    .d(_09859_),
    .o1(_09984_));
 b15nona23ah1n32x5 _18641_ (.a(net496),
    .b(net492),
    .c(net504),
    .d(net500),
    .out0(_09985_));
 b15oai012ah1n08x5 _18642_ (.a(_09984_),
    .b(_09985_),
    .c(_09888_),
    .o1(_09986_));
 b15aoi112ah1n06x5 _18643_ (.a(_09969_),
    .b(_09981_),
    .c(_09986_),
    .d(_09931_),
    .o1(_09987_));
 b15nona23ar1n12x5 _18644_ (.a(_09920_),
    .b(_09943_),
    .c(_09956_),
    .d(_09987_),
    .out0(_09988_));
 b15nandp3al1n04x5 _18645_ (.a(_09899_),
    .b(_09858_),
    .c(_09938_),
    .o1(_09989_));
 b15nona23as1n32x5 _18646_ (.a(net504),
    .b(net500),
    .c(net496),
    .d(net492),
    .out0(_09990_));
 b15oai012al1n02x5 _18647_ (.a(_09989_),
    .b(_09990_),
    .c(_09856_),
    .o1(_09991_));
 b15and002as1n16x5 _18648_ (.a(net505),
    .b(net501),
    .o(_09992_));
 b15nand02aq1n32x5 _18649_ (.a(_09992_),
    .b(_09964_),
    .o1(_09993_));
 b15nanb02as1n24x5 _18650_ (.a(net513),
    .b(net517),
    .out0(_09994_));
 b15zdnd00an1n01x5 FILLER_0_1200 ();
 b15nonb02as1n16x5 _18652_ (.a(net506),
    .b(net507),
    .out0(_09996_));
 b15nand02an1n12x5 _18653_ (.a(_09996_),
    .b(_09951_),
    .o1(_09997_));
 b15oai022ar1n06x5 _18654_ (.a(_09905_),
    .b(_09993_),
    .c(_09994_),
    .d(_09997_),
    .o1(_09998_));
 b15zdnd11an1n04x5 FILLER_0_1196 ();
 b15nonb03ah1n02x5 _18656_ (.a(net511),
    .b(net497),
    .c(net492),
    .out0(_10000_));
 b15oai012ar1n04x5 _18657_ (.a(_10000_),
    .b(_09996_),
    .c(_09858_),
    .o1(_10001_));
 b15nandp2aq1n04x5 _18658_ (.a(_09892_),
    .b(_09868_),
    .o1(_10002_));
 b15nanb03as1n16x5 _18659_ (.a(net502),
    .b(net498),
    .c(net493),
    .out0(_10003_));
 b15oaoi13ar1n08x5 _18660_ (.a(_09916_),
    .b(_10001_),
    .c(_10002_),
    .d(_10003_),
    .o1(_10004_));
 b15nor004as1n03x5 _18661_ (.a(net519),
    .b(_09991_),
    .c(_09998_),
    .d(_10004_),
    .o1(_10005_));
 b15orn002ah1n24x5 _18662_ (.a(net515),
    .b(net510),
    .o(_10006_));
 b15zdnd11an1n04x5 FILLER_0_1188 ();
 b15nandp3aq1n16x5 _18664_ (.a(net501),
    .b(net497),
    .c(net494),
    .o1(_10008_));
 b15nor002aq1n16x5 _18665_ (.a(_10008_),
    .b(_09922_),
    .o1(_10009_));
 b15nor002an1n16x5 _18666_ (.a(_09896_),
    .b(_09925_),
    .o1(_10010_));
 b15aoai13ah1n02x5 _18667_ (.a(_10006_),
    .b(_10009_),
    .c(_10010_),
    .d(_09876_),
    .o1(_10011_));
 b15aoi012ah1n04x5 _18668_ (.a(_10005_),
    .b(_10011_),
    .c(net519),
    .o1(_10012_));
 b15zdnd11an1n04x5 FILLER_0_1179 ();
 b15norp02ah1n24x5 _18670_ (.a(net520),
    .b(net516),
    .o1(_10014_));
 b15andc04aq1n16x5 _18671_ (.a(net505),
    .b(net500),
    .c(net497),
    .d(net492),
    .o(_10015_));
 b15aoi013ar1n02x5 _18672_ (.a(net508),
    .b(_10014_),
    .c(_10015_),
    .d(net513),
    .o1(_10016_));
 b15nand02as1n32x5 _18673_ (.a(net519),
    .b(net517),
    .o1(_10017_));
 b15aoi012ar1n02x5 _18674_ (.a(_10015_),
    .b(_09945_),
    .c(_10017_),
    .o1(_10018_));
 b15zdnd11an1n04x5 FILLER_0_1170 ();
 b15oai013al1n02x5 _18676_ (.a(_10016_),
    .b(_10018_),
    .c(_10014_),
    .d(net513),
    .o1(_10020_));
 b15zdnd11an1n04x5 FILLER_0_1162 ();
 b15nandp2an1n12x5 _18678_ (.a(_09858_),
    .b(_09964_),
    .o1(_10022_));
 b15nonb02ah1n16x5 _18679_ (.a(\u0.tmp_w[1] ),
    .b(net518),
    .out0(_10023_));
 b15nandp2ar1n08x5 _18680_ (.a(net511),
    .b(_10023_),
    .o1(_10024_));
 b15nona23aq1n32x5 _18681_ (.a(\u0.tmp_w[4] ),
    .b(net491),
    .c(net495),
    .d(net499),
    .out0(_10025_));
 b15oai122ah1n08x5 _18682_ (.a(net508),
    .b(_09934_),
    .c(_10022_),
    .d(_10024_),
    .e(_10025_),
    .o1(_10026_));
 b15nandp2ar1n05x5 _18683_ (.a(_09892_),
    .b(_09962_),
    .o1(_10027_));
 b15zdnd00an1n01x5 FILLER_0_1157 ();
 b15oaoi13aq1n03x5 _18685_ (.a(_10023_),
    .b(_10027_),
    .c(_10022_),
    .d(_09892_),
    .o1(_10029_));
 b15nanb02aq1n06x5 _18686_ (.a(net499),
    .b(net513),
    .out0(_10030_));
 b15and002ah1n04x5 _18687_ (.a(\u0.tmp_w[1] ),
    .b(net506),
    .o(_10031_));
 b15nonb02as1n16x5 _18688_ (.a(net495),
    .b(net491),
    .out0(_10032_));
 b15zdnd00an1n02x5 FILLER_0_1155 ();
 b15aoai13an1n08x5 _18690_ (.a(net518),
    .b(_09970_),
    .c(_10031_),
    .d(_10032_),
    .o1(_10034_));
 b15nandp2al1n08x5 _18691_ (.a(net514),
    .b(_09901_),
    .o1(_10035_));
 b15oaoi13ah1n03x5 _18692_ (.a(_10030_),
    .b(_10034_),
    .c(_10035_),
    .d(_09925_),
    .o1(_10036_));
 b15oai013an1n06x5 _18693_ (.a(_10020_),
    .b(_10026_),
    .c(_10029_),
    .d(_10036_),
    .o1(_10037_));
 b15inv020ah1n80x5 _18694_ (.a(net507),
    .o1(_10038_));
 b15zdnd11an1n04x5 FILLER_0_1151 ();
 b15nandp2ah1n08x5 _18696_ (.a(_09967_),
    .b(_09964_),
    .o1(_10040_));
 b15oai012ar1n06x5 _18697_ (.a(_10038_),
    .b(_09887_),
    .c(_10040_),
    .o1(_10041_));
 b15orn003aq1n04x5 _18698_ (.a(net506),
    .b(net495),
    .c(net491),
    .o(_10042_));
 b15nand02aq1n16x5 _18699_ (.a(_09932_),
    .b(net504),
    .o1(_10043_));
 b15nand02an1n48x5 _18700_ (.a(net496),
    .b(net492),
    .o1(_10044_));
 b15oai012ar1n02x5 _18701_ (.a(_10042_),
    .b(_10043_),
    .c(_10044_),
    .o1(_10045_));
 b15norp02ar1n02x5 _18702_ (.a(_10014_),
    .b(_10030_),
    .o1(_10046_));
 b15aoi012ah1n02x5 _18703_ (.a(_10041_),
    .b(_10045_),
    .c(_10046_),
    .o1(_10047_));
 b15nandp3ar1n02x5 _18704_ (.a(_09859_),
    .b(_10014_),
    .c(_10030_),
    .o1(_10048_));
 b15nano22aq1n06x5 _18705_ (.a(net495),
    .b(net491),
    .c(net519),
    .out0(_10049_));
 b15norp03an1n24x5 _18706_ (.a(net500),
    .b(net496),
    .c(net492),
    .o1(_10050_));
 b15aoai13as1n02x5 _18707_ (.a(net517),
    .b(_10049_),
    .c(_10050_),
    .d(_09863_),
    .o1(_10051_));
 b15oai112al1n04x5 _18708_ (.a(_10048_),
    .b(_10051_),
    .c(net513),
    .d(_10044_),
    .o1(_10052_));
 b15nano23an1n16x5 _18709_ (.a(net506),
    .b(net499),
    .c(net495),
    .d(net491),
    .out0(_10053_));
 b15nor002ar1n24x5 _18710_ (.a(_09982_),
    .b(_10044_),
    .o1(_10054_));
 b15ao0022ar1n02x5 _18711_ (.a(net512),
    .b(_10053_),
    .c(_10054_),
    .d(_09932_),
    .o(_10055_));
 b15zdnd11an1n04x5 FILLER_0_1143 ();
 b15aoi022as1n04x5 _18713_ (.a(net505),
    .b(_10052_),
    .c(_10055_),
    .d(net519),
    .o1(_10057_));
 b15aoai13aq1n08x5 _18714_ (.a(_10037_),
    .b(_10047_),
    .c(_10057_),
    .d(net508),
    .o1(_10058_));
 b15nor004as1n12x5 _18715_ (.a(_09912_),
    .b(_09988_),
    .c(_10012_),
    .d(_10058_),
    .o1(_10059_));
 b15xor002aq1n12x5 _18716_ (.a(\u0.w[0][8] ),
    .b(_10059_),
    .out0(_10060_));
 b15xor002ar1n16x5 _18717_ (.a(\u0.w[1][8] ),
    .b(_10060_),
    .out0(_10061_));
 b15xor002ah1n08x5 _18718_ (.a(\u0.w[2][8] ),
    .b(_10061_),
    .out0(_10062_));
 b15xor002ar1n02x5 _18719_ (.a(\u0.tmp_w[8] ),
    .b(_10062_),
    .out0(_10063_));
 b15oai012ar1n02x5 _18720_ (.a(_09850_),
    .b(_10063_),
    .c(net947),
    .o1(_00383_));
 b15inv020aq1n10x5 _18721_ (.a(net128),
    .o1(_10064_));
 b15zdnd11an1n04x5 FILLER_0_1135 ();
 b15zdnd00an1n01x5 FILLER_0_1128 ();
 b15zdnd11an1n04x5 FILLER_0_1124 ();
 b15nonb03as1n12x5 _18725_ (.a(net491),
    .b(net495),
    .c(net499),
    .out0(_10068_));
 b15nand02an1n24x5 _18726_ (.a(_09949_),
    .b(_10068_),
    .o1(_10069_));
 b15oai022ar1n02x5 _18727_ (.a(net507),
    .b(_09984_),
    .c(_10069_),
    .d(_09939_),
    .o1(_10070_));
 b15nanb02as1n24x5 _18728_ (.a(net507),
    .b(\u0.tmp_w[2] ),
    .out0(_10071_));
 b15nand03aq1n12x5 _18729_ (.a(net516),
    .b(net496),
    .c(net492),
    .o1(_10072_));
 b15orn002ar1n24x5 _18730_ (.a(net496),
    .b(net492),
    .o(_10073_));
 b15aoi112al1n08x5 _18731_ (.a(_09983_),
    .b(_10071_),
    .c(_10072_),
    .d(_10073_),
    .o1(_10074_));
 b15orn003an1n02x5 _18732_ (.a(_09915_),
    .b(_10070_),
    .c(_10074_),
    .o(_10075_));
 b15oaoi13ar1n02x5 _18733_ (.a(_09892_),
    .b(_10017_),
    .c(_10074_),
    .d(_09915_),
    .o1(_10076_));
 b15norp02ar1n02x5 _18734_ (.a(net517),
    .b(_09856_),
    .o1(_10077_));
 b15aoi013ar1n02x5 _18735_ (.a(_10077_),
    .b(_09984_),
    .c(_10038_),
    .d(_09892_),
    .o1(_10078_));
 b15oab012al1n03x5 _18736_ (.a(_10076_),
    .b(_10078_),
    .c(net519),
    .out0(_10079_));
 b15oab012ar1n02x5 _18737_ (.a(\u0.tmp_w[4] ),
    .b(_09859_),
    .c(_10049_),
    .out0(_10080_));
 b15mdn022an1n03x5 _18738_ (.a(_10073_),
    .b(_10044_),
    .o1(_10081_),
    .sa(net517));
 b15aoai13al1n04x5 _18739_ (.a(_09910_),
    .b(_10080_),
    .c(_10081_),
    .d(_09888_),
    .o1(_10082_));
 b15zdnd11an1n04x5 FILLER_0_1116 ();
 b15nona22ar1n02x5 _18741_ (.a(net506),
    .b(net491),
    .c(net499),
    .out0(_10084_));
 b15zdnd11an1n04x5 FILLER_0_1108 ();
 b15nanb02ar1n02x5 _18743_ (.a(net499),
    .b(net491),
    .out0(_10086_));
 b15nandp2ah1n12x5 _18744_ (.a(net517),
    .b(net506),
    .o1(_10087_));
 b15oaoi13aq1n02x5 _18745_ (.a(net519),
    .b(_10084_),
    .c(_10086_),
    .d(_10087_),
    .o1(_10088_));
 b15nona22aq1n04x5 _18746_ (.a(net499),
    .b(net491),
    .c(\u0.tmp_w[4] ),
    .out0(_10089_));
 b15oab012ah1n02x5 _18747_ (.a(_10088_),
    .b(_10089_),
    .c(_10017_),
    .out0(_10090_));
 b15nanb02an1n08x5 _18748_ (.a(net507),
    .b(net495),
    .out0(_10091_));
 b15oai112al1n12x5 _18749_ (.a(net513),
    .b(_10082_),
    .c(_10090_),
    .d(_10091_),
    .o1(_10092_));
 b15zdnd11an1n04x5 FILLER_0_1100 ();
 b15zdnd11an1n04x5 FILLER_0_1091 ();
 b15zdnd11an1n04x5 FILLER_0_1082 ();
 b15nor003ah1n02x5 _18753_ (.a(_09932_),
    .b(_09980_),
    .c(_10003_),
    .o1(_10096_));
 b15aoai13as1n03x5 _18754_ (.a(net518),
    .b(_10096_),
    .c(_10053_),
    .d(net507),
    .o1(_10097_));
 b15zdnd11an1n04x5 FILLER_0_1074 ();
 b15aoi022ar1n02x5 _18756_ (.a(_10032_),
    .b(_09910_),
    .c(_09978_),
    .d(_10038_),
    .o1(_10099_));
 b15nonb02an1n12x5 _18757_ (.a(net506),
    .b(net518),
    .out0(_10100_));
 b15nanb02al1n06x5 _18758_ (.a(_10099_),
    .b(_10100_),
    .out0(_10101_));
 b15nandp2ar1n24x5 _18759_ (.a(net507),
    .b(_09907_),
    .o1(_10102_));
 b15nandp3ar1n02x5 _18760_ (.a(_09888_),
    .b(_09868_),
    .c(_09951_),
    .o1(_10103_));
 b15aob012an1n04x5 _18761_ (.a(_09932_),
    .b(_10102_),
    .c(_10103_),
    .out0(_10104_));
 b15nand04ah1n12x5 _18762_ (.a(_09892_),
    .b(_10097_),
    .c(_10101_),
    .d(_10104_),
    .o1(_10105_));
 b15aoi022aq1n12x5 _18763_ (.a(_10075_),
    .b(_10079_),
    .c(_10092_),
    .d(_10105_),
    .o1(_10106_));
 b15nano22al1n24x5 _18764_ (.a(net502),
    .b(net498),
    .c(net493),
    .out0(_10107_));
 b15nand02as1n16x5 _18765_ (.a(_09996_),
    .b(_10107_),
    .o1(_10108_));
 b15norp02ar1n02x5 _18766_ (.a(net513),
    .b(_10108_),
    .o1(_10109_));
 b15orn002ah1n03x5 _18767_ (.a(net504),
    .b(net499),
    .o(_10110_));
 b15norp03ar1n08x5 _18768_ (.a(_10071_),
    .b(_10110_),
    .c(_09925_),
    .o1(_10111_));
 b15nanb02aq1n16x5 _18769_ (.a(net510),
    .b(net509),
    .out0(_10112_));
 b15zdnd00an1n01x5 FILLER_0_1069 ();
 b15aoi012ah1n02x5 _18771_ (.a(_10053_),
    .b(_09951_),
    .c(net512),
    .o1(_10114_));
 b15oai022ar1n02x5 _18772_ (.a(_10112_),
    .b(_09993_),
    .c(_10114_),
    .d(net508),
    .o1(_10115_));
 b15oai013ar1n02x5 _18773_ (.a(net519),
    .b(_10109_),
    .c(_10111_),
    .d(_10115_),
    .o1(_10116_));
 b15nand02as1n12x5 _18774_ (.a(net516),
    .b(net508),
    .o1(_10117_));
 b15nandp3ar1n02x5 _18775_ (.a(_09982_),
    .b(_09887_),
    .c(_09983_),
    .o1(_10118_));
 b15and002an1n08x5 _18776_ (.a(net520),
    .b(net511),
    .o(_10119_));
 b15aoi012ar1n02x5 _18777_ (.a(_10119_),
    .b(_09921_),
    .c(_09871_),
    .o1(_10120_));
 b15aoi112ah1n02x5 _18778_ (.a(_10044_),
    .b(_10117_),
    .c(_10118_),
    .d(_10120_),
    .o1(_10121_));
 b15oai013an1n02x5 _18779_ (.a(_09946_),
    .b(_10022_),
    .c(_09994_),
    .d(net508),
    .o1(_10122_));
 b15oai012ar1n04x5 _18780_ (.a(_10006_),
    .b(_09940_),
    .c(net519),
    .o1(_10123_));
 b15aoi112aq1n04x5 _18781_ (.a(_10121_),
    .b(_10122_),
    .c(_10123_),
    .d(_10009_),
    .o1(_10124_));
 b15norp02an1n04x5 _18782_ (.a(net518),
    .b(_09940_),
    .o1(_10125_));
 b15nanb02ah1n04x5 _18783_ (.a(net494),
    .b(net503),
    .out0(_10126_));
 b15nand02as1n03x5 _18784_ (.a(net511),
    .b(net497),
    .o1(_10127_));
 b15nanb02ah1n24x5 _18785_ (.a(net506),
    .b(net494),
    .out0(_10128_));
 b15orn002as1n04x5 _18786_ (.a(net510),
    .b(net497),
    .o(_10129_));
 b15oai022as1n06x5 _18787_ (.a(_10126_),
    .b(_10127_),
    .c(_10128_),
    .d(_10129_),
    .o1(_10130_));
 b15nand03ah1n06x5 _18788_ (.a(net509),
    .b(net500),
    .c(_10130_),
    .o1(_10131_));
 b15orn003an1n24x5 _18789_ (.a(net501),
    .b(net498),
    .c(net493),
    .o(_10132_));
 b15norp03aq1n02x5 _18790_ (.a(net518),
    .b(_09980_),
    .c(_10132_),
    .o1(_10133_));
 b15aoi013an1n04x5 _18791_ (.a(_10133_),
    .b(_10130_),
    .c(net500),
    .d(net509),
    .o1(_10134_));
 b15oai022aq1n16x5 _18792_ (.a(_10125_),
    .b(_10131_),
    .c(_10134_),
    .d(_10006_),
    .o1(_10135_));
 b15norp03ar1n02x5 _18793_ (.a(net518),
    .b(net512),
    .c(net507),
    .o1(_10136_));
 b15ao0022ar1n03x5 _18794_ (.a(net507),
    .b(_10053_),
    .c(_10136_),
    .d(_09907_),
    .o(_10137_));
 b15nona23aq1n04x5 _18795_ (.a(net502),
    .b(net498),
    .c(net509),
    .d(net506),
    .out0(_10138_));
 b15orn003aq1n03x5 _18796_ (.a(net506),
    .b(net502),
    .c(net498),
    .o(_10139_));
 b15nand03as1n06x5 _18797_ (.a(net506),
    .b(net502),
    .c(net498),
    .o1(_10140_));
 b15aoai13as1n08x5 _18798_ (.a(_10138_),
    .b(_10071_),
    .c(_10139_),
    .d(_10140_),
    .o1(_10141_));
 b15aoi112ah1n06x5 _18799_ (.a(\u0.tmp_w[1] ),
    .b(_10137_),
    .c(_10141_),
    .d(net491),
    .o1(_10142_));
 b15norp02aq1n02x5 _18800_ (.a(net517),
    .b(_10142_),
    .o1(_10143_));
 b15nano23an1n05x5 _18801_ (.a(_10116_),
    .b(_10124_),
    .c(_10135_),
    .d(_10143_),
    .out0(_10144_));
 b15zdnd11an1n04x5 FILLER_0_1065 ();
 b15aoi013ar1n02x5 _18803_ (.a(_09932_),
    .b(net513),
    .c(_09949_),
    .d(_10068_),
    .o1(_10146_));
 b15nandp3ar1n02x5 _18804_ (.a(_09892_),
    .b(_09949_),
    .c(_10068_),
    .o1(_10147_));
 b15nandp2ah1n08x5 _18805_ (.a(_09868_),
    .b(_09978_),
    .o1(_10148_));
 b15aoi013ar1n02x5 _18806_ (.a(_10146_),
    .b(_10147_),
    .c(_10148_),
    .d(_09932_),
    .o1(_10149_));
 b15norp02ar1n02x5 _18807_ (.a(_10025_),
    .b(_10117_),
    .o1(_10150_));
 b15orn003ah1n03x5 _18808_ (.a(net513),
    .b(net504),
    .c(net499),
    .o(_10151_));
 b15aoi112al1n02x5 _18809_ (.a(_09908_),
    .b(_09925_),
    .c(_10151_),
    .d(_09896_),
    .o1(_10152_));
 b15orn003ar1n02x5 _18810_ (.a(net519),
    .b(_10150_),
    .c(_10152_),
    .o(_10153_));
 b15nand03an1n08x5 _18811_ (.a(net513),
    .b(net504),
    .c(net499),
    .o1(_10154_));
 b15oai112ar1n02x5 _18812_ (.a(_10038_),
    .b(net495),
    .c(net491),
    .d(_09932_),
    .o1(_10155_));
 b15oaoi13ar1n02x5 _18813_ (.a(_10154_),
    .b(_10155_),
    .c(_10073_),
    .d(_10038_),
    .o1(_10156_));
 b15oai022ar1n04x5 _18814_ (.a(_09888_),
    .b(_10149_),
    .c(_10153_),
    .d(_10156_),
    .o1(_10157_));
 b15nanb03aq1n02x5 _18815_ (.a(net500),
    .b(net504),
    .c(net513),
    .out0(_10158_));
 b15oaoi13ar1n03x5 _18816_ (.a(net520),
    .b(_10158_),
    .c(_09983_),
    .d(net513),
    .o1(_10159_));
 b15nanb03ar1n04x5 _18817_ (.a(net504),
    .b(net500),
    .c(net516),
    .out0(_10160_));
 b15oaoi13al1n03x5 _18818_ (.a(net513),
    .b(_10160_),
    .c(_09982_),
    .d(net516),
    .o1(_10161_));
 b15oai012an1n06x5 _18819_ (.a(_09859_),
    .b(_10159_),
    .c(_10161_),
    .o1(_10162_));
 b15nandp2ah1n12x5 _18820_ (.a(\u0.tmp_w[0] ),
    .b(net503),
    .o1(_10163_));
 b15nor002ar1n16x5 _18821_ (.a(_10003_),
    .b(_10163_),
    .o1(_10164_));
 b15nona23as1n32x5 _18822_ (.a(net499),
    .b(net495),
    .c(net491),
    .d(net504),
    .out0(_10165_));
 b15nor002aq1n16x5 _18823_ (.a(_09932_),
    .b(_10165_),
    .o1(_10166_));
 b15aoai13an1n06x5 _18824_ (.a(_09892_),
    .b(_10164_),
    .c(_10166_),
    .d(_09888_),
    .o1(_10167_));
 b15aoi012al1n08x5 _18825_ (.a(net511),
    .b(_09880_),
    .c(_09962_),
    .o1(_10168_));
 b15zdnd11an1n04x5 FILLER_0_1057 ();
 b15oai012al1n02x5 _18827_ (.a(net516),
    .b(_09926_),
    .c(net519),
    .o1(_10170_));
 b15nand02al1n02x5 _18828_ (.a(_09926_),
    .b(_10165_),
    .o1(_10171_));
 b15aoi012ar1n04x5 _18829_ (.a(_09892_),
    .b(_10170_),
    .c(_10171_),
    .o1(_10172_));
 b15oai112ah1n06x5 _18830_ (.a(_10162_),
    .b(_10167_),
    .c(_10168_),
    .d(_10172_),
    .o1(_10173_));
 b15zdnd00an1n02x5 FILLER_0_1049 ();
 b15aobi12al1n06x5 _18832_ (.a(_10157_),
    .b(_10173_),
    .c(_10038_),
    .out0(_10175_));
 b15nand02an1n12x5 _18833_ (.a(_10032_),
    .b(_09992_),
    .o1(_10176_));
 b15oaoi13as1n02x5 _18834_ (.a(_09994_),
    .b(_10025_),
    .c(_10176_),
    .d(net520),
    .o1(_10177_));
 b15nandp3an1n03x5 _18835_ (.a(net510),
    .b(_09992_),
    .c(_09964_),
    .o1(_10178_));
 b15oaoi13as1n02x5 _18836_ (.a(_09934_),
    .b(_10178_),
    .c(net511),
    .d(_10176_),
    .o1(_10179_));
 b15nandp2ar1n08x5 _18837_ (.a(_10032_),
    .b(_09871_),
    .o1(_10180_));
 b15nonb02as1n16x5 _18838_ (.a(net518),
    .b(net514),
    .out0(_10181_));
 b15nor004ah1n02x5 _18839_ (.a(_09892_),
    .b(_10180_),
    .c(_10023_),
    .d(_10181_),
    .o1(_10182_));
 b15nor003ah1n04x5 _18840_ (.a(_10177_),
    .b(_10179_),
    .c(_10182_),
    .o1(_10183_));
 b15zdnd11an1n04x5 FILLER_0_1045 ();
 b15nand02aq1n16x5 _18842_ (.a(_09888_),
    .b(net512),
    .o1(_10185_));
 b15oai022as1n02x5 _18843_ (.a(net511),
    .b(_10132_),
    .c(_10185_),
    .d(_09993_),
    .o1(_10186_));
 b15nanb02ar1n02x5 _18844_ (.a(_10142_),
    .b(_10186_),
    .out0(_10187_));
 b15aob012an1n06x5 _18845_ (.a(net508),
    .b(_10183_),
    .c(_10187_),
    .out0(_10188_));
 b15nand04as1n16x5 _18846_ (.a(_10106_),
    .b(_10144_),
    .c(_10175_),
    .d(_10188_),
    .o1(_10189_));
 b15xnr002aq1n12x5 _18847_ (.a(\u0.w[0][9] ),
    .b(_10189_),
    .out0(_10190_));
 b15xor002an1n16x5 _18848_ (.a(\u0.w[1][9] ),
    .b(_10190_),
    .out0(_10191_));
 b15xor002as1n16x5 _18849_ (.a(\u0.w[2][9] ),
    .b(_10191_),
    .out0(_10192_));
 b15xor002al1n02x5 _18850_ (.a(\u0.tmp_w[9] ),
    .b(_10192_),
    .out0(_10193_));
 b15mdn022ar1n02x5 _18851_ (.a(_10064_),
    .b(_10193_),
    .o1(_00384_),
    .sa(net944));
 b15nand02al1n16x5 _18852_ (.a(net947),
    .b(net12),
    .o1(_10194_));
 b15zdnd00an1n02x5 FILLER_0_1039 ();
 b15zdnd11an1n08x5 FILLER_0_1031 ();
 b15zdnd11an1n04x5 FILLER_0_1022 ();
 b15zdnd00an1n01x5 FILLER_0_1015 ();
 b15nano23al1n08x5 _18857_ (.a(net501),
    .b(net492),
    .c(net497),
    .d(net503),
    .out0(_10199_));
 b15nandp3as1n03x5 _18858_ (.a(net514),
    .b(net509),
    .c(_10199_),
    .o1(_10200_));
 b15norp02aq1n04x5 _18859_ (.a(net506),
    .b(net493),
    .o1(_10201_));
 b15and002ah1n04x5 _18860_ (.a(net506),
    .b(net493),
    .o(_10202_));
 b15aoi022ah1n06x5 _18861_ (.a(_09899_),
    .b(_10201_),
    .c(_09876_),
    .d(_10202_),
    .o1(_10203_));
 b15nanb02aq1n24x5 _18862_ (.a(net498),
    .b(net502),
    .out0(_10204_));
 b15oaoi13ar1n08x5 _18863_ (.a(net518),
    .b(_10200_),
    .c(_10203_),
    .d(_10204_),
    .o1(_10205_));
 b15nanb02as1n24x5 _18864_ (.a(net508),
    .b(net520),
    .out0(_10206_));
 b15oai012ah1n02x5 _18865_ (.a(_10107_),
    .b(_10006_),
    .c(_09901_),
    .o1(_10207_));
 b15nonb02as1n16x5 _18866_ (.a(net514),
    .b(net510),
    .out0(_10208_));
 b15zdnd11an1n04x5 FILLER_0_1011 ();
 b15aoi112as1n04x5 _18868_ (.a(_10206_),
    .b(_10207_),
    .c(_10208_),
    .d(_10176_),
    .o1(_10210_));
 b15nandp2aq1n16x5 _18869_ (.a(net503),
    .b(net494),
    .o1(_10211_));
 b15nonb02al1n06x5 _18870_ (.a(net497),
    .b(net501),
    .out0(_10212_));
 b15nonb02an1n12x5 _18871_ (.a(\u0.tmp_w[3] ),
    .b(\u0.tmp_w[0] ),
    .out0(_10213_));
 b15xor002al1n03x5 _18872_ (.a(net501),
    .b(net497),
    .out0(_10214_));
 b15aoi022ar1n02x5 _18873_ (.a(net514),
    .b(_10212_),
    .c(_10213_),
    .d(_10214_),
    .o1(_10215_));
 b15nor003ah1n02x5 _18874_ (.a(_09892_),
    .b(_10211_),
    .c(_10215_),
    .o1(_10216_));
 b15nor002aq1n04x5 _18875_ (.a(net518),
    .b(_09892_),
    .o1(_10217_));
 b15oaoi13aq1n04x5 _18876_ (.a(_09918_),
    .b(_10165_),
    .c(_10217_),
    .d(_10176_),
    .o1(_10218_));
 b15nor004an1n06x5 _18877_ (.a(_10205_),
    .b(_10210_),
    .c(_10216_),
    .d(_10218_),
    .o1(_10219_));
 b15nor002an1n12x5 _18878_ (.a(_09982_),
    .b(_10073_),
    .o1(_10220_));
 b15nandp2al1n12x5 _18879_ (.a(net501),
    .b(net497),
    .o1(_10221_));
 b15nanb03ah1n03x5 _18880_ (.a(\u0.tmp_w[3] ),
    .b(net503),
    .c(net494),
    .out0(_10222_));
 b15orn002ar1n08x5 _18881_ (.a(net503),
    .b(net494),
    .o(_10223_));
 b15oaoi13as1n08x5 _18882_ (.a(_10221_),
    .b(_10222_),
    .c(_10223_),
    .d(_10038_),
    .o1(_10224_));
 b15oab012ar1n02x5 _18883_ (.a(_10017_),
    .b(_10220_),
    .c(_10224_),
    .out0(_10225_));
 b15aoai13aq1n03x5 _18884_ (.a(_09892_),
    .b(_10225_),
    .c(_10224_),
    .d(_10014_),
    .o1(_10226_));
 b15norp03aq1n02x5 _18885_ (.a(net509),
    .b(_09939_),
    .c(_09953_),
    .o1(_10227_));
 b15aoi012al1n04x5 _18886_ (.a(_10227_),
    .b(_10224_),
    .c(_10181_),
    .o1(_10228_));
 b15oai112as1n12x5 _18887_ (.a(_10219_),
    .b(_10226_),
    .c(_10228_),
    .d(_09892_),
    .o1(_10229_));
 b15nand02as1n06x5 _18888_ (.a(net501),
    .b(_09859_),
    .o1(_10230_));
 b15aoi012ar1n02x5 _18889_ (.a(_09901_),
    .b(_10017_),
    .c(net512),
    .o1(_10231_));
 b15aoai13al1n02x5 _18890_ (.a(_09994_),
    .b(net514),
    .c(_09858_),
    .d(_09859_),
    .o1(_10232_));
 b15aoi112aq1n03x5 _18891_ (.a(_10230_),
    .b(_10231_),
    .c(_10232_),
    .d(_09888_),
    .o1(_10233_));
 b15aoai13ar1n02x5 _18892_ (.a(net518),
    .b(_09936_),
    .c(_10208_),
    .d(net503),
    .o1(_10234_));
 b15nor002ar1n06x5 _18893_ (.a(net512),
    .b(net503),
    .o1(_10235_));
 b15aob012ah1n03x5 _18894_ (.a(_10234_),
    .b(_10235_),
    .c(_10023_),
    .out0(_10236_));
 b15aoi012an1n08x5 _18895_ (.a(_10233_),
    .b(_10236_),
    .c(_09977_),
    .o1(_10237_));
 b15norp02ah1n12x5 _18896_ (.a(net514),
    .b(net510),
    .o1(_10238_));
 b15norp02ar1n02x5 _18897_ (.a(_09892_),
    .b(_09939_),
    .o1(_10239_));
 b15aoi022an1n04x5 _18898_ (.a(_10220_),
    .b(_10238_),
    .c(_10224_),
    .d(_10239_),
    .o1(_10240_));
 b15nonb02an1n12x5 _18899_ (.a(net514),
    .b(net503),
    .out0(_10241_));
 b15nandp2ar1n03x5 _18900_ (.a(_10212_),
    .b(_10241_),
    .o1(_10242_));
 b15zdnd00an1n01x5 FILLER_0_1006 ();
 b15nonb02as1n08x5 _18902_ (.a(net501),
    .b(net497),
    .out0(_10244_));
 b15nandp3ar1n02x5 _18903_ (.a(net503),
    .b(_10244_),
    .c(_10238_),
    .o1(_10245_));
 b15aoi112aq1n02x5 _18904_ (.a(\u0.tmp_w[0] ),
    .b(net494),
    .c(_10242_),
    .d(_10245_),
    .o1(_10246_));
 b15and002ar1n02x5 _18905_ (.a(net510),
    .b(net501),
    .o(_10247_));
 b15inv000al1n24x5 _18906_ (.a(net501),
    .o1(_10248_));
 b15aoi012ar1n02x5 _18907_ (.a(_10247_),
    .b(_10238_),
    .c(_10248_),
    .o1(_10249_));
 b15nor003ar1n04x5 _18908_ (.a(_10044_),
    .b(_10163_),
    .c(_10249_),
    .o1(_10250_));
 b15nanb02ah1n12x5 _18909_ (.a(net494),
    .b(net510),
    .out0(_10251_));
 b15oaoi13aq1n02x5 _18910_ (.a(_10251_),
    .b(_10242_),
    .c(_10163_),
    .d(_10204_),
    .o1(_10252_));
 b15nand02aq1n16x5 _18911_ (.a(net505),
    .b(_09938_),
    .o1(_10253_));
 b15oai012ar1n02x5 _18912_ (.a(_10208_),
    .b(net501),
    .c(_09888_),
    .o1(_10254_));
 b15oai012aq1n03x5 _18913_ (.a(\u0.tmp_w[3] ),
    .b(_10253_),
    .c(_10254_),
    .o1(_10255_));
 b15nor004as1n04x5 _18914_ (.a(_10246_),
    .b(_10250_),
    .c(_10252_),
    .d(_10255_),
    .o1(_10256_));
 b15aoi022as1n08x5 _18915_ (.a(_10038_),
    .b(_10237_),
    .c(_10240_),
    .d(_10256_),
    .o1(_10257_));
 b15nor004ar1n08x5 _18916_ (.a(_09888_),
    .b(_09856_),
    .c(_09983_),
    .d(_10073_),
    .o1(_10258_));
 b15aoi112ar1n08x5 _18917_ (.a(_09932_),
    .b(_10258_),
    .c(_09945_),
    .d(_09931_),
    .o1(_10259_));
 b15nor002ah1n12x5 _18918_ (.a(net501),
    .b(net494),
    .o1(_10260_));
 b15nano22ar1n03x5 _18919_ (.a(net501),
    .b(net494),
    .c(net505),
    .out0(_10261_));
 b15aoi022ar1n02x5 _18920_ (.a(net505),
    .b(_10260_),
    .c(_10261_),
    .d(\u0.tmp_w[0] ),
    .o1(_10262_));
 b15orn003al1n02x5 _18921_ (.a(net497),
    .b(_09856_),
    .c(_10262_),
    .o(_10263_));
 b15nanb02as1n24x5 _18922_ (.a(net507),
    .b(net506),
    .out0(_10264_));
 b15aoi112an1n03x5 _18923_ (.a(net512),
    .b(net492),
    .c(_10264_),
    .d(_09922_),
    .o1(_10265_));
 b15aoai13aq1n08x5 _18924_ (.a(_10244_),
    .b(_10265_),
    .c(_10202_),
    .d(_09876_),
    .o1(_10266_));
 b15aoi012ar1n02x5 _18925_ (.a(net515),
    .b(_09967_),
    .c(_09964_),
    .o1(_10267_));
 b15aoi013ah1n02x5 _18926_ (.a(_10259_),
    .b(_10263_),
    .c(_10266_),
    .d(_10267_),
    .o1(_10268_));
 b15and002al1n16x5 _18927_ (.a(net509),
    .b(net505),
    .o(_10269_));
 b15and003ar1n02x5 _18928_ (.a(_10017_),
    .b(_10269_),
    .c(_09978_),
    .o(_10270_));
 b15aoi013al1n03x5 _18929_ (.a(_10270_),
    .b(_10054_),
    .c(_09880_),
    .d(_10038_),
    .o1(_10271_));
 b15oai022ar1n02x5 _18930_ (.a(net514),
    .b(_09856_),
    .c(_09994_),
    .d(\u0.tmp_w[0] ),
    .o1(_10272_));
 b15orn002ah1n16x5 _18931_ (.a(net510),
    .b(\u0.tmp_w[3] ),
    .o(_10273_));
 b15oai012ar1n02x5 _18932_ (.a(_09856_),
    .b(_10273_),
    .c(net514),
    .o1(_10274_));
 b15aoi012ar1n02x5 _18933_ (.a(_10272_),
    .b(_10274_),
    .c(\u0.tmp_w[0] ),
    .o1(_10275_));
 b15oai022ar1n02x5 _18934_ (.a(net510),
    .b(_10271_),
    .c(_10275_),
    .d(_09926_),
    .o1(_10276_));
 b15aoi012al1n08x5 _18935_ (.a(_09970_),
    .b(_10023_),
    .c(_09974_),
    .o1(_10277_));
 b15nor003ah1n02x5 _18936_ (.a(net500),
    .b(_10112_),
    .c(_10277_),
    .o1(_10278_));
 b15nand03al1n08x5 _18937_ (.a(_09949_),
    .b(_10181_),
    .c(_09951_),
    .o1(_10279_));
 b15nonb02aq1n16x5 _18938_ (.a(net501),
    .b(net514),
    .out0(_10280_));
 b15orn003as1n02x5 _18939_ (.a(_10071_),
    .b(_10128_),
    .c(_10280_),
    .o(_10281_));
 b15nand02aq1n24x5 _18940_ (.a(\u0.tmp_w[1] ),
    .b(net511),
    .o1(_10282_));
 b15nand02as1n08x5 _18941_ (.a(_09868_),
    .b(_10050_),
    .o1(_10283_));
 b15oai112al1n16x5 _18942_ (.a(_10279_),
    .b(_10281_),
    .c(_10282_),
    .d(_10283_),
    .o1(_10284_));
 b15nano22al1n02x5 _18943_ (.a(net497),
    .b(net494),
    .c(net503),
    .out0(_10285_));
 b15oai112al1n06x5 _18944_ (.a(_10208_),
    .b(_10285_),
    .c(_10213_),
    .d(_10248_),
    .o1(_10286_));
 b15aoi012ar1n02x5 _18945_ (.a(_10208_),
    .b(_09905_),
    .c(_09888_),
    .o1(_10287_));
 b15aob012ar1n02x5 _18946_ (.a(_10286_),
    .b(_10287_),
    .c(_10009_),
    .out0(_10288_));
 b15nor003an1n02x5 _18947_ (.a(_10181_),
    .b(_10273_),
    .c(_09993_),
    .o1(_10289_));
 b15nor004aq1n06x5 _18948_ (.a(_10278_),
    .b(_10284_),
    .c(_10288_),
    .d(_10289_),
    .o1(_10290_));
 b15aoai13ar1n02x5 _18949_ (.a(net520),
    .b(net510),
    .c(_10264_),
    .d(_10068_),
    .o1(_10291_));
 b15aoi013aq1n03x5 _18950_ (.a(_10291_),
    .b(_10148_),
    .c(_10102_),
    .d(net510),
    .o1(_10292_));
 b15aoi013al1n03x5 _18951_ (.a(_10292_),
    .b(_10224_),
    .c(_10014_),
    .d(_10038_),
    .o1(_10293_));
 b15nona23aq1n08x5 _18952_ (.a(_10268_),
    .b(_10276_),
    .c(_10290_),
    .d(_10293_),
    .out0(_10294_));
 b15norp03ar1n24x5 _18953_ (.a(_10229_),
    .b(_10257_),
    .c(_10294_),
    .o1(_10295_));
 b15xor002as1n06x5 _18954_ (.a(\u0.w[0][10] ),
    .b(_10295_),
    .out0(_10296_));
 b15xor002as1n08x5 _18955_ (.a(\u0.w[1][10] ),
    .b(_10296_),
    .out0(_10297_));
 b15xor002al1n16x5 _18956_ (.a(\u0.w[2][10] ),
    .b(_10297_),
    .out0(_10298_));
 b15xor002ar1n02x5 _18957_ (.a(\u0.tmp_w[10] ),
    .b(_10298_),
    .out0(_10299_));
 b15oai012al1n02x5 _18958_ (.a(_10194_),
    .b(_10299_),
    .c(net945),
    .o1(_00354_));
 b15nand02aq1n12x5 _18959_ (.a(net129),
    .b(net23),
    .o1(_10300_));
 b15zdnd11an1n04x5 FILLER_0_1002 ();
 b15zdnd11an1n04x5 FILLER_0_994 ();
 b15zdnd00an1n01x5 FILLER_0_989 ();
 b15zdnd11an1n04x5 FILLER_0_985 ();
 b15aoi112ar1n02x5 _18964_ (.a(net519),
    .b(_10166_),
    .c(_10010_),
    .d(_09932_),
    .o1(_10305_));
 b15aoi012al1n04x5 _18965_ (.a(_09894_),
    .b(_10151_),
    .c(_10154_),
    .o1(_10306_));
 b15nanb02as1n12x5 _18966_ (.a(\u0.tmp_w[4] ),
    .b(net513),
    .out0(_10307_));
 b15nand02aq1n04x5 _18967_ (.a(net499),
    .b(net491),
    .o1(_10308_));
 b15oai022al1n08x5 _18968_ (.a(net513),
    .b(_10089_),
    .c(_10307_),
    .d(_10308_),
    .o1(_10309_));
 b15nonb02an1n04x5 _18969_ (.a(net517),
    .b(net495),
    .out0(_10310_));
 b15aoi022ah1n06x5 _18970_ (.a(_09932_),
    .b(_10306_),
    .c(_10309_),
    .d(_10310_),
    .o1(_10311_));
 b15norp02ar1n02x5 _18971_ (.a(net517),
    .b(_10165_),
    .o1(_10312_));
 b15aoi012al1n02x5 _18972_ (.a(_10312_),
    .b(_10010_),
    .c(net517),
    .o1(_10313_));
 b15aoi013ar1n04x5 _18973_ (.a(_10305_),
    .b(_10311_),
    .c(_10313_),
    .d(net519),
    .o1(_10314_));
 b15aoi012ar1n02x5 _18974_ (.a(net519),
    .b(_09905_),
    .c(_10010_),
    .o1(_10315_));
 b15aoi012ah1n02x5 _18975_ (.a(_10315_),
    .b(_10311_),
    .c(_09993_),
    .o1(_10316_));
 b15oai022ah1n08x5 _18976_ (.a(net513),
    .b(_10314_),
    .c(_10316_),
    .d(_09945_),
    .o1(_10317_));
 b15nand02aq1n06x5 _18977_ (.a(net511),
    .b(_09915_),
    .o1(_10318_));
 b15orn002aq1n04x5 _18978_ (.a(net501),
    .b(net497),
    .o(_10319_));
 b15oaoi13aq1n03x5 _18979_ (.a(_10126_),
    .b(_10221_),
    .c(_10319_),
    .d(net514),
    .o1(_10320_));
 b15aoi013aq1n08x5 _18980_ (.a(_10320_),
    .b(_10241_),
    .c(_09964_),
    .d(net500),
    .o1(_10321_));
 b15oaoi13aq1n04x5 _18981_ (.a(net518),
    .b(_10318_),
    .c(_10321_),
    .d(net511),
    .o1(_10322_));
 b15nand03aq1n03x5 _18982_ (.a(net518),
    .b(_09859_),
    .c(_10280_),
    .o1(_10323_));
 b15oaoi13ar1n08x5 _18983_ (.a(_10307_),
    .b(_10323_),
    .c(_10044_),
    .d(_10280_),
    .o1(_10324_));
 b15nor004al1n12x5 _18984_ (.a(_10038_),
    .b(_09907_),
    .c(_10322_),
    .d(_10324_),
    .o1(_10325_));
 b15oai112ar1n08x5 _18985_ (.a(_09888_),
    .b(_10043_),
    .c(_10282_),
    .d(net505),
    .o1(_10326_));
 b15oai112al1n12x5 _18986_ (.a(_10050_),
    .b(_10326_),
    .c(_09888_),
    .d(_09936_),
    .o1(_10327_));
 b15aoi012aq1n06x5 _18987_ (.a(net509),
    .b(_10220_),
    .c(_10208_),
    .o1(_10328_));
 b15aoi022an1n16x5 _18988_ (.a(_10317_),
    .b(_10325_),
    .c(_10327_),
    .d(_10328_),
    .o1(_10329_));
 b15zdnd00an1n01x5 FILLER_0_979 ();
 b15oai112ar1n02x5 _18990_ (.a(net514),
    .b(_10185_),
    .c(_10199_),
    .d(net512),
    .o1(_10331_));
 b15nandp2al1n12x5 _18991_ (.a(net518),
    .b(net512),
    .o1(_10332_));
 b15oai012ar1n02x5 _18992_ (.a(_10332_),
    .b(_10164_),
    .c(net512),
    .o1(_10333_));
 b15oai012ah1n02x5 _18993_ (.a(_10331_),
    .b(_10333_),
    .c(net514),
    .o1(_10334_));
 b15oai012al1n08x5 _18994_ (.a(_10334_),
    .b(_10199_),
    .c(_10054_),
    .o1(_10335_));
 b15oai012ar1n03x5 _18995_ (.a(net520),
    .b(_09936_),
    .c(_10208_),
    .o1(_10336_));
 b15aoi012ar1n02x5 _18996_ (.a(_10176_),
    .b(_10024_),
    .c(_10336_),
    .o1(_10337_));
 b15oab012an1n02x5 _18997_ (.a(_10337_),
    .b(_10178_),
    .c(_10181_),
    .out0(_10338_));
 b15aoi012an1n06x5 _18998_ (.a(net509),
    .b(_10335_),
    .c(_10338_),
    .o1(_10339_));
 b15nand03an1n06x5 _18999_ (.a(_09858_),
    .b(_09938_),
    .c(_09916_),
    .o1(_10340_));
 b15nand04as1n02x5 _19000_ (.a(net500),
    .b(_09859_),
    .c(_09876_),
    .d(_10043_),
    .o1(_10341_));
 b15oai112as1n06x5 _19001_ (.a(_10340_),
    .b(_10341_),
    .c(_10273_),
    .d(_09993_),
    .o1(_10342_));
 b15aoai13ar1n02x5 _19002_ (.a(net492),
    .b(_09967_),
    .c(_09992_),
    .d(net508),
    .o1(_10343_));
 b15aoi022aq1n02x5 _19003_ (.a(net508),
    .b(_09858_),
    .c(_09996_),
    .d(_10248_),
    .o1(_10344_));
 b15oai022ar1n02x5 _19004_ (.a(net511),
    .b(_10343_),
    .c(_10344_),
    .d(_10251_),
    .o1(_10345_));
 b15aoai13ah1n02x5 _19005_ (.a(net520),
    .b(_10342_),
    .c(_10345_),
    .d(net497),
    .o1(_10346_));
 b15aoi022an1n04x5 _19006_ (.a(net515),
    .b(_10269_),
    .c(_10006_),
    .d(_09868_),
    .o1(_10347_));
 b15oai013aq1n08x5 _19007_ (.a(_10346_),
    .b(_10347_),
    .c(_10008_),
    .d(net520),
    .o1(_10348_));
 b15norp03ar1n04x5 _19008_ (.a(net515),
    .b(_10008_),
    .c(_09922_),
    .o1(_10349_));
 b15nor002ar1n03x5 _19009_ (.a(\u0.tmp_w[0] ),
    .b(_10349_),
    .o1(_10350_));
 b15oab012ar1n02x5 _19010_ (.a(_10009_),
    .b(_10040_),
    .c(net508),
    .out0(_10351_));
 b15nor003al1n04x5 _19011_ (.a(net511),
    .b(_10350_),
    .c(_10351_),
    .o1(_10352_));
 b15norp02ar1n08x5 _19012_ (.a(net512),
    .b(net499),
    .o1(_10353_));
 b15oai112ar1n04x5 _19013_ (.a(_09964_),
    .b(_10353_),
    .c(_09996_),
    .d(_09949_),
    .o1(_10354_));
 b15nandp2al1n03x5 _19014_ (.a(net502),
    .b(_10032_),
    .o1(_10355_));
 b15nand02as1n12x5 _19015_ (.a(net511),
    .b(_09949_),
    .o1(_10356_));
 b15oai012al1n02x5 _19016_ (.a(\u0.tmp_w[1] ),
    .b(_10355_),
    .c(_10356_),
    .o1(_10357_));
 b15oai022ar1n02x5 _19017_ (.a(_10180_),
    .b(_10206_),
    .c(_10069_),
    .d(net518),
    .o1(_10358_));
 b15nonb03ah1n03x5 _19018_ (.a(_10354_),
    .b(_10357_),
    .c(_10358_),
    .out0(_10359_));
 b15nanb02aq1n12x5 _19019_ (.a(net518),
    .b(net502),
    .out0(_10360_));
 b15nano23ar1n02x5 _19020_ (.a(_10032_),
    .b(_10360_),
    .c(_10307_),
    .d(net507),
    .out0(_10361_));
 b15oai022ar1n02x5 _19021_ (.a(_09860_),
    .b(_10206_),
    .c(_09985_),
    .d(_10185_),
    .o1(_10362_));
 b15norp03aq1n03x5 _19022_ (.a(\u0.tmp_w[1] ),
    .b(_10361_),
    .c(_10362_),
    .o1(_10363_));
 b15oaoi13an1n08x5 _19023_ (.a(_10359_),
    .b(_10363_),
    .c(_10332_),
    .d(_10069_),
    .o1(_10364_));
 b15oai022ar1n02x5 _19024_ (.a(net515),
    .b(_09990_),
    .c(_10002_),
    .d(_09914_),
    .o1(_10365_));
 b15aoi012ar1n02x5 _19025_ (.a(_10356_),
    .b(_10132_),
    .c(_10008_),
    .o1(_10366_));
 b15oab012an1n02x5 _19026_ (.a(net520),
    .b(_10365_),
    .c(_10366_),
    .out0(_10367_));
 b15nandp2ar1n03x5 _19027_ (.a(net514),
    .b(_10248_),
    .o1(_10368_));
 b15aoi022ar1n02x5 _19028_ (.a(net505),
    .b(_09938_),
    .c(_10235_),
    .d(_09859_),
    .o1(_10369_));
 b15oai012al1n02x5 _19029_ (.a(_10027_),
    .b(_10368_),
    .c(_10369_),
    .o1(_10370_));
 b15aoi013an1n02x5 _19030_ (.a(_10367_),
    .b(_10370_),
    .c(_09887_),
    .d(net508),
    .o1(_10371_));
 b15nand02aq1n16x5 _19031_ (.a(_10248_),
    .b(_09964_),
    .o1(_10372_));
 b15norp03as1n04x5 _19032_ (.a(_10264_),
    .b(_10372_),
    .c(_10332_),
    .o1(_10373_));
 b15nanb02aq1n08x5 _19033_ (.a(net503),
    .b(net497),
    .out0(_10374_));
 b15nanb02aq1n12x5 _19034_ (.a(net497),
    .b(net503),
    .out0(_10375_));
 b15oai022ar1n02x5 _19035_ (.a(net509),
    .b(_10374_),
    .c(_10375_),
    .d(_09918_),
    .o1(_10376_));
 b15nandp3ar1n02x5 _19036_ (.a(_10260_),
    .b(_10217_),
    .c(_10376_),
    .o1(_10377_));
 b15oai013aq1n02x5 _19037_ (.a(_10377_),
    .b(_09994_),
    .c(_09914_),
    .d(_09980_),
    .o1(_10378_));
 b15orn003ar1n02x5 _19038_ (.a(_10223_),
    .b(_10273_),
    .c(_10214_),
    .o(_10379_));
 b15nand02al1n12x5 _19039_ (.a(net514),
    .b(_09962_),
    .o1(_10380_));
 b15aoi012aq1n04x5 _19040_ (.a(_10379_),
    .b(_10380_),
    .c(_09888_),
    .o1(_10381_));
 b15and002an1n02x5 _19041_ (.a(_10139_),
    .b(_10140_),
    .o(_10382_));
 b15nanb02as1n12x5 _19042_ (.a(net509),
    .b(net493),
    .out0(_10383_));
 b15aoi012al1n02x5 _19043_ (.a(_09932_),
    .b(_10015_),
    .c(_10185_),
    .o1(_10384_));
 b15nor004aq1n06x5 _19044_ (.a(_10181_),
    .b(_10382_),
    .c(_10383_),
    .d(_10384_),
    .o1(_10385_));
 b15nor004an1n06x5 _19045_ (.a(_10373_),
    .b(_10378_),
    .c(_10381_),
    .d(_10385_),
    .o1(_10386_));
 b15nona23as1n04x5 _19046_ (.a(_10352_),
    .b(_10364_),
    .c(_10371_),
    .d(_10386_),
    .out0(_10387_));
 b15nor004as1n12x5 _19047_ (.a(_10329_),
    .b(_10339_),
    .c(_10348_),
    .d(_10387_),
    .o1(_10388_));
 b15xor002ah1n03x5 _19048_ (.a(\u0.w[0][11] ),
    .b(_10388_),
    .out0(_10389_));
 b15xor002aq1n06x5 _19049_ (.a(\u0.w[1][11] ),
    .b(_10389_),
    .out0(_10390_));
 b15xor003ar1n02x5 _19050_ (.a(\u0.tmp_w[11] ),
    .b(\u0.w[2][11] ),
    .c(_10390_),
    .out0(_10391_));
 b15oai012ar1n02x5 _19051_ (.a(_10300_),
    .b(_10391_),
    .c(net942),
    .o1(_00355_));
 b15nand02ar1n02x5 _19052_ (.a(net944),
    .b(net32),
    .o1(_10392_));
 b15zdnd11an1n04x5 FILLER_0_975 ();
 b15zdnd11an1n04x5 FILLER_0_965 ();
 b15norp03al1n03x5 _19055_ (.a(_09892_),
    .b(net508),
    .c(net492),
    .o1(_10395_));
 b15nand02aq1n04x5 _19056_ (.a(net508),
    .b(net492),
    .o1(_10396_));
 b15norp02ar1n03x5 _19057_ (.a(net513),
    .b(_10396_),
    .o1(_10397_));
 b15oai112al1n08x5 _19058_ (.a(net496),
    .b(_09871_),
    .c(_10395_),
    .d(_10397_),
    .o1(_10398_));
 b15norp02ar1n02x5 _19059_ (.a(_09892_),
    .b(_10165_),
    .o1(_10399_));
 b15norp03ar1n02x5 _19060_ (.a(net513),
    .b(_10110_),
    .c(_09925_),
    .o1(_10400_));
 b15oai112as1n02x5 _19061_ (.a(_09888_),
    .b(_10038_),
    .c(_10399_),
    .d(_10400_),
    .o1(_10401_));
 b15oai022ar1n02x5 _19062_ (.a(net504),
    .b(_09894_),
    .c(_10264_),
    .d(_09925_),
    .o1(_10402_));
 b15norp02ar1n02x5 _19063_ (.a(net500),
    .b(_09994_),
    .o1(_10403_));
 b15aoai13ah1n02x5 _19064_ (.a(net519),
    .b(_10111_),
    .c(_10402_),
    .d(_10403_),
    .o1(_10404_));
 b15aoi013as1n03x5 _19065_ (.a(_10014_),
    .b(_10398_),
    .c(_10401_),
    .d(_10404_),
    .o1(_10405_));
 b15nanb02aq1n04x5 _19066_ (.a(net502),
    .b(net498),
    .out0(_10406_));
 b15oaoi13ar1n08x5 _19067_ (.a(_10383_),
    .b(_10406_),
    .c(net512),
    .d(_10204_),
    .o1(_10407_));
 b15aoai13ah1n08x5 _19068_ (.a(_10100_),
    .b(_10407_),
    .c(net509),
    .d(_09977_),
    .o1(_10408_));
 b15aoi012aq1n02x5 _19069_ (.a(_09932_),
    .b(_09907_),
    .c(_09899_),
    .o1(_10409_));
 b15nandp3ah1n08x5 _19070_ (.a(_10069_),
    .b(_10408_),
    .c(_10409_),
    .o1(_10410_));
 b15oai112ah1n06x5 _19071_ (.a(_09932_),
    .b(_09952_),
    .c(_10108_),
    .d(net519),
    .o1(_10411_));
 b15aoi012aq1n08x5 _19072_ (.a(_10405_),
    .b(_10410_),
    .c(_10411_),
    .o1(_10412_));
 b15nor002an1n03x5 _19073_ (.a(net511),
    .b(_09901_),
    .o1(_10413_));
 b15nand02ar1n02x5 _19074_ (.a(_09951_),
    .b(_10413_),
    .o1(_10414_));
 b15aoi012an1n02x5 _19075_ (.a(net508),
    .b(_09860_),
    .c(_10414_),
    .o1(_10415_));
 b15oaoi13ar1n02x5 _19076_ (.a(net505),
    .b(_10008_),
    .c(_10132_),
    .d(net520),
    .o1(_10416_));
 b15oai012ar1n02x5 _19077_ (.a(_09892_),
    .b(_09897_),
    .c(_10416_),
    .o1(_10417_));
 b15oai012an1n04x5 _19078_ (.a(_10417_),
    .b(_09993_),
    .c(_09888_),
    .o1(_10418_));
 b15aoai13aq1n06x5 _19079_ (.a(_09932_),
    .b(_10415_),
    .c(_10418_),
    .d(_10273_),
    .o1(_10419_));
 b15nandp3ar1n02x5 _19080_ (.a(net508),
    .b(_09858_),
    .c(_09863_),
    .o1(_10420_));
 b15aoi022ar1n02x5 _19081_ (.a(_09899_),
    .b(_09992_),
    .c(_09876_),
    .d(_09967_),
    .o1(_10421_));
 b15oaoi13ah1n03x5 _19082_ (.a(_09894_),
    .b(_10420_),
    .c(_10421_),
    .d(net520),
    .o1(_10422_));
 b15aoai13ar1n04x5 _19083_ (.a(net519),
    .b(_09940_),
    .c(_10238_),
    .d(net508),
    .o1(_10423_));
 b15nand03an1n02x5 _19084_ (.a(net511),
    .b(_09908_),
    .c(_09918_),
    .o1(_10424_));
 b15aoi012al1n04x5 _19085_ (.a(_09985_),
    .b(_10423_),
    .c(_10424_),
    .o1(_10425_));
 b15nand03an1n12x5 _19086_ (.a(_10038_),
    .b(_09858_),
    .c(_09859_),
    .o1(_10426_));
 b15nandp3ar1n02x5 _19087_ (.a(_10269_),
    .b(_09978_),
    .c(_10208_),
    .o1(_10427_));
 b15aoi012aq1n02x5 _19088_ (.a(net520),
    .b(_10426_),
    .c(_10427_),
    .o1(_10428_));
 b15nor004as1n02x5 _19089_ (.a(net508),
    .b(_09983_),
    .c(_10044_),
    .d(_10014_),
    .o1(_10429_));
 b15aoi112aq1n04x5 _19090_ (.a(net513),
    .b(_10429_),
    .c(_09915_),
    .d(net508),
    .o1(_10430_));
 b15nor003ah1n02x5 _19091_ (.a(net504),
    .b(net500),
    .c(net496),
    .o1(_10431_));
 b15and002ar1n02x5 _19092_ (.a(_09916_),
    .b(_10431_),
    .o(_10432_));
 b15oai022ar1n04x5 _19093_ (.a(_10038_),
    .b(_09982_),
    .c(_09983_),
    .d(_10206_),
    .o1(_10433_));
 b15and002ar1n02x5 _19094_ (.a(net516),
    .b(net496),
    .o(_10434_));
 b15aoai13aq1n03x5 _19095_ (.a(net492),
    .b(_10432_),
    .c(_10433_),
    .d(_10434_),
    .o1(_10435_));
 b15aoi022ar1n02x5 _19096_ (.a(net496),
    .b(_09992_),
    .c(_10431_),
    .d(net520),
    .o1(_10436_));
 b15oa0022ah1n02x5 _19097_ (.a(net508),
    .b(_10132_),
    .c(_10360_),
    .d(_10044_),
    .o(_10437_));
 b15oa0022ar1n02x5 _19098_ (.a(_10396_),
    .b(_10436_),
    .c(_10437_),
    .d(_10043_),
    .o(_10438_));
 b15aoi013an1n04x5 _19099_ (.a(_10430_),
    .b(_10435_),
    .c(_10438_),
    .d(_09898_),
    .o1(_10439_));
 b15nor004ah1n06x5 _19100_ (.a(_10422_),
    .b(_10425_),
    .c(_10428_),
    .d(_10439_),
    .o1(_10440_));
 b15oai012ar1n04x5 _19101_ (.a(net520),
    .b(_09867_),
    .c(_10050_),
    .o1(_10441_));
 b15oaoi13ar1n02x5 _19102_ (.a(_10356_),
    .b(_10441_),
    .c(net515),
    .d(_10132_),
    .o1(_10442_));
 b15oai112al1n02x5 _19103_ (.a(_09901_),
    .b(_10050_),
    .c(_10006_),
    .d(net520),
    .o1(_10443_));
 b15aoi112al1n02x5 _19104_ (.a(net508),
    .b(_10119_),
    .c(_10443_),
    .d(_09990_),
    .o1(_10444_));
 b15nandp3ar1n02x5 _19105_ (.a(net510),
    .b(net497),
    .c(net494),
    .o1(_10445_));
 b15oai012al1n02x5 _19106_ (.a(_10445_),
    .b(_10129_),
    .c(net494),
    .o1(_10446_));
 b15aob012ah1n04x5 _19107_ (.a(net515),
    .b(_09967_),
    .c(_10446_),
    .out0(_10447_));
 b15aoi012ar1n02x5 _19108_ (.a(_10442_),
    .b(_10444_),
    .c(_10447_),
    .o1(_10448_));
 b15nand03an1n08x5 _19109_ (.a(net520),
    .b(_09905_),
    .c(_09994_),
    .o1(_10449_));
 b15oaoi13al1n04x5 _19110_ (.a(_10148_),
    .b(_10449_),
    .c(net520),
    .d(_09994_),
    .o1(_10450_));
 b15oai022ar1n02x5 _19111_ (.a(_10008_),
    .b(_09918_),
    .c(_10132_),
    .d(_09908_),
    .o1(_10451_));
 b15nonb02ar1n02x5 _19112_ (.a(_10451_),
    .b(_10163_),
    .out0(_10452_));
 b15aoi012ar1n04x5 _19113_ (.a(_09892_),
    .b(_09939_),
    .c(_09945_),
    .o1(_10453_));
 b15nand03an1n06x5 _19114_ (.a(net492),
    .b(_09910_),
    .c(_10006_),
    .o1(_10454_));
 b15aoi112ar1n08x5 _19115_ (.a(_10453_),
    .b(_10454_),
    .c(_10374_),
    .d(_10375_),
    .o1(_10455_));
 b15norp03as1n04x5 _19116_ (.a(_10450_),
    .b(_10452_),
    .c(_10455_),
    .o1(_10456_));
 b15norp03ar1n02x5 _19117_ (.a(net520),
    .b(_09936_),
    .c(_10208_),
    .o1(_10457_));
 b15aoai13ar1n03x5 _19118_ (.a(_09962_),
    .b(_10457_),
    .c(_10208_),
    .d(net520),
    .o1(_10458_));
 b15aoi022aq1n02x5 _19119_ (.a(_10260_),
    .b(_10413_),
    .c(_10261_),
    .d(_10119_),
    .o1(_10459_));
 b15nandp2ar1n03x5 _19120_ (.a(_09932_),
    .b(net497),
    .o1(_10460_));
 b15oaoi13aq1n04x5 _19121_ (.a(net508),
    .b(_10458_),
    .c(_10459_),
    .d(_10460_),
    .o1(_10461_));
 b15oai112an1n04x5 _19122_ (.a(net520),
    .b(_10160_),
    .c(_10006_),
    .d(_09982_),
    .o1(_10462_));
 b15oai012an1n04x5 _19123_ (.a(_10158_),
    .b(_09983_),
    .c(net516),
    .o1(_10463_));
 b15oai112aq1n08x5 _19124_ (.a(_09859_),
    .b(_10462_),
    .c(_10463_),
    .d(net520),
    .o1(_10464_));
 b15qgbno2an1n10x5 _19125_ (.a(_09888_),
    .b(_09932_),
    .o1(_10465_));
 b15nonb02ar1n02x5 _19126_ (.a(net492),
    .b(net515),
    .out0(_10466_));
 b15oaoi13ar1n02x5 _19127_ (.a(_09936_),
    .b(net520),
    .c(net511),
    .d(_10466_),
    .o1(_10467_));
 b15oa0022al1n02x5 _19128_ (.a(_10465_),
    .b(_10251_),
    .c(_10467_),
    .d(net496),
    .o(_10468_));
 b15oaoi13an1n03x5 _19129_ (.a(_10038_),
    .b(_10464_),
    .c(_10468_),
    .d(_09983_),
    .o1(_10469_));
 b15nano23al1n06x5 _19130_ (.a(_10448_),
    .b(_10456_),
    .c(_10461_),
    .d(_10469_),
    .out0(_10470_));
 b15nand04as1n16x5 _19131_ (.a(_10412_),
    .b(_10419_),
    .c(_10440_),
    .d(_10470_),
    .o1(_10471_));
 b15xnr002as1n16x5 _19132_ (.a(\u0.w[0][12] ),
    .b(_10471_),
    .out0(_10472_));
 b15xor002ah1n12x5 _19133_ (.a(\u0.w[1][12] ),
    .b(_10472_),
    .out0(_10473_));
 b15xor002as1n16x5 _19134_ (.a(\u0.w[2][12] ),
    .b(_10473_),
    .out0(_10474_));
 b15xor002ar1n02x5 _19135_ (.a(net475),
    .b(_10474_),
    .out0(_10475_));
 b15oai012ar1n02x5 _19136_ (.a(_10392_),
    .b(_10475_),
    .c(net943),
    .o1(_00356_));
 b15nand02ar1n02x5 _19137_ (.a(net943),
    .b(net33),
    .o1(_10476_));
 b15zdnd00an1n01x5 FILLER_0_960 ();
 b15zdnd11an1n08x5 FILLER_0_952 ();
 b15zdnd11an1n04x5 FILLER_0_943 ();
 b15aoi012ar1n02x5 _19141_ (.a(net515),
    .b(_09868_),
    .c(_09951_),
    .o1(_10480_));
 b15nand03as1n08x5 _19142_ (.a(_09992_),
    .b(_09876_),
    .c(_09964_),
    .o1(_10481_));
 b15aoi013al1n04x5 _19143_ (.a(_10480_),
    .b(_10481_),
    .c(_09989_),
    .d(net515),
    .o1(_10482_));
 b15oai012as1n03x5 _19144_ (.a(_10355_),
    .b(_10372_),
    .c(_10282_),
    .o1(_10483_));
 b15aoi013aq1n03x5 _19145_ (.a(_10482_),
    .b(_10483_),
    .c(net507),
    .d(_09901_),
    .o1(_10484_));
 b15oai112an1n04x5 _19146_ (.a(net507),
    .b(_10068_),
    .c(_10017_),
    .d(_09901_),
    .o1(_10485_));
 b15aob012ar1n02x5 _19147_ (.a(_09892_),
    .b(_10283_),
    .c(_10485_),
    .out0(_10486_));
 b15aoi012ar1n02x5 _19148_ (.a(_09888_),
    .b(_09876_),
    .c(_09915_),
    .o1(_10487_));
 b15oaoi13ar1n02x5 _19149_ (.a(_10273_),
    .b(_09860_),
    .c(_10372_),
    .d(_10035_),
    .o1(_10488_));
 b15nano22aq1n03x5 _19150_ (.a(_10486_),
    .b(_10487_),
    .c(_10488_),
    .out0(_10489_));
 b15nand02al1n02x5 _19151_ (.a(net513),
    .b(net504),
    .o1(_10490_));
 b15nandp2ar1n02x5 _19152_ (.a(net508),
    .b(_09978_),
    .o1(_10491_));
 b15oaoi13an1n04x5 _19153_ (.a(_10490_),
    .b(_10491_),
    .c(net508),
    .d(_09914_),
    .o1(_10492_));
 b15oai022aq1n02x5 _19154_ (.a(_10038_),
    .b(_09926_),
    .c(_10022_),
    .d(_10273_),
    .o1(_10493_));
 b15nano23as1n06x5 _19155_ (.a(_09888_),
    .b(_10340_),
    .c(_10492_),
    .d(_10493_),
    .out0(_10494_));
 b15aoi022ar1n02x5 _19156_ (.a(_09868_),
    .b(_09951_),
    .c(_10009_),
    .d(net513),
    .o1(_10495_));
 b15nanb02as1n03x5 _19157_ (.a(_10495_),
    .b(net517),
    .out0(_10496_));
 b15aoi022ar1n12x5 _19158_ (.a(_10484_),
    .b(_10489_),
    .c(_10494_),
    .d(_10496_),
    .o1(_10497_));
 b15oai012ar1n02x5 _19159_ (.a(_10038_),
    .b(_09905_),
    .c(_10165_),
    .o1(_10498_));
 b15oai022ar1n02x5 _19160_ (.a(net517),
    .b(_10165_),
    .c(_09985_),
    .d(_09994_),
    .o1(_10499_));
 b15aoi012as1n02x5 _19161_ (.a(_10498_),
    .b(_10499_),
    .c(_09888_),
    .o1(_10500_));
 b15oaoi13an1n02x5 _19162_ (.a(net519),
    .b(_09990_),
    .c(_09925_),
    .d(_09896_),
    .o1(_10501_));
 b15aoi112al1n03x5 _19163_ (.a(net513),
    .b(_10501_),
    .c(_10010_),
    .d(net517),
    .o1(_10502_));
 b15orn003ar1n02x5 _19164_ (.a(_09901_),
    .b(_10248_),
    .c(net491),
    .o(_10503_));
 b15aob012ar1n02x5 _19165_ (.a(_10181_),
    .b(_09990_),
    .c(_10503_),
    .out0(_10504_));
 b15aoi013ar1n02x5 _19166_ (.a(_10502_),
    .b(_10504_),
    .c(_09985_),
    .d(net513),
    .o1(_10505_));
 b15norp02aq1n02x5 _19167_ (.a(net493),
    .b(_10087_),
    .o1(_10506_));
 b15nor002al1n06x5 _19168_ (.a(net512),
    .b(_10406_),
    .o1(_10507_));
 b15aoai13an1n08x5 _19169_ (.a(_10506_),
    .b(_10507_),
    .c(_10244_),
    .d(net518),
    .o1(_10508_));
 b15nand02an1n03x5 _19170_ (.a(_10032_),
    .b(_10100_),
    .o1(_10509_));
 b15aoi012al1n02x5 _19171_ (.a(_10353_),
    .b(_09940_),
    .c(net502),
    .o1(_10510_));
 b15oai112as1n08x5 _19172_ (.a(net507),
    .b(_10508_),
    .c(_10509_),
    .d(_10510_),
    .o1(_10511_));
 b15oab012an1n04x5 _19173_ (.a(_10500_),
    .b(_10505_),
    .c(_10511_),
    .out0(_10512_));
 b15aoi022ar1n12x5 _19174_ (.a(_09859_),
    .b(_10280_),
    .c(_10507_),
    .d(net493),
    .o1(_10513_));
 b15oai022an1n16x5 _19175_ (.a(_09860_),
    .b(_10185_),
    .c(_10513_),
    .d(net503),
    .o1(_10514_));
 b15nandp2ah1n03x5 _19176_ (.a(_09867_),
    .b(_09996_),
    .o1(_10515_));
 b15oai112an1n12x5 _19177_ (.a(_10181_),
    .b(_10515_),
    .c(_10108_),
    .d(net512),
    .o1(_10516_));
 b15aoi013an1n02x5 _19178_ (.a(net518),
    .b(_09936_),
    .c(_09949_),
    .d(_10068_),
    .o1(_10517_));
 b15oaoi13aq1n04x5 _19179_ (.a(_10517_),
    .b(net517),
    .c(net507),
    .d(_09953_),
    .o1(_10518_));
 b15aoi022ar1n04x5 _19180_ (.a(_09892_),
    .b(_09910_),
    .c(_09876_),
    .d(net499),
    .o1(_10519_));
 b15oai012al1n06x5 _19181_ (.a(_09932_),
    .b(_10253_),
    .c(_10519_),
    .o1(_10520_));
 b15nor002as1n02x5 _19182_ (.a(_10071_),
    .b(_10308_),
    .o1(_10521_));
 b15nanb02ar1n03x5 _19183_ (.a(net491),
    .b(net507),
    .out0(_10522_));
 b15aoi013ar1n04x5 _19184_ (.a(_10521_),
    .b(_10522_),
    .c(_10353_),
    .d(_10383_),
    .o1(_10523_));
 b15nand03an1n03x5 _19185_ (.a(\u0.tmp_w[4] ),
    .b(net495),
    .c(_09939_),
    .o1(_10524_));
 b15oai022as1n06x5 _19186_ (.a(_09876_),
    .b(_09926_),
    .c(_10523_),
    .d(_10524_),
    .o1(_10525_));
 b15aoi222as1n12x5 _19187_ (.a(_10038_),
    .b(_10514_),
    .c(_10516_),
    .d(_10518_),
    .e(_10520_),
    .f(_10525_),
    .o1(_10526_));
 b15oaoi13aq1n04x5 _19188_ (.a(_10168_),
    .b(net511),
    .c(_09926_),
    .d(_10465_),
    .o1(_10527_));
 b15oai022ar1n04x5 _19189_ (.a(_09905_),
    .b(_09953_),
    .c(_10003_),
    .d(_10087_),
    .o1(_10528_));
 b15aoai13al1n03x5 _19190_ (.a(_10038_),
    .b(_10527_),
    .c(_10528_),
    .d(_09888_),
    .o1(_10529_));
 b15orn002aq1n08x5 _19191_ (.a(net518),
    .b(net507),
    .o(_10530_));
 b15oai013ar1n02x5 _19192_ (.a(_10485_),
    .b(_10530_),
    .c(_09914_),
    .d(\u0.tmp_w[4] ),
    .o1(_10531_));
 b15aoi022ar1n02x5 _19193_ (.a(_09858_),
    .b(_09859_),
    .c(_10015_),
    .d(_10006_),
    .o1(_10532_));
 b15oaoi13ar1n02x5 _19194_ (.a(_10532_),
    .b(net518),
    .c(net511),
    .d(_09860_),
    .o1(_10533_));
 b15aoi022aq1n02x5 _19195_ (.a(_10208_),
    .b(_10531_),
    .c(_10533_),
    .d(net507),
    .o1(_10534_));
 b15oai112an1n02x5 _19196_ (.a(_09858_),
    .b(_09876_),
    .c(_09964_),
    .d(_10032_),
    .o1(_10535_));
 b15oa0012al1n04x5 _19197_ (.a(_10200_),
    .b(_10535_),
    .c(_09939_),
    .o(_10536_));
 b15oai022ar1n02x5 _19198_ (.a(net511),
    .b(_09980_),
    .c(_10375_),
    .d(_09856_),
    .o1(_10537_));
 b15nandp3aq1n03x5 _19199_ (.a(net492),
    .b(_10280_),
    .c(_10537_),
    .o1(_10538_));
 b15oai112al1n16x5 _19200_ (.a(_10269_),
    .b(_10449_),
    .c(_09892_),
    .d(_09880_),
    .o1(_10539_));
 b15oai112ah1n12x5 _19201_ (.a(_10536_),
    .b(_10538_),
    .c(_10539_),
    .d(_10132_),
    .o1(_10540_));
 b15nandp3ar1n02x5 _19202_ (.a(_09939_),
    .b(_10269_),
    .c(_10107_),
    .o1(_10541_));
 b15aob012aq1n02x5 _19203_ (.a(_09892_),
    .b(_09997_),
    .c(_10541_),
    .out0(_10542_));
 b15nona23al1n05x5 _19204_ (.a(_09894_),
    .b(_10280_),
    .c(_09996_),
    .d(_10368_),
    .out0(_10543_));
 b15oai112as1n08x5 _19205_ (.a(_09935_),
    .b(_10542_),
    .c(_10543_),
    .d(_09892_),
    .o1(_10544_));
 b15nano23as1n08x5 _19206_ (.a(_10529_),
    .b(_10534_),
    .c(_10540_),
    .d(_10544_),
    .out0(_10545_));
 b15nona23as1n32x5 _19207_ (.a(_10497_),
    .b(_10512_),
    .c(_10526_),
    .d(_10545_),
    .out0(_10546_));
 b15xnr002as1n16x5 _19208_ (.a(\u0.w[0][13] ),
    .b(_10546_),
    .out0(_10547_));
 b15xor002ah1n12x5 _19209_ (.a(\u0.w[1][13] ),
    .b(_10547_),
    .out0(_10548_));
 b15xor002as1n16x5 _19210_ (.a(\u0.w[2][13] ),
    .b(_10548_),
    .out0(_10549_));
 b15xor002ar1n02x5 _19211_ (.a(\u0.tmp_w[13] ),
    .b(_10549_),
    .out0(_10550_));
 b15zdnd00an1n01x5 FILLER_0_938 ();
 b15zdnd00an1n02x5 FILLER_0_936 ();
 b15oai012ar1n02x5 _19214_ (.a(_10476_),
    .b(_10550_),
    .c(net943),
    .o1(_00357_));
 b15inv020aq1n08x5 _19215_ (.a(net34),
    .o1(_10553_));
 b15zdnd11an1n04x5 FILLER_0_932 ();
 b15zdnd00an1n02x5 FILLER_0_926 ();
 b15zdnd11an1n16x5 FILLER_0_910 ();
 b15aoi013ar1n02x5 _19219_ (.a(net518),
    .b(\u0.tmp_w[1] ),
    .c(_09867_),
    .d(_09996_),
    .o1(_10557_));
 b15aoai13ah1n02x5 _19220_ (.a(net512),
    .b(_10557_),
    .c(_10515_),
    .d(_10069_),
    .o1(_10558_));
 b15oaoi13ar1n02x5 _19221_ (.a(net518),
    .b(_09922_),
    .c(_10264_),
    .d(\u0.tmp_w[1] ),
    .o1(_10559_));
 b15norp02ar1n02x5 _19222_ (.a(\u0.tmp_w[1] ),
    .b(_09922_),
    .o1(_10560_));
 b15oab012al1n04x5 _19223_ (.a(_10003_),
    .b(_10559_),
    .c(_10560_),
    .out0(_10561_));
 b15nano23al1n05x5 _19224_ (.a(net504),
    .b(net491),
    .c(net499),
    .d(net507),
    .out0(_10562_));
 b15nano23aq1n03x5 _19225_ (.a(net507),
    .b(net499),
    .c(net491),
    .d(net504),
    .out0(_10563_));
 b15oai012ar1n12x5 _19226_ (.a(_10310_),
    .b(_10562_),
    .c(_10563_),
    .o1(_10564_));
 b15oai122ah1n12x5 _19227_ (.a(_10564_),
    .b(_10530_),
    .c(_10165_),
    .d(_10017_),
    .e(_09997_),
    .o1(_10565_));
 b15oai013an1n08x5 _19228_ (.a(_10558_),
    .b(_10561_),
    .c(_10565_),
    .d(net512),
    .o1(_10566_));
 b15aoai13ar1n02x5 _19229_ (.a(net518),
    .b(_10107_),
    .c(_10068_),
    .d(net514),
    .o1(_10567_));
 b15oaoi13aq1n02x5 _19230_ (.a(net503),
    .b(_10567_),
    .c(_10372_),
    .d(_09880_),
    .o1(_10568_));
 b15oai022ar1n08x5 _19231_ (.a(\u0.tmp_w[1] ),
    .b(_09982_),
    .c(_10241_),
    .d(_10360_),
    .o1(_10569_));
 b15aoai13ah1n04x5 _19232_ (.a(_09931_),
    .b(_10568_),
    .c(_10569_),
    .d(_10032_),
    .o1(_10570_));
 b15nandp2an1n05x5 _19233_ (.a(_09858_),
    .b(_09938_),
    .o1(_10571_));
 b15oai122as1n04x5 _19234_ (.a(_10038_),
    .b(_10132_),
    .c(_09892_),
    .d(_10571_),
    .e(net514),
    .o1(_10572_));
 b15and003ar1n02x5 _19235_ (.a(net512),
    .b(net502),
    .c(net491),
    .o(_10573_));
 b15aoi012ar1n02x5 _19236_ (.a(_10573_),
    .b(_10260_),
    .c(_09921_),
    .o1(_10574_));
 b15nor003as1n03x5 _19237_ (.a(net495),
    .b(_10035_),
    .c(_10574_),
    .o1(_10575_));
 b15aoi012ah1n02x5 _19238_ (.a(_10202_),
    .b(_10201_),
    .c(net512),
    .o1(_10576_));
 b15nor003an1n08x5 _19239_ (.a(_10204_),
    .b(_09940_),
    .c(_10576_),
    .o1(_10577_));
 b15oai013an1n04x5 _19240_ (.a(net507),
    .b(_10023_),
    .c(_10132_),
    .d(_10307_),
    .o1(_10578_));
 b15oai013al1n08x5 _19241_ (.a(_10572_),
    .b(_10575_),
    .c(_10577_),
    .d(_10578_),
    .o1(_10579_));
 b15nanb02ar1n08x5 _19242_ (.a(_10206_),
    .b(_10053_),
    .out0(_10580_));
 b15nand03ar1n03x5 _19243_ (.a(net507),
    .b(_10031_),
    .c(_10107_),
    .o1(_10581_));
 b15oaoi13an1n03x5 _19244_ (.a(net512),
    .b(_10580_),
    .c(_10581_),
    .d(net518),
    .o1(_10582_));
 b15nand03aq1n02x5 _19245_ (.a(_09863_),
    .b(_09868_),
    .c(_09951_),
    .o1(_10583_));
 b15nor002ar1n02x5 _19246_ (.a(net507),
    .b(net495),
    .o1(_10584_));
 b15aoi022al1n06x5 _19247_ (.a(net495),
    .b(_09910_),
    .c(_10584_),
    .d(net502),
    .o1(_10585_));
 b15oai013ar1n08x5 _19248_ (.a(_10583_),
    .b(_10585_),
    .c(net518),
    .d(_10128_),
    .o1(_10586_));
 b15nand02al1n04x5 _19249_ (.a(net509),
    .b(net506),
    .o1(_10587_));
 b15nor002an1n06x5 _19250_ (.a(_10587_),
    .b(_10372_),
    .o1(_10588_));
 b15oaoi13al1n08x5 _19251_ (.a(_10582_),
    .b(_09932_),
    .c(_10586_),
    .d(_10588_),
    .o1(_10589_));
 b15nand04as1n16x5 _19252_ (.a(_10566_),
    .b(_10570_),
    .c(_10579_),
    .d(_10589_),
    .o1(_10590_));
 b15oai022as1n02x5 _19253_ (.a(_10038_),
    .b(_10375_),
    .c(_10530_),
    .d(_10374_),
    .o1(_10591_));
 b15oai022al1n04x5 _19254_ (.a(_10071_),
    .b(_10374_),
    .c(_10375_),
    .d(_10112_),
    .o1(_10592_));
 b15aoi022ar1n08x5 _19255_ (.a(_09940_),
    .b(_10591_),
    .c(_10592_),
    .d(_10181_),
    .o1(_10593_));
 b15nanb02an1n02x5 _19256_ (.a(_10593_),
    .b(_10260_),
    .out0(_10594_));
 b15aoi022an1n02x5 _19257_ (.a(net508),
    .b(_09858_),
    .c(_09876_),
    .d(_09967_),
    .o1(_10595_));
 b15oai112ar1n08x5 _19258_ (.a(net519),
    .b(_09946_),
    .c(_10072_),
    .d(_10595_),
    .o1(_10596_));
 b15oai022ah1n06x5 _19259_ (.a(_09918_),
    .b(_10025_),
    .c(_10481_),
    .d(_09932_),
    .o1(_10597_));
 b15oai012ar1n12x5 _19260_ (.a(_10596_),
    .b(_10597_),
    .c(net519),
    .o1(_10598_));
 b15norp03al1n02x5 _19261_ (.a(net510),
    .b(_10014_),
    .c(_09926_),
    .o1(_10599_));
 b15aoai13an1n03x5 _19262_ (.a(_10038_),
    .b(_10599_),
    .c(_09962_),
    .d(_09936_),
    .o1(_10600_));
 b15nor003ar1n06x5 _19263_ (.a(_09901_),
    .b(_09894_),
    .c(_10206_),
    .o1(_10601_));
 b15aoai13as1n02x5 _19264_ (.a(net510),
    .b(_10349_),
    .c(_10601_),
    .d(net515),
    .o1(_10602_));
 b15nand04as1n08x5 _19265_ (.a(_10594_),
    .b(_10598_),
    .c(_10600_),
    .d(_10602_),
    .o1(_10603_));
 b15norp03ar1n02x5 _19266_ (.a(net505),
    .b(_09908_),
    .c(_10204_),
    .o1(_10604_));
 b15aoi012ar1n02x5 _19267_ (.a(_10604_),
    .b(_10269_),
    .c(_10212_),
    .o1(_10605_));
 b15aoi022ar1n08x5 _19268_ (.a(_09916_),
    .b(_10010_),
    .c(_10054_),
    .d(_10213_),
    .o1(_10606_));
 b15oai022ar1n02x5 _19269_ (.a(_10251_),
    .b(_10605_),
    .c(_10606_),
    .d(net510),
    .o1(_10607_));
 b15aoi013ar1n02x5 _19270_ (.a(_09932_),
    .b(_09868_),
    .c(_09978_),
    .d(_10119_),
    .o1(_10608_));
 b15aoi012ar1n02x5 _19271_ (.a(_10608_),
    .b(_10102_),
    .c(_09932_),
    .o1(_10609_));
 b15aoi012ah1n02x5 _19272_ (.a(_10609_),
    .b(_10601_),
    .c(_10248_),
    .o1(_10610_));
 b15aoi012ar1n02x5 _19273_ (.a(_09888_),
    .b(_10038_),
    .c(_09993_),
    .o1(_10611_));
 b15oab012ar1n02x5 _19274_ (.a(net515),
    .b(_10038_),
    .c(_10054_),
    .out0(_10612_));
 b15oai122aq1n04x5 _19275_ (.a(_10611_),
    .b(_09962_),
    .c(_10112_),
    .d(_09892_),
    .e(_10612_),
    .o1(_10613_));
 b15nona23an1n05x5 _19276_ (.a(_10135_),
    .b(_10607_),
    .c(_10610_),
    .d(_10613_),
    .out0(_10614_));
 b15and003ar1n02x5 _19277_ (.a(net503),
    .b(net501),
    .c(net492),
    .o(_10615_));
 b15norp03ar1n03x5 _19278_ (.a(net503),
    .b(net501),
    .c(net492),
    .o1(_10616_));
 b15oai112ar1n08x5 _19279_ (.a(net497),
    .b(_09936_),
    .c(_10615_),
    .d(_10616_),
    .o1(_10617_));
 b15oai112as1n06x5 _19280_ (.a(net518),
    .b(_10617_),
    .c(_10087_),
    .d(_10230_),
    .o1(_10618_));
 b15aoi012aq1n08x5 _19281_ (.a(_10151_),
    .b(_09925_),
    .c(_09894_),
    .o1(_10619_));
 b15aoai13ar1n03x5 _19282_ (.a(_09992_),
    .b(_10000_),
    .c(_09938_),
    .d(_09892_),
    .o1(_10620_));
 b15aoi012ar1n04x5 _19283_ (.a(net515),
    .b(_10040_),
    .c(_10620_),
    .o1(_10621_));
 b15oai013aq1n04x5 _19284_ (.a(_10618_),
    .b(_10619_),
    .c(_10621_),
    .d(net518),
    .o1(_10622_));
 b15norp03aq1n02x5 _19285_ (.a(_09888_),
    .b(_09860_),
    .c(_10006_),
    .o1(_10623_));
 b15aoi112al1n03x5 _19286_ (.a(net509),
    .b(_10623_),
    .c(_10220_),
    .d(net514),
    .o1(_10624_));
 b15norp02an1n03x5 _19287_ (.a(_10127_),
    .b(_10211_),
    .o1(_10625_));
 b15oaoi13aq1n03x5 _19288_ (.a(net497),
    .b(_10126_),
    .c(_10128_),
    .d(_09892_),
    .o1(_10626_));
 b15oai112an1n12x5 _19289_ (.a(_09888_),
    .b(_10248_),
    .c(_10625_),
    .d(_10626_),
    .o1(_10627_));
 b15aoi022aq1n08x5 _19290_ (.a(net509),
    .b(_10622_),
    .c(_10624_),
    .d(_10627_),
    .o1(_10628_));
 b15nor004as1n12x5 _19291_ (.a(_10590_),
    .b(_10603_),
    .c(_10614_),
    .d(_10628_),
    .o1(_10629_));
 b15xor002as1n16x5 _19292_ (.a(\u0.w[0][14] ),
    .b(_10629_),
    .out0(_10630_));
 b15xor002an1n16x5 _19293_ (.a(\u0.w[1][14] ),
    .b(_10630_),
    .out0(_10631_));
 b15xor002as1n16x5 _19294_ (.a(\u0.w[2][14] ),
    .b(_10631_),
    .out0(_10632_));
 b15xor002ar1n02x5 _19295_ (.a(\u0.tmp_w[14] ),
    .b(_10632_),
    .out0(_10633_));
 b15mdn022ar1n02x5 _19296_ (.a(_10553_),
    .b(_10633_),
    .o1(_00358_),
    .sa(net943));
 b15zdnd11an1n04x5 FILLER_0_900 ();
 b15zdnd11an1n04x5 FILLER_0_891 ();
 b15zdnd00an1n01x5 FILLER_0_885 ();
 b15zdnd11an1n04x5 FILLER_0_881 ();
 b15oai022ar1n08x5 _19301_ (.a(net514),
    .b(_10221_),
    .c(_10319_),
    .d(_09994_),
    .o1(_10638_));
 b15nand03ar1n02x5 _19302_ (.a(net493),
    .b(_09868_),
    .c(_10638_),
    .o1(_10639_));
 b15aob012ar1n02x5 _19303_ (.a(_09940_),
    .b(_10102_),
    .c(_10283_),
    .out0(_10640_));
 b15oai112an1n04x5 _19304_ (.a(_10639_),
    .b(_10640_),
    .c(_10006_),
    .d(_10102_),
    .o1(_10641_));
 b15oai012ah1n03x5 _19305_ (.a(_10318_),
    .b(_10006_),
    .c(_10025_),
    .o1(_10642_));
 b15aoi012aq1n02x5 _19306_ (.a(net509),
    .b(_09962_),
    .c(_09892_),
    .o1(_10643_));
 b15nand04an1n08x5 _19307_ (.a(_09932_),
    .b(net510),
    .c(_09967_),
    .d(_09964_),
    .o1(_10644_));
 b15aoai13as1n08x5 _19308_ (.a(_10643_),
    .b(_09888_),
    .c(_10380_),
    .d(_10644_),
    .o1(_10645_));
 b15aoai13ah1n04x5 _19309_ (.a(net518),
    .b(_10641_),
    .c(_10642_),
    .d(_10645_),
    .o1(_10646_));
 b15nand04aq1n03x5 _19310_ (.a(net511),
    .b(net505),
    .c(_09880_),
    .d(_10107_),
    .o1(_10647_));
 b15oai112al1n06x5 _19311_ (.a(net508),
    .b(_10647_),
    .c(_10022_),
    .d(_10465_),
    .o1(_10648_));
 b15nand02ar1n02x5 _19312_ (.a(net520),
    .b(_10282_),
    .o1(_10649_));
 b15aoi012ar1n02x5 _19313_ (.a(_10180_),
    .b(_10649_),
    .c(_10024_),
    .o1(_10650_));
 b15orn002an1n02x5 _19314_ (.a(net514),
    .b(net497),
    .o(_10651_));
 b15aoi112an1n06x5 _19315_ (.a(_09887_),
    .b(_10128_),
    .c(_10651_),
    .d(_10221_),
    .o1(_10652_));
 b15oai013ar1n04x5 _19316_ (.a(_10648_),
    .b(_10650_),
    .c(_10652_),
    .d(net509),
    .o1(_10653_));
 b15oai022ar1n04x5 _19317_ (.a(_10206_),
    .b(_10165_),
    .c(_09985_),
    .d(_10117_),
    .o1(_10654_));
 b15nandp2ar1n02x5 _19318_ (.a(_09892_),
    .b(_10654_),
    .o1(_10655_));
 b15aoi022al1n02x5 _19319_ (.a(_09897_),
    .b(_09916_),
    .c(_10015_),
    .d(_10213_),
    .o1(_10656_));
 b15oai012an1n06x5 _19320_ (.a(_10655_),
    .b(_10656_),
    .c(_09892_),
    .o1(_10657_));
 b15aoai13ar1n02x5 _19321_ (.a(net509),
    .b(net514),
    .c(net512),
    .d(_10054_),
    .o1(_10658_));
 b15aoi012ar1n02x5 _19322_ (.a(_10164_),
    .b(_10235_),
    .c(_09977_),
    .o1(_10659_));
 b15aoi012an1n02x5 _19323_ (.a(_10658_),
    .b(_10659_),
    .c(net514),
    .o1(_10660_));
 b15nonb03aq1n04x5 _19324_ (.a(_10653_),
    .b(_10657_),
    .c(_10660_),
    .out0(_10661_));
 b15nandp3al1n02x5 _19325_ (.a(_10032_),
    .b(_09992_),
    .c(_10213_),
    .o1(_10662_));
 b15oaoi13al1n02x5 _19326_ (.a(net511),
    .b(_10662_),
    .c(_10069_),
    .d(net514),
    .o1(_10663_));
 b15aob012aq1n02x5 _19327_ (.a(_10038_),
    .b(_10220_),
    .c(_10336_),
    .out0(_10664_));
 b15oai012an1n03x5 _19328_ (.a(_10217_),
    .b(_09953_),
    .c(net514),
    .o1(_10665_));
 b15oai012an1n02x5 _19329_ (.a(_09953_),
    .b(_09990_),
    .c(net514),
    .o1(_10666_));
 b15aoi013ah1n03x5 _19330_ (.a(_10663_),
    .b(_10664_),
    .c(_10665_),
    .d(_10666_),
    .o1(_10667_));
 b15oaoi13an1n04x5 _19331_ (.a(_10282_),
    .b(_10426_),
    .c(_09990_),
    .d(_10038_),
    .o1(_10668_));
 b15aoai13al1n06x5 _19332_ (.a(_09880_),
    .b(_10100_),
    .c(net512),
    .d(_09901_),
    .o1(_10669_));
 b15oai013as1n08x5 _19333_ (.a(_10580_),
    .b(_10669_),
    .c(net507),
    .d(_10003_),
    .o1(_10670_));
 b15oai012as1n04x5 _19334_ (.a(_10154_),
    .b(_10110_),
    .c(_09887_),
    .o1(_10671_));
 b15and003an1n04x5 _19335_ (.a(_09938_),
    .b(_09916_),
    .c(_10671_),
    .o(_10672_));
 b15nandp3ar1n02x5 _19336_ (.a(_09867_),
    .b(_09868_),
    .c(_09940_),
    .o1(_10673_));
 b15aoi022ar1n02x5 _19337_ (.a(_10032_),
    .b(_09899_),
    .c(_09964_),
    .d(_10038_),
    .o1(_10674_));
 b15oai013aq1n04x5 _19338_ (.a(_10673_),
    .b(_10674_),
    .c(_10043_),
    .d(_10248_),
    .o1(_10675_));
 b15nor004ah1n08x5 _19339_ (.a(_10668_),
    .b(_10670_),
    .c(_10672_),
    .d(_10675_),
    .o1(_10676_));
 b15oai022an1n02x5 _19340_ (.a(_09994_),
    .b(_10102_),
    .c(_10283_),
    .d(_09905_),
    .o1(_10677_));
 b15aoi013ah1n02x5 _19341_ (.a(_09888_),
    .b(net508),
    .c(_10015_),
    .d(_10238_),
    .o1(_10678_));
 b15nand03ah1n06x5 _19342_ (.a(_10481_),
    .b(_10108_),
    .c(_10678_),
    .o1(_10679_));
 b15norp02aq1n02x5 _19343_ (.a(_10571_),
    .b(_10117_),
    .o1(_10680_));
 b15oai022as1n06x5 _19344_ (.a(net520),
    .b(_10677_),
    .c(_10679_),
    .d(_10680_),
    .o1(_10681_));
 b15norp03ar1n04x5 _19345_ (.a(_09980_),
    .b(_09914_),
    .c(_10332_),
    .o1(_10682_));
 b15aoai13aq1n08x5 _19346_ (.a(net514),
    .b(_10682_),
    .c(_10588_),
    .d(_09921_),
    .o1(_10683_));
 b15nand04aq1n16x5 _19347_ (.a(_10667_),
    .b(_10676_),
    .c(_10681_),
    .d(_10683_),
    .o1(_10684_));
 b15oai022ar1n02x5 _19348_ (.a(net514),
    .b(_10223_),
    .c(_10017_),
    .d(_10211_),
    .o1(_10685_));
 b15oaoi13ar1n02x5 _19349_ (.a(net518),
    .b(_10223_),
    .c(_10211_),
    .d(net514),
    .o1(_10686_));
 b15oab012al1n06x5 _19350_ (.a(_10319_),
    .b(_10685_),
    .c(_10686_),
    .out0(_10687_));
 b15aoi012ar1n02x5 _19351_ (.a(_10100_),
    .b(_10181_),
    .c(_09901_),
    .o1(_10688_));
 b15oai012ah1n04x5 _19352_ (.a(net509),
    .b(_10230_),
    .c(_10688_),
    .o1(_10689_));
 b15oai122ah1n12x5 _19353_ (.a(net512),
    .b(net509),
    .c(_10166_),
    .d(_10687_),
    .e(_10689_),
    .o1(_10690_));
 b15norp02ar1n02x5 _19354_ (.a(_10282_),
    .b(_10025_),
    .o1(_10691_));
 b15aoi013al1n02x5 _19355_ (.a(_10691_),
    .b(_10332_),
    .c(_10031_),
    .d(_09978_),
    .o1(_10692_));
 b15aoi013as1n03x5 _19356_ (.a(_10038_),
    .b(_09858_),
    .c(_10282_),
    .d(_10049_),
    .o1(_10693_));
 b15aob012aq1n04x5 _19357_ (.a(_10645_),
    .b(_10692_),
    .c(_10693_),
    .out0(_10694_));
 b15nanb02an1n03x5 _19358_ (.a(net512),
    .b(net499),
    .out0(_10695_));
 b15oaoi13as1n08x5 _19359_ (.a(_10695_),
    .b(_10042_),
    .c(_10091_),
    .d(_10211_),
    .o1(_10696_));
 b15oai022ah1n02x5 _19360_ (.a(_09980_),
    .b(_09914_),
    .c(_10587_),
    .d(_10372_),
    .o1(_10697_));
 b15aoi012al1n06x5 _19361_ (.a(_10696_),
    .b(_10697_),
    .c(_09892_),
    .o1(_10698_));
 b15aob012ar1n02x5 _19362_ (.a(_09888_),
    .b(_09918_),
    .c(_10696_),
    .out0(_10699_));
 b15aoai13an1n06x5 _19363_ (.a(_10699_),
    .b(_09932_),
    .c(_10206_),
    .d(_10696_),
    .o1(_10700_));
 b15oai112as1n16x5 _19364_ (.a(_10690_),
    .b(_10694_),
    .c(_10698_),
    .d(_10700_),
    .o1(_10701_));
 b15nano23as1n24x5 _19365_ (.a(_10646_),
    .b(_10661_),
    .c(_10684_),
    .d(_10701_),
    .out0(_10702_));
 b15xor002as1n16x5 _19366_ (.a(\u0.w[0][15] ),
    .b(_10702_),
    .out0(_10703_));
 b15xor002ah1n16x5 _19367_ (.a(\u0.w[1][15] ),
    .b(_10703_),
    .out0(_10704_));
 b15xor002as1n16x5 _19368_ (.a(\u0.w[2][15] ),
    .b(_10704_),
    .out0(_10705_));
 b15nanb03ar1n02x5 _19369_ (.a(net943),
    .b(\u0.tmp_w[15] ),
    .c(_10705_),
    .out0(_10706_));
 b15orn003ar1n02x5 _19370_ (.a(net943),
    .b(\u0.tmp_w[15] ),
    .c(_10705_),
    .o(_10707_));
 b15zdnd11an1n32x5 FILLER_0_849 ();
 b15nand02ar1n02x5 _19372_ (.a(net943),
    .b(net35),
    .o1(_10709_));
 b15nand03al1n03x5 _19373_ (.a(_10706_),
    .b(_10707_),
    .c(_10709_),
    .o1(_00359_));
 b15inv040ah1n02x5 _19374_ (.a(net36),
    .o1(_10710_));
 b15zdnd11an1n04x5 FILLER_0_839 ();
 b15zdnd11an1n08x5 FILLER_0_831 ();
 b15zdnd11an1n04x5 FILLER_0_823 ();
 b15zdnd11an1n04x5 FILLER_0_814 ();
 b15zdnd11an1n08x5 FILLER_0_806 ();
 b15zdnd11an1n16x5 FILLER_0_790 ();
 b15zdnd11an1n64x5 FILLER_0_726 ();
 b15and002ar1n24x5 _19382_ (.a(net473),
    .b(net469),
    .o(_10718_));
 b15zdnd00an1n02x5 FILLER_0_716 ();
 b15nonb02as1n16x5 _19384_ (.a(net466),
    .b(net462),
    .out0(_10720_));
 b15nandp2as1n32x5 _19385_ (.a(_10718_),
    .b(_10720_),
    .o1(_10721_));
 b15zdnd11an1n04x5 FILLER_0_712 ();
 b15nand02al1n16x5 _19387_ (.a(net486),
    .b(net480),
    .o1(_10723_));
 b15nonb02as1n16x5 _19388_ (.a(net473),
    .b(net469),
    .out0(_10724_));
 b15norp02ah1n48x5 _19389_ (.a(net468),
    .b(net463),
    .o1(_10725_));
 b15nandp2as1n24x5 _19390_ (.a(_10724_),
    .b(_10725_),
    .o1(_10726_));
 b15zdnd11an1n64x5 FILLER_0_648 ();
 b15inv000an1n56x5 _19392_ (.a(net482),
    .o1(_10728_));
 b15nand02al1n16x5 _19393_ (.a(net485),
    .b(_10728_),
    .o1(_10729_));
 b15oai022ar1n02x5 _19394_ (.a(_10721_),
    .b(_10723_),
    .c(_10726_),
    .d(_10729_),
    .o1(_10730_));
 b15norp02aq1n02x5 _19395_ (.a(net476),
    .b(_10730_),
    .o1(_10731_));
 b15inv020as1n80x5 _19396_ (.a(net489),
    .o1(_10732_));
 b15zdnd11an1n64x5 FILLER_0_584 ();
 b15zdnd11an1n64x5 FILLER_0_520 ();
 b15zdnd11an1n64x5 FILLER_0_456 ();
 b15zdnd11an1n64x5 FILLER_0_392 ();
 b15zdnd11an1n64x5 FILLER_0_328 ();
 b15nona23an1n32x5 _19402_ (.a(net473),
    .b(net467),
    .c(net465),
    .d(net472),
    .out0(_10738_));
 b15zdnd11an1n64x5 FILLER_0_264 ();
 b15nonb02as1n16x5 _19404_ (.a(\u0.tmp_w[9] ),
    .b(net479),
    .out0(_10740_));
 b15norp03an1n02x5 _19405_ (.a(_10732_),
    .b(_10738_),
    .c(_10740_),
    .o1(_10741_));
 b15nano23aq1n24x5 _19406_ (.a(net472),
    .b(net467),
    .c(net465),
    .d(\u0.tmp_w[12] ),
    .out0(_10742_));
 b15zdnd11an1n64x5 FILLER_0_200 ();
 b15zdnd11an1n64x5 FILLER_0_136 ();
 b15nonb02as1n16x5 _19409_ (.a(net485),
    .b(net489),
    .out0(_10745_));
 b15zdnd11an1n64x5 FILLER_0_72 ();
 b15zdnd11an1n64x5 FILLER_0_8 ();
 b15aoi013ar1n04x5 _19412_ (.a(_10741_),
    .b(_10742_),
    .c(_10745_),
    .d(net481),
    .o1(_10748_));
 b15cbf000an1n16x5 clkbuf_opt_1_1_clk (.clk(clknet_opt_1_0_clk),
    .clkout(clknet_opt_1_1_clk));
 b15nor004as1n12x5 _19414_ (.a(net473),
    .b(net472),
    .c(net467),
    .d(net465),
    .o1(_10750_));
 b15nand02ar1n02x5 _19415_ (.a(_10740_),
    .b(_10750_),
    .o1(_10751_));
 b15cbf000an1n16x5 clkbuf_opt_1_0_clk (.clk(clknet_1_1__leaf_clk),
    .clkout(clknet_opt_1_0_clk));
 b15cbf000an1n16x5 clkbuf_1_1__f_clk (.clk(clknet_0_clk),
    .clkout(clknet_1_1__leaf_clk));
 b15norp02ar1n32x5 _19418_ (.a(net473),
    .b(net469),
    .o1(_10754_));
 b15nanb02as1n24x5 _19419_ (.a(net463),
    .b(net468),
    .out0(_10755_));
 b15and002al1n08x5 _19420_ (.a(net483),
    .b(net480),
    .o(_10756_));
 b15oai112al1n06x5 _19421_ (.a(_10754_),
    .b(_10755_),
    .c(_10756_),
    .d(net486),
    .o1(_10757_));
 b15inv000aq1n20x5 _19422_ (.a(net468),
    .o1(_10758_));
 b15nandp2an1n32x5 _19423_ (.a(net487),
    .b(net484),
    .o1(_10759_));
 b15oaoi13al1n02x5 _19424_ (.a(_10728_),
    .b(_10758_),
    .c(net462),
    .d(_10759_),
    .o1(_10760_));
 b15oai012as1n04x5 _19425_ (.a(_10751_),
    .b(_10757_),
    .c(_10760_),
    .o1(_10761_));
 b15cbf000an1n16x5 clkbuf_1_0__f_clk (.clk(clknet_0_clk),
    .clkout(clknet_1_0__leaf_clk));
 b15cbf000an1n16x5 clkbuf_0_clk (.clk(clk),
    .clkout(clknet_0_clk));
 b15nano22ar1n02x5 _19428_ (.a(net469),
    .b(net462),
    .c(net480),
    .out0(_10764_));
 b15nor002al1n24x5 _19429_ (.a(net470),
    .b(net463),
    .o1(_10765_));
 b15nanb02as1n24x5 _19430_ (.a(net485),
    .b(net482),
    .out0(_10766_));
 b15aoi013an1n04x5 _19431_ (.a(_10764_),
    .b(_10765_),
    .c(net486),
    .d(_10766_),
    .o1(_10767_));
 b15orn002ar1n08x5 _19432_ (.a(net486),
    .b(net483),
    .o(_10768_));
 b15and002al1n04x5 _19433_ (.a(_10723_),
    .b(_10768_),
    .o(_10769_));
 b15nand02al1n06x5 _19434_ (.a(net469),
    .b(_10725_),
    .o1(_10770_));
 b15cbf000an1n16x5 clkbuf_leaf_18_clk (.clk(clknet_1_0__leaf_clk),
    .clkout(clknet_leaf_18_clk));
 b15cbf000an1n16x5 clkbuf_leaf_17_clk (.clk(clknet_1_0__leaf_clk),
    .clkout(clknet_leaf_17_clk));
 b15nonb02as1n04x5 _19437_ (.a(net483),
    .b(net466),
    .out0(_10773_));
 b15nand03al1n12x5 _19438_ (.a(net480),
    .b(net462),
    .c(_10773_),
    .o1(_10774_));
 b15cbf000an1n16x5 clkbuf_leaf_16_clk (.clk(clknet_1_0__leaf_clk),
    .clkout(clknet_leaf_16_clk));
 b15oai222ah1n16x5 _19440_ (.a(_10758_),
    .b(_10767_),
    .c(_10769_),
    .d(_10770_),
    .e(_10774_),
    .f(net469),
    .o1(_10776_));
 b15aoi012ar1n12x5 _19441_ (.a(_10761_),
    .b(_10776_),
    .c(net473),
    .o1(_10777_));
 b15aoi013al1n06x5 _19442_ (.a(_10731_),
    .b(_10748_),
    .c(_10777_),
    .d(\u0.tmp_w[11] ),
    .o1(_10778_));
 b15cbf000an1n16x5 clkbuf_leaf_15_clk (.clk(clknet_1_0__leaf_clk),
    .clkout(clknet_leaf_15_clk));
 b15cbf000an1n16x5 clkbuf_leaf_14_clk (.clk(clknet_1_0__leaf_clk),
    .clkout(clknet_leaf_14_clk));
 b15orn002al1n08x5 _19445_ (.a(net480),
    .b(net463),
    .o(_10781_));
 b15cbf000an1n16x5 clkbuf_leaf_13_clk (.clk(clknet_1_0__leaf_clk),
    .clkout(clknet_leaf_13_clk));
 b15nand02al1n12x5 _19447_ (.a(net490),
    .b(net475),
    .o1(_10783_));
 b15cbf000an1n16x5 clkbuf_leaf_12_clk (.clk(clknet_1_0__leaf_clk),
    .clkout(clknet_leaf_12_clk));
 b15nandp2ah1n08x5 _19449_ (.a(net472),
    .b(net467),
    .o1(_10785_));
 b15nand02ah1n32x5 _19450_ (.a(net484),
    .b(net477),
    .o1(_10786_));
 b15orn002ah1n08x5 _19451_ (.a(net472),
    .b(net467),
    .o(_10787_));
 b15oai022ar1n02x5 _19452_ (.a(net477),
    .b(_10785_),
    .c(_10786_),
    .d(_10787_),
    .o1(_10788_));
 b15nanb02ar1n03x5 _19453_ (.a(_10783_),
    .b(_10788_),
    .out0(_10789_));
 b15cbf000an1n16x5 clkbuf_leaf_11_clk (.clk(clknet_1_0__leaf_clk),
    .clkout(clknet_leaf_11_clk));
 b15cbf000an1n16x5 clkbuf_leaf_10_clk (.clk(clknet_1_1__leaf_clk),
    .clkout(clknet_leaf_10_clk));
 b15nanb02aq1n12x5 _19456_ (.a(net474),
    .b(net490),
    .out0(_10792_));
 b15nanb02ar1n02x5 _19457_ (.a(net487),
    .b(net474),
    .out0(_10793_));
 b15oai022ar1n04x5 _19458_ (.a(_10785_),
    .b(_10792_),
    .c(_10793_),
    .d(_10787_),
    .o1(_10794_));
 b15nanb02al1n16x5 _19459_ (.a(net466),
    .b(net474),
    .out0(_10795_));
 b15nonb02ah1n04x5 _19460_ (.a(net466),
    .b(net474),
    .out0(_10796_));
 b15nanb02ah1n03x5 _19461_ (.a(net477),
    .b(net469),
    .out0(_10797_));
 b15norp02ar1n02x5 _19462_ (.a(_10796_),
    .b(_10797_),
    .o1(_10798_));
 b15aoi022ah1n04x5 _19463_ (.a(net477),
    .b(_10794_),
    .c(_10795_),
    .d(_10798_),
    .o1(_10799_));
 b15cbf000an1n16x5 clkbuf_leaf_9_clk (.clk(clknet_1_1__leaf_clk),
    .clkout(clknet_leaf_9_clk));
 b15cbf000an1n16x5 clkbuf_leaf_8_clk (.clk(clknet_1_1__leaf_clk),
    .clkout(clknet_leaf_8_clk));
 b15oaoi13aq1n08x5 _19466_ (.a(_10781_),
    .b(_10789_),
    .c(_10799_),
    .d(net483),
    .o1(_10802_));
 b15cbf000an1n16x5 clkbuf_leaf_7_clk (.clk(clknet_1_1__leaf_clk),
    .clkout(clknet_leaf_7_clk));
 b15nanb02as1n24x5 _19468_ (.a(net473),
    .b(net469),
    .out0(_10804_));
 b15orn002ah1n16x5 _19469_ (.a(net466),
    .b(net462),
    .o(_10805_));
 b15nandp2ar1n24x5 _19470_ (.a(net480),
    .b(net478),
    .o1(_10806_));
 b15norp03ar1n02x5 _19471_ (.a(_10804_),
    .b(_10805_),
    .c(_10806_),
    .o1(_10807_));
 b15orn002aq1n24x5 _19472_ (.a(net482),
    .b(net478),
    .o(_10808_));
 b15norp02as1n04x5 _19473_ (.a(_10732_),
    .b(_10808_),
    .o1(_10809_));
 b15nandp2as1n16x5 _19474_ (.a(net467),
    .b(net465),
    .o1(_10810_));
 b15nor002ar1n12x5 _19475_ (.a(_10810_),
    .b(_10804_),
    .o1(_10811_));
 b15aoai13ar1n02x5 _19476_ (.a(net483),
    .b(_10807_),
    .c(_10809_),
    .d(_10811_),
    .o1(_10812_));
 b15nanb02as1n24x5 _19477_ (.a(net486),
    .b(net483),
    .out0(_10813_));
 b15cbf000an1n16x5 clkbuf_leaf_6_clk (.clk(clknet_1_1__leaf_clk),
    .clkout(clknet_leaf_6_clk));
 b15orn003al1n16x5 _19479_ (.a(net471),
    .b(net468),
    .c(net463),
    .o(_10815_));
 b15orn002al1n08x5 _19480_ (.a(net476),
    .b(net474),
    .o(_10816_));
 b15orn002ah1n03x5 _19481_ (.a(net488),
    .b(net480),
    .o(_10817_));
 b15nor003as1n02x5 _19482_ (.a(_10815_),
    .b(_10816_),
    .c(_10817_),
    .o1(_10818_));
 b15nano23as1n24x5 _19483_ (.a(net473),
    .b(net466),
    .c(net462),
    .d(net469),
    .out0(_10819_));
 b15norp02as1n24x5 _19484_ (.a(net479),
    .b(net476),
    .o1(_10820_));
 b15aoai13ar1n08x5 _19485_ (.a(_10813_),
    .b(_10818_),
    .c(_10819_),
    .d(_10820_),
    .o1(_10821_));
 b15nano23as1n24x5 _19486_ (.a(net473),
    .b(net471),
    .c(net467),
    .d(net465),
    .out0(_10822_));
 b15cbf000an1n16x5 clkbuf_leaf_5_clk (.clk(clknet_1_1__leaf_clk),
    .clkout(clknet_leaf_5_clk));
 b15norp02ah1n32x5 _19488_ (.a(net490),
    .b(\u0.tmp_w[9] ),
    .o1(_10824_));
 b15norp02ar1n02x5 _19489_ (.a(_10808_),
    .b(_10824_),
    .o1(_10825_));
 b15orn002as1n03x5 _19490_ (.a(net485),
    .b(net477),
    .o(_10826_));
 b15aoi012ar1n06x5 _19491_ (.a(_10826_),
    .b(net481),
    .c(net488),
    .o1(_10827_));
 b15orn002ah1n32x5 _19492_ (.a(net475),
    .b(net470),
    .o(_10828_));
 b15nor002ar1n06x5 _19493_ (.a(_10828_),
    .b(_10755_),
    .o1(_10829_));
 b15aoi022ar1n02x5 _19494_ (.a(_10822_),
    .b(_10825_),
    .c(_10827_),
    .d(_10829_),
    .o1(_10830_));
 b15nonb02aq1n16x5 _19495_ (.a(net487),
    .b(net483),
    .out0(_10831_));
 b15nor002as1n02x5 _19496_ (.a(net480),
    .b(_10831_),
    .o1(_10832_));
 b15nonb02as1n16x5 _19497_ (.a(net475),
    .b(net476),
    .out0(_10833_));
 b15nano22as1n24x5 _19498_ (.a(net472),
    .b(net465),
    .c(net467),
    .out0(_10834_));
 b15and002ah1n04x5 _19499_ (.a(_10833_),
    .b(_10834_),
    .o(_10835_));
 b15cbf000an1n16x5 clkbuf_leaf_4_clk (.clk(clknet_1_1__leaf_clk),
    .clkout(clknet_leaf_4_clk));
 b15and003ar1n02x5 _19501_ (.a(net477),
    .b(_10742_),
    .c(_10813_),
    .o(_10837_));
 b15oai012ah1n03x5 _19502_ (.a(_10832_),
    .b(_10835_),
    .c(_10837_),
    .o1(_10838_));
 b15nand04aq1n03x5 _19503_ (.a(_10812_),
    .b(_10821_),
    .c(_10830_),
    .d(_10838_),
    .o1(_10839_));
 b15nand04as1n16x5 _19504_ (.a(\u0.tmp_w[12] ),
    .b(net472),
    .c(net467),
    .d(net465),
    .o1(_10840_));
 b15nor002ah1n02x5 _19505_ (.a(_10840_),
    .b(_10786_),
    .o1(_10841_));
 b15norp03ar1n02x5 _19506_ (.a(_10808_),
    .b(_10804_),
    .c(_10805_),
    .o1(_10842_));
 b15oab012aq1n03x5 _19507_ (.a(net488),
    .b(_10841_),
    .c(_10842_),
    .out0(_10843_));
 b15cbf000an1n16x5 clkbuf_leaf_3_clk (.clk(clknet_opt_1_1_clk),
    .clkout(clknet_leaf_3_clk));
 b15nanb03an1n12x5 _19509_ (.a(net485),
    .b(net482),
    .c(net478),
    .out0(_10845_));
 b15aoi012an1n06x5 _19510_ (.a(net488),
    .b(_10808_),
    .c(_10845_),
    .o1(_10846_));
 b15and002as1n32x5 _19511_ (.a(net466),
    .b(net462),
    .o(_10847_));
 b15nandp3as1n04x5 _19512_ (.a(net488),
    .b(net485),
    .c(net482),
    .o1(_10848_));
 b15nand04ar1n06x5 _19513_ (.a(net478),
    .b(_10847_),
    .c(_10724_),
    .d(_10848_),
    .o1(_10849_));
 b15nonb02as1n16x5 _19514_ (.a(net470),
    .b(net475),
    .out0(_10850_));
 b15nandp2al1n16x5 _19515_ (.a(_10850_),
    .b(_10720_),
    .o1(_10851_));
 b15oaoi13as1n04x5 _19516_ (.a(_10846_),
    .b(_10849_),
    .c(net478),
    .d(_10851_),
    .o1(_10852_));
 b15cbf000an1n16x5 clkbuf_leaf_2_clk (.clk(clknet_1_1__leaf_clk),
    .clkout(clknet_leaf_2_clk));
 b15nand03ar1n08x5 _19518_ (.a(net478),
    .b(_10720_),
    .c(_10848_),
    .o1(_10854_));
 b15aoai13ah1n06x5 _19519_ (.a(net482),
    .b(net485),
    .c(_10720_),
    .d(_10754_),
    .o1(_10855_));
 b15cbf000an1n16x5 clkbuf_leaf_1_clk (.clk(clknet_1_0__leaf_clk),
    .clkout(clknet_leaf_1_clk));
 b15cbf000an1n16x5 clkbuf_leaf_0_clk (.clk(clknet_1_0__leaf_clk),
    .clkout(clknet_leaf_0_clk));
 b15nandp2al1n16x5 _19522_ (.a(net482),
    .b(_10718_),
    .o1(_10858_));
 b15aoi122as1n08x5 _19523_ (.a(_10854_),
    .b(_10855_),
    .c(_10732_),
    .d(_10828_),
    .e(_10858_),
    .o1(_10859_));
 b15nonb02as1n16x5 _19524_ (.a(net485),
    .b(net478),
    .out0(_10860_));
 b15nor002as1n03x5 _19525_ (.a(\u0.tmp_w[12] ),
    .b(net467),
    .o1(_10861_));
 b15and003ar1n02x5 _19526_ (.a(net479),
    .b(net474),
    .c(net468),
    .o(_10862_));
 b15oai112aq1n08x5 _19527_ (.a(_10860_),
    .b(_10765_),
    .c(_10861_),
    .d(_10862_),
    .o1(_10863_));
 b15qgbna2an1n05x5 _19528_ (.o1(_10864_),
    .a(net489),
    .b(net476));
 b15orn002ah1n04x5 _19529_ (.a(_10785_),
    .b(_10864_),
    .o(_10865_));
 b15nonb02al1n12x5 _19530_ (.a(net475),
    .b(net464),
    .out0(_10866_));
 b15nonb02as1n08x5 _19531_ (.a(\u0.tmp_w[15] ),
    .b(net475),
    .out0(_10867_));
 b15aoi022aq1n08x5 _19532_ (.a(_10740_),
    .b(_10866_),
    .c(_10867_),
    .d(net479),
    .o1(_10868_));
 b15nonb02ah1n16x5 _19533_ (.a(net476),
    .b(net474),
    .out0(_10869_));
 b15bfn001as1n64x5 max_length948 (.a(net129),
    .o(net948));
 b15aoi012aq1n04x5 _19535_ (.a(_10869_),
    .b(_10833_),
    .c(net488),
    .o1(_10871_));
 b15nonb02as1n16x5 _19536_ (.a(net481),
    .b(net485),
    .out0(_10872_));
 b15nano22as1n12x5 _19537_ (.a(net468),
    .b(net463),
    .c(net471),
    .out0(_10873_));
 b15nand02ah1n04x5 _19538_ (.a(_10872_),
    .b(_10873_),
    .o1(_10874_));
 b15oai122as1n16x5 _19539_ (.a(_10863_),
    .b(_10865_),
    .c(_10868_),
    .d(_10871_),
    .e(_10874_),
    .o1(_10875_));
 b15nor004an1n12x5 _19540_ (.a(_10843_),
    .b(_10852_),
    .c(_10859_),
    .d(_10875_),
    .o1(_10876_));
 b15nanb02as1n24x5 _19541_ (.a(net468),
    .b(net463),
    .out0(_10877_));
 b15nonb02an1n16x5 _19542_ (.a(net477),
    .b(net479),
    .out0(_10878_));
 b15nand04an1n08x5 _19543_ (.a(_10850_),
    .b(_10877_),
    .c(_10755_),
    .d(_10878_),
    .o1(_10879_));
 b15nonb02aq1n16x5 _19544_ (.a(net475),
    .b(net479),
    .out0(_10880_));
 b15nonb02al1n12x5 _19545_ (.a(net463),
    .b(net470),
    .out0(_10881_));
 b15nonb02aq1n12x5 _19546_ (.a(net479),
    .b(net475),
    .out0(_10882_));
 b15nonb02aq1n08x5 _19547_ (.a(net470),
    .b(net463),
    .out0(_10883_));
 b15aoi022al1n04x5 _19548_ (.a(_10880_),
    .b(_10881_),
    .c(_10882_),
    .d(_10883_),
    .o1(_10884_));
 b15bfn001ah1n48x5 max_length947 (.a(net129),
    .o(net947));
 b15oai013aq1n06x5 _19550_ (.a(_10879_),
    .b(_10884_),
    .c(net477),
    .d(net466),
    .o1(_10886_));
 b15norp02ar1n03x5 _19551_ (.a(net484),
    .b(_10758_),
    .o1(_10887_));
 b15aoai13aq1n06x5 _19552_ (.a(net490),
    .b(_10887_),
    .c(_10879_),
    .d(net484),
    .o1(_10888_));
 b15orn002ar1n08x5 _19553_ (.a(net490),
    .b(net468),
    .o(_10889_));
 b15bfn001ah1n48x5 max_length946 (.a(net948),
    .o(net946));
 b15oai112as1n16x5 _19555_ (.a(_10886_),
    .b(_10888_),
    .c(_10889_),
    .d(net484),
    .o1(_10891_));
 b15nona23ah1n12x5 _19556_ (.a(_10802_),
    .b(_10839_),
    .c(_10876_),
    .d(_10891_),
    .out0(_10892_));
 b15inv040ah1n36x5 _19557_ (.a(net484),
    .o1(_10893_));
 b15bfn001ah1n48x5 wire945 (.a(net946),
    .o(net945));
 b15bfn001as1n32x5 wire944 (.a(net945),
    .o(net944));
 b15norp02as1n03x5 _19560_ (.a(net471),
    .b(_10805_),
    .o1(_10896_));
 b15aoai13aq1n03x5 _19561_ (.a(_10893_),
    .b(_10811_),
    .c(_10896_),
    .d(net488),
    .o1(_10897_));
 b15nandp3ah1n16x5 _19562_ (.a(net475),
    .b(net470),
    .c(net463),
    .o1(_10898_));
 b15orn002ah1n04x5 _19563_ (.a(net471),
    .b(net464),
    .o(_10899_));
 b15oai012al1n02x5 _19564_ (.a(_10898_),
    .b(_10899_),
    .c(\u0.tmp_w[12] ),
    .o1(_10900_));
 b15aoi022as1n04x5 _19565_ (.a(_10745_),
    .b(_10866_),
    .c(_10900_),
    .d(net487),
    .o1(_10901_));
 b15oaoi13ar1n08x5 _19566_ (.a(net476),
    .b(_10897_),
    .c(_10901_),
    .d(net467),
    .o1(_10902_));
 b15nand02an1n32x5 _19567_ (.a(net474),
    .b(net469),
    .o1(_10903_));
 b15nor002aq1n06x5 _19568_ (.a(_10877_),
    .b(_10903_),
    .o1(_10904_));
 b15aoai13as1n08x5 _19569_ (.a(net481),
    .b(_10902_),
    .c(_10904_),
    .d(_10824_),
    .o1(_10905_));
 b15bfn001ah1n48x5 max_length943 (.a(net944),
    .o(net943));
 b15norp02ar1n03x5 _19571_ (.a(_10810_),
    .b(_10808_),
    .o1(_10907_));
 b15bfn001ah1n48x5 wire942 (.a(net946),
    .o(net942));
 b15norp02ar1n02x5 _19573_ (.a(net485),
    .b(_10804_),
    .o1(_10909_));
 b15bfn001as1n24x5 wire941 (.a(net942),
    .o(net941));
 b15aoai13as1n02x5 _19575_ (.a(_10907_),
    .b(_10909_),
    .c(_10724_),
    .d(net485),
    .o1(_10911_));
 b15nano23al1n24x5 _19576_ (.a(net472),
    .b(net465),
    .c(net467),
    .d(net473),
    .out0(_10912_));
 b15nano23as1n24x5 _19577_ (.a(net467),
    .b(net465),
    .c(\u0.tmp_w[12] ),
    .d(net472),
    .out0(_10913_));
 b15nonb03as1n12x5 _19578_ (.a(net485),
    .b(net482),
    .c(net478),
    .out0(_10914_));
 b15aoi022an1n02x5 _19579_ (.a(_10872_),
    .b(_10912_),
    .c(_10913_),
    .d(_10914_),
    .o1(_10915_));
 b15bfn001ah1n48x5 wire940 (.a(net942),
    .o(net940));
 b15aoi012ar1n02x5 _19581_ (.a(_10873_),
    .b(_10725_),
    .c(net471),
    .o1(_10917_));
 b15orn003as1n03x5 _19582_ (.a(net473),
    .b(_10917_),
    .c(_10806_),
    .o(_10918_));
 b15aoi013ar1n04x5 _19583_ (.a(net489),
    .b(_10911_),
    .c(_10915_),
    .d(_10918_),
    .o1(_10919_));
 b15nonb02ah1n16x5 _19584_ (.a(net462),
    .b(net466),
    .out0(_10920_));
 b15nandp2an1n24x5 _19585_ (.a(_10920_),
    .b(_10754_),
    .o1(_10921_));
 b15bfn001ah1n48x5 wire939 (.a(net940),
    .o(net939));
 b15aoi012an1n02x5 _19587_ (.a(\u0.tmp_w[11] ),
    .b(_10921_),
    .c(_10840_),
    .o1(_10923_));
 b15nor002an1n24x5 _19588_ (.a(net483),
    .b(net480),
    .o1(_10924_));
 b15aoi112as1n08x5 _19589_ (.a(net486),
    .b(_10756_),
    .c(_10924_),
    .d(_10921_),
    .o1(_10925_));
 b15bfn001ah1n48x5 wire938 (.a(net939),
    .o(net938));
 b15bfn001ah1n48x5 max_length937 (.a(net938),
    .o(net937));
 b15bfn000as1n32x5 wire936 (.a(net940),
    .o(net936));
 b15nor002al1n12x5 _19593_ (.a(_10877_),
    .b(_10828_),
    .o1(_10929_));
 b15nandp2al1n02x5 _19594_ (.a(net481),
    .b(_10929_),
    .o1(_10930_));
 b15bfn001as1n48x5 load_slew935 (.a(\us00.a[0] ),
    .o(net935));
 b15oaoi13al1n04x5 _19596_ (.a(_10732_),
    .b(_10930_),
    .c(_10840_),
    .d(net481),
    .o1(_10932_));
 b15oaoi13as1n08x5 _19597_ (.a(_10919_),
    .b(_10923_),
    .c(_10925_),
    .d(_10932_),
    .o1(_10933_));
 b15nona23as1n32x5 _19598_ (.a(_10778_),
    .b(_10892_),
    .c(_10905_),
    .d(_10933_),
    .out0(_10934_));
 b15xnr002ah1n08x5 _19599_ (.a(\u0.w[0][16] ),
    .b(_10934_),
    .out0(_10935_));
 b15xor002ah1n03x5 _19600_ (.a(\u0.w[1][16] ),
    .b(_10935_),
    .out0(_10936_));
 b15xor002aq1n02x5 _19601_ (.a(\u0.w[2][16] ),
    .b(_10936_),
    .out0(_10937_));
 b15xor002ar1n02x5 _19602_ (.a(\u0.tmp_w[16] ),
    .b(_10937_),
    .out0(_10938_));
 b15mdn022ar1n02x5 _19603_ (.a(_10710_),
    .b(_10938_),
    .o1(_00360_),
    .sa(net947));
 b15inv020ah1n64x5 _19604_ (.a(\u0.tmp_w[11] ),
    .o1(_10939_));
 b15bfn001as1n64x5 max_length934 (.a(net935),
    .o(net934));
 b15nonb02aq1n16x5 _19606_ (.a(net479),
    .b(net490),
    .out0(_10941_));
 b15nano22aq1n02x5 _19607_ (.a(\u0.tmp_w[12] ),
    .b(net465),
    .c(net467),
    .out0(_10942_));
 b15nand02ar1n02x5 _19608_ (.a(_10941_),
    .b(_10942_),
    .o1(_10943_));
 b15orn002ar1n12x5 _19609_ (.a(net479),
    .b(net475),
    .o(_10944_));
 b15oai112an1n04x5 _19610_ (.a(net472),
    .b(_10943_),
    .c(_10944_),
    .d(_10755_),
    .o1(_10945_));
 b15aoi012ar1n02x5 _19611_ (.a(net472),
    .b(_10725_),
    .c(_10880_),
    .o1(_10946_));
 b15nand02ar1n02x5 _19612_ (.a(net479),
    .b(_10867_),
    .o1(_10947_));
 b15aoai13ar1n02x5 _19613_ (.a(net490),
    .b(_10867_),
    .c(_10866_),
    .d(net479),
    .o1(_10948_));
 b15aoai13as1n02x5 _19614_ (.a(_10946_),
    .b(_10758_),
    .c(_10947_),
    .d(_10948_),
    .o1(_10949_));
 b15nand03as1n06x5 _19615_ (.a(net484),
    .b(_10945_),
    .c(_10949_),
    .o1(_10950_));
 b15bfn001ah1n64x5 max_length933 (.a(\us00.a[0] ),
    .o(net933));
 b15nandp2as1n24x5 _19617_ (.a(net483),
    .b(net482),
    .o1(_10952_));
 b15nandp3ar1n03x5 _19618_ (.a(net488),
    .b(_10952_),
    .c(_10904_),
    .o1(_10953_));
 b15bfn001as1n48x5 load_slew932 (.a(\us00.a[1] ),
    .o(net932));
 b15bfn001ah1n64x5 max_length931 (.a(\us00.a[1] ),
    .o(net931));
 b15bfn001ah1n64x5 wire930 (.a(\us00.a[1] ),
    .o(net930));
 b15nonb02ah1n16x5 _19622_ (.a(net468),
    .b(net470),
    .out0(_10957_));
 b15nandp3ar1n02x5 _19623_ (.a(\u0.tmp_w[12] ),
    .b(_10872_),
    .c(_10957_),
    .o1(_10958_));
 b15nor002an1n06x5 _19624_ (.a(net470),
    .b(net468),
    .o1(_10959_));
 b15and002an1n08x5 _19625_ (.a(net470),
    .b(net466),
    .o(_10960_));
 b15mdn022as1n02x5 _19626_ (.a(_10959_),
    .b(_10960_),
    .o1(_10961_),
    .sa(net474));
 b15oaoi13an1n02x5 _19627_ (.a(net464),
    .b(_10958_),
    .c(_10961_),
    .d(_10893_),
    .o1(_10962_));
 b15aoai13al1n04x5 _19628_ (.a(_10732_),
    .b(_10962_),
    .c(_10913_),
    .d(net479),
    .o1(_10963_));
 b15aoi013an1n03x5 _19629_ (.a(_10939_),
    .b(_10950_),
    .c(_10953_),
    .d(_10963_),
    .o1(_10964_));
 b15nanb03as1n08x5 _19630_ (.a(net468),
    .b(net463),
    .c(net471),
    .out0(_10965_));
 b15nandp2aq1n16x5 _19631_ (.a(net484),
    .b(net474),
    .o1(_10966_));
 b15orn002as1n02x5 _19632_ (.a(_10965_),
    .b(_10966_),
    .o(_10967_));
 b15nand03al1n12x5 _19633_ (.a(net480),
    .b(_10724_),
    .c(_10725_),
    .o1(_10968_));
 b15aoi012aq1n06x5 _19634_ (.a(net487),
    .b(_10967_),
    .c(_10968_),
    .o1(_10969_));
 b15nand02al1n02x5 _19635_ (.a(_10732_),
    .b(_10904_),
    .o1(_10970_));
 b15oaoi13al1n04x5 _19636_ (.a(net479),
    .b(_10970_),
    .c(_10726_),
    .d(\u0.tmp_w[9] ),
    .o1(_10971_));
 b15oaoi13as1n08x5 _19637_ (.a(_10964_),
    .b(_10939_),
    .c(_10969_),
    .d(_10971_),
    .o1(_10972_));
 b15bfn001ah1n64x5 load_slew929 (.a(\us00.a[2] ),
    .o(net929));
 b15nanb02as1n24x5 _19639_ (.a(net482),
    .b(net478),
    .out0(_10974_));
 b15bfn001as1n48x5 wire928 (.a(net929),
    .o(net928));
 b15oai022ar1n02x5 _19641_ (.a(\u0.tmp_w[11] ),
    .b(_10738_),
    .c(_10921_),
    .d(_10974_),
    .o1(_10976_));
 b15nand02al1n02x5 _19642_ (.a(_10893_),
    .b(_10976_),
    .o1(_10977_));
 b15nand02al1n02x5 _19643_ (.a(net478),
    .b(_10929_),
    .o1(_10978_));
 b15oai112ah1n02x5 _19644_ (.a(net489),
    .b(_10977_),
    .c(_10978_),
    .d(_10952_),
    .o1(_10979_));
 b15bfn001ah1n64x5 wire927 (.a(\us00.a[2] ),
    .o(net927));
 b15nanb02ah1n24x5 _19646_ (.a(net476),
    .b(net484),
    .out0(_10981_));
 b15nand03ar1n02x5 _19647_ (.a(_10728_),
    .b(_10981_),
    .c(_10819_),
    .o1(_10982_));
 b15nand03ah1n08x5 _19648_ (.a(net478),
    .b(_10847_),
    .c(_10724_),
    .o1(_10983_));
 b15oai112an1n04x5 _19649_ (.a(_10732_),
    .b(_10982_),
    .c(_10983_),
    .d(_10766_),
    .o1(_10984_));
 b15nandp2ar1n05x5 _19650_ (.a(_10979_),
    .b(_10984_),
    .o1(_10985_));
 b15bfn001as1n48x5 load_slew926 (.a(\us00.a[3] ),
    .o(net926));
 b15nand02ar1n02x5 _19652_ (.a(net485),
    .b(_10750_),
    .o1(_10987_));
 b15nano23as1n24x5 _19653_ (.a(net473),
    .b(net465),
    .c(net467),
    .d(net472),
    .out0(_10988_));
 b15nand02ar1n02x5 _19654_ (.a(_10893_),
    .b(_10988_),
    .o1(_10989_));
 b15oai012ar1n02x5 _19655_ (.a(net482),
    .b(_10750_),
    .c(_10988_),
    .o1(_10990_));
 b15nand04aq1n03x5 _19656_ (.a(\u0.tmp_w[11] ),
    .b(_10987_),
    .c(_10989_),
    .d(_10990_),
    .o1(_10991_));
 b15nanb02as1n24x5 _19657_ (.a(net481),
    .b(net489),
    .out0(_10992_));
 b15nona23as1n32x5 _19658_ (.a(net469),
    .b(net466),
    .c(net462),
    .d(net473),
    .out0(_10993_));
 b15norp03an1n04x5 _19659_ (.a(_10766_),
    .b(_10903_),
    .c(_10755_),
    .o1(_10994_));
 b15aoi012ar1n06x5 _19660_ (.a(_10994_),
    .b(_10988_),
    .c(_10740_),
    .o1(_10995_));
 b15oai222as1n08x5 _19661_ (.a(_10721_),
    .b(_10992_),
    .c(_10993_),
    .d(_10766_),
    .e(net489),
    .f(_10995_),
    .o1(_10996_));
 b15oai012an1n06x5 _19662_ (.a(_10991_),
    .b(_10996_),
    .c(net478),
    .o1(_10997_));
 b15nand02ar1n24x5 _19663_ (.a(_10724_),
    .b(_10720_),
    .o1(_10998_));
 b15bfn001as1n64x5 max_length925 (.a(\us00.a[3] ),
    .o(net925));
 b15oaoi13ar1n08x5 _19665_ (.a(_10723_),
    .b(_10983_),
    .c(_10998_),
    .d(net477),
    .o1(_11000_));
 b15aoi022al1n02x5 _19666_ (.a(_10725_),
    .b(_10880_),
    .c(_10941_),
    .d(_10847_),
    .o1(_11001_));
 b15nor002as1n04x5 _19667_ (.a(_10797_),
    .b(_11001_),
    .o1(_11002_));
 b15bfn001as1n64x5 max_length924 (.a(\us00.a[3] ),
    .o(net924));
 b15nand02an1n24x5 _19669_ (.a(_10847_),
    .b(_10724_),
    .o1(_11004_));
 b15nor003aq1n06x5 _19670_ (.a(net486),
    .b(_10974_),
    .c(_11004_),
    .o1(_11005_));
 b15oai013as1n04x5 _19671_ (.a(net483),
    .b(_11000_),
    .c(_11002_),
    .d(_11005_),
    .o1(_11006_));
 b15and002an1n02x5 _19672_ (.a(_10873_),
    .b(_10833_),
    .o(_11007_));
 b15oai012ah1n02x5 _19673_ (.a(net486),
    .b(_10841_),
    .c(_11007_),
    .o1(_11008_));
 b15nanb02as1n24x5 _19674_ (.a(net478),
    .b(net482),
    .out0(_11009_));
 b15nanb02as1n12x5 _19675_ (.a(net464),
    .b(net470),
    .out0(_11010_));
 b15norp02aq1n03x5 _19676_ (.a(net487),
    .b(_11010_),
    .o1(_11011_));
 b15aoai13as1n08x5 _19677_ (.a(_10796_),
    .b(_11011_),
    .c(_10881_),
    .d(net487),
    .o1(_11012_));
 b15oaoi13aq1n04x5 _19678_ (.a(_11009_),
    .b(_11012_),
    .c(_10921_),
    .d(_10745_),
    .o1(_11013_));
 b15bfn001ah1n64x5 max_length923 (.a(\us00.a[4] ),
    .o(net923));
 b15aoai13al1n06x5 _19680_ (.a(_10809_),
    .b(_10822_),
    .c(net485),
    .d(_10913_),
    .o1(_11015_));
 b15inv000ar1n03x5 _19681_ (.a(_10848_),
    .o1(_11016_));
 b15nand02al1n32x5 _19682_ (.a(_10754_),
    .b(_10720_),
    .o1(_11017_));
 b15oai013al1n08x5 _19683_ (.a(_11015_),
    .b(_11016_),
    .c(_10846_),
    .d(_11017_),
    .o1(_11018_));
 b15nano23ah1n08x5 _19684_ (.a(_11006_),
    .b(_11008_),
    .c(_11013_),
    .d(_11018_),
    .out0(_11019_));
 b15nor002ar1n06x5 _19685_ (.a(net476),
    .b(\u0.tmp_w[12] ),
    .o1(_11020_));
 b15aoi013an1n03x5 _19686_ (.a(net484),
    .b(net472),
    .c(_10725_),
    .d(_11020_),
    .o1(_11021_));
 b15nandp2aq1n02x5 _19687_ (.a(_10725_),
    .b(_11020_),
    .o1(_11022_));
 b15oaoi13as1n08x5 _19688_ (.a(_11021_),
    .b(_11022_),
    .c(_10721_),
    .d(_10974_),
    .o1(_11023_));
 b15oab012an1n04x5 _19689_ (.a(_11023_),
    .b(_10978_),
    .c(_10729_),
    .out0(_11024_));
 b15oai112as1n16x5 _19690_ (.a(_10997_),
    .b(_11019_),
    .c(_11024_),
    .d(net489),
    .o1(_11025_));
 b15nandp2as1n02x5 _19691_ (.a(net490),
    .b(net471),
    .o1(_11026_));
 b15nandp2an1n02x5 _19692_ (.a(_10725_),
    .b(_10833_),
    .o1(_11027_));
 b15aoi012ar1n06x5 _19693_ (.a(_10866_),
    .b(_10867_),
    .c(net484),
    .o1(_11028_));
 b15nand02aq1n04x5 _19694_ (.a(net476),
    .b(net468),
    .o1(_11029_));
 b15oaoi13as1n08x5 _19695_ (.a(_11026_),
    .b(_11027_),
    .c(_11028_),
    .d(_11029_),
    .o1(_11030_));
 b15aoi012ar1n04x5 _19696_ (.a(_10833_),
    .b(_10869_),
    .c(_10732_),
    .o1(_11031_));
 b15nand03aq1n04x5 _19697_ (.a(_10893_),
    .b(net471),
    .c(_10847_),
    .o1(_11032_));
 b15oai022an1n12x5 _19698_ (.a(_10721_),
    .b(_10786_),
    .c(_11031_),
    .d(_11032_),
    .o1(_11033_));
 b15oai012ar1n32x5 _19699_ (.a(net479),
    .b(_11030_),
    .c(_11033_),
    .o1(_11034_));
 b15nandp2aq1n08x5 _19700_ (.a(net477),
    .b(net469),
    .o1(_11035_));
 b15nand03al1n02x5 _19701_ (.a(net473),
    .b(_10847_),
    .c(_10756_),
    .o1(_11036_));
 b15bfn001as1n48x5 max_length922 (.a(\us00.a[4] ),
    .o(net922));
 b15norp02ar1n02x5 _19703_ (.a(net480),
    .b(net473),
    .o1(_11038_));
 b15and002ah1n08x5 _19704_ (.a(net479),
    .b(net475),
    .o(_11039_));
 b15aoi022ar1n02x5 _19705_ (.a(_10847_),
    .b(_11038_),
    .c(_11039_),
    .d(_10725_),
    .o1(_11040_));
 b15and002aq1n03x5 _19706_ (.a(net486),
    .b(net483),
    .o(_11041_));
 b15oaoi13aq1n02x5 _19707_ (.a(_11035_),
    .b(_11036_),
    .c(_11040_),
    .d(_11041_),
    .o1(_11042_));
 b15norp03ar1n02x5 _19708_ (.a(net478),
    .b(net469),
    .c(_11036_),
    .o1(_11043_));
 b15norp02aq1n04x5 _19709_ (.a(_11042_),
    .b(_11043_),
    .o1(_11044_));
 b15nand02an1n02x5 _19710_ (.a(_10750_),
    .b(_10824_),
    .o1(_11045_));
 b15oaoi13an1n08x5 _19711_ (.a(_10808_),
    .b(_11045_),
    .c(_10824_),
    .d(_10851_),
    .o1(_11046_));
 b15norp02as1n16x5 _19712_ (.a(net489),
    .b(net481),
    .o1(_11047_));
 b15norp03ar1n12x5 _19713_ (.a(net473),
    .b(net467),
    .c(net465),
    .o1(_11048_));
 b15aoi022ar1n02x5 _19714_ (.a(_10913_),
    .b(_11047_),
    .c(_11048_),
    .d(net481),
    .o1(_11049_));
 b15nor002an1n02x5 _19715_ (.a(_10826_),
    .b(_11049_),
    .o1(_11050_));
 b15nano23al1n06x5 _19716_ (.a(_11034_),
    .b(_11044_),
    .c(_11046_),
    .d(_11050_),
    .out0(_11051_));
 b15bfn001as1n64x5 wire921 (.a(\us00.a[4] ),
    .o(net921));
 b15oai112al1n04x5 _19718_ (.a(net478),
    .b(_10813_),
    .c(_10822_),
    .d(_10912_),
    .o1(_11053_));
 b15oai013ar1n06x5 _19719_ (.a(_11053_),
    .b(_10813_),
    .c(_10921_),
    .d(net478),
    .o1(_11054_));
 b15nanb02an1n16x5 _19720_ (.a(net485),
    .b(net478),
    .out0(_11055_));
 b15nor003al1n04x5 _19721_ (.a(_10732_),
    .b(_10721_),
    .c(_11055_),
    .o1(_11056_));
 b15aoi112al1n06x5 _19722_ (.a(_11054_),
    .b(_11056_),
    .c(_10860_),
    .d(_11048_),
    .o1(_11057_));
 b15nor003ar1n02x5 _19723_ (.a(_10893_),
    .b(net478),
    .c(_10738_),
    .o1(_11058_));
 b15aoi013as1n03x5 _19724_ (.a(_11058_),
    .b(_10819_),
    .c(net478),
    .d(_10893_),
    .o1(_11059_));
 b15aoai13as1n08x5 _19725_ (.a(_11051_),
    .b(net482),
    .c(_11057_),
    .d(_11059_),
    .o1(_11060_));
 b15nano23as1n24x5 _19726_ (.a(_10972_),
    .b(_10985_),
    .c(_11025_),
    .d(_11060_),
    .out0(_11061_));
 b15xor002al1n12x5 _19727_ (.a(\u0.w[0][17] ),
    .b(_11061_),
    .out0(_11062_));
 b15xnr002as1n06x5 _19728_ (.a(\u0.w[1][17] ),
    .b(_11062_),
    .out0(_11063_));
 b15bfn001ah1n64x5 wire920 (.a(\us00.a[5] ),
    .o(net920));
 b15bfn001as1n64x5 max_length919 (.a(\us00.a[5] ),
    .o(net919));
 b15bfn001as1n48x5 load_slew918 (.a(\us00.a[6] ),
    .o(net918));
 b15xor002ar1n02x5 _19732_ (.a(\u0.tmp_w[17] ),
    .b(\u0.w[2][17] ),
    .out0(_11067_));
 b15xor002ar1n02x5 _19733_ (.a(_11063_),
    .b(_11067_),
    .out0(_11068_));
 b15cmbn22ar1n02x5 _19734_ (.clk1(net37),
    .clk2(_11068_),
    .clkout(_00361_),
    .s(net946));
 b15nand02ah1n03x5 _19735_ (.a(net129),
    .b(net38),
    .o1(_11069_));
 b15bfn001ah1n64x5 load_slew917 (.a(\us00.a[6] ),
    .o(net917));
 b15bfn001as1n64x5 max_length916 (.a(\us00.a[7] ),
    .o(net916));
 b15bfn001as1n64x5 max_length915 (.a(\us00.a[7] ),
    .o(net915));
 b15bfn001as1n64x5 wire914 (.a(\us00.a[7] ),
    .o(net914));
 b15and003ar1n02x5 _19740_ (.a(net483),
    .b(_10873_),
    .c(_10833_),
    .o(_11074_));
 b15nor002an1n08x5 _19741_ (.a(_10939_),
    .b(_10993_),
    .o1(_11075_));
 b15oaoi13ar1n03x5 _19742_ (.a(_11074_),
    .b(net486),
    .c(_11007_),
    .d(_11075_),
    .o1(_11076_));
 b15nanb02an1n03x5 _19743_ (.a(net483),
    .b(net486),
    .out0(_11077_));
 b15aoi012ar1n02x5 _19744_ (.a(_11077_),
    .b(_10903_),
    .c(net480),
    .o1(_11078_));
 b15aob012ar1n02x5 _19745_ (.a(net486),
    .b(net480),
    .c(_10750_),
    .out0(_11079_));
 b15aoi012as1n02x5 _19746_ (.a(_11078_),
    .b(_11079_),
    .c(net483),
    .o1(_11080_));
 b15nor003al1n06x5 _19747_ (.a(net478),
    .b(net466),
    .c(net462),
    .o1(_11081_));
 b15aob012an1n03x5 _19748_ (.a(_11081_),
    .b(_10858_),
    .c(_10828_),
    .out0(_11082_));
 b15oai022ah1n02x5 _19749_ (.a(net480),
    .b(_11076_),
    .c(_11080_),
    .d(_11082_),
    .o1(_11083_));
 b15oai012ar1n02x5 _19750_ (.a(net486),
    .b(_10872_),
    .c(_10860_),
    .o1(_11084_));
 b15oaoi13aq1n03x5 _19751_ (.a(_10721_),
    .b(_11084_),
    .c(_10974_),
    .d(net483),
    .o1(_11085_));
 b15aoai13ar1n02x5 _19752_ (.a(net486),
    .b(net483),
    .c(net480),
    .d(net477),
    .o1(_11086_));
 b15nand04an1n02x5 _19753_ (.a(_10808_),
    .b(_10920_),
    .c(_10718_),
    .d(_11086_),
    .o1(_11087_));
 b15nanb02as1n16x5 _19754_ (.a(net483),
    .b(net474),
    .out0(_11088_));
 b15aoi022aq1n08x5 _19755_ (.a(net477),
    .b(_10881_),
    .c(_10883_),
    .d(_10820_),
    .o1(_11089_));
 b15oai013ah1n03x5 _19756_ (.a(_11087_),
    .b(_11088_),
    .c(_11089_),
    .d(net466),
    .o1(_11090_));
 b15nonb02aq1n04x5 _19757_ (.a(_10838_),
    .b(_11090_),
    .out0(_11091_));
 b15xor002as1n08x5 _19758_ (.a(net479),
    .b(net476),
    .out0(_11092_));
 b15oai022ar1n04x5 _19759_ (.a(_10806_),
    .b(_10750_),
    .c(_11092_),
    .d(net486),
    .o1(_11093_));
 b15oai112ar1n02x5 _19760_ (.a(net477),
    .b(_10750_),
    .c(_10745_),
    .d(net480),
    .o1(_11094_));
 b15aoi022ar1n02x5 _19761_ (.a(net483),
    .b(_11093_),
    .c(_11094_),
    .d(_10921_),
    .o1(_11095_));
 b15nonb02as1n04x5 _19762_ (.a(net467),
    .b(net476),
    .out0(_11096_));
 b15oai112an1n06x5 _19763_ (.a(net464),
    .b(_11096_),
    .c(_10850_),
    .d(_10724_),
    .o1(_11097_));
 b15aoi022aq1n08x5 _19764_ (.a(_10959_),
    .b(_10833_),
    .c(_10869_),
    .d(_10960_),
    .o1(_11098_));
 b15oai013an1n12x5 _19765_ (.a(_11097_),
    .b(_11098_),
    .c(net487),
    .d(net464),
    .o1(_11099_));
 b15aoi012al1n04x5 _19766_ (.a(_11095_),
    .b(_11099_),
    .c(_10756_),
    .o1(_11100_));
 b15nona23ah1n12x5 _19767_ (.a(_11083_),
    .b(_11085_),
    .c(_11091_),
    .d(_11100_),
    .out0(_11101_));
 b15bfn001ah1n80x5 wire913 (.a(\us10.a[0] ),
    .o(net913));
 b15norp03as1n02x5 _19769_ (.a(_10724_),
    .b(_10850_),
    .c(_10729_),
    .o1(_11103_));
 b15oaoi13al1n03x5 _19770_ (.a(_10732_),
    .b(_10858_),
    .c(_10828_),
    .d(net485),
    .o1(_11104_));
 b15oai112al1n08x5 _19771_ (.a(net478),
    .b(_10847_),
    .c(_11103_),
    .d(_11104_),
    .o1(_11105_));
 b15nor002ah1n06x5 _19772_ (.a(_10804_),
    .b(_10805_),
    .o1(_11106_));
 b15nonb02al1n06x5 _19773_ (.a(net481),
    .b(net476),
    .out0(_11107_));
 b15nanb02aq1n12x5 _19774_ (.a(net487),
    .b(net477),
    .out0(_11108_));
 b15aoi012an1n06x5 _19775_ (.a(net480),
    .b(_11108_),
    .c(net483),
    .o1(_11109_));
 b15aoi012al1n02x5 _19776_ (.a(_10732_),
    .b(net476),
    .c(_10952_),
    .o1(_11110_));
 b15oai013an1n06x5 _19777_ (.a(_11106_),
    .b(_11107_),
    .c(_11109_),
    .d(_11110_),
    .o1(_11111_));
 b15nandp3ar1n02x5 _19778_ (.a(_10724_),
    .b(_10914_),
    .c(_10725_),
    .o1(_11112_));
 b15oai013ar1n02x5 _19779_ (.a(_11112_),
    .b(_10878_),
    .c(_10851_),
    .d(net485),
    .o1(_11113_));
 b15nand02al1n04x5 _19780_ (.a(net477),
    .b(net473),
    .o1(_11114_));
 b15oai022al1n02x5 _19781_ (.a(net477),
    .b(_10804_),
    .c(_11114_),
    .d(net471),
    .o1(_11115_));
 b15aoi013al1n03x5 _19782_ (.a(_11113_),
    .b(_11115_),
    .c(net481),
    .d(_10720_),
    .o1(_11116_));
 b15oai112as1n08x5 _19783_ (.a(_11105_),
    .b(_11111_),
    .c(_10732_),
    .d(_11116_),
    .o1(_11117_));
 b15nanb02aq1n06x5 _19784_ (.a(net470),
    .b(net464),
    .out0(_11118_));
 b15norp02ar1n08x5 _19785_ (.a(net475),
    .b(_11118_),
    .o1(_11119_));
 b15orn003ar1n02x5 _19786_ (.a(_10783_),
    .b(_10881_),
    .c(_10883_),
    .o(_11120_));
 b15oaoi13an1n04x5 _19787_ (.a(net479),
    .b(_11120_),
    .c(_10828_),
    .d(net487),
    .o1(_11121_));
 b15oai112as1n16x5 _19788_ (.a(net484),
    .b(net466),
    .c(_11119_),
    .d(_11121_),
    .o1(_11122_));
 b15aoi012ar1n02x5 _19789_ (.a(net476),
    .b(_10740_),
    .c(_10988_),
    .o1(_11123_));
 b15nandp2al1n03x5 _19790_ (.a(net472),
    .b(net464),
    .o1(_11124_));
 b15nanb02ar1n02x5 _19791_ (.a(_11124_),
    .b(_10992_),
    .out0(_11125_));
 b15nonb02aq1n16x5 _19792_ (.a(\u0.tmp_w[12] ),
    .b(\u0.tmp_w[9] ),
    .out0(_11126_));
 b15aoi022ar1n02x5 _19793_ (.a(net488),
    .b(_10861_),
    .c(_11126_),
    .d(net467),
    .o1(_11127_));
 b15oai012aq1n03x5 _19794_ (.a(_11123_),
    .b(_11125_),
    .c(_11127_),
    .o1(_11128_));
 b15nonb02aq1n16x5 _19795_ (.a(net470),
    .b(net468),
    .out0(_11129_));
 b15aoi012ah1n08x5 _19796_ (.a(_10957_),
    .b(_11129_),
    .c(net484),
    .o1(_11130_));
 b15nand02al1n02x5 _19797_ (.a(_10720_),
    .b(_10831_),
    .o1(_11131_));
 b15obai22ah1n02x5 _19798_ (.a(_10867_),
    .b(_11130_),
    .c(_11131_),
    .d(net471),
    .out0(_11132_));
 b15aoi012aq1n06x5 _19799_ (.a(_11128_),
    .b(_11132_),
    .c(net479),
    .o1(_11133_));
 b15oai112an1n06x5 _19800_ (.a(_10729_),
    .b(_10811_),
    .c(net488),
    .d(_10872_),
    .o1(_11134_));
 b15oai013ar1n02x5 _19801_ (.a(net477),
    .b(_10805_),
    .c(_10903_),
    .d(_10723_),
    .o1(_11135_));
 b15nanb02ah1n12x5 _19802_ (.a(\u0.tmp_w[12] ),
    .b(net485),
    .out0(_11136_));
 b15oai022ar1n04x5 _19803_ (.a(_10805_),
    .b(_11088_),
    .c(_11136_),
    .d(_10810_),
    .o1(_11137_));
 b15aoi013an1n03x5 _19804_ (.a(_11135_),
    .b(_11137_),
    .c(_11047_),
    .d(net471),
    .o1(_11138_));
 b15aoi022aq1n12x5 _19805_ (.a(_11122_),
    .b(_11133_),
    .c(_11134_),
    .d(_11138_),
    .o1(_11139_));
 b15oai012ar1n03x5 _19806_ (.a(_10738_),
    .b(_10998_),
    .c(net481),
    .o1(_11140_));
 b15oai022ar1n02x5 _19807_ (.a(_10766_),
    .b(_10738_),
    .c(_10726_),
    .d(net481),
    .o1(_11141_));
 b15aoi022al1n02x5 _19808_ (.a(_10745_),
    .b(_11140_),
    .c(_11141_),
    .d(net489),
    .o1(_11142_));
 b15aoai13ar1n02x5 _19809_ (.a(net489),
    .b(_10740_),
    .c(_10726_),
    .d(_10872_),
    .o1(_11143_));
 b15nand03ar1n02x5 _19810_ (.a(net485),
    .b(_11017_),
    .c(_11004_),
    .o1(_11144_));
 b15oai112ar1n04x5 _19811_ (.a(_10893_),
    .b(_10726_),
    .c(_11047_),
    .d(_11004_),
    .o1(_11145_));
 b15nandp3ar1n04x5 _19812_ (.a(_11143_),
    .b(_11144_),
    .c(_11145_),
    .o1(_11146_));
 b15aoi012as1n04x5 _19813_ (.a(_10939_),
    .b(_11142_),
    .c(_11146_),
    .o1(_11147_));
 b15nor004as1n12x5 _19814_ (.a(_11101_),
    .b(_11117_),
    .c(_11139_),
    .d(_11147_),
    .o1(_11148_));
 b15xor002an1n08x5 _19815_ (.a(\u0.w[0][18] ),
    .b(_11148_),
    .out0(_11149_));
 b15xor002ar1n08x5 _19816_ (.a(\u0.w[1][18] ),
    .b(_11149_),
    .out0(_11150_));
 b15xor002aq1n02x5 _19817_ (.a(\u0.w[2][18] ),
    .b(_11150_),
    .out0(_11151_));
 b15xor002ar1n02x5 _19818_ (.a(\u0.tmp_w[18] ),
    .b(_11151_),
    .out0(_11152_));
 b15oai012ar1n02x5 _19819_ (.a(_11069_),
    .b(_11152_),
    .c(net946),
    .o1(_00362_));
 b15inv020as1n05x5 _19820_ (.a(net39),
    .o1(_11153_));
 b15bfn001as1n64x5 max_length912 (.a(net913),
    .o(net912));
 b15bfn001ah1n64x5 max_length911 (.a(net912),
    .o(net911));
 b15bfn001as1n48x5 max_length910 (.a(net911),
    .o(net910));
 b15norp02ar1n02x5 _19824_ (.a(_10952_),
    .b(_11114_),
    .o1(_11157_));
 b15nona22aq1n02x5 _19825_ (.a(net477),
    .b(\u0.tmp_w[12] ),
    .c(net481),
    .out0(_11158_));
 b15oai012aq1n02x5 _19826_ (.a(_11158_),
    .b(_11114_),
    .c(net481),
    .o1(_11159_));
 b15aoai13aq1n04x5 _19827_ (.a(_10834_),
    .b(_11157_),
    .c(_11159_),
    .d(_10824_),
    .o1(_11160_));
 b15nona23aq1n16x5 _19828_ (.a(net473),
    .b(net469),
    .c(net466),
    .d(net462),
    .out0(_11161_));
 b15nand03aq1n03x5 _19829_ (.a(net478),
    .b(_11161_),
    .c(_10993_),
    .o1(_11162_));
 b15bfn001as1n48x5 wire909 (.a(\us10.a[1] ),
    .o(net909));
 b15oai013ar1n04x5 _19831_ (.a(_10939_),
    .b(_10828_),
    .c(_10755_),
    .d(_11041_),
    .o1(_11164_));
 b15nand03al1n08x5 _19832_ (.a(net480),
    .b(_11162_),
    .c(_11164_),
    .o1(_11165_));
 b15aoai13al1n03x5 _19833_ (.a(_10817_),
    .b(_10835_),
    .c(net477),
    .d(_10750_),
    .o1(_11166_));
 b15aoi012al1n02x5 _19834_ (.a(_10732_),
    .b(_10766_),
    .c(_10835_),
    .o1(_11167_));
 b15oai112ah1n06x5 _19835_ (.a(_11160_),
    .b(_11165_),
    .c(_11166_),
    .d(_11167_),
    .o1(_11168_));
 b15norp02aq1n02x5 _19836_ (.a(_10903_),
    .b(_10755_),
    .o1(_11169_));
 b15nandp3al1n03x5 _19837_ (.a(_10939_),
    .b(_11169_),
    .c(_10831_),
    .o1(_11170_));
 b15aoi022an1n04x5 _19838_ (.a(_10860_),
    .b(_11169_),
    .c(_10829_),
    .d(net477),
    .o1(_11171_));
 b15oai112ar1n12x5 _19839_ (.a(net480),
    .b(_11170_),
    .c(_11171_),
    .d(net488),
    .o1(_11172_));
 b15oai022ar1n02x5 _19840_ (.a(net477),
    .b(_10840_),
    .c(_10786_),
    .d(_10738_),
    .o1(_11173_));
 b15nand02al1n02x5 _19841_ (.a(_10732_),
    .b(_11173_),
    .o1(_11174_));
 b15oai112al1n08x5 _19842_ (.a(_10728_),
    .b(_11174_),
    .c(_10840_),
    .d(_10981_),
    .o1(_11175_));
 b15oai122aq1n08x5 _19843_ (.a(_10732_),
    .b(_10721_),
    .c(_10974_),
    .d(_10826_),
    .e(_10921_),
    .o1(_11176_));
 b15aoai13al1n03x5 _19844_ (.a(net478),
    .b(_10994_),
    .c(_10750_),
    .d(_10740_),
    .o1(_11177_));
 b15nand02al1n03x5 _19845_ (.a(_10820_),
    .b(_10929_),
    .o1(_11178_));
 b15aoai13al1n04x5 _19846_ (.a(_11107_),
    .b(_11106_),
    .c(net485),
    .d(_10822_),
    .o1(_11179_));
 b15nand04an1n08x5 _19847_ (.a(net488),
    .b(_11177_),
    .c(_11178_),
    .d(_11179_),
    .o1(_11180_));
 b15aoi122an1n06x5 _19848_ (.a(_11168_),
    .b(_11172_),
    .c(_11175_),
    .d(_11176_),
    .e(_11180_),
    .o1(_11181_));
 b15nand02an1n02x5 _19849_ (.a(_10822_),
    .b(_10941_),
    .o1(_11182_));
 b15nandp2ar1n02x5 _19850_ (.a(net488),
    .b(_10939_),
    .o1(_11183_));
 b15nandp2as1n05x5 _19851_ (.a(_10850_),
    .b(_10725_),
    .o1(_11184_));
 b15oai112ar1n08x5 _19852_ (.a(_10893_),
    .b(_11182_),
    .c(_11183_),
    .d(_11184_),
    .o1(_11185_));
 b15oai022ar1n02x5 _19853_ (.a(_10939_),
    .b(_10840_),
    .c(_10815_),
    .d(_11158_),
    .o1(_11186_));
 b15and002al1n02x5 _19854_ (.a(_10732_),
    .b(_11186_),
    .o(_11187_));
 b15nonb02aq1n03x5 _19855_ (.a(net478),
    .b(net489),
    .out0(_11188_));
 b15aoi022al1n02x5 _19856_ (.a(_10820_),
    .b(_10742_),
    .c(_11188_),
    .d(_10929_),
    .o1(_11189_));
 b15oai112aq1n08x5 _19857_ (.a(net485),
    .b(_11189_),
    .c(_10998_),
    .d(_10732_),
    .o1(_11190_));
 b15nor002an1n08x5 _19858_ (.a(net471),
    .b(_10877_),
    .o1(_11191_));
 b15oai012al1n08x5 _19859_ (.a(_11191_),
    .b(_10869_),
    .c(_10833_),
    .o1(_11192_));
 b15and002al1n03x5 _19860_ (.a(net476),
    .b(net474),
    .o(_11193_));
 b15aoi022aq1n08x5 _19861_ (.a(_11020_),
    .b(_11129_),
    .c(_11193_),
    .d(_10957_),
    .o1(_11194_));
 b15aob012an1n06x5 _19862_ (.a(net464),
    .b(_11092_),
    .c(_10732_),
    .out0(_11195_));
 b15oai022al1n16x5 _19863_ (.a(net479),
    .b(_11192_),
    .c(_11194_),
    .d(_11195_),
    .o1(_11196_));
 b15oai013ar1n08x5 _19864_ (.a(_11185_),
    .b(_11187_),
    .c(_11190_),
    .d(_11196_),
    .o1(_11197_));
 b15aoi012ar1n02x5 _19865_ (.a(_10811_),
    .b(_10742_),
    .c(_10808_),
    .o1(_11198_));
 b15oai112ar1n02x5 _19866_ (.a(net488),
    .b(_10981_),
    .c(_10742_),
    .d(_10766_),
    .o1(_11199_));
 b15aoi012ar1n02x5 _19867_ (.a(_11107_),
    .b(_10878_),
    .c(net485),
    .o1(_11200_));
 b15aoai13ar1n03x5 _19868_ (.a(_11200_),
    .b(net485),
    .c(net477),
    .d(_10811_),
    .o1(_11201_));
 b15oaoi13ah1n03x5 _19869_ (.a(_11198_),
    .b(_11199_),
    .c(_11201_),
    .d(net488),
    .o1(_11202_));
 b15aob012an1n06x5 _19870_ (.a(_10795_),
    .b(_10796_),
    .c(_10939_),
    .out0(_11203_));
 b15nand04as1n06x5 _19871_ (.a(_10765_),
    .b(_10832_),
    .c(_11108_),
    .d(_11203_),
    .o1(_11204_));
 b15inv000aq1n20x5 _19872_ (.a(net475),
    .o1(_11205_));
 b15oai112as1n02x5 _19873_ (.a(_10873_),
    .b(_10827_),
    .c(_10817_),
    .d(_11205_),
    .o1(_11206_));
 b15aoi112ar1n02x5 _19874_ (.a(_10815_),
    .b(_11088_),
    .c(_11009_),
    .d(net486),
    .o1(_11207_));
 b15nanb02al1n16x5 _19875_ (.a(net471),
    .b(\u0.tmp_w[12] ),
    .out0(_11208_));
 b15nanb02an1n03x5 _19876_ (.a(net481),
    .b(net471),
    .out0(_11209_));
 b15oai022al1n02x5 _19877_ (.a(_10728_),
    .b(_11208_),
    .c(_10816_),
    .d(_11209_),
    .o1(_11210_));
 b15aoi013an1n03x5 _19878_ (.a(_11207_),
    .b(_11210_),
    .c(net486),
    .d(_10720_),
    .o1(_11211_));
 b15aoai13al1n03x5 _19879_ (.a(net477),
    .b(_10819_),
    .c(_10813_),
    .d(_10913_),
    .o1(_11212_));
 b15nand04al1n08x5 _19880_ (.a(_11204_),
    .b(_11206_),
    .c(_11211_),
    .d(_11212_),
    .o1(_11213_));
 b15nor003al1n03x5 _19881_ (.a(net480),
    .b(_10813_),
    .c(_10993_),
    .o1(_11214_));
 b15nor002as1n04x5 _19882_ (.a(net480),
    .b(_10993_),
    .o1(_11215_));
 b15norp03aq1n08x5 _19883_ (.a(_10728_),
    .b(_10804_),
    .c(_10805_),
    .o1(_11216_));
 b15oaoi13as1n04x5 _19884_ (.a(_11214_),
    .b(_10831_),
    .c(_11215_),
    .d(_11216_),
    .o1(_11217_));
 b15norp03al1n02x5 _19885_ (.a(net483),
    .b(_10810_),
    .c(_10804_),
    .o1(_11218_));
 b15norp02ar1n02x5 _19886_ (.a(_10840_),
    .b(_10759_),
    .o1(_11219_));
 b15oai022ar1n02x5 _19887_ (.a(_10810_),
    .b(_10804_),
    .c(_10840_),
    .d(net483),
    .o1(_11220_));
 b15aoi112ah1n02x5 _19888_ (.a(_11218_),
    .b(_11219_),
    .c(_11220_),
    .d(_10732_),
    .o1(_11221_));
 b15oai022ah1n06x5 _19889_ (.a(_10939_),
    .b(_11217_),
    .c(_11221_),
    .d(_11009_),
    .o1(_11222_));
 b15nor003aq1n06x5 _19890_ (.a(_11202_),
    .b(_11213_),
    .c(_11222_),
    .o1(_11223_));
 b15nor003ar1n02x5 _19891_ (.a(_11205_),
    .b(_10981_),
    .c(_11010_),
    .o1(_11224_));
 b15orn002aq1n04x5 _19892_ (.a(net484),
    .b(net475),
    .o(_11225_));
 b15oaoi13ar1n02x5 _19893_ (.a(_10939_),
    .b(_10898_),
    .c(_11225_),
    .d(_10899_),
    .o1(_11226_));
 b15oai012an1n02x5 _19894_ (.a(net468),
    .b(_11224_),
    .c(_11226_),
    .o1(_11227_));
 b15oaoi13as1n04x5 _19895_ (.a(net479),
    .b(_11227_),
    .c(_10816_),
    .d(_10815_),
    .o1(_11228_));
 b15aoi012al1n02x5 _19896_ (.a(_11039_),
    .b(_10944_),
    .c(net484),
    .o1(_11229_));
 b15nand02an1n02x5 _19897_ (.a(net476),
    .b(_10834_),
    .o1(_11230_));
 b15nand03al1n06x5 _19898_ (.a(net484),
    .b(net479),
    .c(net475),
    .o1(_11231_));
 b15aob012al1n03x5 _19899_ (.a(_10873_),
    .b(_10944_),
    .c(_11231_),
    .out0(_11232_));
 b15oai022an1n08x5 _19900_ (.a(_11229_),
    .b(_11230_),
    .c(_11232_),
    .d(net476),
    .o1(_11233_));
 b15nand03al1n03x5 _19901_ (.a(net479),
    .b(_10833_),
    .c(_11191_),
    .o1(_11234_));
 b15norp02ar1n02x5 _19902_ (.a(net476),
    .b(_10815_),
    .o1(_11235_));
 b15aoi013ah1n02x5 _19903_ (.a(_11235_),
    .b(_11191_),
    .c(net476),
    .d(net479),
    .o1(_11236_));
 b15oai012al1n06x5 _19904_ (.a(_11234_),
    .b(_11236_),
    .c(_11225_),
    .o1(_11237_));
 b15oai013as1n12x5 _19905_ (.a(net490),
    .b(_11228_),
    .c(_11233_),
    .d(_11237_),
    .o1(_11238_));
 b15nand04as1n16x5 _19906_ (.a(_11181_),
    .b(_11197_),
    .c(_11223_),
    .d(_11238_),
    .o1(_11239_));
 b15xnr002al1n12x5 _19907_ (.a(\u0.w[0][19] ),
    .b(_11239_),
    .out0(_11240_));
 b15xor002ah1n04x5 _19908_ (.a(\u0.w[1][19] ),
    .b(_11240_),
    .out0(_11241_));
 b15xor002al1n04x5 _19909_ (.a(\u0.w[2][19] ),
    .b(_11241_),
    .out0(_11242_));
 b15xor002al1n02x5 _19910_ (.a(\u0.tmp_w[19] ),
    .b(_11242_),
    .out0(_11243_));
 b15mdn022ar1n02x5 _19911_ (.a(_11153_),
    .b(_11243_),
    .o1(_00363_),
    .sa(net946));
 b15nand02ar1n02x5 _19912_ (.a(net939),
    .b(net41),
    .o1(_11244_));
 b15bfn001as1n48x5 load_slew908 (.a(net909),
    .o(net908));
 b15bfn001ah1n64x5 max_length907 (.a(net909),
    .o(net907));
 b15bfn001as1n48x5 max_length906 (.a(net909),
    .o(net906));
 b15nandp3al1n08x5 _19916_ (.a(net480),
    .b(_10768_),
    .c(_10783_),
    .o1(_11248_));
 b15oai012aq1n06x5 _19917_ (.a(_11136_),
    .b(_11126_),
    .c(_10732_),
    .o1(_11249_));
 b15oai112al1n12x5 _19918_ (.a(_10896_),
    .b(_11248_),
    .c(_11249_),
    .d(net481),
    .o1(_11250_));
 b15norp02ar1n02x5 _19919_ (.a(_10804_),
    .b(_10992_),
    .o1(_11251_));
 b15nanb02aq1n08x5 _19920_ (.a(net489),
    .b(net481),
    .out0(_11252_));
 b15oai022ar1n02x5 _19921_ (.a(net481),
    .b(_10804_),
    .c(_11252_),
    .d(_11208_),
    .o1(_11253_));
 b15aoai13ah1n02x5 _19922_ (.a(_10847_),
    .b(_11251_),
    .c(_11253_),
    .d(net485),
    .o1(_11254_));
 b15aoi012ah1n04x5 _19923_ (.a(net476),
    .b(_11250_),
    .c(_11254_),
    .o1(_11255_));
 b15and002ar1n08x5 _19924_ (.a(net482),
    .b(net478),
    .o(_11256_));
 b15aoi122aq1n08x5 _19925_ (.a(_10732_),
    .b(_11256_),
    .c(_10750_),
    .d(_10988_),
    .e(_10914_),
    .o1(_11257_));
 b15norp02ar1n02x5 _19926_ (.a(net478),
    .b(_10822_),
    .o1(_11258_));
 b15and002ar1n02x5 _19927_ (.a(_10728_),
    .b(_11055_),
    .o(_11259_));
 b15aoi022ar1n04x5 _19928_ (.a(_10847_),
    .b(_10718_),
    .c(_10822_),
    .d(_10845_),
    .o1(_11260_));
 b15oai013ar1n03x5 _19929_ (.a(_11257_),
    .b(_11258_),
    .c(_11259_),
    .d(_11260_),
    .o1(_11261_));
 b15oai022aq1n06x5 _19930_ (.a(_11184_),
    .b(_11055_),
    .c(_11009_),
    .d(_11017_),
    .o1(_11262_));
 b15nor002aq1n02x5 _19931_ (.a(_11259_),
    .b(_11260_),
    .o1(_11263_));
 b15oai012aq1n08x5 _19932_ (.a(_10732_),
    .b(_10728_),
    .c(_10860_),
    .o1(_11264_));
 b15aoai13aq1n06x5 _19933_ (.a(_11261_),
    .b(_11262_),
    .c(_11263_),
    .d(_11264_),
    .o1(_11265_));
 b15oai012ar1n06x5 _19934_ (.a(_10858_),
    .b(_10974_),
    .c(_10828_),
    .o1(_11266_));
 b15and002al1n04x5 _19935_ (.a(net474),
    .b(net464),
    .o(_11267_));
 b15nandp2ar1n08x5 _19936_ (.a(_10820_),
    .b(_11267_),
    .o1(_11268_));
 b15norp03ar1n08x5 _19937_ (.a(net477),
    .b(net475),
    .c(net468),
    .o1(_11269_));
 b15nand02ah1n02x5 _19938_ (.a(net475),
    .b(net468),
    .o1(_11270_));
 b15oab012ah1n06x5 _19939_ (.a(_11269_),
    .b(_10974_),
    .c(_11270_),
    .out0(_11271_));
 b15oai022ar1n24x5 _19940_ (.a(_11130_),
    .b(_11268_),
    .c(_11271_),
    .d(_11010_),
    .o1(_11272_));
 b15aoi022ar1n12x5 _19941_ (.a(_10720_),
    .b(_11266_),
    .c(_11272_),
    .d(_10759_),
    .o1(_11273_));
 b15oai013aq1n02x5 _19942_ (.a(_10732_),
    .b(net478),
    .c(_10952_),
    .d(_10993_),
    .o1(_11274_));
 b15aoi013ah1n04x5 _19943_ (.a(_11274_),
    .b(_10750_),
    .c(net478),
    .d(_10893_),
    .o1(_11275_));
 b15oai112as1n16x5 _19944_ (.a(_11265_),
    .b(_11273_),
    .c(_11275_),
    .d(_11257_),
    .o1(_11276_));
 b15nor004al1n02x5 _19945_ (.a(net471),
    .b(_10755_),
    .c(_10941_),
    .d(_11088_),
    .o1(_11277_));
 b15aoi013aq1n03x5 _19946_ (.a(_11277_),
    .b(_10882_),
    .c(_11191_),
    .d(_10813_),
    .o1(_11278_));
 b15and002aq1n03x5 _19947_ (.a(_10939_),
    .b(_11278_),
    .o(_11279_));
 b15oai022aq1n02x5 _19948_ (.a(_10729_),
    .b(_10921_),
    .c(_10721_),
    .d(net485),
    .o1(_11280_));
 b15aoai13an1n08x5 _19949_ (.a(_10732_),
    .b(_11280_),
    .c(_10913_),
    .d(net481),
    .o1(_11281_));
 b15aoai13ar1n02x5 _19950_ (.a(\u0.tmp_w[9] ),
    .b(_10929_),
    .c(_10904_),
    .d(_11047_),
    .o1(_11282_));
 b15aoai13al1n02x5 _19951_ (.a(net485),
    .b(_10941_),
    .c(_10993_),
    .d(_10728_),
    .o1(_11283_));
 b15oai022as1n06x5 _19952_ (.a(_10810_),
    .b(_10804_),
    .c(_10924_),
    .d(_10993_),
    .o1(_11284_));
 b15oai112al1n06x5 _19953_ (.a(_11283_),
    .b(_11284_),
    .c(_11252_),
    .d(_10988_),
    .o1(_11285_));
 b15and003ar1n03x5 _19954_ (.a(net476),
    .b(_11282_),
    .c(_11285_),
    .o(_11286_));
 b15xor002ar1n02x5 _19955_ (.a(net479),
    .b(net468),
    .out0(_11287_));
 b15nand02aq1n02x5 _19956_ (.a(_10867_),
    .b(_11287_),
    .o1(_11288_));
 b15aoi022ah1n02x5 _19957_ (.a(_10725_),
    .b(_10880_),
    .c(_10867_),
    .d(net479),
    .o1(_11289_));
 b15oaoi13as1n04x5 _19958_ (.a(\u0.tmp_w[13] ),
    .b(_11288_),
    .c(_11289_),
    .d(net484),
    .o1(_11290_));
 b15aoai13an1n08x5 _19959_ (.a(net488),
    .b(_11290_),
    .c(_11126_),
    .d(_10834_),
    .o1(_11291_));
 b15aoi022al1n12x5 _19960_ (.a(_11279_),
    .b(_11281_),
    .c(_11286_),
    .d(_11291_),
    .o1(_11292_));
 b15oai022ar1n02x5 _19961_ (.a(_10912_),
    .b(_10742_),
    .c(_10974_),
    .d(net489),
    .o1(_11293_));
 b15aob012ar1n02x5 _19962_ (.a(_10742_),
    .b(_11252_),
    .c(_10992_),
    .out0(_11294_));
 b15nandp3ar1n02x5 _19963_ (.a(_10912_),
    .b(_11252_),
    .c(_10992_),
    .o1(_11295_));
 b15aoi013ar1n02x5 _19964_ (.a(_11293_),
    .b(_11294_),
    .c(_11295_),
    .d(net485),
    .o1(_11296_));
 b15oai012ar1n02x5 _19965_ (.a(_10728_),
    .b(_10912_),
    .c(_10732_),
    .o1(_11297_));
 b15aoi022as1n02x5 _19966_ (.a(_10851_),
    .b(_11047_),
    .c(_11297_),
    .d(_10939_),
    .o1(_11298_));
 b15oai012an1n04x5 _19967_ (.a(_11296_),
    .b(_11298_),
    .c(net485),
    .o1(_11299_));
 b15nandp3ar1n02x5 _19968_ (.a(_10834_),
    .b(_11107_),
    .c(_11126_),
    .o1(_11300_));
 b15aoi022al1n04x5 _19969_ (.a(_10820_),
    .b(_10957_),
    .c(_11129_),
    .d(net476),
    .o1(_11301_));
 b15oai013as1n02x5 _19970_ (.a(_11300_),
    .b(_11301_),
    .c(_11136_),
    .d(net464),
    .o1(_11302_));
 b15nand02al1n02x5 _19971_ (.a(net489),
    .b(_11302_),
    .o1(_11303_));
 b15norp02aq1n08x5 _19972_ (.a(\u0.tmp_w[12] ),
    .b(net465),
    .o1(_11304_));
 b15nona23as1n02x5 _19973_ (.a(net472),
    .b(_11304_),
    .c(net467),
    .d(\u0.tmp_w[9] ),
    .out0(_11305_));
 b15nonb02al1n06x5 _19974_ (.a(net490),
    .b(net465),
    .out0(_11306_));
 b15oaoi13ah1n04x5 _19975_ (.a(_11305_),
    .b(net479),
    .c(_11205_),
    .d(_11306_),
    .o1(_11307_));
 b15norp02ar1n02x5 _19976_ (.a(_10726_),
    .b(_11252_),
    .o1(_11308_));
 b15oai012al1n03x5 _19977_ (.a(net476),
    .b(_11307_),
    .c(_11308_),
    .o1(_11309_));
 b15nandp2ar1n03x5 _19978_ (.a(_10893_),
    .b(_10913_),
    .o1(_11310_));
 b15oai122al1n04x5 _19979_ (.a(_10728_),
    .b(_11004_),
    .c(_10864_),
    .d(_11310_),
    .e(net476),
    .o1(_11311_));
 b15oai022ah1n04x5 _19980_ (.a(_11124_),
    .b(_10792_),
    .c(_10966_),
    .d(_10899_),
    .o1(_11312_));
 b15aoi022ar1n08x5 _19981_ (.a(net476),
    .b(_11106_),
    .c(_11096_),
    .d(_11312_),
    .o1(_11313_));
 b15aob012as1n03x5 _19982_ (.a(_11311_),
    .b(_11313_),
    .c(net481),
    .out0(_11314_));
 b15nand04aq1n08x5 _19983_ (.a(_11299_),
    .b(_11303_),
    .c(_11309_),
    .d(_11314_),
    .o1(_11315_));
 b15nor004as1n12x5 _19984_ (.a(_11255_),
    .b(_11276_),
    .c(_11292_),
    .d(_11315_),
    .o1(_11316_));
 b15xor002as1n16x5 _19985_ (.a(\u0.w[0][20] ),
    .b(_11316_),
    .out0(_11317_));
 b15xor002ah1n16x5 _19986_ (.a(\u0.w[1][20] ),
    .b(_11317_),
    .out0(_11318_));
 b15xor002al1n03x5 _19987_ (.a(\u0.w[2][20] ),
    .b(_11318_),
    .out0(_11319_));
 b15xor002ar1n02x5 _19988_ (.a(\u0.tmp_w[20] ),
    .b(_11319_),
    .out0(_11320_));
 b15oai012ar1n02x5 _19989_ (.a(_11244_),
    .b(_11320_),
    .c(net939),
    .o1(_00365_));
 b15inv040as1n12x5 _19990_ (.a(net42),
    .o1(_11321_));
 b15bfn001ah1n64x5 wire905 (.a(net906),
    .o(net905));
 b15bfn001as1n64x5 wire904 (.a(\us10.a[2] ),
    .o(net904));
 b15bfn001as1n64x5 max_length903 (.a(net904),
    .o(net903));
 b15norp02ar1n02x5 _19994_ (.a(_10808_),
    .b(_10815_),
    .o1(_11325_));
 b15aob012ar1n02x5 _19995_ (.a(net486),
    .b(_11088_),
    .c(_11136_),
    .out0(_11326_));
 b15nor004ar1n02x5 _19996_ (.a(_10877_),
    .b(_10833_),
    .c(_10869_),
    .d(_11209_),
    .o1(_11327_));
 b15aoi022aq1n02x5 _19997_ (.a(_11249_),
    .b(_11325_),
    .c(_11326_),
    .d(_11327_),
    .o1(_11328_));
 b15nandp2al1n02x5 _19998_ (.a(_10893_),
    .b(_11081_),
    .o1(_11329_));
 b15and003al1n03x5 _19999_ (.a(net483),
    .b(net466),
    .c(net462),
    .o(_11330_));
 b15aoi012al1n04x5 _20000_ (.a(_11081_),
    .b(_11330_),
    .c(net478),
    .o1(_11331_));
 b15oaoi13an1n08x5 _20001_ (.a(_10804_),
    .b(_11329_),
    .c(_11331_),
    .d(_10992_),
    .o1(_11332_));
 b15aoai13an1n03x5 _20002_ (.a(_10847_),
    .b(_10724_),
    .c(_10850_),
    .d(_10893_),
    .o1(_11333_));
 b15aoai13an1n03x5 _20003_ (.a(_10732_),
    .b(net485),
    .c(_10847_),
    .d(_10850_),
    .o1(_11334_));
 b15aoi112an1n06x5 _20004_ (.a(net478),
    .b(_11333_),
    .c(_11334_),
    .d(net482),
    .o1(_11335_));
 b15nand02al1n02x5 _20005_ (.a(_10914_),
    .b(_10819_),
    .o1(_11336_));
 b15oaoi13as1n04x5 _20006_ (.a(_10732_),
    .b(_11336_),
    .c(_10845_),
    .d(_10726_),
    .o1(_11337_));
 b15aoi012ar1n06x5 _20007_ (.a(_11161_),
    .b(_11264_),
    .c(_10808_),
    .o1(_11338_));
 b15nor004as1n12x5 _20008_ (.a(_11332_),
    .b(_11335_),
    .c(_11337_),
    .d(_11338_),
    .o1(_11339_));
 b15oai022ar1n02x5 _20009_ (.a(_10944_),
    .b(_11118_),
    .c(_11010_),
    .d(_10966_),
    .o1(_11340_));
 b15and003as1n02x5 _20010_ (.a(net476),
    .b(_10758_),
    .c(_11340_),
    .o(_11341_));
 b15aoi112ar1n03x5 _20011_ (.a(_10728_),
    .b(net476),
    .c(_11017_),
    .d(_10967_),
    .o1(_11342_));
 b15oai012al1n06x5 _20012_ (.a(net487),
    .b(_11341_),
    .c(_11342_),
    .o1(_11343_));
 b15nandp2aq1n02x5 _20013_ (.a(net471),
    .b(_11188_),
    .o1(_11344_));
 b15aoai13al1n02x5 _20014_ (.a(net481),
    .b(_11048_),
    .c(_10847_),
    .d(net473),
    .o1(_11345_));
 b15oaoi13aq1n04x5 _20015_ (.a(_11344_),
    .b(_11345_),
    .c(_10966_),
    .d(_10810_),
    .o1(_11346_));
 b15nand03al1n03x5 _20016_ (.a(_10847_),
    .b(_10724_),
    .c(_10813_),
    .o1(_11347_));
 b15nandp3al1n03x5 _20017_ (.a(net485),
    .b(_10920_),
    .c(_10754_),
    .o1(_11348_));
 b15aoi013ah1n03x5 _20018_ (.a(_10974_),
    .b(_11184_),
    .c(_11347_),
    .d(_11348_),
    .o1(_11349_));
 b15nor004as1n08x5 _20019_ (.a(_10859_),
    .b(_11046_),
    .c(_11346_),
    .d(_11349_),
    .o1(_11350_));
 b15nand04an1n08x5 _20020_ (.a(_11328_),
    .b(_11339_),
    .c(_11343_),
    .d(_11350_),
    .o1(_11351_));
 b15aoi022ar1n12x5 _20021_ (.a(net485),
    .b(_10920_),
    .c(_10720_),
    .d(net486),
    .o1(_11352_));
 b15oai122ah1n16x5 _20022_ (.a(net478),
    .b(_10805_),
    .c(_10858_),
    .d(_11352_),
    .e(_10804_),
    .o1(_11353_));
 b15aoi022ar1n02x5 _20023_ (.a(net483),
    .b(_10819_),
    .c(_10831_),
    .d(_10988_),
    .o1(_11354_));
 b15aoai13ar1n02x5 _20024_ (.a(_10732_),
    .b(_10819_),
    .c(_10988_),
    .d(net483),
    .o1(_11355_));
 b15aoi012ar1n02x5 _20025_ (.a(net480),
    .b(_11354_),
    .c(_11355_),
    .o1(_11356_));
 b15aoi112an1n02x5 _20026_ (.a(net464),
    .b(_11039_),
    .c(_10787_),
    .d(_10745_),
    .o1(_11357_));
 b15nand03an1n08x5 _20027_ (.a(net474),
    .b(net469),
    .c(net466),
    .o1(_11358_));
 b15oai012an1n02x5 _20028_ (.a(_11358_),
    .b(_10831_),
    .c(_10787_),
    .o1(_11359_));
 b15aoi112aq1n03x5 _20029_ (.a(_11353_),
    .b(_11356_),
    .c(_11357_),
    .d(_11359_),
    .o1(_11360_));
 b15aoai13ar1n02x5 _20030_ (.a(_10732_),
    .b(_10728_),
    .c(_10721_),
    .d(net483),
    .o1(_11361_));
 b15oaoi13ar1n02x5 _20031_ (.a(_10740_),
    .b(_10840_),
    .c(_10721_),
    .d(_10872_),
    .o1(_11362_));
 b15nand02an1n02x5 _20032_ (.a(_11361_),
    .b(_11362_),
    .o1(_11363_));
 b15oai112al1n02x5 _20033_ (.a(_10872_),
    .b(_10959_),
    .c(_11267_),
    .d(_11304_),
    .o1(_11364_));
 b15aoi022ar1n02x5 _20034_ (.a(_10765_),
    .b(_10882_),
    .c(_11267_),
    .d(_10924_),
    .o1(_11365_));
 b15oai112as1n02x5 _20035_ (.a(_10939_),
    .b(_11364_),
    .c(_11365_),
    .d(_10889_),
    .o1(_11366_));
 b15oai012al1n02x5 _20036_ (.a(_10903_),
    .b(_10828_),
    .c(_10732_),
    .o1(_11367_));
 b15aoi013an1n03x5 _20037_ (.a(_11366_),
    .b(_11367_),
    .c(_10920_),
    .d(_10740_),
    .o1(_11368_));
 b15aoi012al1n02x5 _20038_ (.a(_10813_),
    .b(_10738_),
    .c(net480),
    .o1(_11369_));
 b15oai013an1n08x5 _20039_ (.a(_11369_),
    .b(_10829_),
    .c(_10822_),
    .d(net480),
    .o1(_11370_));
 b15aoi013ah1n04x5 _20040_ (.a(_11360_),
    .b(_11363_),
    .c(_11368_),
    .d(_11370_),
    .o1(_11371_));
 b15nandp2ar1n04x5 _20041_ (.a(net484),
    .b(_10796_),
    .o1(_11372_));
 b15aoai13ar1n08x5 _20042_ (.a(net462),
    .b(_11035_),
    .c(_11372_),
    .d(_10795_),
    .o1(_11373_));
 b15aoi022ar1n02x5 _20043_ (.a(_10939_),
    .b(_10850_),
    .c(_10959_),
    .d(_11193_),
    .o1(_11374_));
 b15mdn022ar1n03x5 _20044_ (.a(_10957_),
    .b(_11129_),
    .o1(_11375_),
    .sa(net474));
 b15oai022ah1n02x5 _20045_ (.a(_10893_),
    .b(_11374_),
    .c(_11375_),
    .d(net476),
    .o1(_11376_));
 b15oai112ah1n06x5 _20046_ (.a(_10732_),
    .b(_11373_),
    .c(_11376_),
    .d(net464),
    .o1(_11377_));
 b15nanb03al1n03x5 _20047_ (.a(\u0.tmp_w[12] ),
    .b(net465),
    .c(net476),
    .out0(_11378_));
 b15nona22ar1n02x5 _20048_ (.a(net476),
    .b(net465),
    .c(\u0.tmp_w[12] ),
    .out0(_11379_));
 b15aoi012aq1n04x5 _20049_ (.a(_10787_),
    .b(_11378_),
    .c(_11379_),
    .o1(_11380_));
 b15aob012an1n03x5 _20050_ (.a(_11310_),
    .b(_11380_),
    .c(\u0.tmp_w[9] ),
    .out0(_11381_));
 b15aoi022ah1n08x5 _20051_ (.a(_10824_),
    .b(_11380_),
    .c(_11381_),
    .d(net489),
    .o1(_11382_));
 b15aoi022ar1n06x5 _20052_ (.a(net476),
    .b(_10834_),
    .c(_11096_),
    .d(_10765_),
    .o1(_11383_));
 b15oai112as1n08x5 _20053_ (.a(_11377_),
    .b(_11382_),
    .c(_11383_),
    .d(_11088_),
    .o1(_11384_));
 b15aoi112as1n08x5 _20054_ (.a(_11351_),
    .b(_11371_),
    .c(_11384_),
    .d(net481),
    .o1(_11385_));
 b15xor002as1n16x5 _20055_ (.a(\u0.w[0][21] ),
    .b(_11385_),
    .out0(_11386_));
 b15xor002as1n16x5 _20056_ (.a(\u0.w[1][21] ),
    .b(_11386_),
    .out0(_11387_));
 b15xor002as1n12x5 _20057_ (.a(\u0.w[2][21] ),
    .b(_11387_),
    .out0(_11388_));
 b15xor002an1n02x5 _20058_ (.a(net443),
    .b(_11388_),
    .out0(_11389_));
 b15bfn001as1n64x5 max_length902 (.a(net903),
    .o(net902));
 b15mdn022ar1n02x5 _20060_ (.a(_11321_),
    .b(_11389_),
    .o1(_00366_),
    .sa(net936));
 b15nand02ar1n02x5 _20061_ (.a(net939),
    .b(net43),
    .o1(_11391_));
 b15bfn001as1n48x5 wire901 (.a(net903),
    .o(net901));
 b15bfn001as1n64x5 wire900 (.a(\us10.a[3] ),
    .o(net900));
 b15bfn001as1n64x5 max_length899 (.a(net900),
    .o(net899));
 b15bfn001as1n64x5 max_length898 (.a(net900),
    .o(net898));
 b15nonb03ar1n02x5 _20066_ (.a(net467),
    .b(net465),
    .c(\u0.tmp_w[12] ),
    .out0(_11396_));
 b15oai112ah1n02x5 _20067_ (.a(net472),
    .b(_10820_),
    .c(_10942_),
    .d(_11396_),
    .o1(_11397_));
 b15nand04ar1n03x5 _20068_ (.a(net479),
    .b(net476),
    .c(_10847_),
    .d(_10724_),
    .o1(_11398_));
 b15nand02ar1n02x5 _20069_ (.a(_10820_),
    .b(_10913_),
    .o1(_11399_));
 b15aoai13an1n02x5 _20070_ (.a(_11397_),
    .b(\u0.tmp_w[9] ),
    .c(_11398_),
    .d(_11399_),
    .o1(_11400_));
 b15nand02an1n12x5 _20071_ (.a(net476),
    .b(_10988_),
    .o1(_11401_));
 b15nandp3ar1n02x5 _20072_ (.a(\u0.tmp_w[9] ),
    .b(_10939_),
    .c(_10913_),
    .o1(_11402_));
 b15oai112aq1n02x5 _20073_ (.a(_11401_),
    .b(_11402_),
    .c(\u0.tmp_w[9] ),
    .d(_11017_),
    .o1(_11403_));
 b15aoai13an1n03x5 _20074_ (.a(net488),
    .b(_11400_),
    .c(_11403_),
    .d(net479),
    .o1(_11404_));
 b15nano22al1n03x5 _20075_ (.a(net487),
    .b(_10840_),
    .c(_10819_),
    .out0(_11405_));
 b15aoai13aq1n04x5 _20076_ (.a(_10847_),
    .b(_10724_),
    .c(_10718_),
    .d(net483),
    .o1(_11406_));
 b15aoi112ar1n08x5 _20077_ (.a(_11009_),
    .b(_11405_),
    .c(_11406_),
    .d(_10732_),
    .o1(_11407_));
 b15oai022al1n02x5 _20078_ (.a(net476),
    .b(_10787_),
    .c(_10785_),
    .d(\u0.tmp_w[9] ),
    .o1(_11408_));
 b15oai012al1n02x5 _20079_ (.a(_10939_),
    .b(_10742_),
    .c(\u0.tmp_w[9] ),
    .o1(_11409_));
 b15oai012ar1n02x5 _20080_ (.a(_10864_),
    .b(_10750_),
    .c(net476),
    .o1(_11410_));
 b15aoi022an1n04x5 _20081_ (.a(_11047_),
    .b(_11409_),
    .c(_11410_),
    .d(net481),
    .o1(_11411_));
 b15aoi013ar1n03x5 _20082_ (.a(_11407_),
    .b(_11408_),
    .c(_11411_),
    .d(_11304_),
    .o1(_11412_));
 b15nandp3al1n02x5 _20083_ (.a(net476),
    .b(_10765_),
    .c(_10889_),
    .o1(_11413_));
 b15oai012as1n04x5 _20084_ (.a(_11413_),
    .b(_10965_),
    .c(net476),
    .o1(_11414_));
 b15aoai13an1n08x5 _20085_ (.a(_10893_),
    .b(_11075_),
    .c(_11414_),
    .d(_10880_),
    .o1(_11415_));
 b15aoi022ar1n02x5 _20086_ (.a(net485),
    .b(_10912_),
    .c(_10834_),
    .d(_11126_),
    .o1(_11416_));
 b15oai022as1n02x5 _20087_ (.a(_10738_),
    .b(_10786_),
    .c(_11416_),
    .d(_10732_),
    .o1(_11417_));
 b15nand02ah1n02x5 _20088_ (.a(net481),
    .b(_11417_),
    .o1(_11418_));
 b15nand04ah1n08x5 _20089_ (.a(_11404_),
    .b(_11412_),
    .c(_11415_),
    .d(_11418_),
    .o1(_11419_));
 b15orn002ar1n02x5 _20090_ (.a(net480),
    .b(net466),
    .o(_11420_));
 b15nona23ar1n02x5 _20091_ (.a(net486),
    .b(net469),
    .c(net462),
    .d(net473),
    .out0(_11421_));
 b15nona22ar1n05x5 _20092_ (.a(net473),
    .b(net462),
    .c(net469),
    .out0(_11422_));
 b15oaoi13as1n03x5 _20093_ (.a(_11420_),
    .b(_11421_),
    .c(_11422_),
    .d(_11077_),
    .o1(_11423_));
 b15oaoi13ar1n08x5 _20094_ (.a(_11423_),
    .b(net483),
    .c(_11215_),
    .d(_11216_),
    .o1(_11424_));
 b15aoi112ah1n03x5 _20095_ (.a(net490),
    .b(_10965_),
    .c(_11225_),
    .d(_11231_),
    .o1(_11425_));
 b15and003as1n02x5 _20096_ (.a(net484),
    .b(net471),
    .c(_10725_),
    .o(_11426_));
 b15aoi112ar1n06x5 _20097_ (.a(net490),
    .b(net471),
    .c(_10877_),
    .d(_10755_),
    .o1(_11427_));
 b15oaoi13as1n08x5 _20098_ (.a(_11425_),
    .b(_10869_),
    .c(_11426_),
    .d(_11427_),
    .o1(_11428_));
 b15oai022aq1n06x5 _20099_ (.a(net477),
    .b(_11424_),
    .c(_11428_),
    .d(_11256_),
    .o1(_11429_));
 b15oai012ar1n02x5 _20100_ (.a(_10759_),
    .b(_10766_),
    .c(net486),
    .o1(_11430_));
 b15aoai13ar1n02x5 _20101_ (.a(_11088_),
    .b(net480),
    .c(_10732_),
    .d(_11205_),
    .o1(_11431_));
 b15aoi022ar1n02x5 _20102_ (.a(_10822_),
    .b(_11430_),
    .c(_11431_),
    .d(_10834_),
    .o1(_11432_));
 b15aoi012aq1n02x5 _20103_ (.a(net484),
    .b(_11118_),
    .c(_11010_),
    .o1(_11433_));
 b15norp02ar1n03x5 _20104_ (.a(_10792_),
    .b(_11118_),
    .o1(_11434_));
 b15oai112ah1n08x5 _20105_ (.a(_10758_),
    .b(_10882_),
    .c(_11433_),
    .d(_11434_),
    .o1(_11435_));
 b15aoai13ar1n02x5 _20106_ (.a(_10913_),
    .b(_10924_),
    .c(_10952_),
    .d(_10732_),
    .o1(_11436_));
 b15aoi013ar1n02x5 _20107_ (.a(_10939_),
    .b(_11432_),
    .c(_11435_),
    .d(_11436_),
    .o1(_11437_));
 b15norp02ar1n02x5 _20108_ (.a(_10860_),
    .b(_10992_),
    .o1(_11438_));
 b15nand04ar1n02x5 _20109_ (.a(net477),
    .b(_10718_),
    .c(_10720_),
    .d(_10768_),
    .o1(_11439_));
 b15oaoi13aq1n02x5 _20110_ (.a(_11438_),
    .b(_11439_),
    .c(net477),
    .d(_10726_),
    .o1(_11440_));
 b15norp02ar1n02x5 _20111_ (.a(net483),
    .b(net466),
    .o1(_11441_));
 b15nor004an1n02x5 _20112_ (.a(net464),
    .b(_11208_),
    .c(_10806_),
    .d(_11441_),
    .o1(_11442_));
 b15oai112al1n06x5 _20113_ (.a(_10960_),
    .b(_10869_),
    .c(_10728_),
    .d(net464),
    .o1(_11443_));
 b15oab012al1n03x5 _20114_ (.a(net479),
    .b(net464),
    .c(net487),
    .out0(_11444_));
 b15oaoi13ah1n04x5 _20115_ (.a(_11443_),
    .b(_10759_),
    .c(net484),
    .d(_11444_),
    .o1(_11445_));
 b15nor004aq1n04x5 _20116_ (.a(_11005_),
    .b(_11440_),
    .c(_11442_),
    .d(_11445_),
    .o1(_11446_));
 b15nona23ah1n08x5 _20117_ (.a(_11429_),
    .b(_11437_),
    .c(_11446_),
    .d(_10821_),
    .out0(_11447_));
 b15nor002ah1n03x5 _20118_ (.a(\u0.tmp_w[9] ),
    .b(_10840_),
    .o1(_11448_));
 b15aoai13ah1n03x5 _20119_ (.a(_11047_),
    .b(_11448_),
    .c(\u0.tmp_w[9] ),
    .d(_10750_),
    .o1(_11449_));
 b15and002ar1n02x5 _20120_ (.a(_10893_),
    .b(_10750_),
    .o(_11450_));
 b15oaoi13al1n04x5 _20121_ (.a(_11450_),
    .b(net489),
    .c(_10750_),
    .d(_11448_),
    .o1(_11451_));
 b15oai112ar1n16x5 _20122_ (.a(net476),
    .b(_11449_),
    .c(_11451_),
    .d(_10728_),
    .o1(_11452_));
 b15nor002as1n03x5 _20123_ (.a(net484),
    .b(net474),
    .o1(_11453_));
 b15aoi013ah1n02x5 _20124_ (.a(net477),
    .b(_10960_),
    .c(_10781_),
    .d(_11453_),
    .o1(_11454_));
 b15mdn022aq1n02x5 _20125_ (.a(_10881_),
    .b(_10883_),
    .o1(_11455_),
    .sa(_10728_));
 b15oai013ah1n03x5 _20126_ (.a(_11454_),
    .b(_11455_),
    .c(_11270_),
    .d(_10759_),
    .o1(_11456_));
 b15nano23aq1n02x5 _20127_ (.a(net484),
    .b(net463),
    .c(net470),
    .d(net475),
    .out0(_11457_));
 b15aoai13as1n04x5 _20128_ (.a(net490),
    .b(_11457_),
    .c(_10883_),
    .d(net475),
    .o1(_11458_));
 b15aob012an1n02x5 _20129_ (.a(_11458_),
    .b(_11119_),
    .c(_10824_),
    .out0(_11459_));
 b15aoi013as1n04x5 _20130_ (.a(_11456_),
    .b(_11459_),
    .c(_10728_),
    .d(_10758_),
    .o1(_11460_));
 b15nandp3ar1n02x5 _20131_ (.a(net474),
    .b(_10847_),
    .c(_10924_),
    .o1(_11461_));
 b15aoai13ar1n02x5 _20132_ (.a(_10882_),
    .b(_10920_),
    .c(net483),
    .d(_10720_),
    .o1(_11462_));
 b15aoi012al1n02x5 _20133_ (.a(net469),
    .b(_11461_),
    .c(_11462_),
    .o1(_11463_));
 b15aoi013ar1n06x5 _20134_ (.a(_11463_),
    .b(_10880_),
    .c(_10720_),
    .d(net469),
    .o1(_11464_));
 b15oai012as1n12x5 _20135_ (.a(_11460_),
    .b(_11464_),
    .c(net487),
    .o1(_11465_));
 b15aoi112as1n08x5 _20136_ (.a(_11419_),
    .b(_11447_),
    .c(_11452_),
    .d(_11465_),
    .o1(_11466_));
 b15xor002as1n16x5 _20137_ (.a(\u0.w[0][22] ),
    .b(_11466_),
    .out0(_11467_));
 b15xor002as1n16x5 _20138_ (.a(\u0.w[1][22] ),
    .b(_11467_),
    .out0(_11468_));
 b15xor002ah1n04x5 _20139_ (.a(\u0.w[2][22] ),
    .b(_11468_),
    .out0(_11469_));
 b15xor002ar1n02x5 _20140_ (.a(\u0.tmp_w[22] ),
    .b(_11469_),
    .out0(_11470_));
 b15oai012ar1n02x5 _20141_ (.a(_11391_),
    .b(_11470_),
    .c(net939),
    .o1(_00367_));
 b15inv000al1n10x5 _20142_ (.a(net44),
    .o1(_11471_));
 b15bfn001as1n64x5 max_length897 (.a(net898),
    .o(net897));
 b15bfn001ah1n64x5 wire896 (.a(\us10.a[4] ),
    .o(net896));
 b15bfn001as1n64x5 load_slew895 (.a(net896),
    .o(net895));
 b15bfn001as1n64x5 max_length894 (.a(net895),
    .o(net894));
 b15norp03ar1n02x5 _20147_ (.a(net466),
    .b(_10804_),
    .c(_11108_),
    .o1(_11476_));
 b15oai022an1n08x5 _20148_ (.a(_10804_),
    .b(_10981_),
    .c(_11055_),
    .d(_11208_),
    .o1(_11477_));
 b15and002al1n03x5 _20149_ (.a(net480),
    .b(net466),
    .o(_11478_));
 b15aoai13al1n02x5 _20150_ (.a(net462),
    .b(_11476_),
    .c(_11477_),
    .d(_11478_),
    .o1(_11479_));
 b15oai012al1n03x5 _20151_ (.a(_10939_),
    .b(_11161_),
    .c(_10952_),
    .o1(_11480_));
 b15nandp2ar1n03x5 _20152_ (.a(net480),
    .b(net463),
    .o1(_11481_));
 b15oai022as1n02x5 _20153_ (.a(_10828_),
    .b(_11481_),
    .c(_10781_),
    .d(_10903_),
    .o1(_11482_));
 b15aoi013al1n02x5 _20154_ (.a(_11480_),
    .b(_11482_),
    .c(net466),
    .d(net487),
    .o1(_11483_));
 b15xor002an1n04x5 _20155_ (.a(net483),
    .b(net480),
    .out0(_11484_));
 b15oai022ar1n02x5 _20156_ (.a(net480),
    .b(_10813_),
    .c(_11484_),
    .d(_10732_),
    .o1(_11485_));
 b15nand02al1n03x5 _20157_ (.a(_10819_),
    .b(_11485_),
    .o1(_11486_));
 b15aoi013an1n02x5 _20158_ (.a(_10939_),
    .b(_10759_),
    .c(_10750_),
    .d(net480),
    .o1(_11487_));
 b15aoai13ar1n04x5 _20159_ (.a(_11479_),
    .b(_11483_),
    .c(_11486_),
    .d(_11487_),
    .o1(_11488_));
 b15norp02ar1n02x5 _20160_ (.a(_10804_),
    .b(_10974_),
    .o1(_11489_));
 b15nanb03ar1n02x5 _20161_ (.a(net487),
    .b(net466),
    .c(net462),
    .out0(_11490_));
 b15oai013al1n02x5 _20162_ (.a(_11490_),
    .b(_10720_),
    .c(_10920_),
    .d(_10893_),
    .o1(_11491_));
 b15oai122ah1n02x5 _20163_ (.a(_10808_),
    .b(_10806_),
    .c(_10893_),
    .d(_11484_),
    .e(_10732_),
    .o1(_11492_));
 b15aoi022ar1n02x5 _20164_ (.a(_11489_),
    .b(_11491_),
    .c(_11492_),
    .d(_10742_),
    .o1(_11493_));
 b15oai013ar1n03x5 _20165_ (.a(_11358_),
    .b(_10831_),
    .c(_10828_),
    .d(net466),
    .o1(_11494_));
 b15aoi012ar1n02x5 _20166_ (.a(net487),
    .b(net483),
    .c(net474),
    .o1(_11495_));
 b15aoi013ar1n02x5 _20167_ (.a(_11495_),
    .b(_11136_),
    .c(_11088_),
    .d(net487),
    .o1(_11496_));
 b15aoi022ar1n04x5 _20168_ (.a(_10813_),
    .b(_11494_),
    .c(_11496_),
    .d(_10957_),
    .o1(_11497_));
 b15oai013as1n02x5 _20169_ (.a(_11493_),
    .b(_11497_),
    .c(net462),
    .d(_11009_),
    .o1(_11498_));
 b15nanb02an1n04x5 _20170_ (.a(_11217_),
    .b(net478),
    .out0(_11499_));
 b15nandp3ar1n02x5 _20171_ (.a(_10728_),
    .b(_10847_),
    .c(_10850_),
    .o1(_11500_));
 b15oaoi13ah1n02x5 _20172_ (.a(net487),
    .b(_11500_),
    .c(_10968_),
    .d(net483),
    .o1(_11501_));
 b15aoi022ah1n04x5 _20173_ (.a(_10732_),
    .b(_10834_),
    .c(_11306_),
    .d(_10957_),
    .o1(_11502_));
 b15nor003an1n12x5 _20174_ (.a(net484),
    .b(_10944_),
    .c(_11502_),
    .o1(_11503_));
 b15nanb03ar1n02x5 _20175_ (.a(net469),
    .b(net462),
    .c(net473),
    .out0(_11504_));
 b15aoi112al1n02x5 _20176_ (.a(net466),
    .b(_10952_),
    .c(_11422_),
    .d(_11504_),
    .o1(_11505_));
 b15and003ar1n02x5 _20177_ (.a(_10847_),
    .b(_10850_),
    .c(_10924_),
    .o(_11506_));
 b15nand04ah1n03x5 _20178_ (.a(net480),
    .b(_10724_),
    .c(_10725_),
    .d(_11041_),
    .o1(_11507_));
 b15nor003ar1n02x5 _20179_ (.a(net482),
    .b(net466),
    .c(net462),
    .o1(_11508_));
 b15oai112ah1n04x5 _20180_ (.a(_10724_),
    .b(_10759_),
    .c(_11330_),
    .d(_11508_),
    .o1(_11509_));
 b15nona23aq1n08x5 _20181_ (.a(_11505_),
    .b(_11506_),
    .c(_11507_),
    .d(_11509_),
    .out0(_11510_));
 b15oai013aq1n06x5 _20182_ (.a(_10939_),
    .b(_11501_),
    .c(_11503_),
    .d(_11510_),
    .o1(_11511_));
 b15nona23ar1n12x5 _20183_ (.a(_11488_),
    .b(_11498_),
    .c(_11499_),
    .d(_11511_),
    .out0(_11512_));
 b15oai022ar1n02x5 _20184_ (.a(_11161_),
    .b(_10806_),
    .c(_10786_),
    .d(_11004_),
    .o1(_11513_));
 b15aoi012ar1n02x5 _20185_ (.a(_10808_),
    .b(_10998_),
    .c(_10993_),
    .o1(_11514_));
 b15nano22ar1n02x5 _20186_ (.a(net469),
    .b(net462),
    .c(net477),
    .out0(_11515_));
 b15aoai13aq1n02x5 _20187_ (.a(_11478_),
    .b(_11515_),
    .c(net477),
    .d(_10765_),
    .o1(_11516_));
 b15nanb03ar1n02x5 _20188_ (.a(net462),
    .b(_10878_),
    .c(_11129_),
    .out0(_11517_));
 b15aoi012ah1n02x5 _20189_ (.a(net474),
    .b(_11516_),
    .c(_11517_),
    .o1(_11518_));
 b15oai013ar1n03x5 _20190_ (.a(net486),
    .b(_11513_),
    .c(_11514_),
    .d(_11518_),
    .o1(_11519_));
 b15aoai13al1n02x5 _20191_ (.a(net486),
    .b(_10835_),
    .c(_11075_),
    .d(net483),
    .o1(_11520_));
 b15oai012ar1n06x5 _20192_ (.a(_11520_),
    .b(_11401_),
    .c(_10768_),
    .o1(_11521_));
 b15aob012ah1n04x5 _20193_ (.a(_11519_),
    .b(_11521_),
    .c(net480),
    .out0(_11522_));
 b15norp02ar1n02x5 _20194_ (.a(net462),
    .b(_10806_),
    .o1(_11523_));
 b15aoi012ar1n02x5 _20195_ (.a(_10795_),
    .b(net470),
    .c(net487),
    .o1(_11524_));
 b15oai112ar1n04x5 _20196_ (.a(_11523_),
    .b(_11524_),
    .c(net469),
    .d(_10813_),
    .o1(_11525_));
 b15oai112ah1n06x5 _20197_ (.a(_10893_),
    .b(_10834_),
    .c(_10869_),
    .d(_10833_),
    .o1(_11526_));
 b15norp03ah1n03x5 _20198_ (.a(net462),
    .b(_10795_),
    .c(_10974_),
    .o1(_11527_));
 b15aobi12ar1n02x5 _20199_ (.a(_11526_),
    .b(_11527_),
    .c(net483),
    .out0(_11528_));
 b15norp02ar1n02x5 _20200_ (.a(_10773_),
    .b(_11478_),
    .o1(_11529_));
 b15nor003ah1n03x5 _20201_ (.a(_10898_),
    .b(_11108_),
    .c(_11529_),
    .o1(_11530_));
 b15nonb03an1n02x5 _20202_ (.a(net470),
    .b(net463),
    .c(net480),
    .out0(_11531_));
 b15and003ar1n02x5 _20203_ (.a(net477),
    .b(net475),
    .c(net468),
    .o(_11532_));
 b15oai112al1n06x5 _20204_ (.a(_10759_),
    .b(_11531_),
    .c(_11532_),
    .d(_11269_),
    .o1(_11533_));
 b15aob012ar1n02x5 _20205_ (.a(net466),
    .b(_11481_),
    .c(_10781_),
    .out0(_11534_));
 b15oai013as1n02x5 _20206_ (.a(_11533_),
    .b(_11534_),
    .c(_10828_),
    .d(_10786_),
    .o1(_11535_));
 b15nano23ar1n06x5 _20207_ (.a(_11525_),
    .b(_11528_),
    .c(_11530_),
    .d(_11535_),
    .out0(_11536_));
 b15oai013ah1n03x5 _20208_ (.a(_10974_),
    .b(_11009_),
    .c(_10732_),
    .d(net466),
    .o1(_11537_));
 b15aoi013ar1n06x5 _20209_ (.a(_11527_),
    .b(_11537_),
    .c(net462),
    .d(_11453_),
    .o1(_11538_));
 b15oai112aq1n16x5 _20210_ (.a(_11034_),
    .b(_11536_),
    .c(_11538_),
    .d(net469),
    .o1(_11539_));
 b15aoi012ar1n02x5 _20211_ (.a(_10773_),
    .b(_10831_),
    .c(net466),
    .o1(_11540_));
 b15norp03al1n02x5 _20212_ (.a(_10939_),
    .b(_10898_),
    .c(_11540_),
    .o1(_11541_));
 b15oaoi13ar1n02x5 _20213_ (.a(net487),
    .b(_11358_),
    .c(_10828_),
    .d(net484),
    .o1(_11542_));
 b15aoai13an1n02x5 _20214_ (.a(net462),
    .b(_11542_),
    .c(_11126_),
    .d(_10960_),
    .o1(_11543_));
 b15oaoi13aq1n04x5 _20215_ (.a(net477),
    .b(_11543_),
    .c(_11458_),
    .d(net466),
    .o1(_11544_));
 b15oab012ar1n06x5 _20216_ (.a(net480),
    .b(_11541_),
    .c(_11544_),
    .out0(_11545_));
 b15nor004as1n12x5 _20217_ (.a(_11512_),
    .b(_11522_),
    .c(_11539_),
    .d(_11545_),
    .o1(_11546_));
 b15xor002an1n06x5 _20218_ (.a(\u0.w[0][23] ),
    .b(_11546_),
    .out0(_11547_));
 b15xor002ah1n03x5 _20219_ (.a(\u0.w[1][23] ),
    .b(_11547_),
    .out0(_11548_));
 b15xor002ar1n08x5 _20220_ (.a(\u0.w[2][23] ),
    .b(net391),
    .out0(_11549_));
 b15xor002ar1n03x5 _20221_ (.a(\u0.tmp_w[23] ),
    .b(_11549_),
    .out0(_11550_));
 b15mdn022ar1n02x5 _20222_ (.a(_11471_),
    .b(_11550_),
    .o1(_00368_),
    .sa(net940));
 b15nand02ar1n12x5 _20223_ (.a(net129),
    .b(net45),
    .o1(_11551_));
 b15bfn001as1n64x5 max_length893 (.a(\us10.a[5] ),
    .o(net893));
 b15bfn001as1n64x5 max_length892 (.a(\us10.a[5] ),
    .o(net892));
 b15bfn001ah1n64x5 load_slew891 (.a(\us10.a[6] ),
    .o(net891));
 b15bfn001as1n48x5 max_length890 (.a(\us10.a[6] ),
    .o(net890));
 b15nanb02as1n24x5 _20228_ (.a(net449),
    .b(net447),
    .out0(_11556_));
 b15bfn001ah1n64x5 max_length889 (.a(\us10.a[6] ),
    .o(net889));
 b15bfn001as1n80x5 wire888 (.a(\us10.a[7] ),
    .o(net888));
 b15nona22as1n32x5 _20231_ (.a(\u0.tmp_w[22] ),
    .b(net435),
    .c(net443),
    .out0(_11559_));
 b15bfn001ah1n64x5 load_slew887 (.a(net888),
    .o(net887));
 b15norp02al1n02x5 _20233_ (.a(_11556_),
    .b(_11559_),
    .o1(_11561_));
 b15bfn001ah1n64x5 wire886 (.a(net888),
    .o(net886));
 b15bfn001as1n48x5 load_slew885 (.a(\us20.a[0] ),
    .o(net885));
 b15orn003as1n12x5 _20236_ (.a(net443),
    .b(net439),
    .c(net433),
    .o(_11564_));
 b15nandp2an1n48x5 _20237_ (.a(net449),
    .b(\u0.tmp_w[20] ),
    .o1(_11565_));
 b15bfn001ah1n64x5 load_slew884 (.a(\us20.a[0] ),
    .o(net884));
 b15norp02as1n04x5 _20239_ (.a(_11564_),
    .b(_11565_),
    .o1(_11567_));
 b15bfn001ah1n48x5 max_length883 (.a(net885),
    .o(net883));
 b15aoai13ar1n02x5 _20241_ (.a(net460),
    .b(_11561_),
    .c(_11567_),
    .d(net455),
    .o1(_11569_));
 b15bfn001as1n48x5 max_length882 (.a(net883),
    .o(net882));
 b15nor002as1n24x5 _20243_ (.a(net461),
    .b(net456),
    .o1(_11571_));
 b15aoi022ar1n02x5 _20244_ (.a(net455),
    .b(_11561_),
    .c(_11567_),
    .d(_11571_),
    .o1(_11572_));
 b15aoi012aq1n02x5 _20245_ (.a(net454),
    .b(_11569_),
    .c(_11572_),
    .o1(_11573_));
 b15nonb02as1n16x5 _20246_ (.a(net454),
    .b(net448),
    .out0(_11574_));
 b15nanb02as1n24x5 _20247_ (.a(net433),
    .b(net439),
    .out0(_11575_));
 b15bfn001as1n64x5 load_slew881 (.a(\us20.a[1] ),
    .o(net881));
 b15bfn001ah1n64x5 max_length880 (.a(\us20.a[1] ),
    .o(net880));
 b15bfn001ah1n64x5 load_slew879 (.a(net880),
    .o(net879));
 b15inv000ah1n80x5 _20251_ (.a(net459),
    .o1(_11579_));
 b15bfn001as1n48x5 load_slew878 (.a(\us20.a[2] ),
    .o(net878));
 b15aoi012ar1n02x5 _20253_ (.a(_11575_),
    .b(net444),
    .c(_11579_),
    .o1(_11581_));
 b15bfn001ah1n64x5 max_length877 (.a(net878),
    .o(net877));
 b15bfn001as1n48x5 max_length876 (.a(net878),
    .o(net876));
 b15nanb03an1n04x5 _20256_ (.a(net435),
    .b(net447),
    .c(net457),
    .out0(_11584_));
 b15bfn001ah1n64x5 wire875 (.a(\us20.a[2] ),
    .o(net875));
 b15nanb02al1n16x5 _20258_ (.a(net447),
    .b(net435),
    .out0(_11586_));
 b15bfn001as1n64x5 max_length874 (.a(\us20.a[3] ),
    .o(net874));
 b15oai012al1n06x5 _20260_ (.a(_11584_),
    .b(_11586_),
    .c(net457),
    .o1(_11588_));
 b15norp02ar1n02x5 _20261_ (.a(net460),
    .b(net439),
    .o1(_11589_));
 b15aoai13ar1n02x5 _20262_ (.a(net443),
    .b(_11581_),
    .c(_11588_),
    .d(_11589_),
    .o1(_11590_));
 b15nonb02aq1n12x5 _20263_ (.a(net455),
    .b(net447),
    .out0(_11591_));
 b15bfn001as1n64x5 max_length873 (.a(net874),
    .o(net873));
 b15norp03as1n24x5 _20265_ (.a(net441),
    .b(net439),
    .c(net433),
    .o1(_11593_));
 b15aob012as1n02x5 _20266_ (.a(_11590_),
    .b(_11591_),
    .c(_11593_),
    .out0(_11594_));
 b15aoi012as1n06x5 _20267_ (.a(_11573_),
    .b(_11574_),
    .c(_11594_),
    .o1(_11595_));
 b15bfn001as1n64x5 max_length872 (.a(net874),
    .o(net872));
 b15nanb02as1n24x5 _20269_ (.a(net438),
    .b(\u0.tmp_w[23] ),
    .out0(_11597_));
 b15bfn001as1n48x5 load_slew871 (.a(\us20.a[4] ),
    .o(net871));
 b15nor003ah1n02x5 _20271_ (.a(net451),
    .b(net440),
    .c(_11597_),
    .o1(_11599_));
 b15bfn001ah1n64x5 load_slew870 (.a(\us20.a[4] ),
    .o(net870));
 b15qgbin1an1n40x5 _20273_ (.a(net444),
    .o1(_11601_));
 b15nandp2al1n24x5 _20274_ (.a(\u0.tmp_w[18] ),
    .b(_11601_),
    .o1(_11602_));
 b15inv000as1n80x5 _20275_ (.a(net452),
    .o1(_11603_));
 b15nandp2aq1n04x5 _20276_ (.a(_11603_),
    .b(net445),
    .o1(_11604_));
 b15bfn001as1n64x5 max_length869 (.a(\us20.a[5] ),
    .o(net869));
 b15nanb02as1n24x5 _20278_ (.a(net461),
    .b(net456),
    .out0(_11606_));
 b15oai022aq1n02x5 _20279_ (.a(net456),
    .b(_11602_),
    .c(_11604_),
    .d(_11606_),
    .o1(_11607_));
 b15oaoi13as1n02x5 _20280_ (.a(_11579_),
    .b(_11602_),
    .c(_11604_),
    .d(net456),
    .o1(_11608_));
 b15oai012ah1n06x5 _20281_ (.a(_11599_),
    .b(_11607_),
    .c(_11608_),
    .o1(_11609_));
 b15bfn001as1n64x5 max_length868 (.a(\us20.a[5] ),
    .o(net868));
 b15bfn001as1n48x5 load_slew867 (.a(net869),
    .o(net867));
 b15bfn001as1n64x5 max_length866 (.a(\us20.a[6] ),
    .o(net866));
 b15nonb02aq1n16x5 _20285_ (.a(net444),
    .b(net448),
    .out0(_11613_));
 b15nonb02as1n16x5 _20286_ (.a(\u0.tmp_w[18] ),
    .b(net456),
    .out0(_11614_));
 b15bfn001as1n48x5 max_length865 (.a(net866),
    .o(net865));
 b15nano22ah1n12x5 _20288_ (.a(net437),
    .b(net434),
    .c(net440),
    .out0(_11616_));
 b15nand04an1n02x5 _20289_ (.a(net461),
    .b(_11613_),
    .c(_11614_),
    .d(_11616_),
    .o1(_11617_));
 b15nonb02as1n16x5 _20290_ (.a(net456),
    .b(net461),
    .out0(_11618_));
 b15nonb02aq1n12x5 _20291_ (.a(\u0.tmp_w[16] ),
    .b(net456),
    .out0(_11619_));
 b15aoi022ar1n02x5 _20292_ (.a(_11613_),
    .b(_11618_),
    .c(_11619_),
    .d(_11565_),
    .o1(_11620_));
 b15bfn001as1n64x5 max_length864 (.a(\us20.a[7] ),
    .o(net864));
 b15oai013ar1n02x5 _20294_ (.a(_11617_),
    .b(_11620_),
    .c(_11603_),
    .d(_11564_),
    .o1(_11622_));
 b15and002aq1n12x5 _20295_ (.a(net453),
    .b(net450),
    .o(_11623_));
 b15nor004as1n12x5 _20296_ (.a(net446),
    .b(net442),
    .c(net438),
    .d(net436),
    .o1(_11624_));
 b15bfn001as1n48x5 wire863 (.a(net864),
    .o(net863));
 b15nandp3ar1n02x5 _20298_ (.a(net455),
    .b(_11623_),
    .c(_11624_),
    .o1(_11626_));
 b15bfn001ah1n64x5 load_slew862 (.a(\us30.a[0] ),
    .o(net862));
 b15orn002an1n24x5 _20300_ (.a(net453),
    .b(net451),
    .o(_11628_));
 b15nona22as1n24x5 _20301_ (.a(net442),
    .b(net438),
    .c(net436),
    .out0(_11629_));
 b15oai013al1n02x5 _20302_ (.a(_11626_),
    .b(_11628_),
    .c(_11629_),
    .d(net445),
    .o1(_11630_));
 b15bfn001ah1n64x5 load_slew861 (.a(net862),
    .o(net861));
 b15bfn001as1n48x5 wire860 (.a(net862),
    .o(net860));
 b15aoi012al1n02x5 _20305_ (.a(_11622_),
    .b(_11630_),
    .c(_11579_),
    .o1(_11633_));
 b15bfn001ah1n64x5 max_length859 (.a(\us30.a[1] ),
    .o(net859));
 b15nanb02as1n24x5 _20307_ (.a(net450),
    .b(net453),
    .out0(_11635_));
 b15nor004ar1n02x5 _20308_ (.a(net461),
    .b(net445),
    .c(_11559_),
    .d(_11635_),
    .o1(_11636_));
 b15nona22as1n16x5 _20309_ (.a(net443),
    .b(net435),
    .c(net439),
    .out0(_11637_));
 b15nor002al1n12x5 _20310_ (.a(_11565_),
    .b(_11637_),
    .o1(_11638_));
 b15bfn001ah1n64x5 max_length858 (.a(net859),
    .o(net858));
 b15bfn001as1n48x5 max_length857 (.a(net859),
    .o(net857));
 b15aoai13ar1n03x5 _20313_ (.a(net455),
    .b(_11636_),
    .c(_11638_),
    .d(net461),
    .o1(_11641_));
 b15bfn001as1n64x5 max_length856 (.a(\us30.a[2] ),
    .o(net856));
 b15nandp2as1n48x5 _20315_ (.a(net444),
    .b(net441),
    .o1(_11643_));
 b15nor002as1n24x5 _20316_ (.a(_11575_),
    .b(_11643_),
    .o1(_11644_));
 b15bfn001as1n64x5 max_length855 (.a(\us30.a[2] ),
    .o(net855));
 b15nand02as1n48x5 _20318_ (.a(\u0.tmp_w[18] ),
    .b(net451),
    .o1(_11646_));
 b15bfn001ah1n64x5 load_slew854 (.a(net855),
    .o(net854));
 b15oai022an1n02x5 _20320_ (.a(net456),
    .b(_11628_),
    .c(_11646_),
    .d(_11606_),
    .o1(_11648_));
 b15nanb02as1n24x5 _20321_ (.a(\u0.tmp_w[18] ),
    .b(net456),
    .out0(_11649_));
 b15bfn001ah1n64x5 wire853 (.a(net855),
    .o(net853));
 b15oaoi13as1n02x5 _20323_ (.a(_11579_),
    .b(_11649_),
    .c(_11646_),
    .d(net456),
    .o1(_11651_));
 b15oai012ar1n08x5 _20324_ (.a(_11644_),
    .b(_11648_),
    .c(_11651_),
    .o1(_11652_));
 b15nandp2as1n04x5 _20325_ (.a(net457),
    .b(net450),
    .o1(_11653_));
 b15bfn001as1n64x5 max_length852 (.a(\us30.a[3] ),
    .o(net852));
 b15orn002ah1n08x5 _20327_ (.a(net458),
    .b(net446),
    .o(_11655_));
 b15oai112an1n08x5 _20328_ (.a(net461),
    .b(_11653_),
    .c(_11655_),
    .d(_11559_),
    .o1(_11656_));
 b15norp02al1n16x5 _20329_ (.a(net454),
    .b(net444),
    .o1(_11657_));
 b15bfn001as1n48x5 load_slew851 (.a(\us30.a[3] ),
    .o(net851));
 b15bfn001as1n64x5 max_length850 (.a(net851),
    .o(net850));
 b15nand03al1n12x5 _20332_ (.a(net448),
    .b(net437),
    .c(net434),
    .o1(_11660_));
 b15orn002al1n16x5 _20333_ (.a(net439),
    .b(net434),
    .o(_11661_));
 b15bfn001as1n64x5 max_length849 (.a(\us30.a[4] ),
    .o(net849));
 b15aoai13al1n08x5 _20335_ (.a(_11660_),
    .b(_11661_),
    .c(net448),
    .d(_11571_),
    .o1(_11663_));
 b15nand04an1n16x5 _20336_ (.a(net441),
    .b(_11656_),
    .c(_11657_),
    .d(_11663_),
    .o1(_11664_));
 b15xor002as1n16x5 _20337_ (.a(net458),
    .b(net452),
    .out0(_11665_));
 b15inv000ah1n64x5 _20338_ (.a(net449),
    .o1(_11666_));
 b15nonb02as1n16x5 _20339_ (.a(net458),
    .b(net453),
    .out0(_11667_));
 b15bfn001as1n64x5 max_length848 (.a(\us30.a[4] ),
    .o(net848));
 b15bfn001ah1n48x5 load_slew847 (.a(\us30.a[5] ),
    .o(net847));
 b15bfn001as1n48x5 load_slew846 (.a(net847),
    .o(net846));
 b15nona23ah1n32x5 _20343_ (.a(net446),
    .b(net438),
    .c(net436),
    .d(net442),
    .out0(_11671_));
 b15norp03ar1n02x5 _20344_ (.a(_11666_),
    .b(_11667_),
    .c(_11671_),
    .o1(_11672_));
 b15nand04as1n16x5 _20345_ (.a(net446),
    .b(net442),
    .c(net438),
    .d(net436),
    .o1(_11673_));
 b15and002an1n16x5 _20346_ (.a(net460),
    .b(net454),
    .o(_11674_));
 b15norp03an1n02x5 _20347_ (.a(net450),
    .b(_11673_),
    .c(_11674_),
    .o1(_11675_));
 b15oai022an1n02x5 _20348_ (.a(net461),
    .b(_11665_),
    .c(_11672_),
    .d(_11675_),
    .o1(_11676_));
 b15nand04as1n06x5 _20349_ (.a(_11641_),
    .b(_11652_),
    .c(_11664_),
    .d(_11676_),
    .o1(_11677_));
 b15inv020an1n28x5 _20350_ (.a(net434),
    .o1(_11678_));
 b15norp02as1n08x5 _20351_ (.a(net456),
    .b(net445),
    .o1(_11679_));
 b15bfn001ah1n64x5 load_slew845 (.a(\us30.a[6] ),
    .o(net845));
 b15nor004as1n02x5 _20353_ (.a(net460),
    .b(net451),
    .c(net440),
    .d(net437),
    .o1(_11681_));
 b15bfn001as1n48x5 load_slew844 (.a(\us30.a[6] ),
    .o(net844));
 b15and003ar1n02x5 _20355_ (.a(net451),
    .b(net440),
    .c(net437),
    .o(_11683_));
 b15oai112aq1n08x5 _20356_ (.a(_11678_),
    .b(_11679_),
    .c(_11681_),
    .d(_11683_),
    .o1(_11684_));
 b15nona23as1n32x5 _20357_ (.a(net446),
    .b(net436),
    .c(net438),
    .d(net442),
    .out0(_11685_));
 b15nandp2al1n12x5 _20358_ (.a(net460),
    .b(net451),
    .o1(_11686_));
 b15oaoi13as1n08x5 _20359_ (.a(net454),
    .b(_11684_),
    .c(_11685_),
    .d(_11686_),
    .o1(_11687_));
 b15nano23al1n08x5 _20360_ (.a(_11609_),
    .b(_11633_),
    .c(_11677_),
    .d(_11687_),
    .out0(_11688_));
 b15inv020aq1n32x5 _20361_ (.a(net440),
    .o1(_11689_));
 b15bfn001ah1n64x5 load_slew843 (.a(\us30.a[7] ),
    .o(net843));
 b15nonb02ah1n08x5 _20363_ (.a(net439),
    .b(net444),
    .out0(_11691_));
 b15nand04al1n02x5 _20364_ (.a(net450),
    .b(net434),
    .c(_11614_),
    .d(_11691_),
    .o1(_11692_));
 b15nandp2as1n24x5 _20365_ (.a(net458),
    .b(net446),
    .o1(_11693_));
 b15norp02ah1n32x5 _20366_ (.a(net460),
    .b(net454),
    .o1(_11694_));
 b15norp02ar1n02x5 _20367_ (.a(_11693_),
    .b(_11694_),
    .o1(_11695_));
 b15inv040as1n60x5 _20368_ (.a(net458),
    .o1(_11696_));
 b15bfn001ah1n64x5 wire842 (.a(\us01.a[0] ),
    .o(net842));
 b15bfn001ah1n64x5 max_length841 (.a(net842),
    .o(net841));
 b15nor002as1n04x5 _20371_ (.a(net460),
    .b(net444),
    .o1(_11699_));
 b15oaoi13an1n02x5 _20372_ (.a(_11695_),
    .b(_11696_),
    .c(_11603_),
    .d(_11699_),
    .o1(_11700_));
 b15oai013aq1n03x5 _20373_ (.a(_11692_),
    .b(_11700_),
    .c(net450),
    .d(_11575_),
    .o1(_11701_));
 b15nandp2ar1n08x5 _20374_ (.a(_11689_),
    .b(_11701_),
    .o1(_11702_));
 b15bfn001as1n48x5 load_slew840 (.a(\us01.a[0] ),
    .o(net840));
 b15nonb03ah1n03x5 _20376_ (.a(net436),
    .b(net438),
    .c(net442),
    .out0(_11704_));
 b15nand02ar1n32x5 _20377_ (.a(net455),
    .b(net454),
    .o1(_11705_));
 b15nanb02ah1n08x5 _20378_ (.a(net446),
    .b(net459),
    .out0(_11706_));
 b15aob012as1n03x5 _20379_ (.a(_11704_),
    .b(_11705_),
    .c(_11706_),
    .out0(_11707_));
 b15xnr002ar1n02x5 _20380_ (.a(net452),
    .b(net442),
    .out0(_11708_));
 b15bfn001ah1n64x5 wire839 (.a(\us01.a[1] ),
    .o(net839));
 b15nor003ah1n08x5 _20382_ (.a(\u0.tmp_w[20] ),
    .b(net438),
    .c(\u0.tmp_w[23] ),
    .o1(_11710_));
 b15xor002al1n03x5 _20383_ (.a(net459),
    .b(net452),
    .out0(_11711_));
 b15oai112as1n02x5 _20384_ (.a(_11708_),
    .b(_11710_),
    .c(net458),
    .d(_11711_),
    .o1(_11712_));
 b15nandp2ar1n16x5 _20385_ (.a(net445),
    .b(_11616_),
    .o1(_11713_));
 b15bfn001as1n64x5 max_length838 (.a(net839),
    .o(net838));
 b15oai112an1n06x5 _20387_ (.a(_11707_),
    .b(_11712_),
    .c(_11713_),
    .d(net452),
    .o1(_11715_));
 b15nona23as1n32x5 _20388_ (.a(net438),
    .b(\u0.tmp_w[23] ),
    .c(\u0.tmp_w[20] ),
    .d(net443),
    .out0(_11716_));
 b15bfn001ah1n48x5 load_slew837 (.a(net839),
    .o(net837));
 b15oai122aq1n08x5 _20390_ (.a(net459),
    .b(net458),
    .c(_11713_),
    .d(_11716_),
    .e(_11603_),
    .o1(_11718_));
 b15nanb03as1n16x5 _20391_ (.a(net443),
    .b(net438),
    .c(\u0.tmp_w[23] ),
    .out0(_11719_));
 b15oai122aq1n08x5 _20392_ (.a(_11579_),
    .b(_11693_),
    .c(_11719_),
    .d(_11716_),
    .e(net458),
    .o1(_11720_));
 b15aoai13an1n08x5 _20393_ (.a(net449),
    .b(_11715_),
    .c(_11718_),
    .d(_11720_),
    .o1(_11721_));
 b15nandp2as1n24x5 _20394_ (.a(net439),
    .b(net434),
    .o1(_11722_));
 b15oai013al1n02x5 _20395_ (.a(_11661_),
    .b(_11722_),
    .c(net460),
    .d(net444),
    .o1(_11723_));
 b15bfn001as1n48x5 load_slew836 (.a(net838),
    .o(net836));
 b15norp03an1n02x5 _20397_ (.a(net450),
    .b(net441),
    .c(_11649_),
    .o1(_11725_));
 b15nand04an1n02x5 _20398_ (.a(_11666_),
    .b(net434),
    .c(_11614_),
    .d(_11691_),
    .o1(_11726_));
 b15nonb02ah1n12x5 _20399_ (.a(net437),
    .b(net435),
    .out0(_11727_));
 b15nonb02as1n06x5 _20400_ (.a(net435),
    .b(net437),
    .out0(_11728_));
 b15nonb02al1n16x5 _20401_ (.a(net444),
    .b(net455),
    .out0(_11729_));
 b15aoi022ar1n02x5 _20402_ (.a(_11727_),
    .b(_11591_),
    .c(_11728_),
    .d(_11729_),
    .o1(_11730_));
 b15nanb02as1n24x5 _20403_ (.a(net459),
    .b(net452),
    .out0(_11731_));
 b15oai013as1n03x5 _20404_ (.a(_11726_),
    .b(_11730_),
    .c(_11731_),
    .d(_11666_),
    .o1(_11732_));
 b15aoi022as1n04x5 _20405_ (.a(_11723_),
    .b(_11725_),
    .c(_11732_),
    .d(net441),
    .o1(_11733_));
 b15nand03as1n04x5 _20406_ (.a(net455),
    .b(net444),
    .c(net441),
    .o1(_11734_));
 b15orn002al1n32x5 _20407_ (.a(net444),
    .b(net441),
    .o(_11735_));
 b15bfn001as1n64x5 max_length835 (.a(\us01.a[2] ),
    .o(net835));
 b15oaoi13ar1n04x5 _20409_ (.a(_11660_),
    .b(_11734_),
    .c(_11603_),
    .d(_11735_),
    .o1(_11737_));
 b15nor003ah1n02x5 _20410_ (.a(_11693_),
    .b(_11628_),
    .c(_11719_),
    .o1(_11738_));
 b15norp02ar1n48x5 _20411_ (.a(net458),
    .b(net449),
    .o1(_11739_));
 b15bfn001as1n64x5 max_length834 (.a(\us01.a[2] ),
    .o(net834));
 b15nanb02as1n24x5 _20413_ (.a(net445),
    .b(net440),
    .out0(_11741_));
 b15nor002as1n24x5 _20414_ (.a(_11741_),
    .b(_11722_),
    .o1(_11742_));
 b15aoi112al1n03x5 _20415_ (.a(_11737_),
    .b(_11738_),
    .c(_11739_),
    .d(_11742_),
    .o1(_11743_));
 b15norp03ah1n03x5 _20416_ (.a(_11559_),
    .b(_11635_),
    .c(_11655_),
    .o1(_11744_));
 b15nanb02ar1n24x5 _20417_ (.a(net435),
    .b(net441),
    .out0(_11745_));
 b15orn002ah1n08x5 _20418_ (.a(net448),
    .b(net444),
    .o(_11746_));
 b15norp02ar1n02x5 _20419_ (.a(_11745_),
    .b(_11746_),
    .o1(_11747_));
 b15nanb02as1n24x5 _20420_ (.a(net454),
    .b(net448),
    .out0(_11748_));
 b15nanb02ah1n16x5 _20421_ (.a(net435),
    .b(net447),
    .out0(_11749_));
 b15aoi112al1n06x5 _20422_ (.a(net443),
    .b(_11748_),
    .c(_11586_),
    .d(_11749_),
    .o1(_11750_));
 b15oaoi13al1n03x5 _20423_ (.a(_11744_),
    .b(net439),
    .c(_11747_),
    .d(_11750_),
    .o1(_11751_));
 b15mdn022aq1n04x5 _20424_ (.a(_11743_),
    .b(_11751_),
    .o1(_11752_),
    .sa(_11579_));
 b15nandp3ar1n02x5 _20425_ (.a(net460),
    .b(net443),
    .c(net435),
    .o1(_11753_));
 b15nanb03aq1n06x5 _20426_ (.a(net447),
    .b(net439),
    .c(net448),
    .out0(_11754_));
 b15bfn001as1n48x5 load_slew833 (.a(\us01.a[2] ),
    .o(net833));
 b15oaoi13ah1n02x5 _20428_ (.a(_11753_),
    .b(_11754_),
    .c(_11556_),
    .d(net439),
    .o1(_11756_));
 b15norp02as1n16x5 _20429_ (.a(_11597_),
    .b(_11643_),
    .o1(_11757_));
 b15aoai13ar1n03x5 _20430_ (.a(net454),
    .b(_11756_),
    .c(_11757_),
    .d(_11739_),
    .o1(_11758_));
 b15bfn001as1n64x5 max_length832 (.a(\us01.a[3] ),
    .o(net832));
 b15nanb02as1n24x5 _20432_ (.a(\u0.tmp_w[20] ),
    .b(net449),
    .out0(_11760_));
 b15bfn001as1n48x5 load_slew831 (.a(\us01.a[3] ),
    .o(net831));
 b15oai012ar1n08x5 _20434_ (.a(net454),
    .b(_11637_),
    .c(_11760_),
    .o1(_11762_));
 b15norp03ar1n08x5 _20435_ (.a(_11637_),
    .b(_11694_),
    .c(_11760_),
    .o1(_11763_));
 b15bfn001as1n48x5 wire830 (.a(net832),
    .o(net830));
 b15nor003al1n08x5 _20437_ (.a(net448),
    .b(_11597_),
    .c(_11643_),
    .o1(_11765_));
 b15and002an1n16x5 _20438_ (.a(net455),
    .b(net454),
    .o(_11766_));
 b15oaoi13aq1n04x5 _20439_ (.a(_11766_),
    .b(_11696_),
    .c(_11637_),
    .d(_11760_),
    .o1(_11767_));
 b15oai122as1n16x5 _20440_ (.a(_11762_),
    .b(_11763_),
    .c(_11765_),
    .d(_11579_),
    .e(_11767_),
    .o1(_11768_));
 b15bfn001as1n64x5 max_length829 (.a(\us01.a[4] ),
    .o(net829));
 b15nandp3as1n24x5 _20442_ (.a(net441),
    .b(net438),
    .c(net435),
    .o1(_11770_));
 b15nor002aq1n03x5 _20443_ (.a(_11565_),
    .b(_11770_),
    .o1(_11771_));
 b15nanb02aq1n24x5 _20444_ (.a(net449),
    .b(net458),
    .out0(_11772_));
 b15norp02ah1n12x5 _20445_ (.a(_11579_),
    .b(_11772_),
    .o1(_11773_));
 b15aoi012ah1n06x5 _20446_ (.a(_11771_),
    .b(_11773_),
    .c(_11742_),
    .o1(_11774_));
 b15oai112al1n08x5 _20447_ (.a(_11758_),
    .b(_11768_),
    .c(net454),
    .d(_11774_),
    .o1(_11775_));
 b15nano23an1n08x5 _20448_ (.a(_11721_),
    .b(_11733_),
    .c(_11752_),
    .d(_11775_),
    .out0(_11776_));
 b15nand04as1n16x5 _20449_ (.a(_11595_),
    .b(_11688_),
    .c(_11702_),
    .d(_11776_),
    .o1(_11777_));
 b15xor002aq1n06x5 _20450_ (.a(\u0.r0.out[24] ),
    .b(\u0.w[0][24] ),
    .out0(_11778_));
 b15qgbxo2an1n10x5 _20451_ (.a(_11777_),
    .b(_11778_),
    .out0(_11779_));
 b15xnr002al1n08x5 _20452_ (.a(\u0.w[1][24] ),
    .b(_11779_),
    .out0(_11780_));
 b15qgbxo2an1n05x5 _20453_ (.a(\u0.w[2][24] ),
    .b(_11780_),
    .out0(_11781_));
 b15xor002ar1n02x5 _20454_ (.a(\u0.tmp_w[24] ),
    .b(_11781_),
    .out0(_11782_));
 b15oai012ar1n02x5 _20455_ (.a(_11551_),
    .b(_11782_),
    .c(net945),
    .o1(_00369_));
 b15bfn001ah1n64x5 wire828 (.a(net829),
    .o(net828));
 b15nand02al1n08x5 _20457_ (.a(net129),
    .b(net46),
    .o1(_11784_));
 b15xnr002aq1n04x5 _20458_ (.a(\u0.r0.out[25] ),
    .b(\u0.w[0][25] ),
    .out0(_11785_));
 b15nanb02ah1n16x5 _20459_ (.a(net453),
    .b(net459),
    .out0(_11786_));
 b15nanb03as1n16x5 _20460_ (.a(net439),
    .b(net433),
    .c(net443),
    .out0(_11787_));
 b15nor003ar1n02x5 _20461_ (.a(_11786_),
    .b(_11760_),
    .c(_11787_),
    .o1(_11788_));
 b15aoi012al1n02x5 _20462_ (.a(_11788_),
    .b(_11667_),
    .c(_11624_),
    .o1(_11789_));
 b15norp02aq1n04x5 _20463_ (.a(net451),
    .b(_11649_),
    .o1(_11790_));
 b15nona23aq1n24x5 _20464_ (.a(net442),
    .b(net438),
    .c(net436),
    .d(net446),
    .out0(_11791_));
 b15oai012an1n02x5 _20465_ (.a(_11671_),
    .b(_11791_),
    .c(\u0.tmp_w[16] ),
    .o1(_11792_));
 b15oai022al1n02x5 _20466_ (.a(_11559_),
    .b(_11628_),
    .c(_11646_),
    .d(_11719_),
    .o1(_11793_));
 b15nor002ar1n02x5 _20467_ (.a(net446),
    .b(_11619_),
    .o1(_11794_));
 b15aoi022ar1n06x5 _20468_ (.a(_11790_),
    .b(_11792_),
    .c(_11793_),
    .d(_11794_),
    .o1(_11795_));
 b15nor002ah1n06x5 _20469_ (.a(_11661_),
    .b(_11643_),
    .o1(_11796_));
 b15aoi012ar1n02x5 _20470_ (.a(_11624_),
    .b(_11796_),
    .c(_11579_),
    .o1(_11797_));
 b15oai112aq1n08x5 _20471_ (.a(_11789_),
    .b(_11795_),
    .c(_11646_),
    .d(_11797_),
    .o1(_11798_));
 b15nandp3ar1n02x5 _20472_ (.a(net456),
    .b(net451),
    .c(net440),
    .o1(_11799_));
 b15orn002aq1n04x5 _20473_ (.a(net451),
    .b(net440),
    .o(_11800_));
 b15oai012aq1n04x5 _20474_ (.a(_11799_),
    .b(_11800_),
    .c(net456),
    .o1(_11801_));
 b15nand04ar1n12x5 _20475_ (.a(net445),
    .b(_11727_),
    .c(_11694_),
    .d(_11801_),
    .o1(_11802_));
 b15nanb03aq1n03x5 _20476_ (.a(net437),
    .b(net435),
    .c(net445),
    .out0(_11803_));
 b15aoi112ah1n04x5 _20477_ (.a(_11646_),
    .b(_11803_),
    .c(net440),
    .d(_11606_),
    .o1(_11804_));
 b15nanb02aq1n12x5 _20478_ (.a(net451),
    .b(net461),
    .out0(_11805_));
 b15oai022as1n02x5 _20479_ (.a(net440),
    .b(_11565_),
    .c(_11741_),
    .d(_11805_),
    .o1(_11806_));
 b15bfn001as1n64x5 max_length827 (.a(\us01.a[5] ),
    .o(net827));
 b15aoi013as1n03x5 _20481_ (.a(_11804_),
    .b(_11806_),
    .c(_11728_),
    .d(_11696_),
    .o1(_11808_));
 b15nand02ar1n12x5 _20482_ (.a(_11696_),
    .b(net440),
    .o1(_11809_));
 b15bfn001ah1n64x5 wire826 (.a(\us01.a[5] ),
    .o(net826));
 b15norp03as1n02x5 _20484_ (.a(net445),
    .b(_11597_),
    .c(_11748_),
    .o1(_11811_));
 b15mdn022an1n03x5 _20485_ (.a(_11661_),
    .b(_11722_),
    .o1(_11812_),
    .sa(net451));
 b15and002ah1n16x5 _20486_ (.a(net452),
    .b(\u0.tmp_w[20] ),
    .o(_11813_));
 b15aoi012ar1n06x5 _20487_ (.a(_11811_),
    .b(_11812_),
    .c(_11813_),
    .o1(_11814_));
 b15oai112al1n16x5 _20488_ (.a(_11802_),
    .b(_11808_),
    .c(_11809_),
    .d(_11814_),
    .o1(_11815_));
 b15aoi012aq1n02x5 _20489_ (.a(net450),
    .b(_11685_),
    .c(_11667_),
    .o1(_11816_));
 b15aoai13an1n03x5 _20490_ (.a(net461),
    .b(_11766_),
    .c(_11685_),
    .d(_11603_),
    .o1(_11817_));
 b15nor002as1n03x5 _20491_ (.a(net454),
    .b(_11571_),
    .o1(_11818_));
 b15oai112aq1n12x5 _20492_ (.a(_11816_),
    .b(_11817_),
    .c(_11624_),
    .d(_11818_),
    .o1(_11819_));
 b15bfn001as1n64x5 max_length825 (.a(\us01.a[6] ),
    .o(net825));
 b15nandp2an1n12x5 _20494_ (.a(net443),
    .b(net439),
    .o1(_11821_));
 b15nano23as1n05x5 _20495_ (.a(_11584_),
    .b(_11586_),
    .c(_11821_),
    .d(_11731_),
    .out0(_11822_));
 b15aoai13ah1n06x5 _20496_ (.a(_11666_),
    .b(_11822_),
    .c(_11757_),
    .d(_11618_),
    .o1(_11823_));
 b15aoi012ar1n02x5 _20497_ (.a(_11635_),
    .b(_11719_),
    .c(_11716_),
    .o1(_11824_));
 b15oai012al1n02x5 _20498_ (.a(_11643_),
    .b(_11735_),
    .c(net454),
    .o1(_11825_));
 b15and002ah1n04x5 _20499_ (.a(net455),
    .b(net450),
    .o(_11826_));
 b15and002ah1n16x5 _20500_ (.a(net438),
    .b(net436),
    .o(_11827_));
 b15qgbao4an1n05x5 _20501_ (.o1(_11828_),
    .a(_11824_),
    .b(_11825_),
    .c(_11826_),
    .d(_11827_));
 b15oai112ah1n12x5 _20502_ (.a(_11819_),
    .b(_11823_),
    .c(_11828_),
    .d(_11579_),
    .o1(_11829_));
 b15nor003ah1n06x5 _20503_ (.a(_11798_),
    .b(_11815_),
    .c(_11829_),
    .o1(_11830_));
 b15qgbno2an1n10x5 _20504_ (.a(_11575_),
    .b(_11735_),
    .o1(_11831_));
 b15aob012al1n02x5 _20505_ (.a(_11579_),
    .b(_11628_),
    .c(_11831_),
    .out0(_11832_));
 b15nano23as1n24x5 _20506_ (.a(net446),
    .b(net438),
    .c(net436),
    .d(net442),
    .out0(_11833_));
 b15qgbna2an1n10x5 _20507_ (.a(_11666_),
    .b(_11833_),
    .o1(_11834_));
 b15and003ar1n02x5 _20508_ (.a(net459),
    .b(net457),
    .c(_11834_),
    .o(_11835_));
 b15aoai13ar1n04x5 _20509_ (.a(net453),
    .b(_11835_),
    .c(_11571_),
    .d(net450),
    .o1(_11836_));
 b15nor002aq1n03x5 _20510_ (.a(net441),
    .b(_11575_),
    .o1(_11837_));
 b15nand04ar1n06x5 _20511_ (.a(net457),
    .b(net453),
    .c(_11613_),
    .d(_11837_),
    .o1(_11838_));
 b15nano22al1n24x5 _20512_ (.a(net442),
    .b(net438),
    .c(net436),
    .out0(_11839_));
 b15nanb02al1n06x5 _20513_ (.a(_11565_),
    .b(_11839_),
    .out0(_11840_));
 b15orn002ah1n12x5 _20514_ (.a(net456),
    .b(\u0.tmp_w[18] ),
    .o(_11841_));
 b15oai012al1n06x5 _20515_ (.a(_11838_),
    .b(_11840_),
    .c(_11841_),
    .o1(_11842_));
 b15oai112ah1n06x5 _20516_ (.a(_11832_),
    .b(_11836_),
    .c(_11842_),
    .d(_11831_),
    .o1(_11843_));
 b15aoai13al1n02x5 _20517_ (.a(net459),
    .b(_11644_),
    .c(_11742_),
    .d(net458),
    .o1(_11844_));
 b15aoi022al1n02x5 _20518_ (.a(net458),
    .b(_11644_),
    .c(_11742_),
    .d(_11571_),
    .o1(_11845_));
 b15aoi012aq1n04x5 _20519_ (.a(_11646_),
    .b(_11844_),
    .c(_11845_),
    .o1(_11846_));
 b15nor004as1n03x5 _20520_ (.a(net450),
    .b(_11575_),
    .c(_11643_),
    .d(_11786_),
    .o1(_11847_));
 b15norp02ah1n04x5 _20521_ (.a(_11846_),
    .b(_11847_),
    .o1(_11848_));
 b15nonb02ah1n08x5 _20522_ (.a(net444),
    .b(net439),
    .out0(_11849_));
 b15oai012ah1n04x5 _20523_ (.a(_11800_),
    .b(_11686_),
    .c(_11689_),
    .o1(_11850_));
 b15aoi013ah1n06x5 _20524_ (.a(net456),
    .b(net434),
    .c(_11849_),
    .d(_11850_),
    .o1(_11851_));
 b15aoi112ar1n02x5 _20525_ (.a(_11696_),
    .b(_11771_),
    .c(_11616_),
    .d(_11613_),
    .o1(_11852_));
 b15oai012as1n03x5 _20526_ (.a(net453),
    .b(_11851_),
    .c(_11852_),
    .o1(_11853_));
 b15nanb02aq1n24x5 _20527_ (.a(net438),
    .b(net442),
    .out0(_11854_));
 b15norp02an1n02x5 _20528_ (.a(_11854_),
    .b(_11565_),
    .o1(_11855_));
 b15nanb02al1n16x5 _20529_ (.a(net442),
    .b(net438),
    .out0(_11856_));
 b15nor003ar1n03x5 _20530_ (.a(net446),
    .b(_11856_),
    .c(_11772_),
    .o1(_11857_));
 b15oai112aq1n08x5 _20531_ (.a(net459),
    .b(net436),
    .c(_11855_),
    .d(_11857_),
    .o1(_11858_));
 b15bfn001as1n64x5 max_length824 (.a(\us01.a[6] ),
    .o(net824));
 b15nor002an1n06x5 _20533_ (.a(_11601_),
    .b(_11564_),
    .o1(_11860_));
 b15oai012ar1n02x5 _20534_ (.a(net457),
    .b(_11716_),
    .c(_11579_),
    .o1(_11861_));
 b15xor002an1n16x5 _20535_ (.a(net441),
    .b(net439),
    .out0(_11862_));
 b15nano22aq1n02x5 _20536_ (.a(_11678_),
    .b(_11862_),
    .c(_11565_),
    .out0(_11863_));
 b15aoi022as1n04x5 _20537_ (.a(_11739_),
    .b(_11860_),
    .c(_11861_),
    .d(_11863_),
    .o1(_11864_));
 b15oai022ar1n02x5 _20538_ (.a(_11601_),
    .b(_11854_),
    .c(_11655_),
    .d(_11856_),
    .o1(_11865_));
 b15aoi013an1n03x5 _20539_ (.a(_11638_),
    .b(_11865_),
    .c(_11666_),
    .d(net436),
    .o1(_11866_));
 b15oai112al1n12x5 _20540_ (.a(_11858_),
    .b(_11864_),
    .c(net459),
    .d(_11866_),
    .o1(_11867_));
 b15oai012ar1n12x5 _20541_ (.a(_11853_),
    .b(_11867_),
    .c(net453),
    .o1(_11868_));
 b15nand04ah1n12x5 _20542_ (.a(_11830_),
    .b(_11843_),
    .c(_11848_),
    .d(_11868_),
    .o1(_11869_));
 b15and002aq1n12x5 _20543_ (.a(net441),
    .b(net439),
    .o(_11870_));
 b15norp02as1n12x5 _20544_ (.a(net443),
    .b(net439),
    .o1(_11871_));
 b15aoi012ar1n02x5 _20545_ (.a(_11870_),
    .b(_11871_),
    .c(net461),
    .o1(_11872_));
 b15nona22al1n05x5 _20546_ (.a(net453),
    .b(net445),
    .c(net435),
    .out0(_11873_));
 b15oai122as1n02x5 _20547_ (.a(_11696_),
    .b(_11731_),
    .c(_11713_),
    .d(_11872_),
    .e(_11873_),
    .o1(_11874_));
 b15nand02ah1n06x5 _20548_ (.a(_11657_),
    .b(_11839_),
    .o1(_11875_));
 b15nona22as1n02x5 _20549_ (.a(net439),
    .b(net434),
    .c(net444),
    .out0(_11876_));
 b15nanb02an1n06x5 _20550_ (.a(net460),
    .b(net434),
    .out0(_11877_));
 b15oai013al1n12x5 _20551_ (.a(_11876_),
    .b(_11877_),
    .c(_11849_),
    .d(_11691_),
    .o1(_11878_));
 b15nand02an1n16x5 _20552_ (.a(net444),
    .b(net439),
    .o1(_11879_));
 b15oai012aq1n03x5 _20553_ (.a(_11879_),
    .b(_11597_),
    .c(net444),
    .o1(_11880_));
 b15aoi022ah1n08x5 _20554_ (.a(_11603_),
    .b(_11878_),
    .c(_11880_),
    .d(_11674_),
    .o1(_11881_));
 b15oai112al1n06x5 _20555_ (.a(net457),
    .b(_11875_),
    .c(_11881_),
    .d(net441),
    .o1(_11882_));
 b15nandp2al1n04x5 _20556_ (.a(_11874_),
    .b(_11882_),
    .o1(_11883_));
 b15bfn001as1n64x5 max_length823 (.a(\us01.a[7] ),
    .o(net823));
 b15nanb02ah1n16x5 _20558_ (.a(net458),
    .b(net453),
    .out0(_11885_));
 b15nonb02ar1n12x5 _20559_ (.a(net437),
    .b(net440),
    .out0(_11886_));
 b15nand02as1n04x5 _20560_ (.a(net445),
    .b(_11886_),
    .o1(_11887_));
 b15norp02ar1n02x5 _20561_ (.a(net447),
    .b(_11821_),
    .o1(_11888_));
 b15aoi012ar1n02x5 _20562_ (.a(_11888_),
    .b(_11871_),
    .c(net447),
    .o1(_11889_));
 b15oai022aq1n02x5 _20563_ (.a(_11885_),
    .b(_11887_),
    .c(_11889_),
    .d(_11696_),
    .o1(_11890_));
 b15aoi022aq1n08x5 _20564_ (.a(_11603_),
    .b(_11742_),
    .c(_11890_),
    .d(_11678_),
    .o1(_11891_));
 b15oai112as1n16x5 _20565_ (.a(net448),
    .b(_11883_),
    .c(_11891_),
    .d(net461),
    .o1(_11892_));
 b15nor002ah1n12x5 _20566_ (.a(net446),
    .b(_11629_),
    .o1(_11893_));
 b15norp02ar1n16x5 _20567_ (.a(net446),
    .b(_11559_),
    .o1(_11894_));
 b15norp03ar1n02x5 _20568_ (.a(\u0.tmp_w[17] ),
    .b(_11893_),
    .c(_11894_),
    .o1(_11895_));
 b15oai012ar1n02x5 _20569_ (.a(\u0.tmp_w[16] ),
    .b(net446),
    .c(_11629_),
    .o1(_11896_));
 b15oai013ar1n02x5 _20570_ (.a(_11896_),
    .b(_11742_),
    .c(_11894_),
    .d(\u0.tmp_w[16] ),
    .o1(_11897_));
 b15aoi112ar1n02x5 _20571_ (.a(_11603_),
    .b(_11895_),
    .c(_11897_),
    .d(\u0.tmp_w[17] ),
    .o1(_11898_));
 b15aoi022ar1n02x5 _20572_ (.a(_11893_),
    .b(_11667_),
    .c(_11813_),
    .d(_11593_),
    .o1(_11899_));
 b15oai012ar1n02x5 _20573_ (.a(_11579_),
    .b(_11696_),
    .c(_11716_),
    .o1(_11900_));
 b15nor002ar1n24x5 _20574_ (.a(_11601_),
    .b(_11719_),
    .o1(_11901_));
 b15oai012al1n02x5 _20575_ (.a(_11900_),
    .b(_11796_),
    .c(_11901_),
    .o1(_11902_));
 b15oai022an1n02x5 _20576_ (.a(\u0.tmp_w[16] ),
    .b(_11899_),
    .c(_11902_),
    .d(\u0.tmp_w[18] ),
    .o1(_11903_));
 b15orn003al1n04x5 _20577_ (.a(net451),
    .b(_11898_),
    .c(_11903_),
    .o(_11904_));
 b15aoi012al1n12x5 _20578_ (.a(_11869_),
    .b(_11892_),
    .c(_11904_),
    .o1(_11905_));
 b15xor002aq1n06x5 _20579_ (.a(_11785_),
    .b(_11905_),
    .out0(_11906_));
 b15xnr002as1n04x5 _20580_ (.a(\u0.w[1][25] ),
    .b(_11906_),
    .out0(_11907_));
 b15xor002ar1n02x5 _20581_ (.a(\u0.tmp_w[25] ),
    .b(\u0.w[2][25] ),
    .out0(_11908_));
 b15xor002ar1n02x5 _20582_ (.a(_11907_),
    .b(_11908_),
    .out0(_11909_));
 b15oai012al1n02x5 _20583_ (.a(_11784_),
    .b(_11909_),
    .c(net945),
    .o1(_00370_));
 b15nand02ar1n02x5 _20584_ (.a(net946),
    .b(net47),
    .o1(_11910_));
 b15and003ar1n02x5 _20585_ (.a(_11603_),
    .b(_11644_),
    .c(_11773_),
    .o(_11911_));
 b15orn002ah1n08x5 _20586_ (.a(_11629_),
    .b(_11746_),
    .o(_11912_));
 b15nano23ah1n24x5 _20587_ (.a(net443),
    .b(net435),
    .c(net439),
    .d(net447),
    .out0(_11913_));
 b15nor002aq1n08x5 _20588_ (.a(net450),
    .b(_11571_),
    .o1(_11914_));
 b15nand02ar1n02x5 _20589_ (.a(_11913_),
    .b(_11914_),
    .o1(_11915_));
 b15nanb02ah1n08x5 _20590_ (.a(net458),
    .b(net451),
    .out0(_11916_));
 b15oai112as1n02x5 _20591_ (.a(_11912_),
    .b(_11915_),
    .c(_11791_),
    .d(_11916_),
    .o1(_11917_));
 b15aoi012al1n04x5 _20592_ (.a(_11911_),
    .b(_11917_),
    .c(\u0.tmp_w[18] ),
    .o1(_11918_));
 b15norp02as1n08x5 _20593_ (.a(_11722_),
    .b(_11643_),
    .o1(_11919_));
 b15oai022al1n04x5 _20594_ (.a(net453),
    .b(_11854_),
    .c(_11885_),
    .d(_11856_),
    .o1(_11920_));
 b15norp02ar1n02x5 _20595_ (.a(net446),
    .b(net436),
    .o1(_11921_));
 b15aoi022an1n02x5 _20596_ (.a(_11667_),
    .b(_11919_),
    .c(_11920_),
    .d(_11921_),
    .o1(_11922_));
 b15norp02aq1n02x5 _20597_ (.a(_11805_),
    .b(_11922_),
    .o1(_11923_));
 b15nonb02ah1n16x5 _20598_ (.a(net450),
    .b(net444),
    .out0(_11924_));
 b15nand02as1n16x5 _20599_ (.a(_11924_),
    .b(_11839_),
    .o1(_11925_));
 b15nand02an1n32x5 _20600_ (.a(net461),
    .b(net453),
    .o1(_11926_));
 b15oaoi13an1n03x5 _20601_ (.a(net457),
    .b(_11912_),
    .c(_11925_),
    .d(_11926_),
    .o1(_11927_));
 b15nonb02ar1n12x5 _20602_ (.a(net449),
    .b(net453),
    .out0(_11928_));
 b15norp03ah1n03x5 _20603_ (.a(\u0.tmp_w[16] ),
    .b(_11574_),
    .c(_11928_),
    .o1(_11929_));
 b15oai012ar1n03x5 _20604_ (.a(_11757_),
    .b(_11790_),
    .c(_11929_),
    .o1(_11930_));
 b15aoi022aq1n08x5 _20605_ (.a(_11871_),
    .b(_11606_),
    .c(_11870_),
    .d(net457),
    .o1(_11931_));
 b15nandp2an1n08x5 _20606_ (.a(net446),
    .b(net436),
    .o1(_11932_));
 b15oai013an1n03x5 _20607_ (.a(_11930_),
    .b(_11931_),
    .c(_11748_),
    .d(_11932_),
    .o1(_11933_));
 b15norp03ar1n08x5 _20608_ (.a(_11923_),
    .b(_11927_),
    .c(_11933_),
    .o1(_11934_));
 b15nand03al1n02x5 _20609_ (.a(_11606_),
    .b(_11623_),
    .c(_11624_),
    .o1(_11935_));
 b15nanb02al1n06x5 _20610_ (.a(net459),
    .b(net451),
    .out0(_11936_));
 b15orn002al1n04x5 _20611_ (.a(net446),
    .b(net436),
    .o(_11937_));
 b15oa0022al1n04x5 _20612_ (.a(net451),
    .b(_11932_),
    .c(_11936_),
    .d(_11937_),
    .o(_11938_));
 b15inv000ar1n24x5 _20613_ (.a(net439),
    .o1(_11939_));
 b15nand02ah1n08x5 _20614_ (.a(_11689_),
    .b(_11939_),
    .o1(_11940_));
 b15oai013ah1n04x5 _20615_ (.a(_11935_),
    .b(_11938_),
    .c(_11649_),
    .d(_11940_),
    .o1(_11941_));
 b15oaoi13an1n04x5 _20616_ (.a(_11926_),
    .b(_11673_),
    .c(_11671_),
    .d(net456),
    .o1(_11942_));
 b15norp03an1n03x5 _20617_ (.a(\u0.tmp_w[18] ),
    .b(net446),
    .c(_11629_),
    .o1(_11943_));
 b15oaoi13an1n04x5 _20618_ (.a(_11941_),
    .b(net451),
    .c(_11942_),
    .d(_11943_),
    .o1(_11944_));
 b15aoi012ar1n02x5 _20619_ (.a(net442),
    .b(_11635_),
    .c(_11649_),
    .o1(_11945_));
 b15nor002ah1n06x5 _20620_ (.a(net459),
    .b(_11666_),
    .o1(_11946_));
 b15aoai13ar1n02x5 _20621_ (.a(_11827_),
    .b(_11945_),
    .c(_11946_),
    .d(_11667_),
    .o1(_11947_));
 b15oaoi13as1n02x5 _20622_ (.a(net446),
    .b(_11947_),
    .c(_11635_),
    .d(_11559_),
    .o1(_11948_));
 b15aoi122aq1n02x5 _20623_ (.a(\u0.tmp_w[16] ),
    .b(_11919_),
    .c(_11739_),
    .d(_11928_),
    .e(_11894_),
    .o1(_11949_));
 b15orn003ar1n02x5 _20624_ (.a(_11770_),
    .b(_11760_),
    .c(_11841_),
    .o(_11950_));
 b15aoi013ar1n04x5 _20625_ (.a(_11949_),
    .b(_11950_),
    .c(_11912_),
    .d(\u0.tmp_w[16] ),
    .o1(_11951_));
 b15nor002aq1n06x5 _20626_ (.a(_11696_),
    .b(net443),
    .o1(_11952_));
 b15aoai13an1n08x5 _20627_ (.a(_11952_),
    .b(_11710_),
    .c(_11827_),
    .d(net446),
    .o1(_11953_));
 b15and002as1n03x5 _20628_ (.a(net461),
    .b(net456),
    .o(_11954_));
 b15nor003aq1n03x5 _20629_ (.a(net437),
    .b(_11678_),
    .c(_11954_),
    .o1(_11955_));
 b15aoi012al1n08x5 _20630_ (.a(_11955_),
    .b(_11727_),
    .c(net461),
    .o1(_11956_));
 b15oaoi13as1n02x5 _20631_ (.a(_11635_),
    .b(_11953_),
    .c(_11956_),
    .d(_11643_),
    .o1(_11957_));
 b15nor003aq1n06x5 _20632_ (.a(_11948_),
    .b(_11951_),
    .c(_11957_),
    .o1(_11958_));
 b15nand04ar1n16x5 _20633_ (.a(_11918_),
    .b(_11934_),
    .c(_11944_),
    .d(_11958_),
    .o1(_11959_));
 b15nonb02an1n08x5 _20634_ (.a(net445),
    .b(net440),
    .out0(_11960_));
 b15aoai13ah1n03x5 _20635_ (.a(net460),
    .b(_11679_),
    .c(_11960_),
    .d(net456),
    .o1(_11961_));
 b15aoi012ar1n02x5 _20636_ (.a(net437),
    .b(_11809_),
    .c(_11961_),
    .o1(_11962_));
 b15norp02ar1n02x5 _20637_ (.a(_11606_),
    .b(_11735_),
    .o1(_11963_));
 b15oab012ar1n02x5 _20638_ (.a(net435),
    .b(_11962_),
    .c(_11963_),
    .out0(_11964_));
 b15orn002an1n08x5 _20639_ (.a(net461),
    .b(net456),
    .o(_11965_));
 b15aoai13ar1n02x5 _20640_ (.a(_11603_),
    .b(_11964_),
    .c(_11901_),
    .d(_11965_),
    .o1(_11966_));
 b15nandp2al1n03x5 _20641_ (.a(\u0.tmp_w[18] ),
    .b(_11618_),
    .o1(_11967_));
 b15nand02an1n16x5 _20642_ (.a(net445),
    .b(_11593_),
    .o1(_11968_));
 b15oaoi13aq1n03x5 _20643_ (.a(net451),
    .b(_11966_),
    .c(_11967_),
    .d(_11968_),
    .o1(_11969_));
 b15oai012ar1n02x5 _20644_ (.a(_11579_),
    .b(_11841_),
    .c(_11925_),
    .o1(_11970_));
 b15bfn001as1n48x5 load_slew822 (.a(\us01.a[7] ),
    .o(net822));
 b15oai022ar1n02x5 _20646_ (.a(_11685_),
    .b(_11646_),
    .c(_11760_),
    .d(_11787_),
    .o1(_11972_));
 b15aoi012ar1n02x5 _20647_ (.a(_11970_),
    .b(_11972_),
    .c(net455),
    .o1(_11973_));
 b15bfn001as1n64x5 max_length821 (.a(\us11.a[0] ),
    .o(net821));
 b15nandp3ar1n03x5 _20649_ (.a(_11666_),
    .b(_11665_),
    .c(_11833_),
    .o1(_11975_));
 b15oaoi13ar1n02x5 _20650_ (.a(_11685_),
    .b(_11635_),
    .c(_11666_),
    .d(_11649_),
    .o1(_11976_));
 b15and002as1n04x5 _20651_ (.a(net449),
    .b(net435),
    .o(_11977_));
 b15obai22ar1n16x5 _20652_ (.a(_11977_),
    .b(net441),
    .c(net448),
    .d(_11745_),
    .out0(_11978_));
 b15aoi013al1n03x5 _20653_ (.a(_11976_),
    .b(_11978_),
    .c(_11679_),
    .d(net437),
    .o1(_11979_));
 b15aoi013aq1n04x5 _20654_ (.a(_11973_),
    .b(_11975_),
    .c(_11979_),
    .d(net461),
    .o1(_11980_));
 b15nor003ah1n02x5 _20655_ (.a(net459),
    .b(_11556_),
    .c(_11559_),
    .o1(_11981_));
 b15aoai13an1n06x5 _20656_ (.a(net458),
    .b(_11981_),
    .c(_11936_),
    .d(_11742_),
    .o1(_11982_));
 b15nanb02as1n24x5 _20657_ (.a(_11741_),
    .b(_11827_),
    .out0(_11983_));
 b15oaoi13an1n08x5 _20658_ (.a(_11603_),
    .b(_11982_),
    .c(_11983_),
    .d(_11916_),
    .o1(_11984_));
 b15oab012ar1n02x5 _20659_ (.a(_11926_),
    .b(_11796_),
    .c(_11833_),
    .out0(_11985_));
 b15nor003ah1n03x5 _20660_ (.a(_11696_),
    .b(_11575_),
    .c(_11735_),
    .o1(_11986_));
 b15aoi012an1n02x5 _20661_ (.a(_11985_),
    .b(_11986_),
    .c(_11786_),
    .o1(_11987_));
 b15norp03ar1n02x5 _20662_ (.a(\u0.tmp_w[18] ),
    .b(_11618_),
    .c(_11968_),
    .o1(_11988_));
 b15aoi012al1n02x5 _20663_ (.a(_11988_),
    .b(_11644_),
    .c(_11619_),
    .o1(_11989_));
 b15nonb02ah1n03x5 _20664_ (.a(net440),
    .b(net437),
    .out0(_11990_));
 b15rm6013eq1n12x5 _20665_ (.a(net460),
    .b(net455),
    .c(_11678_),
    .carryb(_11991_));
 b15oai012an1n03x5 _20666_ (.a(_11809_),
    .b(_11606_),
    .c(net440),
    .o1(_11992_));
 b15aoi022aq1n06x5 _20667_ (.a(_11990_),
    .b(_11991_),
    .c(_11992_),
    .d(_11727_),
    .o1(_11993_));
 b15oai112ah1n06x5 _20668_ (.a(_11987_),
    .b(_11989_),
    .c(_11604_),
    .d(_11993_),
    .o1(_11994_));
 b15aoi112ah1n04x5 _20669_ (.a(_11980_),
    .b(_11984_),
    .c(net451),
    .d(_11994_),
    .o1(_11995_));
 b15nonb03as1n12x5 _20670_ (.a(net441),
    .b(net437),
    .c(net434),
    .out0(_11996_));
 b15nandp3al1n02x5 _20671_ (.a(_11613_),
    .b(_11996_),
    .c(_11674_),
    .o1(_11997_));
 b15oai013ah1n03x5 _20672_ (.a(_11997_),
    .b(_11770_),
    .c(_11556_),
    .d(_11603_),
    .o1(_11998_));
 b15nanb02an1n16x5 _20673_ (.a(net441),
    .b(net434),
    .out0(_11999_));
 b15oai012ah1n04x5 _20674_ (.a(_11999_),
    .b(_11745_),
    .c(net454),
    .o1(_12000_));
 b15aoi013aq1n08x5 _20675_ (.a(_11998_),
    .b(_12000_),
    .c(_11924_),
    .d(_11939_),
    .o1(_12001_));
 b15nanb02ar1n12x5 _20676_ (.a(net440),
    .b(net445),
    .out0(_12002_));
 b15oaoi13al1n02x5 _20677_ (.a(_12002_),
    .b(_11722_),
    .c(net455),
    .d(_11661_),
    .o1(_12003_));
 b15aoi013aq1n04x5 _20678_ (.a(_12003_),
    .b(_11996_),
    .c(_11591_),
    .d(net460),
    .o1(_12004_));
 b15aoai13ar1n02x5 _20679_ (.a(net451),
    .b(\u0.tmp_w[18] ),
    .c(_11901_),
    .d(_11965_),
    .o1(_12005_));
 b15oai022ar1n04x5 _20680_ (.a(net456),
    .b(_12001_),
    .c(_12004_),
    .d(_12005_),
    .o1(_12006_));
 b15aoi013aq1n02x5 _20681_ (.a(_11667_),
    .b(_11968_),
    .c(_12001_),
    .d(_11614_),
    .o1(_12007_));
 b15oai012al1n06x5 _20682_ (.a(_12006_),
    .b(_12007_),
    .c(_11579_),
    .o1(_12008_));
 b15nona23an1n16x5 _20683_ (.a(_11959_),
    .b(_11969_),
    .c(_11995_),
    .d(_12008_),
    .out0(_12009_));
 b15xor002ah1n08x5 _20684_ (.a(\u0.r0.out[26] ),
    .b(\u0.w[0][26] ),
    .out0(_12010_));
 b15xor002as1n08x5 _20685_ (.a(_12009_),
    .b(_12010_),
    .out0(_12011_));
 b15xnr002an1n08x5 _20686_ (.a(\u0.w[1][26] ),
    .b(_12011_),
    .out0(_12012_));
 b15xor003ar1n02x5 _20687_ (.a(\u0.tmp_w[26] ),
    .b(\u0.w[2][26] ),
    .c(_12012_),
    .out0(_12013_));
 b15oai012ar1n03x5 _20688_ (.a(_11910_),
    .b(_12013_),
    .c(net946),
    .o1(_00371_));
 b15nand02as1n12x5 _20689_ (.a(net129),
    .b(net48),
    .o1(_12014_));
 b15oai013ar1n02x5 _20690_ (.a(_11579_),
    .b(net457),
    .c(_11635_),
    .d(_11671_),
    .o1(_12015_));
 b15norp02as1n03x5 _20691_ (.a(_11629_),
    .b(_11760_),
    .o1(_12016_));
 b15aoi012an1n02x5 _20692_ (.a(_12015_),
    .b(_12016_),
    .c(net457),
    .o1(_12017_));
 b15nandp2ar1n02x5 _20693_ (.a(net457),
    .b(_11833_),
    .o1(_12018_));
 b15aoi012ar1n04x5 _20694_ (.a(net450),
    .b(_11875_),
    .c(_12018_),
    .o1(_12019_));
 b15oai012ar1n04x5 _20695_ (.a(\u0.tmp_w[16] ),
    .b(_11671_),
    .c(_11772_),
    .o1(_12020_));
 b15aoi112aq1n03x5 _20696_ (.a(_12019_),
    .b(_12020_),
    .c(_11614_),
    .d(_12016_),
    .o1(_12021_));
 b15nandp2al1n12x5 _20697_ (.a(_11996_),
    .b(_11679_),
    .o1(_12022_));
 b15oaoi13an1n08x5 _20698_ (.a(_12017_),
    .b(_12021_),
    .c(_11646_),
    .d(_12022_),
    .o1(_12023_));
 b15oaoi13ar1n04x5 _20699_ (.a(_11660_),
    .b(_11735_),
    .c(_11643_),
    .d(_11674_),
    .o1(_12024_));
 b15oaoi13an1n04x5 _20700_ (.a(_11722_),
    .b(_11734_),
    .c(net455),
    .d(_11735_),
    .o1(_12025_));
 b15oai013an1n12x5 _20701_ (.a(_12024_),
    .b(_12025_),
    .c(_11766_),
    .d(net460),
    .o1(_12026_));
 b15orn002ar1n02x5 _20702_ (.a(net456),
    .b(net440),
    .o(_12027_));
 b15orn002ah1n08x5 _20703_ (.a(net445),
    .b(net437),
    .o(_12028_));
 b15oaoi13ar1n02x5 _20704_ (.a(_12027_),
    .b(_12028_),
    .c(_11603_),
    .d(_11879_),
    .o1(_12029_));
 b15nonb02al1n03x5 _20705_ (.a(net445),
    .b(net454),
    .out0(_12030_));
 b15aoi012ar1n02x5 _20706_ (.a(_12029_),
    .b(_11870_),
    .c(_12030_),
    .o1(_12031_));
 b15and003ar1n03x5 _20707_ (.a(net456),
    .b(net444),
    .c(net434),
    .o(_12032_));
 b15aoi022ah1n08x5 _20708_ (.a(_11593_),
    .b(_11699_),
    .c(_11862_),
    .d(_12032_),
    .o1(_12033_));
 b15oai122aq1n16x5 _20709_ (.a(net451),
    .b(_11983_),
    .c(_11841_),
    .d(_12033_),
    .e(_11603_),
    .o1(_12034_));
 b15nona22aq1n05x5 _20710_ (.a(_12031_),
    .b(_11877_),
    .c(_12034_),
    .out0(_12035_));
 b15oai022ar1n02x5 _20711_ (.a(_11603_),
    .b(_11716_),
    .c(_11746_),
    .d(_11719_),
    .o1(_12036_));
 b15nand02ar1n02x5 _20712_ (.a(_11571_),
    .b(_12036_),
    .o1(_12037_));
 b15nona23al1n32x5 _20713_ (.a(net446),
    .b(net442),
    .c(net438),
    .d(net436),
    .out0(_12038_));
 b15norp03ar1n02x5 _20714_ (.a(net450),
    .b(_11786_),
    .c(_12038_),
    .o1(_12039_));
 b15aoi013an1n02x5 _20715_ (.a(_12039_),
    .b(_11739_),
    .c(_11674_),
    .d(_11624_),
    .o1(_12040_));
 b15aoi012ar1n02x5 _20716_ (.a(_11638_),
    .b(_11860_),
    .c(_11571_),
    .o1(_12041_));
 b15oai022ar1n02x5 _20717_ (.a(net450),
    .b(_11671_),
    .c(_11760_),
    .d(_11629_),
    .o1(_12042_));
 b15nor002ah1n16x5 _20718_ (.a(net458),
    .b(net452),
    .o1(_12043_));
 b15oaoi13al1n02x5 _20719_ (.a(_11791_),
    .b(_11579_),
    .c(_11574_),
    .d(_12043_),
    .o1(_12044_));
 b15aoai13al1n02x5 _20720_ (.a(_11603_),
    .b(_11739_),
    .c(_11826_),
    .d(net461),
    .o1(_12045_));
 b15aoi022ar1n02x5 _20721_ (.a(_11667_),
    .b(_12042_),
    .c(_12044_),
    .d(_12045_),
    .o1(_12046_));
 b15andc04as1n04x5 _20722_ (.a(_12037_),
    .b(_12040_),
    .c(_12041_),
    .d(_12046_),
    .o(_12047_));
 b15nor004an1n02x5 _20723_ (.a(net460),
    .b(net450),
    .c(net434),
    .d(_11735_),
    .o1(_12048_));
 b15mdn022al1n04x5 _20724_ (.a(_11603_),
    .b(_11766_),
    .o1(_12049_),
    .sa(net437));
 b15obai22ah1n06x5 _20725_ (.a(_12048_),
    .b(_12049_),
    .c(_11705_),
    .d(_11925_),
    .out0(_12050_));
 b15xor002as1n12x5 _20726_ (.a(net460),
    .b(net456),
    .out0(_12051_));
 b15nor003as1n04x5 _20727_ (.a(_11678_),
    .b(_11643_),
    .c(_12051_),
    .o1(_12052_));
 b15nandp2ar1n02x5 _20728_ (.a(net437),
    .b(_11574_),
    .o1(_12053_));
 b15oai012al1n06x5 _20729_ (.a(_12053_),
    .b(_11748_),
    .c(net437),
    .o1(_12054_));
 b15aoi022aq1n02x5 _20730_ (.a(_11574_),
    .b(_11960_),
    .c(_11924_),
    .d(net440),
    .o1(_12055_));
 b15oai022ah1n06x5 _20731_ (.a(_11649_),
    .b(_11968_),
    .c(_12055_),
    .d(_11575_),
    .o1(_12056_));
 b15aoi122al1n08x5 _20732_ (.a(_12050_),
    .b(_12052_),
    .c(_12054_),
    .d(net460),
    .e(_12056_),
    .o1(_12057_));
 b15nand04ah1n16x5 _20733_ (.a(_12026_),
    .b(_12035_),
    .c(_12047_),
    .d(_12057_),
    .o1(_12058_));
 b15nand02ah1n02x5 _20734_ (.a(net440),
    .b(net434),
    .o1(_12059_));
 b15mdn022al1n02x5 _20735_ (.a(_11691_),
    .b(_11849_),
    .o1(_12060_),
    .sa(_11603_));
 b15norp02as1n03x5 _20736_ (.a(net437),
    .b(net434),
    .o1(_12061_));
 b15aoi022ar1n04x5 _20737_ (.a(net444),
    .b(_11827_),
    .c(_11657_),
    .d(_12061_),
    .o1(_12062_));
 b15nand02ar1n02x5 _20738_ (.a(net455),
    .b(_11689_),
    .o1(_12063_));
 b15oai022as1n02x5 _20739_ (.a(_12059_),
    .b(_12060_),
    .c(_12062_),
    .d(_12063_),
    .o1(_12064_));
 b15aoi012ah1n06x5 _20740_ (.a(_12034_),
    .b(_12064_),
    .c(net460),
    .o1(_12065_));
 b15oai022al1n02x5 _20741_ (.a(_11693_),
    .b(_11821_),
    .c(_11706_),
    .d(_11940_),
    .o1(_12066_));
 b15aoi013al1n03x5 _20742_ (.a(net450),
    .b(net435),
    .c(_12066_),
    .d(_11603_),
    .o1(_12067_));
 b15aoi012ar1n04x5 _20743_ (.a(_11894_),
    .b(_11901_),
    .c(_11885_),
    .o1(_12068_));
 b15nandp2aq1n03x5 _20744_ (.a(\u0.tmp_w[16] ),
    .b(_11649_),
    .o1(_12069_));
 b15oaoi13ar1n08x5 _20745_ (.a(_12065_),
    .b(_12067_),
    .c(_12068_),
    .d(_12069_),
    .o1(_12070_));
 b15nandp2an1n03x5 _20746_ (.a(net461),
    .b(net443),
    .o1(_12071_));
 b15nor002aq1n03x5 _20747_ (.a(_11575_),
    .b(_12071_),
    .o1(_12072_));
 b15oai012ar1n02x5 _20748_ (.a(_11885_),
    .b(_11649_),
    .c(_11601_),
    .o1(_12073_));
 b15aoi012al1n04x5 _20749_ (.a(_11694_),
    .b(_11614_),
    .c(net461),
    .o1(_12074_));
 b15aoi022ar1n02x5 _20750_ (.a(_12072_),
    .b(_12073_),
    .c(_12074_),
    .d(_11757_),
    .o1(_12075_));
 b15nor004ar1n03x5 _20751_ (.a(net461),
    .b(_11741_),
    .c(_11722_),
    .d(_12043_),
    .o1(_12076_));
 b15oai022ar1n02x5 _20752_ (.a(_11655_),
    .b(_11770_),
    .c(_11705_),
    .d(_11716_),
    .o1(_12077_));
 b15aoi112aq1n02x5 _20753_ (.a(net450),
    .b(_12076_),
    .c(_12077_),
    .d(net461),
    .o1(_12078_));
 b15orn002aq1n12x5 _20754_ (.a(net441),
    .b(net434),
    .o(_12079_));
 b15oaoi13an1n04x5 _20755_ (.a(_11601_),
    .b(_11939_),
    .c(_11614_),
    .d(_11694_),
    .o1(_12080_));
 b15nanb02as1n02x5 _20756_ (.a(net455),
    .b(net439),
    .out0(_12081_));
 b15aoi013al1n06x5 _20757_ (.a(net444),
    .b(_12081_),
    .c(net460),
    .d(_11603_),
    .o1(_12082_));
 b15oai012an1n06x5 _20758_ (.a(net439),
    .b(_11618_),
    .c(_11614_),
    .o1(_12083_));
 b15aoi112ah1n08x5 _20759_ (.a(_12079_),
    .b(_12080_),
    .c(_12082_),
    .d(_12083_),
    .o1(_12084_));
 b15orn003ar1n02x5 _20760_ (.a(_11575_),
    .b(_11643_),
    .c(_11731_),
    .o(_12085_));
 b15aoi012al1n04x5 _20761_ (.a(_11696_),
    .b(_11875_),
    .c(_12085_),
    .o1(_12086_));
 b15nano23al1n08x5 _20762_ (.a(_12075_),
    .b(_12078_),
    .c(_12084_),
    .d(_12086_),
    .out0(_12087_));
 b15oai012ar1n02x5 _20763_ (.a(\u0.tmp_w[16] ),
    .b(_11696_),
    .c(_11983_),
    .o1(_12088_));
 b15oai112an1n04x5 _20764_ (.a(net454),
    .b(_12088_),
    .c(_11831_),
    .d(_11742_),
    .o1(_12089_));
 b15nona23ar1n02x5 _20765_ (.a(net445),
    .b(net437),
    .c(net435),
    .d(net456),
    .out0(_12090_));
 b15oai013ar1n04x5 _20766_ (.a(_12090_),
    .b(_11954_),
    .c(_11575_),
    .d(_11601_),
    .o1(_12091_));
 b15and003ar1n02x5 _20767_ (.a(net440),
    .b(_11694_),
    .c(_12091_),
    .o(_12092_));
 b15nor003ar1n06x5 _20768_ (.a(_11575_),
    .b(_11735_),
    .c(_11841_),
    .o1(_12093_));
 b15aoi013ar1n02x5 _20769_ (.a(_12093_),
    .b(_12091_),
    .c(net440),
    .d(\u0.tmp_w[18] ),
    .o1(_12094_));
 b15oab012ah1n04x5 _20770_ (.a(_12092_),
    .b(_12094_),
    .c(_11579_),
    .out0(_12095_));
 b15aoi013an1n04x5 _20771_ (.a(_12087_),
    .b(_12089_),
    .c(_12095_),
    .d(net451),
    .o1(_12096_));
 b15nor004as1n12x5 _20772_ (.a(_12023_),
    .b(_12058_),
    .c(_12070_),
    .d(_12096_),
    .o1(_12097_));
 b15xnr002ar1n16x5 _20773_ (.a(\u0.r0.out[27] ),
    .b(\u0.w[0][27] ),
    .out0(_12098_));
 b15xor002as1n06x5 _20774_ (.a(_12097_),
    .b(_12098_),
    .out0(_12099_));
 b15xnr002ar1n12x5 _20775_ (.a(\u0.w[1][27] ),
    .b(_12099_),
    .out0(_12100_));
 b15xor002aq1n08x5 _20776_ (.a(\u0.w[2][27] ),
    .b(_12100_),
    .out0(_12101_));
 b15xor002ar1n02x5 _20777_ (.a(\u0.tmp_w[27] ),
    .b(_12101_),
    .out0(_12102_));
 b15oai012ar1n02x5 _20778_ (.a(_12014_),
    .b(_12102_),
    .c(net942),
    .o1(_00372_));
 b15nand02ar1n02x5 _20779_ (.a(net944),
    .b(net49),
    .o1(_12103_));
 b15xor002an1n16x5 _20780_ (.a(\u0.r0.out[28] ),
    .b(\u0.w[0][28] ),
    .out0(_12104_));
 b15aoi122ar1n02x5 _20781_ (.a(net459),
    .b(_11696_),
    .c(_11624_),
    .d(_11813_),
    .e(_11593_),
    .o1(_12105_));
 b15nand02ar1n02x5 _20782_ (.a(net452),
    .b(_11624_),
    .o1(_12106_));
 b15nandp3ar1n02x5 _20783_ (.a(net446),
    .b(_11593_),
    .c(_12043_),
    .o1(_12107_));
 b15aoi013an1n02x5 _20784_ (.a(_12105_),
    .b(_12106_),
    .c(_12107_),
    .d(net459),
    .o1(_12108_));
 b15nand02ar1n02x5 _20785_ (.a(_11833_),
    .b(_12043_),
    .o1(_12109_));
 b15oai112ar1n04x5 _20786_ (.a(_11666_),
    .b(_12109_),
    .c(_12038_),
    .d(_11731_),
    .o1(_12110_));
 b15nand02as1n02x5 _20787_ (.a(net459),
    .b(_11667_),
    .o1(_12111_));
 b15oaoi13an1n02x5 _20788_ (.a(_11685_),
    .b(_12111_),
    .c(_11665_),
    .d(net459),
    .o1(_12112_));
 b15oai022ah1n02x5 _20789_ (.a(_11666_),
    .b(_12108_),
    .c(_12110_),
    .d(_12112_),
    .o1(_12113_));
 b15nand02ar1n02x5 _20790_ (.a(net449),
    .b(_11871_),
    .o1(_12114_));
 b15nanb03as1n04x5 _20791_ (.a(net449),
    .b(net443),
    .c(net439),
    .out0(_12115_));
 b15aoi112al1n02x5 _20792_ (.a(net447),
    .b(_11926_),
    .c(_12114_),
    .d(_12115_),
    .o1(_12116_));
 b15nand02ar1n02x5 _20793_ (.a(_11579_),
    .b(\u0.tmp_w[22] ),
    .o1(_12117_));
 b15oai022an1n02x5 _20794_ (.a(\u0.tmp_w[22] ),
    .b(_11760_),
    .c(_12117_),
    .d(_11556_),
    .o1(_12118_));
 b15aoai13as1n03x5 _20795_ (.a(net435),
    .b(_12116_),
    .c(_12118_),
    .d(_11952_),
    .o1(_12119_));
 b15nor003aq1n03x5 _20796_ (.a(_11559_),
    .b(_11646_),
    .c(_11729_),
    .o1(_12120_));
 b15nand02al1n06x5 _20797_ (.a(net460),
    .b(_11678_),
    .o1(_12121_));
 b15aoi012ar1n04x5 _20798_ (.a(_12121_),
    .b(net437),
    .c(net455),
    .o1(_12122_));
 b15aoi013an1n08x5 _20799_ (.a(_12120_),
    .b(_12122_),
    .c(_11960_),
    .d(_11574_),
    .o1(_12123_));
 b15aoi012aq1n06x5 _20800_ (.a(_11754_),
    .b(_11999_),
    .c(_11745_),
    .o1(_12124_));
 b15oai022ar1n02x5 _20801_ (.a(_11685_),
    .b(_11731_),
    .c(_12038_),
    .d(_11649_),
    .o1(_12125_));
 b15aoai13an1n02x5 _20802_ (.a(_12124_),
    .b(_12125_),
    .c(_11705_),
    .d(net459),
    .o1(_12126_));
 b15nand04an1n06x5 _20803_ (.a(_12113_),
    .b(_12119_),
    .c(_12123_),
    .d(_12126_),
    .o1(_12127_));
 b15oaoi13aq1n08x5 _20804_ (.a(_11579_),
    .b(_11996_),
    .c(_11729_),
    .d(_11591_),
    .o1(_12128_));
 b15nor004an1n02x5 _20805_ (.a(net445),
    .b(_11559_),
    .c(_11748_),
    .d(_12128_),
    .o1(_12129_));
 b15norp02ar1n02x5 _20806_ (.a(net459),
    .b(net435),
    .o1(_12130_));
 b15oai112ar1n04x5 _20807_ (.a(_11871_),
    .b(_11813_),
    .c(_11977_),
    .d(_12130_),
    .o1(_12131_));
 b15oai112ar1n04x5 _20808_ (.a(_11696_),
    .b(_12131_),
    .c(_11713_),
    .d(_11628_),
    .o1(_12132_));
 b15aoi013aq1n02x5 _20809_ (.a(_11696_),
    .b(_11666_),
    .c(_11913_),
    .d(_11674_),
    .o1(_12133_));
 b15nand03an1n02x5 _20810_ (.a(_11556_),
    .b(_11694_),
    .c(_11760_),
    .o1(_12134_));
 b15oai012an1n06x5 _20811_ (.a(_12133_),
    .b(_12134_),
    .c(_11787_),
    .o1(_12135_));
 b15nano23as1n16x5 _20812_ (.a(net446),
    .b(net436),
    .c(net438),
    .d(net442),
    .out0(_12136_));
 b15aoi012ar1n02x5 _20813_ (.a(_12136_),
    .b(_11628_),
    .c(_11833_),
    .o1(_12137_));
 b15oaoi13ar1n02x5 _20814_ (.a(net459),
    .b(_11628_),
    .c(_11646_),
    .d(_11833_),
    .o1(_12138_));
 b15aoi012ar1n02x5 _20815_ (.a(_11926_),
    .b(_12136_),
    .c(net448),
    .o1(_12139_));
 b15aoi112an1n02x5 _20816_ (.a(_12137_),
    .b(_12138_),
    .c(_12139_),
    .d(_11834_),
    .o1(_12140_));
 b15oai022ar1n02x5 _20817_ (.a(_12129_),
    .b(_12132_),
    .c(_12135_),
    .d(_12140_),
    .o1(_12141_));
 b15norp02ar1n02x5 _20818_ (.a(net459),
    .b(_11854_),
    .o1(_12142_));
 b15oai012aq1n08x5 _20819_ (.a(_11937_),
    .b(_11649_),
    .c(_11932_),
    .o1(_12143_));
 b15aoi022ar1n06x5 _20820_ (.a(_11813_),
    .b(_11839_),
    .c(_12142_),
    .d(_12143_),
    .o1(_12144_));
 b15oai022ar1n02x5 _20821_ (.a(net459),
    .b(_11575_),
    .c(_11597_),
    .d(_11926_),
    .o1(_12145_));
 b15aoai13ar1n02x5 _20822_ (.a(net441),
    .b(_11710_),
    .c(_12145_),
    .d(net446),
    .o1(_12146_));
 b15nand02as1n02x5 _20823_ (.a(_11616_),
    .b(_11657_),
    .o1(_12147_));
 b15aoai13ar1n02x5 _20824_ (.a(_12144_),
    .b(net458),
    .c(_12146_),
    .d(_12147_),
    .o1(_12148_));
 b15aob012as1n02x5 _20825_ (.a(_12141_),
    .b(_12148_),
    .c(_11666_),
    .out0(_12149_));
 b15oai013aq1n02x5 _20826_ (.a(_11696_),
    .b(_11741_),
    .c(_11722_),
    .d(_11748_),
    .o1(_12150_));
 b15norp02aq1n02x5 _20827_ (.a(_11635_),
    .b(_11735_),
    .o1(_12151_));
 b15aoi013as1n04x5 _20828_ (.a(_12150_),
    .b(_12151_),
    .c(_12121_),
    .d(_11939_),
    .o1(_12152_));
 b15nandp2ar1n02x5 _20829_ (.a(_11579_),
    .b(_11603_),
    .o1(_12153_));
 b15oai012ar1n02x5 _20830_ (.a(net457),
    .b(_12153_),
    .c(_11912_),
    .o1(_12154_));
 b15oai022ar1n02x5 _20831_ (.a(_11666_),
    .b(_11713_),
    .c(_11983_),
    .d(_11628_),
    .o1(_12155_));
 b15oab012aq1n03x5 _20832_ (.a(_12152_),
    .b(_12154_),
    .c(_12155_),
    .out0(_12156_));
 b15aoi012ar1n02x5 _20833_ (.a(_11671_),
    .b(_11885_),
    .c(_11579_),
    .o1(_12157_));
 b15oai112ah1n02x5 _20834_ (.a(net448),
    .b(_12111_),
    .c(_12157_),
    .d(_11644_),
    .o1(_12158_));
 b15nand02ar1n02x5 _20835_ (.a(net454),
    .b(net440),
    .o1(_12159_));
 b15oai012ah1n03x5 _20836_ (.a(_12159_),
    .b(_11649_),
    .c(net440),
    .o1(_12160_));
 b15nand04aq1n12x5 _20837_ (.a(_12061_),
    .b(_11613_),
    .c(_11606_),
    .d(_12160_),
    .o1(_12161_));
 b15aoi022ar1n08x5 _20838_ (.a(_11837_),
    .b(_11924_),
    .c(_11914_),
    .d(_11624_),
    .o1(_12162_));
 b15oai112as1n06x5 _20839_ (.a(_12158_),
    .b(_12161_),
    .c(_12162_),
    .d(net453),
    .o1(_12163_));
 b15aoi022an1n06x5 _20840_ (.a(_11696_),
    .b(_11919_),
    .c(_11831_),
    .d(_11666_),
    .o1(_12164_));
 b15oai022as1n08x5 _20841_ (.a(_11565_),
    .b(_11770_),
    .c(_12164_),
    .d(net459),
    .o1(_12165_));
 b15aoi112al1n08x5 _20842_ (.a(_12156_),
    .b(_12163_),
    .c(_12165_),
    .d(net453),
    .o1(_12166_));
 b15nand02as1n03x5 _20843_ (.a(_11913_),
    .b(_11739_),
    .o1(_12167_));
 b15oaoi13aq1n03x5 _20844_ (.a(net453),
    .b(_12167_),
    .c(_12128_),
    .d(_11666_),
    .o1(_12168_));
 b15nand02ar1n02x5 _20845_ (.a(net453),
    .b(_11871_),
    .o1(_12169_));
 b15oaoi13an1n03x5 _20846_ (.a(_11586_),
    .b(_12169_),
    .c(_11821_),
    .d(net453),
    .o1(_12170_));
 b15nor003an1n08x5 _20847_ (.a(_11575_),
    .b(_11735_),
    .c(_11649_),
    .o1(_12171_));
 b15orn003ar1n04x5 _20848_ (.a(net448),
    .b(_12170_),
    .c(_12171_),
    .o(_12172_));
 b15nano23as1n06x5 _20849_ (.a(net438),
    .b(net436),
    .c(\u0.tmp_w[18] ),
    .d(net442),
    .out0(_12173_));
 b15aoi013ah1n06x5 _20850_ (.a(_12173_),
    .b(net436),
    .c(net442),
    .d(_11696_),
    .o1(_12174_));
 b15oai122as1n16x5 _20851_ (.a(net450),
    .b(_11602_),
    .c(_11770_),
    .d(_12174_),
    .e(_11601_),
    .o1(_12175_));
 b15aoai13aq1n08x5 _20852_ (.a(net459),
    .b(_12168_),
    .c(_12172_),
    .d(_12175_),
    .o1(_12176_));
 b15nona23aq1n24x5 _20853_ (.a(_12127_),
    .b(_12149_),
    .c(_12166_),
    .d(_12176_),
    .out0(_12177_));
 b15xor002as1n12x5 _20854_ (.a(_12104_),
    .b(_12177_),
    .out0(_12178_));
 b15xnr002an1n16x5 _20855_ (.a(\u0.w[1][28] ),
    .b(_12178_),
    .out0(_12179_));
 b15xor002as1n16x5 _20856_ (.a(\u0.w[2][28] ),
    .b(_12179_),
    .out0(_12180_));
 b15xor002ar1n02x5 _20857_ (.a(\u0.tmp_w[28] ),
    .b(_12180_),
    .out0(_12181_));
 b15oai012ar1n02x5 _20858_ (.a(_12103_),
    .b(_12181_),
    .c(net944),
    .o1(_00373_));
 b15nand02ar1n02x5 _20859_ (.a(net943),
    .b(net50),
    .o1(_12182_));
 b15xor002an1n12x5 _20860_ (.a(\u0.r0.out[29] ),
    .b(\u0.w[0][29] ),
    .out0(_12183_));
 b15nandp2an1n05x5 _20861_ (.a(net461),
    .b(net455),
    .o1(_12184_));
 b15aoi012ar1n02x5 _20862_ (.a(_11716_),
    .b(_12184_),
    .c(_11603_),
    .o1(_12185_));
 b15aoi112aq1n02x5 _20863_ (.a(_11666_),
    .b(_12185_),
    .c(_11894_),
    .d(_11603_),
    .o1(_12186_));
 b15oai022an1n02x5 _20864_ (.a(net445),
    .b(_11854_),
    .c(_11887_),
    .d(_12043_),
    .o1(_12187_));
 b15oab012as1n04x5 _20865_ (.a(net436),
    .b(_11711_),
    .c(_11696_),
    .out0(_12188_));
 b15aoi122aq1n04x5 _20866_ (.a(net450),
    .b(_11644_),
    .c(_11766_),
    .d(_12187_),
    .e(_12188_),
    .o1(_12189_));
 b15aoi012ar1n02x5 _20867_ (.a(_11689_),
    .b(net435),
    .c(_12184_),
    .o1(_12190_));
 b15aoi112al1n02x5 _20868_ (.a(_12028_),
    .b(_12190_),
    .c(_11991_),
    .d(_11689_),
    .o1(_12191_));
 b15aoai13al1n04x5 _20869_ (.a(_11603_),
    .b(_12191_),
    .c(_11644_),
    .d(_11619_),
    .o1(_12192_));
 b15aoi012aq1n04x5 _20870_ (.a(_12186_),
    .b(_12189_),
    .c(_12192_),
    .o1(_12193_));
 b15aoi022aq1n04x5 _20871_ (.a(net448),
    .b(_11710_),
    .c(_11739_),
    .d(_12136_),
    .o1(_12194_));
 b15oai012ar1n02x5 _20872_ (.a(_11719_),
    .b(_11559_),
    .c(net453),
    .o1(_12195_));
 b15aoi022as1n04x5 _20873_ (.a(_11623_),
    .b(_11839_),
    .c(_12195_),
    .d(_11666_),
    .o1(_12196_));
 b15oaoi13ah1n08x5 _20874_ (.a(net459),
    .b(_12194_),
    .c(_12196_),
    .d(_11693_),
    .o1(_12197_));
 b15aoi022an1n02x5 _20875_ (.a(net454),
    .b(_11691_),
    .c(_11849_),
    .d(net456),
    .o1(_12198_));
 b15oai013al1n04x5 _20876_ (.a(_11925_),
    .b(_12198_),
    .c(net434),
    .d(_11800_),
    .o1(_12199_));
 b15nandp2as1n08x5 _20877_ (.a(net460),
    .b(_12199_),
    .o1(_12200_));
 b15nano23aq1n08x5 _20878_ (.a(net438),
    .b(net436),
    .c(net446),
    .d(net442),
    .out0(_12201_));
 b15aoi112aq1n04x5 _20879_ (.a(net451),
    .b(_12173_),
    .c(_12201_),
    .d(_11619_),
    .o1(_12202_));
 b15aoai13as1n03x5 _20880_ (.a(_11618_),
    .b(_12201_),
    .c(_11913_),
    .d(\u0.tmp_w[18] ),
    .o1(_12203_));
 b15aoi012al1n04x5 _20881_ (.a(_11614_),
    .b(_11649_),
    .c(\u0.tmp_w[16] ),
    .o1(_12204_));
 b15oai112ar1n16x5 _20882_ (.a(_12202_),
    .b(_12203_),
    .c(_12204_),
    .d(_11673_),
    .o1(_12205_));
 b15aoai13aq1n04x5 _20883_ (.a(net451),
    .b(_11967_),
    .c(_11968_),
    .d(_11983_),
    .o1(_12206_));
 b15nand03al1n03x5 _20884_ (.a(net445),
    .b(_11593_),
    .c(_11614_),
    .o1(_12207_));
 b15oaoi13an1n04x5 _20885_ (.a(_11579_),
    .b(_12207_),
    .c(_11983_),
    .d(_11649_),
    .o1(_12208_));
 b15nand02an1n04x5 _20886_ (.a(_12030_),
    .b(_12051_),
    .o1(_12209_));
 b15oaoi13aq1n08x5 _20887_ (.a(_11629_),
    .b(_12209_),
    .c(_12051_),
    .d(_11602_),
    .o1(_12210_));
 b15oai013aq1n12x5 _20888_ (.a(_12205_),
    .b(_12206_),
    .c(_12208_),
    .d(_12210_),
    .o1(_12211_));
 b15oaoi13ar1n02x5 _20889_ (.a(_11565_),
    .b(_11787_),
    .c(_12079_),
    .d(net454),
    .o1(_12212_));
 b15oai012an1n04x5 _20890_ (.a(_12212_),
    .b(_11665_),
    .c(_11579_),
    .o1(_12213_));
 b15nor003as1n02x5 _20891_ (.a(net461),
    .b(_11673_),
    .c(_12043_),
    .o1(_12214_));
 b15aoai13as1n02x5 _20892_ (.a(net450),
    .b(_12214_),
    .c(_11818_),
    .d(_11893_),
    .o1(_12215_));
 b15norp02al1n02x5 _20893_ (.a(net461),
    .b(net450),
    .o1(_12216_));
 b15aoai13al1n06x5 _20894_ (.a(_12216_),
    .b(_12171_),
    .c(_11860_),
    .d(_11614_),
    .o1(_12217_));
 b15norp03an1n02x5 _20895_ (.a(_11575_),
    .b(_11686_),
    .c(_11643_),
    .o1(_12218_));
 b15aoai13al1n03x5 _20896_ (.a(_11614_),
    .b(_12218_),
    .c(_11666_),
    .d(_12136_),
    .o1(_12219_));
 b15nand04an1n08x5 _20897_ (.a(_12213_),
    .b(_12215_),
    .c(_12217_),
    .d(_12219_),
    .o1(_12220_));
 b15nor004ah1n02x5 _20898_ (.a(net434),
    .b(_11618_),
    .c(_11748_),
    .d(_11879_),
    .o1(_12221_));
 b15norp02ar1n03x5 _20899_ (.a(net450),
    .b(_11705_),
    .o1(_12222_));
 b15and002ar1n02x5 _20900_ (.a(net460),
    .b(net444),
    .o(_12223_));
 b15ao0022aq1n02x5 _20901_ (.a(_11727_),
    .b(_11699_),
    .c(_12223_),
    .d(_11728_),
    .o(_12224_));
 b15aoai13as1n04x5 _20902_ (.a(net441),
    .b(_12221_),
    .c(_12222_),
    .d(_12224_),
    .o1(_12225_));
 b15nor004an1n02x5 _20903_ (.a(_11618_),
    .b(_11999_),
    .c(_11748_),
    .d(_11879_),
    .o1(_12226_));
 b15nand02ar1n02x5 _20904_ (.a(_11616_),
    .b(_11924_),
    .o1(_12227_));
 b15oab012ah1n02x5 _20905_ (.a(_12226_),
    .b(_12227_),
    .c(_12074_),
    .out0(_12228_));
 b15nano23ar1n02x5 _20906_ (.a(_11745_),
    .b(_11999_),
    .c(_11653_),
    .d(_12028_),
    .out0(_12229_));
 b15aoi013an1n03x5 _20907_ (.a(_12229_),
    .b(_11739_),
    .c(_11742_),
    .d(_11926_),
    .o1(_12230_));
 b15nand04as1n08x5 _20908_ (.a(_11819_),
    .b(_12225_),
    .c(_12228_),
    .d(_12230_),
    .o1(_12231_));
 b15nano23al1n12x5 _20909_ (.a(_11768_),
    .b(_12211_),
    .c(_12220_),
    .d(_12231_),
    .out0(_12232_));
 b15nona23an1n32x5 _20910_ (.a(_12193_),
    .b(_12197_),
    .c(_12200_),
    .d(_12232_),
    .out0(_12233_));
 b15xor002as1n16x5 _20911_ (.a(_12183_),
    .b(_12233_),
    .out0(_12234_));
 b15xnr002as1n16x5 _20912_ (.a(\u0.w[1][29] ),
    .b(_12234_),
    .out0(_12235_));
 b15xor002as1n16x5 _20913_ (.a(\u0.w[2][29] ),
    .b(_12235_),
    .out0(_12236_));
 b15xor002ar1n02x5 _20914_ (.a(\u0.tmp_w[29] ),
    .b(_12236_),
    .out0(_12237_));
 b15oai012ar1n02x5 _20915_ (.a(_12182_),
    .b(_12237_),
    .c(net943),
    .o1(_00374_));
 b15nand02ar1n02x5 _20916_ (.a(net938),
    .b(net52),
    .o1(_12238_));
 b15xor002as1n06x5 _20917_ (.a(\u0.r0.out[30] ),
    .b(\u0.w[0][30] ),
    .out0(_12239_));
 b15oai112ah1n06x5 _20918_ (.a(_11579_),
    .b(_12167_),
    .c(_11748_),
    .d(_11713_),
    .o1(_12240_));
 b15oai012al1n06x5 _20919_ (.a(_11834_),
    .b(_11983_),
    .c(_11653_),
    .o1(_12241_));
 b15aoi022ar1n02x5 _20920_ (.a(net448),
    .b(_11871_),
    .c(_11613_),
    .d(_11870_),
    .o1(_12242_));
 b15nor003al1n03x5 _20921_ (.a(_11603_),
    .b(_11678_),
    .c(_12242_),
    .o1(_12243_));
 b15nor003aq1n02x5 _20922_ (.a(_11885_),
    .b(_11637_),
    .c(_11760_),
    .o1(_12244_));
 b15norp03aq1n02x5 _20923_ (.a(_11556_),
    .b(_11719_),
    .c(_11649_),
    .o1(_12245_));
 b15nor004ah1n04x5 _20924_ (.a(_12241_),
    .b(_12243_),
    .c(_12244_),
    .d(_12245_),
    .o1(_12246_));
 b15aoi012an1n04x5 _20925_ (.a(_11765_),
    .b(_11567_),
    .c(_11696_),
    .o1(_12247_));
 b15oai112ah1n12x5 _20926_ (.a(net461),
    .b(_12246_),
    .c(_12247_),
    .d(net454),
    .o1(_12248_));
 b15nand02al1n16x5 _20927_ (.a(_12240_),
    .b(_12248_),
    .o1(_12249_));
 b15oai012aq1n02x5 _20928_ (.a(_11932_),
    .b(_11937_),
    .c(_11696_),
    .o1(_12250_));
 b15nor002al1n02x5 _20929_ (.a(_11856_),
    .b(_11731_),
    .o1(_12251_));
 b15oai022ar1n02x5 _20930_ (.a(net453),
    .b(_11716_),
    .c(_12038_),
    .d(_11665_),
    .o1(_12252_));
 b15aoi022ar1n02x5 _20931_ (.a(_12250_),
    .b(_12251_),
    .c(_12252_),
    .d(net459),
    .o1(_12253_));
 b15aoi012ar1n02x5 _20932_ (.a(_11579_),
    .b(_11685_),
    .c(_12022_),
    .o1(_12254_));
 b15norp02ar1n02x5 _20933_ (.a(net458),
    .b(_11685_),
    .o1(_12255_));
 b15oai012ar1n02x5 _20934_ (.a(_11603_),
    .b(_12254_),
    .c(_12255_),
    .o1(_12256_));
 b15aob012aq1n04x5 _20935_ (.a(_11666_),
    .b(_12253_),
    .c(_12256_),
    .out0(_12257_));
 b15oai013al1n02x5 _20936_ (.a(net455),
    .b(_11629_),
    .c(_11628_),
    .d(_11706_),
    .o1(_12258_));
 b15oaoi13ah1n03x5 _20937_ (.a(_12258_),
    .b(_11894_),
    .c(_11574_),
    .d(_11928_),
    .o1(_12259_));
 b15oai013ar1n02x5 _20938_ (.a(_11696_),
    .b(net444),
    .c(_11559_),
    .d(_11646_),
    .o1(_12260_));
 b15oai022ar1n02x5 _20939_ (.a(_11565_),
    .b(_12059_),
    .c(_12079_),
    .d(_11746_),
    .o1(_12261_));
 b15aoi013an1n02x5 _20940_ (.a(_12260_),
    .b(_12261_),
    .c(_11674_),
    .d(net437),
    .o1(_12262_));
 b15oa0012as1n03x5 _20941_ (.a(_12262_),
    .b(_11685_),
    .c(_11635_),
    .o(_12263_));
 b15norp03an1n02x5 _20942_ (.a(_11689_),
    .b(_11575_),
    .c(_11602_),
    .o1(_12264_));
 b15oai022al1n02x5 _20943_ (.a(net450),
    .b(_11940_),
    .c(_11565_),
    .d(_11821_),
    .o1(_12265_));
 b15aoi013ah1n03x5 _20944_ (.a(_12264_),
    .b(_12265_),
    .c(_11603_),
    .d(net435),
    .o1(_12266_));
 b15oaoi13ar1n08x5 _20945_ (.a(_12259_),
    .b(_12263_),
    .c(_12266_),
    .d(\u0.tmp_w[16] ),
    .o1(_12267_));
 b15aoai13as1n02x5 _20946_ (.a(_11694_),
    .b(_12016_),
    .c(_11839_),
    .d(_11613_),
    .o1(_12268_));
 b15oai012ar1n02x5 _20947_ (.a(_11624_),
    .b(_11965_),
    .c(net454),
    .o1(_12269_));
 b15oai012aq1n03x5 _20948_ (.a(_12269_),
    .b(_11983_),
    .c(net457),
    .o1(_12270_));
 b15aoi012ah1n04x5 _20949_ (.a(_11941_),
    .b(_12270_),
    .c(_11666_),
    .o1(_12271_));
 b15norp03al1n03x5 _20950_ (.a(_11556_),
    .b(_11719_),
    .c(_12153_),
    .o1(_12272_));
 b15norp03ar1n04x5 _20951_ (.a(net453),
    .b(_11556_),
    .c(_11854_),
    .o1(_12273_));
 b15nor003aq1n03x5 _20952_ (.a(net445),
    .b(_11646_),
    .c(_11862_),
    .o1(_12274_));
 b15oaoi13an1n04x5 _20953_ (.a(_12272_),
    .b(net435),
    .c(_12273_),
    .d(_12274_),
    .o1(_12275_));
 b15oai112ah1n08x5 _20954_ (.a(_12268_),
    .b(_12271_),
    .c(net457),
    .d(_12275_),
    .o1(_12276_));
 b15nanb02ar1n02x5 _20955_ (.a(_11786_),
    .b(_11772_),
    .out0(_12277_));
 b15oai022ar1n02x5 _20956_ (.a(_11564_),
    .b(_11556_),
    .c(_11571_),
    .d(_11840_),
    .o1(_12278_));
 b15aoi012ar1n02x5 _20957_ (.a(_11687_),
    .b(_12277_),
    .c(_12278_),
    .o1(_12279_));
 b15aoi112ar1n02x5 _20958_ (.a(_12002_),
    .b(_11916_),
    .c(_11575_),
    .d(_11597_),
    .o1(_12280_));
 b15oab012ar1n02x5 _20959_ (.a(_12280_),
    .b(_11912_),
    .c(_11731_),
    .out0(_12281_));
 b15oai112al1n02x5 _20960_ (.a(_11616_),
    .b(_11924_),
    .c(_12043_),
    .d(_11579_),
    .o1(_12282_));
 b15oai112ah1n04x5 _20961_ (.a(_11705_),
    .b(_12282_),
    .c(_11787_),
    .d(_11565_),
    .o1(_12283_));
 b15nand02ar1n02x5 _20962_ (.a(net448),
    .b(_11593_),
    .o1(_12284_));
 b15oaoi13an1n03x5 _20963_ (.a(_11601_),
    .b(_12284_),
    .c(_11770_),
    .d(net448),
    .o1(_12285_));
 b15oai012ar1n08x5 _20964_ (.a(_12283_),
    .b(_12285_),
    .c(_11705_),
    .o1(_12286_));
 b15nandp3ah1n03x5 _20965_ (.a(_12279_),
    .b(_12281_),
    .c(_12286_),
    .o1(_12287_));
 b15aoi112ah1n03x5 _20966_ (.a(net439),
    .b(_12071_),
    .c(_11586_),
    .d(_11749_),
    .o1(_12288_));
 b15aoi112aq1n08x5 _20967_ (.a(_11696_),
    .b(_12288_),
    .c(_11913_),
    .d(net453),
    .o1(_12289_));
 b15oai022ar1n02x5 _20968_ (.a(net453),
    .b(_11671_),
    .c(_11731_),
    .d(_11716_),
    .o1(_12290_));
 b15norp02an1n02x5 _20969_ (.a(net457),
    .b(_12290_),
    .o1(_12291_));
 b15nor003aq1n06x5 _20970_ (.a(_11666_),
    .b(_12289_),
    .c(_12291_),
    .o1(_12292_));
 b15nor004aq1n12x5 _20971_ (.a(_12267_),
    .b(_12276_),
    .c(_12287_),
    .d(_12292_),
    .o1(_12293_));
 b15aoi122aq1n02x5 _20972_ (.a(net453),
    .b(_11739_),
    .c(_11833_),
    .d(_11946_),
    .e(_11831_),
    .o1(_12294_));
 b15aoi012al1n02x5 _20973_ (.a(_11638_),
    .b(_11644_),
    .c(_11773_),
    .o1(_12295_));
 b15nor004ar1n02x5 _20974_ (.a(net459),
    .b(_11597_),
    .c(_11643_),
    .d(_11772_),
    .o1(_12296_));
 b15aoai13an1n08x5 _20975_ (.a(_11729_),
    .b(_11990_),
    .c(net451),
    .d(_11886_),
    .o1(_12297_));
 b15oai013ar1n02x5 _20976_ (.a(_12297_),
    .b(_11772_),
    .c(_11854_),
    .d(net446),
    .o1(_12298_));
 b15aoi013an1n02x5 _20977_ (.a(_12296_),
    .b(_12298_),
    .c(net436),
    .d(net459),
    .o1(_12299_));
 b15aoi013al1n03x5 _20978_ (.a(_12294_),
    .b(_12295_),
    .c(_12299_),
    .d(net453),
    .o1(_12300_));
 b15inv040as1n02x5 _20979_ (.a(_12300_),
    .o1(_12301_));
 b15nand04as1n16x5 _20980_ (.a(_12249_),
    .b(_12257_),
    .c(_12293_),
    .d(_12301_),
    .o1(_12302_));
 b15xor002as1n16x5 _20981_ (.a(_12239_),
    .b(_12302_),
    .out0(_12303_));
 b15xnr002ah1n16x5 _20982_ (.a(\u0.w[1][30] ),
    .b(_12303_),
    .out0(_12304_));
 b15xor003al1n02x5 _20983_ (.a(\u0.tmp_w[30] ),
    .b(\u0.w[2][30] ),
    .c(_12304_),
    .out0(_12305_));
 b15bfn001as1n64x5 max_length820 (.a(\us11.a[0] ),
    .o(net820));
 b15oai012ar1n02x5 _20985_ (.a(_12238_),
    .b(_12305_),
    .c(net938),
    .o1(_00376_));
 b15nand02ar1n02x5 _20986_ (.a(net943),
    .b(net53),
    .o1(_12307_));
 b15aoi012ar1n04x5 _20987_ (.a(_11849_),
    .b(_11691_),
    .c(_11826_),
    .o1(_12308_));
 b15nanb02an1n04x5 _20988_ (.a(_11805_),
    .b(_11665_),
    .out0(_12309_));
 b15oai013as1n04x5 _20989_ (.a(net454),
    .b(_11601_),
    .c(_11564_),
    .d(_11618_),
    .o1(_12310_));
 b15nona23ah1n12x5 _20990_ (.a(_12079_),
    .b(_12308_),
    .c(_12309_),
    .d(_12310_),
    .out0(_12311_));
 b15nanb02al1n04x5 _20991_ (.a(net458),
    .b(net459),
    .out0(_12312_));
 b15norp03ar1n02x5 _20992_ (.a(_11854_),
    .b(_12312_),
    .c(_11760_),
    .o1(_12313_));
 b15oai022as1n02x5 _20993_ (.a(_12002_),
    .b(_11916_),
    .c(_11772_),
    .d(_11741_),
    .o1(_12314_));
 b15aoai13an1n02x5 _20994_ (.a(net453),
    .b(_12313_),
    .c(_12314_),
    .d(_11827_),
    .o1(_12315_));
 b15oaoi13as1n08x5 _20995_ (.a(_12115_),
    .b(_11873_),
    .c(_11749_),
    .d(_11603_),
    .o1(_12316_));
 b15norp03an1n08x5 _20996_ (.a(_11565_),
    .b(_11614_),
    .c(_11637_),
    .o1(_12317_));
 b15norp02ah1n04x5 _20997_ (.a(_12316_),
    .b(_12317_),
    .o1(_12318_));
 b15nand02ar1n02x5 _20998_ (.a(_11696_),
    .b(_11666_),
    .o1(_12319_));
 b15oai112al1n06x5 _20999_ (.a(_12311_),
    .b(_12315_),
    .c(_12318_),
    .d(_12319_),
    .o1(_12320_));
 b15orn003ah1n02x5 _21000_ (.a(_11846_),
    .b(_11847_),
    .c(_12320_),
    .o(_12321_));
 b15aob012an1n02x5 _21001_ (.a(_11840_),
    .b(_11739_),
    .c(_11893_),
    .out0(_12322_));
 b15aoi122an1n04x5 _21002_ (.a(net453),
    .b(_11893_),
    .c(_11773_),
    .d(_12322_),
    .e(_11579_),
    .o1(_12323_));
 b15oai022an1n02x5 _21003_ (.a(_11696_),
    .b(_11565_),
    .c(_11655_),
    .d(net449),
    .o1(_12324_));
 b15nand03ar1n08x5 _21004_ (.a(net459),
    .b(_11704_),
    .c(_12324_),
    .o1(_12325_));
 b15nand02ar1n02x5 _21005_ (.a(_11696_),
    .b(_11624_),
    .o1(_12326_));
 b15aoai13ar1n02x5 _21006_ (.a(_11579_),
    .b(_11624_),
    .c(_12136_),
    .d(_11696_),
    .o1(_12327_));
 b15aoi012ar1n02x5 _21007_ (.a(_11666_),
    .b(_12326_),
    .c(_12327_),
    .o1(_12328_));
 b15nanb02an1n02x5 _21008_ (.a(_11879_),
    .b(_12051_),
    .out0(_12329_));
 b15oaoi13as1n08x5 _21009_ (.a(_12079_),
    .b(_12329_),
    .c(_12028_),
    .d(_12051_),
    .o1(_12330_));
 b15aoi012as1n02x5 _21010_ (.a(_12328_),
    .b(_12330_),
    .c(_11666_),
    .o1(_12331_));
 b15aoi013al1n06x5 _21011_ (.a(_12323_),
    .b(_12325_),
    .c(_12331_),
    .d(net452),
    .o1(_12332_));
 b15oaoi13al1n03x5 _21012_ (.a(_12093_),
    .b(\u0.tmp_w[18] ),
    .c(_11757_),
    .d(_11986_),
    .o1(_12333_));
 b15nor002as1n04x5 _21013_ (.a(_11805_),
    .b(_12333_),
    .o1(_12334_));
 b15aoai13ar1n03x5 _21014_ (.a(_11919_),
    .b(_11929_),
    .c(_12043_),
    .d(\u0.tmp_w[16] ),
    .o1(_12335_));
 b15norp03ar1n03x5 _21015_ (.a(_11999_),
    .b(_11667_),
    .c(_11760_),
    .o1(_12336_));
 b15aoai13as1n02x5 _21016_ (.a(_12336_),
    .b(_11603_),
    .c(_11965_),
    .d(_12201_),
    .o1(_12337_));
 b15norp02aq1n04x5 _21017_ (.a(_11693_),
    .b(_11597_),
    .o1(_12338_));
 b15nor003ah1n04x5 _21018_ (.a(net446),
    .b(_11575_),
    .c(_12312_),
    .o1(_12339_));
 b15oai112al1n16x5 _21019_ (.a(net442),
    .b(_11928_),
    .c(_12338_),
    .d(_12339_),
    .o1(_12340_));
 b15nand03aq1n08x5 _21020_ (.a(_12335_),
    .b(_12337_),
    .c(_12340_),
    .o1(_12341_));
 b15oaoi13ar1n02x5 _21021_ (.a(net451),
    .b(net454),
    .c(_12184_),
    .d(_11685_),
    .o1(_12342_));
 b15aoai13ar1n02x5 _21022_ (.a(_11685_),
    .b(_11965_),
    .c(_12038_),
    .d(_11671_),
    .o1(_12343_));
 b15aob012aq1n06x5 _21023_ (.a(_11664_),
    .b(_12342_),
    .c(_12343_),
    .out0(_12344_));
 b15norp03ah1n02x5 _21024_ (.a(_11760_),
    .b(_11954_),
    .c(_11787_),
    .o1(_12345_));
 b15oai022an1n02x5 _21025_ (.a(net451),
    .b(_11597_),
    .c(_11748_),
    .d(_11575_),
    .o1(_12346_));
 b15aoi013as1n04x5 _21026_ (.a(_12345_),
    .b(_12346_),
    .c(net440),
    .d(_11729_),
    .o1(_12347_));
 b15aoi022as1n04x5 _21027_ (.a(_11614_),
    .b(_11919_),
    .c(_11901_),
    .d(_11618_),
    .o1(_12348_));
 b15aoi022as1n06x5 _21028_ (.a(_11796_),
    .b(_11946_),
    .c(_12201_),
    .d(_11914_),
    .o1(_12349_));
 b15oai122al1n16x5 _21029_ (.a(_12347_),
    .b(_12348_),
    .c(net451),
    .d(_11603_),
    .e(_12349_),
    .o1(_12350_));
 b15nor004ah1n12x5 _21030_ (.a(_12334_),
    .b(_12341_),
    .c(_12344_),
    .d(_12350_),
    .o1(_12351_));
 b15oai013aq1n04x5 _21031_ (.a(_11685_),
    .b(_11643_),
    .c(net461),
    .d(_11597_),
    .o1(_12352_));
 b15oai022as1n02x5 _21032_ (.a(_11603_),
    .b(_11746_),
    .c(_11748_),
    .d(_11601_),
    .o1(_12353_));
 b15aoi022an1n12x5 _21033_ (.a(_11623_),
    .b(_12352_),
    .c(_12353_),
    .d(_11996_),
    .o1(_12354_));
 b15nandp2ar1n02x5 _21034_ (.a(_11574_),
    .b(_12136_),
    .o1(_12355_));
 b15nor002ar1n03x5 _21035_ (.a(_11666_),
    .b(_11791_),
    .o1(_12356_));
 b15oai013al1n03x5 _21036_ (.a(_11694_),
    .b(_12356_),
    .c(_12316_),
    .d(_12317_),
    .o1(_12357_));
 b15aoi013as1n03x5 _21037_ (.a(_11696_),
    .b(_12354_),
    .c(_12355_),
    .d(_12357_),
    .o1(_12358_));
 b15norp03al1n02x5 _21038_ (.a(net452),
    .b(_11556_),
    .c(_11597_),
    .o1(_12359_));
 b15norp03ar1n02x5 _21039_ (.a(net446),
    .b(_11575_),
    .c(_11646_),
    .o1(_12360_));
 b15oai012ar1n04x5 _21040_ (.a(_11689_),
    .b(_12359_),
    .c(_12360_),
    .o1(_12361_));
 b15nand03aq1n03x5 _21041_ (.a(net457),
    .b(net450),
    .c(_11901_),
    .o1(_12362_));
 b15oaoi13al1n02x5 _21042_ (.a(_11749_),
    .b(_11854_),
    .c(_11856_),
    .d(net453),
    .o1(_12363_));
 b15oab012ah1n02x5 _21043_ (.a(_12363_),
    .b(_11770_),
    .c(_11602_),
    .out0(_12364_));
 b15oai112ah1n08x5 _21044_ (.a(_12361_),
    .b(_12362_),
    .c(_12364_),
    .d(net450),
    .o1(_12365_));
 b15nandp2al1n02x5 _21045_ (.a(_11603_),
    .b(_12356_),
    .o1(_12366_));
 b15aoi012al1n04x5 _21046_ (.a(_11667_),
    .b(_12318_),
    .c(_12366_),
    .o1(_12367_));
 b15oaoi13ah1n08x5 _21047_ (.a(_12358_),
    .b(net459),
    .c(_12365_),
    .d(_12367_),
    .o1(_12368_));
 b15nona23ah1n16x5 _21048_ (.a(_12321_),
    .b(_12332_),
    .c(_12351_),
    .d(_12368_),
    .out0(_12369_));
 b15xnr002an1n16x5 _21049_ (.a(\u0.r0.out[31] ),
    .b(\u0.w[0][31] ),
    .out0(_12370_));
 b15xor002as1n16x5 _21050_ (.a(_12369_),
    .b(_12370_),
    .out0(_12371_));
 b15xor002ah1n12x5 _21051_ (.a(\u0.w[1][31] ),
    .b(_12371_),
    .out0(_12372_));
 b15xor002as1n16x5 _21052_ (.a(\u0.w[2][31] ),
    .b(_12372_),
    .out0(_12373_));
 b15xor002ar1n02x5 _21053_ (.a(net406),
    .b(_12373_),
    .out0(_12374_));
 b15oai012ar1n02x5 _21054_ (.a(_12307_),
    .b(_12374_),
    .c(net943),
    .o1(_00377_));
 b15nandp2aq1n03x5 _21055_ (.a(net129),
    .b(net54),
    .o1(_12375_));
 b15oai012al1n02x5 _21056_ (.a(_12375_),
    .b(_05078_),
    .c(net948),
    .o1(_00321_));
 b15nand02ar1n02x5 _21057_ (.a(net944),
    .b(net55),
    .o1(_12376_));
 b15oai012ar1n02x5 _21058_ (.a(_12376_),
    .b(_06590_),
    .c(net944),
    .o1(_00332_));
 b15nand02ar1n02x5 _21059_ (.a(net942),
    .b(net56),
    .o1(_12377_));
 b15oai012ar1n03x5 _21060_ (.a(_12377_),
    .b(_07621_),
    .c(net942),
    .o1(_00343_));
 b15bfn001as1n48x5 max_length819 (.a(\us11.a[0] ),
    .o(net819));
 b15nand02ar1n02x5 _21062_ (.a(net948),
    .b(net57),
    .o1(_12379_));
 b15oai012ar1n02x5 _21063_ (.a(_12379_),
    .b(_08739_),
    .c(net948),
    .o1(_00346_));
 b15nand02ar1n02x5 _21064_ (.a(net940),
    .b(net58),
    .o1(_12380_));
 b15oai012ar1n02x5 _21065_ (.a(_12380_),
    .b(_09443_),
    .c(net940),
    .o1(_00347_));
 b15nand02ar1n02x5 _21066_ (.a(net937),
    .b(net59),
    .o1(_12381_));
 b15oai012ar1n02x5 _21067_ (.a(_12381_),
    .b(_09694_),
    .c(net937),
    .o1(_00348_));
 b15nand02ar1n02x5 _21068_ (.a(net937),
    .b(net60),
    .o1(_12382_));
 b15oai012ar1n02x5 _21069_ (.a(_12382_),
    .b(_09775_),
    .c(net937),
    .o1(_00349_));
 b15nand02ar1n02x5 _21070_ (.a(net938),
    .b(net61),
    .o1(_12383_));
 b15oai012ar1n02x5 _21071_ (.a(_12383_),
    .b(_09848_),
    .c(net938),
    .o1(_00350_));
 b15nand02ar1n02x5 _21072_ (.a(net948),
    .b(net63),
    .o1(_12384_));
 b15bfn001ah1n64x5 max_length818 (.a(\us11.a[1] ),
    .o(net818));
 b15oai012ar1n02x5 _21074_ (.a(_12384_),
    .b(_10062_),
    .c(net948),
    .o1(_00351_));
 b15nandp2ar1n02x5 _21075_ (.a(net945),
    .b(net64),
    .o1(_12386_));
 b15oai012ar1n02x5 _21076_ (.a(_12386_),
    .b(_10192_),
    .c(net945),
    .o1(_00352_));
 b15nandp2al1n12x5 _21077_ (.a(net129),
    .b(net65),
    .o1(_12387_));
 b15oai012ar1n02x5 _21078_ (.a(_12387_),
    .b(_10298_),
    .c(net942),
    .o1(_00322_));
 b15nand02ar1n16x5 _21079_ (.a(net129),
    .b(net66),
    .o1(_12388_));
 b15xor002ar1n02x5 _21080_ (.a(\u0.w[2][11] ),
    .b(_10390_),
    .out0(_12389_));
 b15oai012ar1n02x5 _21081_ (.a(_12388_),
    .b(_12389_),
    .c(net942),
    .o1(_00323_));
 b15nand02an1n04x5 _21082_ (.a(net940),
    .b(net67),
    .o1(_12390_));
 b15oai012ar1n02x5 _21083_ (.a(_12390_),
    .b(_10474_),
    .c(net940),
    .o1(_00324_));
 b15bfn001as1n48x5 max_length817 (.a(\us11.a[1] ),
    .o(net817));
 b15nand02ar1n02x5 _21085_ (.a(net939),
    .b(net68),
    .o1(_12392_));
 b15oai012ar1n02x5 _21086_ (.a(_12392_),
    .b(_10549_),
    .c(net939),
    .o1(_00325_));
 b15nand02ar1n02x5 _21087_ (.a(net937),
    .b(net69),
    .o1(_12393_));
 b15oai012ar1n02x5 _21088_ (.a(_12393_),
    .b(_10632_),
    .c(net937),
    .o1(_00326_));
 b15nand02ar1n02x5 _21089_ (.a(net940),
    .b(net70),
    .o1(_12394_));
 b15oai012ar1n02x5 _21090_ (.a(_12394_),
    .b(_10705_),
    .c(net940),
    .o1(_00327_));
 b15nand02ar1n02x5 _21091_ (.a(net947),
    .b(net71),
    .o1(_12395_));
 b15oai012ar1n02x5 _21092_ (.a(_12395_),
    .b(_10937_),
    .c(net947),
    .o1(_00328_));
 b15nandp2ar1n05x5 _21093_ (.a(net129),
    .b(net72),
    .o1(_12396_));
 b15and002ar1n02x5 _21094_ (.a(\u0.w[2][17] ),
    .b(_11063_),
    .o(_12397_));
 b15norp02ar1n02x5 _21095_ (.a(\u0.w[2][17] ),
    .b(_11063_),
    .o1(_12398_));
 b15bfn001ah1n48x5 max_length816 (.a(net817),
    .o(net816));
 b15oai013ar1n02x5 _21097_ (.a(_12396_),
    .b(_12397_),
    .c(_12398_),
    .d(net946),
    .o1(_00329_));
 b15nandp2al1n04x5 _21098_ (.a(net129),
    .b(net74),
    .o1(_12400_));
 b15oai012al1n02x5 _21099_ (.a(_12400_),
    .b(_11151_),
    .c(net946),
    .o1(_00330_));
 b15nandp2ar1n08x5 _21100_ (.a(net948),
    .b(net75),
    .o1(_12401_));
 b15bfn001ah1n64x5 load_slew815 (.a(net816),
    .o(net815));
 b15oai012ar1n02x5 _21102_ (.a(_12401_),
    .b(_11242_),
    .c(net946),
    .o1(_00331_));
 b15nand02ar1n02x5 _21103_ (.a(net939),
    .b(net76),
    .o1(_12403_));
 b15oai012al1n02x5 _21104_ (.a(_12403_),
    .b(_11319_),
    .c(net939),
    .o1(_00333_));
 b15nand02ar1n02x5 _21105_ (.a(net939),
    .b(net77),
    .o1(_12404_));
 b15oai012ar1n02x5 _21106_ (.a(_12404_),
    .b(_11388_),
    .c(net939),
    .o1(_00334_));
 b15nand02ar1n02x5 _21107_ (.a(net939),
    .b(net78),
    .o1(_12405_));
 b15oai012ar1n02x5 _21108_ (.a(_12405_),
    .b(_11469_),
    .c(net939),
    .o1(_00335_));
 b15nand02ar1n02x5 _21109_ (.a(net940),
    .b(net79),
    .o1(_12406_));
 b15oai012ar1n02x5 _21110_ (.a(_12406_),
    .b(_11549_),
    .c(net940),
    .o1(_00336_));
 b15inv000ah1n05x5 _21111_ (.a(net80),
    .o1(_12407_));
 b15mdn022al1n03x5 _21112_ (.a(_12407_),
    .b(_11781_),
    .o1(_00337_),
    .sa(net945));
 b15bfn001ah1n64x5 wire814 (.a(\us11.a[2] ),
    .o(net814));
 b15nandp2as1n04x5 _21114_ (.a(net129),
    .b(net81),
    .o1(_12409_));
 b15xor002ar1n02x5 _21115_ (.a(\u0.w[2][25] ),
    .b(_11907_),
    .out0(_12410_));
 b15oai012ar1n02x5 _21116_ (.a(_12409_),
    .b(_12410_),
    .c(net945),
    .o1(_00338_));
 b15nanb03ar1n02x5 _21117_ (.a(net946),
    .b(\u0.w[2][26] ),
    .c(_12012_),
    .out0(_12411_));
 b15orn003ar1n02x5 _21118_ (.a(net946),
    .b(\u0.w[2][26] ),
    .c(_12012_),
    .o(_12412_));
 b15nandp2ar1n08x5 _21119_ (.a(net947),
    .b(net82),
    .o1(_12413_));
 b15nandp3ar1n02x5 _21120_ (.a(_12411_),
    .b(_12412_),
    .c(_12413_),
    .o1(_00339_));
 b15inv000ah1n08x5 _21121_ (.a(net83),
    .o1(_12414_));
 b15mdn022ar1n02x5 _21122_ (.a(_12414_),
    .b(_12101_),
    .o1(_00340_),
    .sa(net942));
 b15nand02al1n02x5 _21123_ (.a(net941),
    .b(net85),
    .o1(_12415_));
 b15oai012ar1n02x5 _21124_ (.a(_12415_),
    .b(_12180_),
    .c(net942),
    .o1(_00341_));
 b15nand02ar1n02x5 _21125_ (.a(net938),
    .b(net86),
    .o1(_12416_));
 b15oai012ar1n02x5 _21126_ (.a(_12416_),
    .b(_12236_),
    .c(net938),
    .o1(_00342_));
 b15inv040ah1n02x5 _21127_ (.a(net87),
    .o1(_12417_));
 b15xor002ar1n03x5 _21128_ (.a(\u0.w[2][30] ),
    .b(_12304_),
    .out0(_12418_));
 b15mdn022ar1n02x5 _21129_ (.a(_12417_),
    .b(_12418_),
    .o1(_00344_),
    .sa(net938));
 b15nand02ar1n02x5 _21130_ (.a(net938),
    .b(net88),
    .o1(_12419_));
 b15oai012ar1n02x5 _21131_ (.a(_12419_),
    .b(_12373_),
    .c(net938),
    .o1(_00345_));
 b15inv040as1n02x5 _21132_ (.a(net89),
    .o1(_12420_));
 b15mdn022al1n03x5 _21133_ (.a(_12420_),
    .b(_05067_),
    .o1(_00289_),
    .sa(net948));
 b15inv040ah1n05x5 _21134_ (.a(net90),
    .o1(_12421_));
 b15mdn022ar1n02x5 _21135_ (.a(_12421_),
    .b(_06579_),
    .o1(_00300_),
    .sa(net944));
 b15inv000as1n08x5 _21136_ (.a(net91),
    .o1(_12422_));
 b15mdn022ar1n02x5 _21137_ (.a(_12422_),
    .b(_07610_),
    .o1(_00311_),
    .sa(net942));
 b15inv040ah1n02x5 _21138_ (.a(net92),
    .o1(_12423_));
 b15mdn022al1n02x5 _21139_ (.a(_12423_),
    .b(_08728_),
    .o1(_00314_),
    .sa(net946));
 b15inv040al1n10x5 _21140_ (.a(net93),
    .o1(_12424_));
 b15mdn022an1n02x5 _21141_ (.a(_12424_),
    .b(_09442_),
    .o1(_00315_),
    .sa(net940));
 b15inv040aq1n06x5 _21142_ (.a(net94),
    .o1(_12425_));
 b15bfn001as1n64x5 max_length813 (.a(net814),
    .o(net813));
 b15mdn022ar1n02x5 _21144_ (.a(_12425_),
    .b(_09693_),
    .o1(_00316_),
    .sa(net939));
 b15inv040as1n05x5 _21145_ (.a(net96),
    .o1(_12427_));
 b15mdn022ar1n02x5 _21146_ (.a(_12427_),
    .b(_09774_),
    .o1(_00317_),
    .sa(net939));
 b15inv020ah1n12x5 _21147_ (.a(net97),
    .o1(_12428_));
 b15mdn022al1n03x5 _21148_ (.a(_12428_),
    .b(_09847_),
    .o1(_00318_),
    .sa(net940));
 b15inv040ah1n02x5 _21149_ (.a(net98),
    .o1(_12429_));
 b15mdn022ar1n02x5 _21150_ (.a(_12429_),
    .b(_10061_),
    .o1(_00319_),
    .sa(net948));
 b15inv040an1n06x5 _21151_ (.a(net99),
    .o1(_12430_));
 b15mdn022ar1n02x5 _21152_ (.a(_12430_),
    .b(_10191_),
    .o1(_00320_),
    .sa(net945));
 b15inv040ah1n05x5 _21153_ (.a(net100),
    .o1(_12431_));
 b15mdn022al1n03x5 _21154_ (.a(_12431_),
    .b(_10297_),
    .o1(_00290_),
    .sa(net945));
 b15nandp2al1n12x5 _21155_ (.a(net129),
    .b(net101),
    .o1(_12432_));
 b15oai012ar1n02x5 _21156_ (.a(_12432_),
    .b(_10390_),
    .c(net942),
    .o1(_00291_));
 b15inv000al1n16x5 _21157_ (.a(net102),
    .o1(_12433_));
 b15mdn022ar1n03x5 _21158_ (.a(_12433_),
    .b(_10473_),
    .o1(_00292_),
    .sa(net940));
 b15inv040an1n08x5 _21159_ (.a(net103),
    .o1(_12434_));
 b15mdn022ar1n03x5 _21160_ (.a(_12434_),
    .b(_10548_),
    .o1(_00293_),
    .sa(net939));
 b15inv000as1n08x5 _21161_ (.a(net104),
    .o1(_12435_));
 b15mdn022ar1n02x5 _21162_ (.a(_12435_),
    .b(_10631_),
    .o1(_00294_),
    .sa(net940));
 b15inv000as1n10x5 _21163_ (.a(net105),
    .o1(_12436_));
 b15mdn022ar1n03x5 _21164_ (.a(_12436_),
    .b(_10704_),
    .o1(_00295_),
    .sa(net940));
 b15inv040ah1n02x5 _21165_ (.a(net107),
    .o1(_12437_));
 b15bfn001ah1n64x5 load_slew812 (.a(net814),
    .o(net812));
 b15mdn022ar1n02x5 _21167_ (.a(_12437_),
    .b(_10936_),
    .o1(_00296_),
    .sa(net947));
 b15bfn001as1n64x5 max_length811 (.a(net813),
    .o(net811));
 b15bfn001ah1n64x5 max_length810 (.a(\us11.a[3] ),
    .o(net810));
 b15norp02ar1n02x5 _21170_ (.a(net946),
    .b(_11063_),
    .o1(_12441_));
 b15inv040ah1n02x5 _21171_ (.a(net108),
    .o1(_12442_));
 b15bfn001as1n48x5 load_slew809 (.a(\us11.a[3] ),
    .o(net809));
 b15aoi012ar1n02x5 _21173_ (.a(_12441_),
    .b(_12442_),
    .c(net946),
    .o1(_00297_));
 b15inv000as1n02x5 _21174_ (.a(net109),
    .o1(_12444_));
 b15mdn022ar1n02x5 _21175_ (.a(_12444_),
    .b(_11150_),
    .o1(_00298_),
    .sa(net946));
 b15inv040ah1n02x5 _21176_ (.a(net110),
    .o1(_12445_));
 b15mdn022ar1n02x5 _21177_ (.a(_12445_),
    .b(_11241_),
    .o1(_00299_),
    .sa(net945));
 b15inv020as1n24x5 _21178_ (.a(net111),
    .o1(_12446_));
 b15mdn022ar1n02x5 _21179_ (.a(_12446_),
    .b(_11318_),
    .o1(_00301_),
    .sa(net940));
 b15inv000al1n20x5 _21180_ (.a(net112),
    .o1(_12447_));
 b15mdn022ar1n02x5 _21181_ (.a(_12447_),
    .b(_11387_),
    .o1(_00302_),
    .sa(net936));
 b15inv000as1n02x5 _21182_ (.a(net113),
    .o1(_12448_));
 b15mdn022ar1n02x5 _21183_ (.a(_12448_),
    .b(_11468_),
    .o1(_00303_),
    .sa(net936));
 b15inv040ah1n05x5 _21184_ (.a(net114),
    .o1(_12449_));
 b15mdn022al1n02x5 _21185_ (.a(_12449_),
    .b(net391),
    .o1(_00304_),
    .sa(net945));
 b15nand02al1n12x5 _21186_ (.a(net129),
    .b(net115),
    .o1(_12450_));
 b15bfn001as1n48x5 load_slew808 (.a(net809),
    .o(net808));
 b15oai012ar1n03x5 _21188_ (.a(_12450_),
    .b(_11780_),
    .c(net945),
    .o1(_00305_));
 b15nand02ah1n06x5 _21189_ (.a(net129),
    .b(net116),
    .o1(_12452_));
 b15oai012ar1n02x5 _21190_ (.a(_12452_),
    .b(_11907_),
    .c(net945),
    .o1(_00306_));
 b15nand02an1n08x5 _21191_ (.a(net947),
    .b(net118),
    .o1(_12453_));
 b15oai012ar1n02x5 _21192_ (.a(_12453_),
    .b(_12012_),
    .c(net946),
    .o1(_00307_));
 b15nandp2ar1n16x5 _21193_ (.a(net129),
    .b(net119),
    .o1(_12454_));
 b15oai012ar1n02x5 _21194_ (.a(_12454_),
    .b(_12100_),
    .c(net942),
    .o1(_00308_));
 b15nandp2al1n16x5 _21195_ (.a(net129),
    .b(net120),
    .o1(_12455_));
 b15oai012ar1n02x5 _21196_ (.a(_12455_),
    .b(_12179_),
    .c(net942),
    .o1(_00309_));
 b15bfn001as1n32x5 wire807 (.a(\us11.a[4] ),
    .o(net807));
 b15nand02ar1n02x5 _21198_ (.a(net940),
    .b(net121),
    .o1(_12457_));
 b15oai012ar1n02x5 _21199_ (.a(_12457_),
    .b(_12235_),
    .c(net940),
    .o1(_00310_));
 b15nand02ar1n02x5 _21200_ (.a(net940),
    .b(net122),
    .o1(_12458_));
 b15oai012al1n02x5 _21201_ (.a(_12458_),
    .b(_12304_),
    .c(net940),
    .o1(_00312_));
 b15nand02ar1n02x5 _21202_ (.a(net938),
    .b(net123),
    .o1(_12459_));
 b15oai012an1n02x5 _21203_ (.a(_12459_),
    .b(_12372_),
    .c(net938),
    .o1(_00313_));
 b15nandp2ar1n05x5 _21204_ (.a(net129),
    .b(net124),
    .o1(_12460_));
 b15oai012ar1n02x5 _21205_ (.a(_12460_),
    .b(_05056_),
    .c(net948),
    .o1(_00257_));
 b15nand02ar1n02x5 _21206_ (.a(net944),
    .b(net125),
    .o1(_12461_));
 b15oai012ar1n02x5 _21207_ (.a(_12461_),
    .b(_06568_),
    .c(net944),
    .o1(_00268_));
 b15nandp2ar1n16x5 _21208_ (.a(net129),
    .b(net126),
    .o1(_12462_));
 b15bfn001ah1n64x5 load_slew806 (.a(net807),
    .o(net806));
 b15oai012ar1n02x5 _21210_ (.a(_12462_),
    .b(_07599_),
    .c(net942),
    .o1(_00279_));
 b15nand02ar1n02x5 _21211_ (.a(net948),
    .b(net127),
    .o1(_12464_));
 b15oai012ar1n02x5 _21212_ (.a(_12464_),
    .b(_08717_),
    .c(net948),
    .o1(_00282_));
 b15nand02aq1n16x5 _21213_ (.a(net129),
    .b(net2),
    .o1(_12465_));
 b15oai012ar1n02x5 _21214_ (.a(_12465_),
    .b(_09441_),
    .c(net941),
    .o1(_00283_));
 b15nand02aq1n16x5 _21215_ (.a(net129),
    .b(net3),
    .o1(_12466_));
 b15oai012ar1n02x5 _21216_ (.a(_12466_),
    .b(_09692_),
    .c(net941),
    .o1(_00284_));
 b15nand02ar1n02x5 _21217_ (.a(net939),
    .b(net4),
    .o1(_12467_));
 b15oai012ar1n02x5 _21218_ (.a(_12467_),
    .b(_09773_),
    .c(net939),
    .o1(_00285_));
 b15bfn001ah1n64x5 load_slew805 (.a(net807),
    .o(net805));
 b15nand02ar1n02x5 _21220_ (.a(net940),
    .b(net5),
    .o1(_12469_));
 b15oai012ar1n02x5 _21221_ (.a(_12469_),
    .b(_09846_),
    .c(net940),
    .o1(_00286_));
 b15nand02an1n04x5 _21222_ (.a(net129),
    .b(net6),
    .o1(_12470_));
 b15oai012ar1n02x5 _21223_ (.a(_12470_),
    .b(_10060_),
    .c(net946),
    .o1(_00287_));
 b15nand02al1n12x5 _21224_ (.a(net947),
    .b(net7),
    .o1(_12471_));
 b15oai012ar1n02x5 _21225_ (.a(_12471_),
    .b(_10190_),
    .c(net946),
    .o1(_00288_));
 b15nandp2ar1n12x5 _21226_ (.a(net129),
    .b(net8),
    .o1(_12472_));
 b15oai012ar1n02x5 _21227_ (.a(_12472_),
    .b(_10296_),
    .c(net945),
    .o1(_00258_));
 b15nand02as1n12x5 _21228_ (.a(net129),
    .b(net9),
    .o1(_12473_));
 b15oai012ar1n02x5 _21229_ (.a(_12473_),
    .b(_10389_),
    .c(net942),
    .o1(_00259_));
 b15nand02aq1n16x5 _21230_ (.a(net129),
    .b(net10),
    .o1(_12474_));
 b15bfn001ah1n64x5 max_length804 (.a(net805),
    .o(net804));
 b15oai012ar1n02x5 _21232_ (.a(_12474_),
    .b(_10472_),
    .c(net941),
    .o1(_00260_));
 b15nandp2al1n24x5 _21233_ (.a(net129),
    .b(net11),
    .o1(_12476_));
 b15oai012ar1n02x5 _21234_ (.a(_12476_),
    .b(_10547_),
    .c(net941),
    .o1(_00261_));
 b15nand02an1n16x5 _21235_ (.a(net129),
    .b(net13),
    .o1(_12477_));
 b15oai012ar1n02x5 _21236_ (.a(_12477_),
    .b(_10630_),
    .c(net941),
    .o1(_00262_));
 b15nandp2an1n16x5 _21237_ (.a(net129),
    .b(net14),
    .o1(_12478_));
 b15oai012ar1n02x5 _21238_ (.a(_12478_),
    .b(_10703_),
    .c(net941),
    .o1(_00263_));
 b15nandp2al1n04x5 _21239_ (.a(net947),
    .b(net15),
    .o1(_12479_));
 b15oai012ar1n02x5 _21240_ (.a(_12479_),
    .b(_10935_),
    .c(net946),
    .o1(_00264_));
 b15bfn001as1n64x5 max_length803 (.a(\us11.a[5] ),
    .o(net803));
 b15nandp2ar1n02x5 _21242_ (.a(net946),
    .b(net16),
    .o1(_12481_));
 b15oai012ar1n02x5 _21243_ (.a(_12481_),
    .b(_11062_),
    .c(net946),
    .o1(_00265_));
 b15nandp2ah1n03x5 _21244_ (.a(net947),
    .b(net17),
    .o1(_12482_));
 b15oai012ar1n02x5 _21245_ (.a(_12482_),
    .b(_11149_),
    .c(net946),
    .o1(_00266_));
 b15nandp2aq1n02x5 _21246_ (.a(net946),
    .b(net18),
    .o1(_12483_));
 b15oai012ar1n02x5 _21247_ (.a(_12483_),
    .b(_11240_),
    .c(net946),
    .o1(_00267_));
 b15nandp2as1n08x5 _21248_ (.a(net947),
    .b(net19),
    .o1(_12484_));
 b15oai012ar1n02x5 _21249_ (.a(_12484_),
    .b(_11317_),
    .c(net945),
    .o1(_00269_));
 b15qgbna2an1n10x5 _21250_ (.a(net947),
    .b(net20),
    .o1(_12485_));
 b15oai012ar1n02x5 _21251_ (.a(_12485_),
    .b(_11386_),
    .c(net945),
    .o1(_00270_));
 b15nand02ar1n16x5 _21252_ (.a(net129),
    .b(net21),
    .o1(_12486_));
 b15bfn001ah1n64x5 max_length802 (.a(net803),
    .o(net802));
 b15oai012ar1n02x5 _21254_ (.a(_12486_),
    .b(_11467_),
    .c(net945),
    .o1(_00271_));
 b15nandp2ar1n12x5 _21255_ (.a(net947),
    .b(net22),
    .o1(_12488_));
 b15oai012ar1n02x5 _21256_ (.a(_12488_),
    .b(_11547_),
    .c(net945),
    .o1(_00272_));
 b15norp02ar1n02x5 _21257_ (.a(net945),
    .b(_11779_),
    .o1(_12489_));
 b15inv000as1n02x5 _21258_ (.a(net24),
    .o1(_12490_));
 b15aoi012ar1n02x5 _21259_ (.a(_12489_),
    .b(_12490_),
    .c(net945),
    .o1(_00273_));
 b15norp02ar1n02x5 _21260_ (.a(net945),
    .b(_11906_),
    .o1(_12491_));
 b15inv040ah1n02x5 _21261_ (.a(net25),
    .o1(_12492_));
 b15aoi012ar1n02x5 _21262_ (.a(_12491_),
    .b(_12492_),
    .c(net945),
    .o1(_00274_));
 b15norp02aq1n04x5 _21263_ (.a(net946),
    .b(_12011_),
    .o1(_12493_));
 b15inv040ah1n02x5 _21264_ (.a(net26),
    .o1(_12494_));
 b15aoi012ar1n02x5 _21265_ (.a(_12493_),
    .b(_12494_),
    .c(net946),
    .o1(_00275_));
 b15nor002ah1n02x5 _21266_ (.a(net942),
    .b(_12099_),
    .o1(_12495_));
 b15inv000as1n06x5 _21267_ (.a(net27),
    .o1(_12496_));
 b15aoi012ar1n02x5 _21268_ (.a(_12495_),
    .b(_12496_),
    .c(net942),
    .o1(_00276_));
 b15norp02ar1n02x5 _21269_ (.a(net942),
    .b(_12178_),
    .o1(_12497_));
 b15inv040as1n04x5 _21270_ (.a(net28),
    .o1(_12498_));
 b15aoi012ar1n02x5 _21271_ (.a(_12497_),
    .b(_12498_),
    .c(net942),
    .o1(_00277_));
 b15norp02ar1n02x5 _21272_ (.a(net942),
    .b(_12234_),
    .o1(_12499_));
 b15inv000ah1n08x5 _21273_ (.a(net29),
    .o1(_12500_));
 b15aoi012ar1n02x5 _21274_ (.a(_12499_),
    .b(_12500_),
    .c(net942),
    .o1(_00278_));
 b15norp02ar1n02x5 _21275_ (.a(net942),
    .b(_12303_),
    .o1(_12501_));
 b15inv040ah1n05x5 _21276_ (.a(net30),
    .o1(_12502_));
 b15aoi012ar1n02x5 _21277_ (.a(_12501_),
    .b(_12502_),
    .c(net942),
    .o1(_00280_));
 b15inv020as1n08x5 _21278_ (.a(net31),
    .o1(_12503_));
 b15mdn022ar1n02x5 _21279_ (.a(_12503_),
    .b(_12371_),
    .o1(_00281_),
    .sa(net942));
 b15norp03al1n03x5 _21280_ (.a(\dcnt[1] ),
    .b(\dcnt[2] ),
    .c(\dcnt[3] ),
    .o1(_12504_));
 b15nano22ar1n02x5 _21281_ (.a(\dcnt[0] ),
    .b(_12504_),
    .c(net947),
    .out0(_00000_));
 b15inv000aq1n12x5 _21282_ (.a(\text_in_r[0] ),
    .o1(_12505_));
 b15bfn001as1n64x5 max_length801 (.a(\us11.a[6] ),
    .o(net801));
 b15bfn001as1n64x5 max_length800 (.a(\us11.a[6] ),
    .o(net800));
 b15bfn001as1n48x5 load_slew799 (.a(net800),
    .o(net799));
 b15bfn001ah1n64x5 load_slew798 (.a(\us11.a[7] ),
    .o(net798));
 b15bfn001as1n48x5 load_slew797 (.a(\us11.a[7] ),
    .o(net797));
 b15inv000an1n64x5 _21288_ (.a(net640),
    .o1(_12511_));
 b15bfn001ah1n64x5 max_length796 (.a(\us21.a[0] ),
    .o(net796));
 b15bfn001ah1n64x5 max_length795 (.a(\us21.a[0] ),
    .o(net795));
 b15bfn001as1n48x5 max_length794 (.a(net795),
    .o(net794));
 b15inv040ar1n48x5 _21292_ (.a(\us03.a[2] ),
    .o1(_12515_));
 b15bfn001ah1n80x5 wire793 (.a(\us21.a[1] ),
    .o(net793));
 b15bfn001as1n64x5 max_length792 (.a(net793),
    .o(net792));
 b15bfn001as1n48x5 max_length791 (.a(net792),
    .o(net791));
 b15nonb02aq1n16x5 _21296_ (.a(net625),
    .b(net622),
    .out0(_12519_));
 b15bfn001ah1n64x5 max_length790 (.a(net793),
    .o(net790));
 b15bfn001ah1n64x5 wire789 (.a(\us21.a[2] ),
    .o(net789));
 b15bfn001as1n64x5 load_slew788 (.a(net789),
    .o(net788));
 b15norp02as1n32x5 _21300_ (.a(net626),
    .b(net629),
    .o1(_12523_));
 b15nand02as1n24x5 _21301_ (.a(_12519_),
    .b(_12523_),
    .o1(_12524_));
 b15oai012as1n03x5 _21302_ (.a(_12511_),
    .b(_12515_),
    .c(_12524_),
    .o1(_12525_));
 b15bfn001as1n64x5 max_length787 (.a(net788),
    .o(net787));
 b15bfn001ah1n48x5 max_length786 (.a(net787),
    .o(net786));
 b15bfn001ah1n48x5 max_length785 (.a(net787),
    .o(net785));
 b15bfn001as1n48x5 wire784 (.a(\us21.a[3] ),
    .o(net784));
 b15bfn001ah1n64x5 max_length783 (.a(net784),
    .o(net783));
 b15oai012al1n06x5 _21308_ (.a(\us03.a[0] ),
    .b(net636),
    .c(_12524_),
    .o1(_12531_));
 b15bfn001as1n48x5 load_slew782 (.a(net784),
    .o(net782));
 b15bfn001as1n48x5 max_length781 (.a(net782),
    .o(net781));
 b15bfn001ah1n64x5 max_length780 (.a(net783),
    .o(net780));
 b15bfn001ah1n64x5 load_slew779 (.a(\us21.a[4] ),
    .o(net779));
 b15bfn001ah1n64x5 load_slew778 (.a(\us21.a[4] ),
    .o(net778));
 b15bfn001ah1n64x5 max_length777 (.a(net778),
    .o(net777));
 b15nonb03as1n12x5 _21315_ (.a(\us03.a[7] ),
    .b(net624),
    .c(\us03.a[4] ),
    .out0(_12538_));
 b15bfn001as1n64x5 max_length776 (.a(\us21.a[5] ),
    .o(net776));
 b15bfn001as1n64x5 max_length775 (.a(\us21.a[5] ),
    .o(net775));
 b15norp02ah1n04x5 _21318_ (.a(\us03.a[2] ),
    .b(\us03.a[5] ),
    .o1(_12541_));
 b15nandp2as1n12x5 _21319_ (.a(_12538_),
    .b(_12541_),
    .o1(_12542_));
 b15aoi012ar1n04x5 _21320_ (.a(\us03.a[1] ),
    .b(_12524_),
    .c(_12542_),
    .o1(_12543_));
 b15oai112ah1n12x5 _21321_ (.a(\us03.a[3] ),
    .b(_12525_),
    .c(_12531_),
    .d(_12543_),
    .o1(_12544_));
 b15inv040as1n40x5 _21322_ (.a(net632),
    .o1(_12545_));
 b15bfn001ah1n64x5 wire774 (.a(net775),
    .o(net774));
 b15nandp2an1n32x5 _21324_ (.a(net626),
    .b(net628),
    .o1(_12547_));
 b15bfn001as1n48x5 load_slew773 (.a(\us21.a[6] ),
    .o(net773));
 b15nanb02as1n24x5 _21326_ (.a(net624),
    .b(net621),
    .out0(_12549_));
 b15norp02ar1n48x5 _21327_ (.a(_12547_),
    .b(_12549_),
    .o1(_12550_));
 b15nonb02ah1n16x5 _21328_ (.a(\us03.a[2] ),
    .b(\us03.a[0] ),
    .out0(_12551_));
 b15nandp2ah1n48x5 _21329_ (.a(\us03.a[7] ),
    .b(net623),
    .o1(_12552_));
 b15nanb02as1n24x5 _21330_ (.a(net627),
    .b(net628),
    .out0(_12553_));
 b15nor002as1n32x5 _21331_ (.a(_12552_),
    .b(_12553_),
    .o1(_12554_));
 b15bfn001ah1n64x5 wire772 (.a(\us21.a[6] ),
    .o(net772));
 b15bfn001as1n64x5 max_length771 (.a(net773),
    .o(net771));
 b15bfn001ah1n64x5 load_slew770 (.a(\us21.a[7] ),
    .o(net770));
 b15bfn001as1n64x5 max_length769 (.a(net770),
    .o(net769));
 b15bfn001as1n48x5 load_slew768 (.a(\us21.a[7] ),
    .o(net768));
 b15aoi122an1n06x5 _21337_ (.a(_12545_),
    .b(_12550_),
    .c(_12551_),
    .d(_12554_),
    .e(\us03.a[0] ),
    .o1(_12560_));
 b15bfn001as1n48x5 load_slew767 (.a(\us31.a[0] ),
    .o(net767));
 b15bfn001as1n48x5 load_slew766 (.a(\us31.a[0] ),
    .o(net766));
 b15and002as1n16x5 _21340_ (.a(net626),
    .b(net629),
    .o(_12563_));
 b15nonb02as1n16x5 _21341_ (.a(net622),
    .b(net625),
    .out0(_12564_));
 b15nandp2an1n16x5 _21342_ (.a(_12563_),
    .b(_12564_),
    .o1(_12565_));
 b15nona23as1n32x5 _21343_ (.a(net629),
    .b(net625),
    .c(net622),
    .d(net626),
    .out0(_12566_));
 b15bfn001as1n64x5 max_length765 (.a(net766),
    .o(net765));
 b15oaoi13an1n02x5 _21345_ (.a(_12515_),
    .b(_12565_),
    .c(_12566_),
    .d(net640),
    .o1(_12568_));
 b15nanb02as1n24x5 _21346_ (.a(net621),
    .b(net623),
    .out0(_12569_));
 b15norp02an1n32x5 _21347_ (.a(_12569_),
    .b(_12547_),
    .o1(_12570_));
 b15aoi112as1n02x5 _21348_ (.a(net632),
    .b(_12568_),
    .c(_12570_),
    .d(_12515_),
    .o1(_12571_));
 b15bfn001as1n48x5 load_slew764 (.a(net766),
    .o(net764));
 b15bfn001as1n64x5 max_length763 (.a(\us31.a[1] ),
    .o(net763));
 b15bfn001as1n64x5 max_length762 (.a(\us31.a[1] ),
    .o(net762));
 b15bfn001ah1n64x5 max_length761 (.a(net762),
    .o(net761));
 b15oai013an1n08x5 _21353_ (.a(_12544_),
    .b(_12560_),
    .c(_12571_),
    .d(\us03.a[1] ),
    .o1(_12576_));
 b15nor002ar1n24x5 _21354_ (.a(_12545_),
    .b(_12566_),
    .o1(_12577_));
 b15bfn001as1n48x5 load_slew760 (.a(net762),
    .o(net760));
 b15and002aq1n04x5 _21356_ (.a(net640),
    .b(net633),
    .o(_12579_));
 b15orn002ah1n24x5 _21357_ (.a(net641),
    .b(net634),
    .o(_12580_));
 b15inv000aq1n56x5 _21358_ (.a(net637),
    .o1(_12581_));
 b15aoi012ah1n02x5 _21359_ (.a(_12579_),
    .b(_12580_),
    .c(_12581_),
    .o1(_12582_));
 b15bfn001ah1n64x5 wire759 (.a(\us31.a[2] ),
    .o(net759));
 b15nand02aq1n24x5 _21361_ (.a(net640),
    .b(net630),
    .o1(_12584_));
 b15bfn001as1n64x5 max_length758 (.a(net759),
    .o(net758));
 b15nonb02as1n16x5 _21363_ (.a(net626),
    .b(net629),
    .out0(_12586_));
 b15and002aq1n32x5 _21364_ (.a(net621),
    .b(net623),
    .o(_12587_));
 b15bfn001as1n48x5 wire757 (.a(\us31.a[2] ),
    .o(net757));
 b15nand03al1n12x5 _21366_ (.a(net636),
    .b(_12586_),
    .c(_12587_),
    .o1(_12589_));
 b15obai22ah1n06x5 _21367_ (.a(_12577_),
    .b(_12582_),
    .c(_12584_),
    .d(_12589_),
    .out0(_12590_));
 b15orn002ah1n32x5 _21368_ (.a(net630),
    .b(net636),
    .o(_12591_));
 b15bfn001as1n48x5 load_slew756 (.a(\us31.a[3] ),
    .o(net756));
 b15nor002ah1n24x5 _21370_ (.a(net622),
    .b(net625),
    .o1(_12593_));
 b15nandp2ar1n24x5 _21371_ (.a(_12586_),
    .b(_12593_),
    .o1(_12594_));
 b15and002aq1n16x5 _21372_ (.a(\us03.a[1] ),
    .b(net640),
    .o(_12595_));
 b15nor003an1n06x5 _21373_ (.a(_12591_),
    .b(_12594_),
    .c(_12595_),
    .o1(_12596_));
 b15nano23as1n24x5 _21374_ (.a(net629),
    .b(net625),
    .c(net622),
    .d(\us03.a[5] ),
    .out0(_12597_));
 b15nano22ah1n12x5 _21375_ (.a(net637),
    .b(net633),
    .c(net630),
    .out0(_12598_));
 b15and002ah1n04x5 _21376_ (.a(_12597_),
    .b(_12598_),
    .o(_12599_));
 b15nand02ar1n48x5 _21377_ (.a(_12564_),
    .b(_12523_),
    .o1(_12600_));
 b15nandp2ah1n32x5 _21378_ (.a(net630),
    .b(net633),
    .o1(_12601_));
 b15bfn001as1n64x5 max_length755 (.a(net756),
    .o(net755));
 b15norp02ar1n32x5 _21380_ (.a(\us03.a[1] ),
    .b(\us03.a[0] ),
    .o1(_12603_));
 b15norp03as1n04x5 _21381_ (.a(_12600_),
    .b(_12601_),
    .c(_12603_),
    .o1(_12604_));
 b15nor004as1n12x5 _21382_ (.a(_12590_),
    .b(_12596_),
    .c(_12599_),
    .d(_12604_),
    .o1(_12605_));
 b15nor002ar1n12x5 _21383_ (.a(net639),
    .b(\us03.a[5] ),
    .o1(_12606_));
 b15bfn001as1n64x5 max_length754 (.a(net755),
    .o(net754));
 b15bfn001as1n64x5 max_length753 (.a(\us31.a[4] ),
    .o(net753));
 b15bfn001as1n64x5 wire752 (.a(\us31.a[4] ),
    .o(net752));
 b15nonb03as1n12x5 _21387_ (.a(net624),
    .b(net621),
    .c(net628),
    .out0(_12610_));
 b15nano23ah1n24x5 _21388_ (.a(net627),
    .b(net624),
    .c(\us03.a[7] ),
    .d(\us03.a[4] ),
    .out0(_12611_));
 b15aoi022an1n06x5 _21389_ (.a(_12606_),
    .b(_12610_),
    .c(_12611_),
    .d(_12580_),
    .o1(_12612_));
 b15nona23as1n32x5 _21390_ (.a(net628),
    .b(net621),
    .c(net624),
    .d(net626),
    .out0(_12613_));
 b15aoi012ah1n02x5 _21391_ (.a(_12612_),
    .b(_12613_),
    .c(_12579_),
    .o1(_12614_));
 b15nanb02as1n24x5 _21392_ (.a(net640),
    .b(net637),
    .out0(_12615_));
 b15bfn001as1n48x5 load_slew751 (.a(\us31.a[5] ),
    .o(net751));
 b15nonb02al1n16x5 _21394_ (.a(net629),
    .b(net626),
    .out0(_12617_));
 b15oai112ar1n02x5 _21395_ (.a(net636),
    .b(_12593_),
    .c(_12617_),
    .d(_12586_),
    .o1(_12618_));
 b15nand02an1n24x5 _21396_ (.a(_12587_),
    .b(_12617_),
    .o1(_12619_));
 b15oaoi13ar1n02x5 _21397_ (.a(_12615_),
    .b(_12618_),
    .c(net636),
    .d(_12619_),
    .o1(_12620_));
 b15nor003aq1n02x5 _21398_ (.a(net632),
    .b(_12614_),
    .c(_12620_),
    .o1(_12621_));
 b15bfn001ah1n64x5 max_length750 (.a(net751),
    .o(net750));
 b15nandp2aq1n03x5 _21400_ (.a(_12586_),
    .b(_12587_),
    .o1(_12623_));
 b15oaoi13ar1n02x5 _21401_ (.a(net636),
    .b(_12619_),
    .c(_12623_),
    .d(net640),
    .o1(_12624_));
 b15oai022ar1n02x5 _21402_ (.a(net640),
    .b(_12619_),
    .c(_12623_),
    .d(net636),
    .o1(_12625_));
 b15aoi012as1n02x5 _21403_ (.a(_12624_),
    .b(_12625_),
    .c(\us03.a[1] ),
    .o1(_12626_));
 b15aoai13an1n06x5 _21404_ (.a(_12605_),
    .b(_12621_),
    .c(_12626_),
    .d(net632),
    .o1(_12627_));
 b15bfn001as1n64x5 wire749 (.a(\us31.a[5] ),
    .o(net749));
 b15nanb02ah1n24x5 _21406_ (.a(net631),
    .b(net639),
    .out0(_12629_));
 b15bfn001ah1n64x5 load_slew748 (.a(\us31.a[6] ),
    .o(net748));
 b15bfn001ah1n64x5 load_slew747 (.a(\us31.a[6] ),
    .o(net747));
 b15nor002an1n06x5 _21409_ (.a(\us03.a[4] ),
    .b(\us03.a[7] ),
    .o1(_12632_));
 b15bfn001ah1n64x5 load_slew746 (.a(net747),
    .o(net746));
 b15bfn001ah1n64x5 wire745 (.a(\us31.a[7] ),
    .o(net745));
 b15nonb02aq1n03x5 _21412_ (.a(\us03.a[2] ),
    .b(\us03.a[5] ),
    .out0(_12635_));
 b15nonb02ar1n16x5 _21413_ (.a(net627),
    .b(\us03.a[2] ),
    .out0(_12636_));
 b15and002al1n04x5 _21414_ (.a(\us03.a[4] ),
    .b(\us03.a[7] ),
    .o(_12637_));
 b15aoi022ah1n02x5 _21415_ (.a(_12632_),
    .b(_12635_),
    .c(_12636_),
    .d(_12637_),
    .o1(_12638_));
 b15norp03an1n08x5 _21416_ (.a(net624),
    .b(_12629_),
    .c(_12638_),
    .o1(_12639_));
 b15bfn001ah1n64x5 load_slew744 (.a(\us31.a[7] ),
    .o(net744));
 b15nonb02an1n16x5 _21418_ (.a(net627),
    .b(net631),
    .out0(_12641_));
 b15nand02an1n03x5 _21419_ (.a(\us03.a[4] ),
    .b(_12641_),
    .o1(_12642_));
 b15nor002al1n24x5 _21420_ (.a(net640),
    .b(net633),
    .o1(_12643_));
 b15aoi022ah1n06x5 _21421_ (.a(_12519_),
    .b(_12579_),
    .c(_12643_),
    .d(_12564_),
    .o1(_12644_));
 b15nano23an1n12x5 _21422_ (.a(net626),
    .b(net629),
    .c(net622),
    .d(net625),
    .out0(_12645_));
 b15nonb02as1n16x5 _21423_ (.a(net631),
    .b(net634),
    .out0(_12646_));
 b15bfn001ah1n64x5 max_length743 (.a(\us02.a[0] ),
    .o(net743));
 b15nandp2ah1n05x5 _21425_ (.a(_12645_),
    .b(_12646_),
    .o1(_12648_));
 b15orn002aq1n24x5 _21426_ (.a(net637),
    .b(net640),
    .o(_12649_));
 b15oai022as1n08x5 _21427_ (.a(_12642_),
    .b(_12644_),
    .c(_12648_),
    .d(_12649_),
    .o1(_12650_));
 b15nonb02an1n12x5 _21428_ (.a(net631),
    .b(net627),
    .out0(_12651_));
 b15aoi022ar1n04x5 _21429_ (.a(_12587_),
    .b(_12641_),
    .c(_12651_),
    .d(_12593_),
    .o1(_12652_));
 b15bfn001as1n48x5 max_length742 (.a(\us02.a[0] ),
    .o(net742));
 b15nanb02as1n16x5 _21431_ (.a(net642),
    .b(net631),
    .out0(_12654_));
 b15bfn001ah1n64x5 load_slew741 (.a(net743),
    .o(net741));
 b15oai112ah1n02x5 _21433_ (.a(_12581_),
    .b(_12654_),
    .c(_12591_),
    .d(_12511_),
    .o1(_12656_));
 b15nandp2aq1n32x5 _21434_ (.a(\us03.a[0] ),
    .b(\us03.a[2] ),
    .o1(_12657_));
 b15orn002ar1n12x5 _21435_ (.a(net640),
    .b(net630),
    .o(_12658_));
 b15nandp3al1n03x5 _21436_ (.a(net638),
    .b(_12657_),
    .c(_12658_),
    .o1(_12659_));
 b15aoi112ar1n04x5 _21437_ (.a(\us03.a[4] ),
    .b(_12652_),
    .c(_12656_),
    .d(_12659_),
    .o1(_12660_));
 b15nor003ar1n06x5 _21438_ (.a(_12639_),
    .b(_12650_),
    .c(_12660_),
    .o1(_12661_));
 b15inv000ar1n32x5 _21439_ (.a(net628),
    .o1(_12662_));
 b15bfn001ah1n64x5 wire740 (.a(\us02.a[0] ),
    .o(net740));
 b15nona23ar1n08x5 _21441_ (.a(net631),
    .b(net623),
    .c(net621),
    .d(net634),
    .out0(_12664_));
 b15norp02ar1n08x5 _21442_ (.a(_12662_),
    .b(_12664_),
    .o1(_12665_));
 b15nonb02ar1n12x5 _21443_ (.a(net628),
    .b(net623),
    .out0(_12666_));
 b15nand02ar1n02x5 _21444_ (.a(net635),
    .b(_12666_),
    .o1(_12667_));
 b15bfn001ah1n64x5 load_slew739 (.a(\us02.a[1] ),
    .o(net739));
 b15nanb02al1n12x5 _21446_ (.a(net628),
    .b(net623),
    .out0(_12669_));
 b15oai012as1n04x5 _21447_ (.a(_12667_),
    .b(_12669_),
    .c(net635),
    .o1(_12670_));
 b15inv020aq1n16x5 _21448_ (.a(\us03.a[7] ),
    .o1(_12671_));
 b15bfn001as1n48x5 load_slew738 (.a(net739),
    .o(net738));
 b15aoi013aq1n08x5 _21450_ (.a(_12665_),
    .b(_12670_),
    .c(_12671_),
    .d(net631),
    .o1(_12673_));
 b15bfn001ah1n48x5 max_length737 (.a(\us02.a[1] ),
    .o(net737));
 b15nand02as1n06x5 _21452_ (.a(net642),
    .b(\us03.a[5] ),
    .o1(_12675_));
 b15bfn001ah1n64x5 load_slew736 (.a(\us02.a[2] ),
    .o(net736));
 b15nona23as1n32x5 _21454_ (.a(net622),
    .b(net625),
    .c(net626),
    .d(net629),
    .out0(_12677_));
 b15bfn001as1n48x5 load_slew735 (.a(net736),
    .o(net735));
 b15oai022ar1n06x5 _21456_ (.a(_12511_),
    .b(_12600_),
    .c(_12615_),
    .d(_12677_),
    .o1(_12679_));
 b15aoi012al1n06x5 _21457_ (.a(net632),
    .b(net634),
    .c(_12679_),
    .o1(_12680_));
 b15bfn001ah1n64x5 max_length734 (.a(net736),
    .o(net734));
 b15bfn001as1n48x5 max_length733 (.a(net734),
    .o(net733));
 b15nandp2as1n24x5 _21460_ (.a(net638),
    .b(net634),
    .o1(_12683_));
 b15nandp2as1n24x5 _21461_ (.a(_12617_),
    .b(_12593_),
    .o1(_12684_));
 b15nandp2al1n08x5 _21462_ (.a(_12515_),
    .b(_12603_),
    .o1(_12685_));
 b15oai122aq1n16x5 _21463_ (.a(net632),
    .b(_12594_),
    .c(_12683_),
    .d(_12684_),
    .e(_12685_),
    .o1(_12686_));
 b15nonb02ah1n16x5 _21464_ (.a(net623),
    .b(net628),
    .out0(_12687_));
 b15nandp3ar1n08x5 _21465_ (.a(net627),
    .b(_12551_),
    .c(_12687_),
    .o1(_12688_));
 b15nanb02as1n24x5 _21466_ (.a(net633),
    .b(net641),
    .out0(_12689_));
 b15bfn001ah1n64x5 load_slew732 (.a(\us02.a[3] ),
    .o(net732));
 b15bfn001ah1n64x5 load_slew731 (.a(net732),
    .o(net731));
 b15nanb02al1n12x5 _21469_ (.a(net623),
    .b(net628),
    .out0(_12692_));
 b15oai013ah1n06x5 _21470_ (.a(_12688_),
    .b(_12689_),
    .c(net627),
    .d(_12692_),
    .o1(_12693_));
 b15bfn001as1n48x5 load_slew730 (.a(\us02.a[3] ),
    .o(net730));
 b15aoi013ah1n06x5 _21472_ (.a(_12686_),
    .b(_12693_),
    .c(_12671_),
    .d(net639),
    .o1(_12695_));
 b15oai122as1n16x5 _21473_ (.a(_12661_),
    .b(_12673_),
    .c(_12675_),
    .d(_12680_),
    .e(_12695_),
    .o1(_12696_));
 b15nano23as1n24x5 _21474_ (.a(net629),
    .b(net622),
    .c(net625),
    .d(\us03.a[5] ),
    .out0(_12697_));
 b15bfn001as1n48x5 wire729 (.a(net730),
    .o(net729));
 b15aoai13ar1n02x5 _21476_ (.a(_12581_),
    .b(_12597_),
    .c(_12697_),
    .d(net640),
    .o1(_12699_));
 b15nonb02as1n16x5 _21477_ (.a(net639),
    .b(net642),
    .out0(_12700_));
 b15aoi022ar1n02x5 _21478_ (.a(net640),
    .b(_12597_),
    .c(_12700_),
    .d(_12697_),
    .o1(_12701_));
 b15aoi012ah1n02x5 _21479_ (.a(_12591_),
    .b(_12699_),
    .c(_12701_),
    .o1(_12702_));
 b15bfn001as1n64x5 max_length728 (.a(\us02.a[4] ),
    .o(net728));
 b15nandp3al1n03x5 _21481_ (.a(_12545_),
    .b(_12519_),
    .c(_12563_),
    .o1(_12704_));
 b15nand03ar1n08x5 _21482_ (.a(net638),
    .b(_12538_),
    .c(_12651_),
    .o1(_12705_));
 b15aoi012ar1n02x5 _21483_ (.a(net633),
    .b(_12704_),
    .c(_12705_),
    .o1(_12706_));
 b15nonb02as1n16x5 _21484_ (.a(net633),
    .b(net630),
    .out0(_12707_));
 b15bfn001as1n64x5 max_length727 (.a(\us02.a[4] ),
    .o(net727));
 b15nandp2aq1n05x5 _21486_ (.a(_12581_),
    .b(_12707_),
    .o1(_12709_));
 b15xnr002an1n16x5 _21487_ (.a(net622),
    .b(net625),
    .out0(_12710_));
 b15nand02ar1n02x5 _21488_ (.a(_12617_),
    .b(_12710_),
    .o1(_12711_));
 b15aoi012an1n02x5 _21489_ (.a(_12709_),
    .b(_12711_),
    .c(_12594_),
    .o1(_12712_));
 b15oaoi13ar1n03x5 _21490_ (.a(_12702_),
    .b(net640),
    .c(_12706_),
    .d(_12712_),
    .o1(_12713_));
 b15nona23as1n32x5 _21491_ (.a(\us03.a[5] ),
    .b(\us03.a[7] ),
    .c(net625),
    .d(\us03.a[4] ),
    .out0(_12714_));
 b15bfn001ah1n64x5 load_slew726 (.a(net728),
    .o(net726));
 b15norp02ar1n02x5 _21493_ (.a(_12714_),
    .b(_12584_),
    .o1(_12716_));
 b15orn002aq1n32x5 _21494_ (.a(net621),
    .b(net623),
    .o(_12717_));
 b15norp02aq1n48x5 _21495_ (.a(_12553_),
    .b(_12717_),
    .o1(_12718_));
 b15bfn001as1n48x5 load_slew725 (.a(net728),
    .o(net725));
 b15norp02as1n16x5 _21497_ (.a(net630),
    .b(net636),
    .o1(_12720_));
 b15aoai13an1n02x5 _21498_ (.a(net637),
    .b(_12716_),
    .c(_12718_),
    .d(_12720_),
    .o1(_12721_));
 b15and002an1n12x5 _21499_ (.a(net631),
    .b(net627),
    .o(_12722_));
 b15nonb02an1n16x5 _21500_ (.a(net628),
    .b(net621),
    .out0(_12723_));
 b15and003al1n12x5 _21501_ (.a(net623),
    .b(_12722_),
    .c(_12723_),
    .o(_12724_));
 b15nanb03as1n16x5 _21502_ (.a(net638),
    .b(net641),
    .c(net634),
    .out0(_12725_));
 b15xor002ah1n12x5 _21503_ (.a(net641),
    .b(net633),
    .out0(_12726_));
 b15aob012aq1n04x5 _21504_ (.a(_12725_),
    .b(_12726_),
    .c(net638),
    .out0(_12727_));
 b15bfn001ah1n64x5 load_slew724 (.a(\us02.a[5] ),
    .o(net724));
 b15norp02aq1n03x5 _21506_ (.a(net638),
    .b(net628),
    .o1(_12729_));
 b15nanb03an1n02x5 _21507_ (.a(net634),
    .b(net627),
    .c(net631),
    .out0(_12730_));
 b15oai022aq1n06x5 _21508_ (.a(net627),
    .b(_12664_),
    .c(_12730_),
    .d(_12569_),
    .o1(_12731_));
 b15aoi022as1n12x5 _21509_ (.a(_12724_),
    .b(_12727_),
    .c(_12729_),
    .d(_12731_),
    .o1(_12732_));
 b15bfn001ah1n64x5 wire723 (.a(\us02.a[5] ),
    .o(net723));
 b15and003ar1n02x5 _21511_ (.a(net632),
    .b(net622),
    .c(net625),
    .o(_12734_));
 b15aoai13ar1n02x5 _21512_ (.a(_12734_),
    .b(_12563_),
    .c(_12523_),
    .d(_12580_),
    .o1(_12735_));
 b15and003ar1n12x5 _21513_ (.a(_12662_),
    .b(_12587_),
    .c(_12606_),
    .o(_12736_));
 b15bfn001ah1n64x5 wire722 (.a(net723),
    .o(net722));
 b15nandp2aq1n04x5 _21515_ (.a(net636),
    .b(_12615_),
    .o1(_12738_));
 b15oab012ah1n02x5 _21516_ (.a(_12735_),
    .b(_12736_),
    .c(_12738_),
    .out0(_12739_));
 b15norp03ar1n02x5 _21517_ (.a(net626),
    .b(net629),
    .c(net625),
    .o1(_12740_));
 b15aoi112ar1n02x5 _21518_ (.a(net632),
    .b(net636),
    .c(net622),
    .d(net640),
    .o1(_12741_));
 b15oai112ah1n02x5 _21519_ (.a(_12740_),
    .b(_12741_),
    .c(net637),
    .d(net622),
    .o1(_12742_));
 b15nona22as1n02x5 _21520_ (.a(net622),
    .b(net625),
    .c(net626),
    .out0(_12743_));
 b15nanb02ar1n02x5 _21521_ (.a(net629),
    .b(net640),
    .out0(_12744_));
 b15nandp2aq1n05x5 _21522_ (.a(net637),
    .b(net629),
    .o1(_12745_));
 b15nona23aq1n02x5 _21523_ (.a(_12601_),
    .b(_12743_),
    .c(_12744_),
    .d(_12745_),
    .out0(_12746_));
 b15nanb03as1n16x5 _21524_ (.a(net636),
    .b(net630),
    .c(net640),
    .out0(_12747_));
 b15oai112ah1n04x5 _21525_ (.a(_12742_),
    .b(_12746_),
    .c(_12714_),
    .d(_12747_),
    .o1(_12748_));
 b15nano23ah1n06x5 _21526_ (.a(_12721_),
    .b(_12732_),
    .c(_12739_),
    .d(_12748_),
    .out0(_12749_));
 b15nona23as1n32x5 _21527_ (.a(net626),
    .b(net625),
    .c(net622),
    .d(net629),
    .out0(_12750_));
 b15nand02ah1n24x5 _21528_ (.a(\us03.a[1] ),
    .b(\us03.a[3] ),
    .o1(_12751_));
 b15nor004as1n12x5 _21529_ (.a(\us03.a[5] ),
    .b(\us03.a[4] ),
    .c(\us03.a[7] ),
    .d(net624),
    .o1(_12752_));
 b15nandp2aq1n04x5 _21530_ (.a(net640),
    .b(_12752_),
    .o1(_12753_));
 b15orn002aq1n12x5 _21531_ (.a(net639),
    .b(net631),
    .o(_12754_));
 b15oai022ar1n04x5 _21532_ (.a(_12750_),
    .b(_12751_),
    .c(_12753_),
    .d(_12754_),
    .o1(_12755_));
 b15nandp2aq1n02x5 _21533_ (.a(net636),
    .b(_12755_),
    .o1(_12756_));
 b15bfn001ah1n64x5 load_slew721 (.a(\us02.a[6] ),
    .o(net721));
 b15bfn001ah1n64x5 load_slew720 (.a(net721),
    .o(net720));
 b15bfn001ah1n64x5 load_slew719 (.a(net721),
    .o(net719));
 b15nand04as1n16x5 _21537_ (.a(net626),
    .b(net629),
    .c(net622),
    .d(net625),
    .o1(_12760_));
 b15norp03ar1n02x5 _21538_ (.a(_12515_),
    .b(_12649_),
    .c(_12760_),
    .o1(_12761_));
 b15ornc04as1n24x5 _21539_ (.a(\us03.a[5] ),
    .b(net629),
    .c(\us03.a[7] ),
    .d(net625),
    .o(_12762_));
 b15nor002ah1n06x5 _21540_ (.a(_12649_),
    .b(_12762_),
    .o1(_12763_));
 b15and003ar1n02x5 _21541_ (.a(_12563_),
    .b(_12649_),
    .c(_12710_),
    .o(_12764_));
 b15oaoi13ar1n02x5 _21542_ (.a(_12761_),
    .b(_12515_),
    .c(_12763_),
    .d(_12764_),
    .o1(_12765_));
 b15nanb02as1n24x5 _21543_ (.a(net628),
    .b(net627),
    .out0(_12766_));
 b15bfn001as1n64x5 wire718 (.a(\us02.a[7] ),
    .o(net718));
 b15bfn001ah1n64x5 load_slew717 (.a(net718),
    .o(net717));
 b15nor003ar1n06x5 _21546_ (.a(_12766_),
    .b(_12584_),
    .c(_12717_),
    .o1(_12769_));
 b15nor003as1n03x5 _21547_ (.a(_12545_),
    .b(_12766_),
    .c(_12717_),
    .o1(_12770_));
 b15nona23as1n32x5 _21548_ (.a(net626),
    .b(net628),
    .c(net621),
    .d(net624),
    .out0(_12771_));
 b15nor002ar1n04x5 _21549_ (.a(_12658_),
    .b(_12771_),
    .o1(_12772_));
 b15oaoi13ar1n08x5 _21550_ (.a(_12769_),
    .b(net637),
    .c(_12770_),
    .d(_12772_),
    .o1(_12773_));
 b15oa0022ah1n03x5 _21551_ (.a(net632),
    .b(_12765_),
    .c(_12773_),
    .d(net636),
    .o(_12774_));
 b15nand04al1n08x5 _21552_ (.a(_12713_),
    .b(_12749_),
    .c(_12756_),
    .d(_12774_),
    .o1(_12775_));
 b15ornc04as1n24x5 _21553_ (.a(_12576_),
    .b(_12627_),
    .c(_12696_),
    .d(_12775_),
    .o(_12776_));
 b15bfn001ah1n64x5 load_slew716 (.a(\us02.a[7] ),
    .o(net716));
 b15bfn001as1n64x5 load_slew715 (.a(\us12.a[0] ),
    .o(net715));
 b15bfn001as1n64x5 max_length714 (.a(net715),
    .o(net714));
 b15bfn001ah1n48x5 wire713 (.a(net715),
    .o(net713));
 b15bfn001as1n48x5 load_slew712 (.a(\us12.a[1] ),
    .o(net712));
 b15inv000ar1n56x5 _21559_ (.a(net905),
    .o1(_12782_));
 b15bfn001ah1n64x5 wire711 (.a(\us12.a[1] ),
    .o(net711));
 b15bfn001ah1n64x5 max_length710 (.a(net712),
    .o(net710));
 b15bfn001ah1n64x5 max_length709 (.a(\us12.a[2] ),
    .o(net709));
 b15bfn001as1n48x5 load_slew708 (.a(\us12.a[2] ),
    .o(net708));
 b15bfn001ah1n48x5 load_slew707 (.a(net708),
    .o(net707));
 b15bfn001as1n64x5 max_length706 (.a(net709),
    .o(net706));
 b15nano23as1n24x5 _21566_ (.a(net895),
    .b(net891),
    .c(net888),
    .d(\us10.a[5] ),
    .out0(_12789_));
 b15nandp2al1n12x5 _21567_ (.a(net897),
    .b(_12789_),
    .o1(_12790_));
 b15nor002al1n03x5 _21568_ (.a(_12782_),
    .b(_12790_),
    .o1(_12791_));
 b15bfn001ah1n64x5 wire705 (.a(\us12.a[3] ),
    .o(net705));
 b15bfn001as1n64x5 max_length704 (.a(net705),
    .o(net704));
 b15bfn001as1n64x5 max_length703 (.a(net705),
    .o(net703));
 b15bfn001ah1n48x5 max_length702 (.a(net705),
    .o(net702));
 b15and002as1n32x5 _21573_ (.a(\us10.a[5] ),
    .b(net895),
    .o(_12796_));
 b15bfn001ah1n48x5 max_length701 (.a(net705),
    .o(net701));
 b15norp02as1n48x5 _21575_ (.a(net888),
    .b(net891),
    .o1(_12798_));
 b15bfn001as1n64x5 max_length700 (.a(\us12.a[4] ),
    .o(net700));
 b15nandp2as1n24x5 _21577_ (.a(_12796_),
    .b(_12798_),
    .o1(_12800_));
 b15bfn001ah1n64x5 wire699 (.a(\us12.a[4] ),
    .o(net699));
 b15bfn001ah1n64x5 wire698 (.a(\us12.a[5] ),
    .o(net698));
 b15oaoi13an1n03x5 _21580_ (.a(net902),
    .b(_12790_),
    .c(_12800_),
    .d(net897),
    .o1(_12803_));
 b15bfn001as1n64x5 max_length697 (.a(net698),
    .o(net697));
 b15bfn001ah1n64x5 wire696 (.a(net698),
    .o(net696));
 b15bfn001as1n64x5 max_length695 (.a(\us12.a[6] ),
    .o(net695));
 b15bfn001ah1n64x5 wire694 (.a(\us12.a[6] ),
    .o(net694));
 b15bfn001ah1n64x5 load_slew693 (.a(\us12.a[7] ),
    .o(net693));
 b15bfn001ah1n64x5 load_slew692 (.a(net693),
    .o(net692));
 b15bfn001as1n64x5 max_length691 (.a(net693),
    .o(net691));
 b15and002al1n16x5 _21588_ (.a(net892),
    .b(net887),
    .o(_12811_));
 b15bfn001ah1n64x5 max_length690 (.a(\us22.a[0] ),
    .o(net690));
 b15bfn001as1n48x5 wire689 (.a(net690),
    .o(net689));
 b15bfn001ah1n64x5 load_slew688 (.a(\us22.a[0] ),
    .o(net688));
 b15bfn001ah1n64x5 load_slew687 (.a(\us22.a[1] ),
    .o(net687));
 b15bfn001ah1n64x5 load_slew686 (.a(net687),
    .o(net686));
 b15bfn001ah1n64x5 load_slew685 (.a(\us22.a[1] ),
    .o(net685));
 b15aoi012al1n04x5 _21595_ (.a(net899),
    .b(net902),
    .c(net908),
    .o1(_12818_));
 b15nand03as1n08x5 _21596_ (.a(net890),
    .b(_12811_),
    .c(_12818_),
    .o1(_12819_));
 b15inv040ah1n40x5 _21597_ (.a(net902),
    .o1(_12820_));
 b15bfn001ah1n48x5 load_slew684 (.a(net685),
    .o(net684));
 b15nonb02as1n16x5 _21599_ (.a(\us10.a[5] ),
    .b(net895),
    .out0(_12822_));
 b15bfn001as1n48x5 max_length683 (.a(\us22.a[2] ),
    .o(net683));
 b15bfn001ah1n64x5 load_slew682 (.a(net683),
    .o(net682));
 b15andc04as1n16x5 _21602_ (.a(net893),
    .b(net896),
    .c(net886),
    .d(\us10.a[6] ),
    .o(_12825_));
 b15bfn001as1n64x5 load_slew681 (.a(net682),
    .o(net681));
 b15orn002ar1n32x5 _21604_ (.a(net905),
    .b(net902),
    .o(_12827_));
 b15oai022ar1n02x5 _21605_ (.a(_12820_),
    .b(_12822_),
    .c(_12825_),
    .d(_12827_),
    .o1(_12828_));
 b15nor002an1n02x5 _21606_ (.a(_12819_),
    .b(_12828_),
    .o1(_12829_));
 b15oai013ah1n06x5 _21607_ (.a(net910),
    .b(_12791_),
    .c(_12803_),
    .d(_12829_),
    .o1(_12830_));
 b15bfn001as1n48x5 wire680 (.a(net683),
    .o(net680));
 b15inv000as1n24x5 _21609_ (.a(net895),
    .o1(_12832_));
 b15bfn001as1n64x5 max_length679 (.a(\us22.a[3] ),
    .o(net679));
 b15bfn001as1n48x5 load_slew678 (.a(net679),
    .o(net678));
 b15bfn001as1n64x5 max_length677 (.a(net678),
    .o(net677));
 b15bfn001as1n64x5 max_length676 (.a(\us22.a[4] ),
    .o(net676));
 b15nandp2ar1n02x5 _21614_ (.a(_12832_),
    .b(net908),
    .o1(_12837_));
 b15oai012al1n06x5 _21615_ (.a(_12837_),
    .b(_12827_),
    .c(_12832_),
    .o1(_12838_));
 b15oai013an1n12x5 _21616_ (.a(_12830_),
    .b(_12838_),
    .c(_12819_),
    .d(net910),
    .o1(_12839_));
 b15bfn001as1n48x5 max_length675 (.a(\us22.a[4] ),
    .o(net675));
 b15bfn001as1n64x5 max_length674 (.a(\us22.a[5] ),
    .o(net674));
 b15bfn001ah1n64x5 max_length673 (.a(\us22.a[5] ),
    .o(net673));
 b15bfn001ah1n64x5 load_slew672 (.a(\us22.a[6] ),
    .o(net672));
 b15nandp3al1n04x5 _21621_ (.a(net908),
    .b(net902),
    .c(net899),
    .o1(_12844_));
 b15bfn001as1n48x5 load_slew671 (.a(\us22.a[6] ),
    .o(net671));
 b15bfn001as1n64x5 max_length670 (.a(\us22.a[7] ),
    .o(net670));
 b15bfn001ah1n64x5 load_slew669 (.a(net670),
    .o(net669));
 b15nonb02as1n16x5 _21625_ (.a(net891),
    .b(net888),
    .out0(_12848_));
 b15bfn001as1n64x5 wire668 (.a(\us32.a[0] ),
    .o(net668));
 b15aoai13as1n04x5 _21627_ (.a(_12844_),
    .b(net899),
    .c(_12796_),
    .d(_12848_),
    .o1(_12850_));
 b15inv000as1n80x5 _21628_ (.a(net897),
    .o1(_12851_));
 b15bfn001as1n48x5 max_length667 (.a(net668),
    .o(net667));
 b15oai112an1n04x5 _21630_ (.a(_12796_),
    .b(_12848_),
    .c(_12827_),
    .d(_12851_),
    .o1(_12853_));
 b15bfn001as1n48x5 max_length666 (.a(net668),
    .o(net666));
 b15bfn001ah1n64x5 max_length665 (.a(\us32.a[1] ),
    .o(net665));
 b15bfn001ah1n64x5 load_slew664 (.a(\us32.a[1] ),
    .o(net664));
 b15nona23as1n32x5 _21634_ (.a(net893),
    .b(net896),
    .c(net886),
    .d(net889),
    .out0(_12857_));
 b15aoi022as1n06x5 _21635_ (.a(net910),
    .b(_12850_),
    .c(_12853_),
    .d(_12857_),
    .o1(_12858_));
 b15bfn001ah1n64x5 max_length663 (.a(net664),
    .o(net663));
 b15bfn001ah1n64x5 wire662 (.a(\us32.a[2] ),
    .o(net662));
 b15bfn001as1n64x5 max_length661 (.a(net662),
    .o(net661));
 b15aoai13ar1n04x5 _21639_ (.a(_12820_),
    .b(net899),
    .c(_12857_),
    .d(net906),
    .o1(_12862_));
 b15nonb02as1n16x5 _21640_ (.a(net904),
    .b(net900),
    .out0(_12863_));
 b15inv020ar1n40x5 _21641_ (.a(net891),
    .o1(_12864_));
 b15nandp2ah1n12x5 _21642_ (.a(net892),
    .b(net894),
    .o1(_12865_));
 b15bfn001ah1n64x5 max_length660 (.a(net661),
    .o(net660));
 b15orn002aq1n04x5 _21644_ (.a(net886),
    .b(net903),
    .o(_12867_));
 b15bfn001as1n64x5 max_length659 (.a(net661),
    .o(net659));
 b15nand02ah1n06x5 _21646_ (.a(net887),
    .b(net904),
    .o1(_12869_));
 b15orn002ah1n16x5 _21647_ (.a(net893),
    .b(net896),
    .o(_12870_));
 b15oa0022ar1n06x5 _21648_ (.a(_12865_),
    .b(_12867_),
    .c(_12869_),
    .d(_12870_),
    .o(_12871_));
 b15oaoi13an1n03x5 _21649_ (.a(_12863_),
    .b(_12782_),
    .c(_12864_),
    .d(_12871_),
    .o1(_12872_));
 b15aoai13ar1n06x5 _21650_ (.a(_12858_),
    .b(net910),
    .c(_12862_),
    .d(_12872_),
    .o1(_12873_));
 b15nonb02as1n16x5 _21651_ (.a(net888),
    .b(net891),
    .out0(_12874_));
 b15nandp2ah1n24x5 _21652_ (.a(_12796_),
    .b(_12874_),
    .o1(_12875_));
 b15bfn001ah1n64x5 wire658 (.a(\us32.a[3] ),
    .o(net658));
 b15nonb02as1n16x5 _21654_ (.a(net908),
    .b(net913),
    .out0(_12877_));
 b15bfn001as1n48x5 wire657 (.a(net658),
    .o(net657));
 b15nanb02as1n24x5 _21656_ (.a(net909),
    .b(net913),
    .out0(_12879_));
 b15bfn001as1n64x5 max_length656 (.a(net658),
    .o(net656));
 b15and002aq1n32x5 _21658_ (.a(net887),
    .b(net891),
    .o(_12881_));
 b15bfn001ah1n64x5 load_slew655 (.a(net656),
    .o(net655));
 b15nonb02as1n16x5 _21660_ (.a(net896),
    .b(net893),
    .out0(_12883_));
 b15bfn001ah1n64x5 load_slew654 (.a(\us32.a[4] ),
    .o(net654));
 b15nandp2ar1n12x5 _21662_ (.a(_12881_),
    .b(_12883_),
    .o1(_12885_));
 b15oai022ah1n04x5 _21663_ (.a(_12875_),
    .b(_12877_),
    .c(_12879_),
    .d(_12885_),
    .o1(_12886_));
 b15bfn001ah1n64x5 load_slew653 (.a(\us32.a[4] ),
    .o(net653));
 b15bfn001as1n64x5 load_slew652 (.a(net653),
    .o(net652));
 b15bfn001as1n64x5 max_length651 (.a(\us32.a[5] ),
    .o(net651));
 b15bfn001as1n64x5 max_length650 (.a(\us32.a[5] ),
    .o(net650));
 b15bfn001ah1n64x5 wire649 (.a(net650),
    .o(net649));
 b15nano22al1n03x5 _21669_ (.a(net895),
    .b(net909),
    .c(\us10.a[5] ),
    .out0(_12892_));
 b15nano22ah1n03x5 _21670_ (.a(\us10.a[5] ),
    .b(net913),
    .c(net895),
    .out0(_12893_));
 b15oai112al1n12x5 _21671_ (.a(net904),
    .b(_12874_),
    .c(_12892_),
    .d(_12893_),
    .o1(_12894_));
 b15bfn001ah1n64x5 wire648 (.a(\us32.a[6] ),
    .o(net648));
 b15oai012as1n04x5 _21673_ (.a(_12894_),
    .b(_12885_),
    .c(net904),
    .o1(_12896_));
 b15bfn001as1n64x5 max_length647 (.a(net648),
    .o(net647));
 b15bfn001as1n64x5 max_length646 (.a(net647),
    .o(net646));
 b15aoi022ar1n12x5 _21676_ (.a(_12863_),
    .b(_12886_),
    .c(_12896_),
    .d(net900),
    .o1(_12899_));
 b15nand02aq1n08x5 _21677_ (.a(net912),
    .b(net899),
    .o1(_12900_));
 b15aoi012ar1n02x5 _21678_ (.a(_12820_),
    .b(_12900_),
    .c(net906),
    .o1(_12901_));
 b15nandp2aq1n03x5 _21679_ (.a(net899),
    .b(_12825_),
    .o1(_12902_));
 b15bfn001as1n64x5 max_length645 (.a(\us32.a[7] ),
    .o(net645));
 b15nanb02as1n24x5 _21681_ (.a(net910),
    .b(net905),
    .out0(_12904_));
 b15bfn001as1n64x5 max_length644 (.a(\us32.a[7] ),
    .o(net644));
 b15oai112an1n04x5 _21683_ (.a(_12851_),
    .b(_12789_),
    .c(_12904_),
    .d(net903),
    .o1(_12906_));
 b15aoi012aq1n04x5 _21684_ (.a(_12901_),
    .b(_12902_),
    .c(_12906_),
    .o1(_12907_));
 b15nor002ar1n24x5 _21685_ (.a(net904),
    .b(net900),
    .o1(_12908_));
 b15nor004as1n12x5 _21686_ (.a(net893),
    .b(net896),
    .c(net886),
    .d(net889),
    .o1(_12909_));
 b15nor002ah1n32x5 _21687_ (.a(net913),
    .b(net908),
    .o1(_12910_));
 b15nandp3ar1n12x5 _21688_ (.o1(_12911_),
    .a(_12908_),
    .b(_12909_),
    .c(_12910_));
 b15nonb02as1n16x5 _21689_ (.a(net904),
    .b(net913),
    .out0(_12912_));
 b15nandp2al1n32x5 _21690_ (.a(net908),
    .b(net902),
    .o1(_12913_));
 b15bfn001ah1n64x5 wire643 (.a(net644),
    .o(net643));
 b15aoi012al1n06x5 _21692_ (.a(_12912_),
    .b(_12913_),
    .c(net910),
    .o1(_12915_));
 b15norp02as1n48x5 _21693_ (.a(\us10.a[5] ),
    .b(net895),
    .o1(_12916_));
 b15nandp2ar1n48x5 _21694_ (.a(_12916_),
    .b(_12848_),
    .o1(_12917_));
 b15bfn001as1n48x5 max_length642 (.a(\us03.a[0] ),
    .o(net642));
 b15oai013as1n12x5 _21696_ (.a(_12911_),
    .b(_12915_),
    .c(_12917_),
    .d(_12851_),
    .o1(_12919_));
 b15bfn001as1n64x5 max_length641 (.a(net642),
    .o(net641));
 b15bfn001ah1n64x5 wire640 (.a(\us03.a[0] ),
    .o(net640));
 b15nonb02as1n16x5 _21699_ (.a(net913),
    .b(net908),
    .out0(_12922_));
 b15bfn001ah1n64x5 max_length639 (.a(\us03.a[1] ),
    .o(net639));
 b15nandp3ah1n16x5 _21701_ (.a(net901),
    .b(_12822_),
    .c(_12798_),
    .o1(_12924_));
 b15bfn001as1n48x5 max_length638 (.a(\us03.a[1] ),
    .o(net638));
 b15bfn001ah1n64x5 load_slew637 (.a(net638),
    .o(net637));
 b15nand04aq1n04x5 _21704_ (.a(_12820_),
    .b(_12883_),
    .c(_12904_),
    .d(_12798_),
    .o1(_12927_));
 b15aoi112ah1n04x5 _21705_ (.a(_12851_),
    .b(_12922_),
    .c(_12924_),
    .d(_12927_),
    .o1(_12928_));
 b15nanb03ar1n16x5 _21706_ (.a(net892),
    .b(net895),
    .c(net888),
    .out0(_12929_));
 b15bfn001ah1n64x5 max_length636 (.a(\us03.a[2] ),
    .o(net636));
 b15nand02as1n12x5 _21708_ (.a(net889),
    .b(net898),
    .o1(_12931_));
 b15orn002ar1n32x5 _21709_ (.a(net903),
    .b(net899),
    .o(_12932_));
 b15bfn001ah1n64x5 max_length635 (.a(net636),
    .o(net635));
 b15oaoi13as1n08x5 _21711_ (.a(_12929_),
    .b(_12931_),
    .c(_12932_),
    .d(net889),
    .o1(_12934_));
 b15and002ar1n03x5 _21712_ (.a(_12922_),
    .b(_12934_),
    .o(_12935_));
 b15nor004ah1n08x5 _21713_ (.a(_12907_),
    .b(_12919_),
    .c(_12928_),
    .d(_12935_),
    .o1(_12936_));
 b15bfn001as1n48x5 load_slew634 (.a(net635),
    .o(net634));
 b15nanb02al1n12x5 _21715_ (.a(net891),
    .b(net913),
    .out0(_12938_));
 b15oai012ar1n02x5 _21716_ (.a(\us10.a[5] ),
    .b(net908),
    .c(net904),
    .o1(_12939_));
 b15nonb02as1n16x5 _21717_ (.a(net888),
    .b(net895),
    .out0(_12940_));
 b15bfn001ah1n64x5 max_length633 (.a(net636),
    .o(net633));
 b15nona23ar1n04x5 _21719_ (.a(_12851_),
    .b(_12938_),
    .c(_12939_),
    .d(_12940_),
    .out0(_12942_));
 b15bfn001ah1n64x5 max_length632 (.a(\us03.a[3] ),
    .o(net632));
 b15bfn001as1n48x5 max_length631 (.a(\us03.a[3] ),
    .o(net631));
 b15nonb03ar1n03x5 _21722_ (.a(net900),
    .b(net904),
    .c(net888),
    .out0(_12945_));
 b15xor002ar1n04x5 _21723_ (.a(net891),
    .b(net909),
    .out0(_12946_));
 b15bfn001ah1n64x5 load_slew630 (.a(net632),
    .o(net630));
 b15oai112ah1n06x5 _21725_ (.a(_12822_),
    .b(_12945_),
    .c(_12946_),
    .d(net913),
    .o1(_12948_));
 b15nand02ah1n16x5 _21726_ (.a(_12864_),
    .b(_12796_),
    .o1(_12949_));
 b15inv000as1n64x5 _21727_ (.a(net910),
    .o1(_12950_));
 b15bfn001as1n64x5 max_length629 (.a(\us03.a[4] ),
    .o(net629));
 b15aoai13as1n02x5 _21729_ (.a(_12908_),
    .b(net908),
    .c(_12950_),
    .d(net887),
    .o1(_12952_));
 b15oai112as1n08x5 _21730_ (.a(_12942_),
    .b(_12948_),
    .c(_12949_),
    .d(_12952_),
    .o1(_12953_));
 b15nanb02aq1n24x5 _21731_ (.a(net907),
    .b(net898),
    .out0(_12954_));
 b15bfn001as1n48x5 load_slew628 (.a(\us03.a[4] ),
    .o(net628));
 b15nanb02aq1n12x5 _21733_ (.a(net889),
    .b(net886),
    .out0(_12956_));
 b15nor002aq1n16x5 _21734_ (.a(_12870_),
    .b(_12956_),
    .o1(_12957_));
 b15oai112ar1n02x5 _21735_ (.a(net902),
    .b(_12954_),
    .c(_12900_),
    .d(_12957_),
    .o1(_12958_));
 b15nano23as1n24x5 _21736_ (.a(net893),
    .b(net889),
    .c(net886),
    .d(net896),
    .out0(_12959_));
 b15nanb02ah1n24x5 _21737_ (.a(net898),
    .b(net907),
    .out0(_12960_));
 b15aoi012ar1n02x5 _21738_ (.a(_12959_),
    .b(_12957_),
    .c(_12960_),
    .o1(_12961_));
 b15oab012aq1n03x5 _21739_ (.a(_12953_),
    .b(_12958_),
    .c(_12961_),
    .out0(_12962_));
 b15nand04as1n12x5 _21740_ (.a(_12873_),
    .b(_12899_),
    .c(_12936_),
    .d(_12962_),
    .o1(_12963_));
 b15and002ar1n08x5 _21741_ (.a(net901),
    .b(net898),
    .o(_12964_));
 b15bfn001as1n48x5 load_slew627 (.a(\us03.a[5] ),
    .o(net627));
 b15nandp3ar1n02x5 _21743_ (.a(net911),
    .b(_12964_),
    .c(_12909_),
    .o1(_12966_));
 b15oai112al1n02x5 _21744_ (.a(_12782_),
    .b(_12966_),
    .c(_12917_),
    .d(_12932_),
    .o1(_12967_));
 b15nonb02as1n16x5 _21745_ (.a(net897),
    .b(net901),
    .out0(_12968_));
 b15bfn001ah1n64x5 load_slew626 (.a(\us03.a[5] ),
    .o(net626));
 b15nand02ar1n02x5 _21747_ (.a(_12968_),
    .b(_12909_),
    .o1(_12970_));
 b15and002al1n32x5 _21748_ (.a(net912),
    .b(net903),
    .o(_12971_));
 b15bfn001as1n64x5 wire625 (.a(\us03.a[6] ),
    .o(net625));
 b15nandp2ah1n12x5 _21750_ (.a(_12883_),
    .b(_12798_),
    .o1(_12973_));
 b15oai013an1n02x5 _21751_ (.a(_12970_),
    .b(_12971_),
    .c(net898),
    .d(_12973_),
    .o1(_12974_));
 b15oai012ah1n04x5 _21752_ (.a(_12967_),
    .b(_12974_),
    .c(_12782_),
    .o1(_12975_));
 b15bfn001as1n64x5 max_length624 (.a(net625),
    .o(net624));
 b15nanb02as1n02x5 _21754_ (.a(net906),
    .b(net886),
    .out0(_12977_));
 b15oa0022aq1n02x5 _21755_ (.a(net886),
    .b(_12960_),
    .c(_12977_),
    .d(_12851_),
    .o(_12978_));
 b15nor002ar1n03x5 _21756_ (.a(_12949_),
    .b(_12978_),
    .o1(_12979_));
 b15aoi022ah1n08x5 _21757_ (.a(net906),
    .b(_12934_),
    .c(_12979_),
    .d(net902),
    .o1(_12980_));
 b15oai012aq1n08x5 _21758_ (.a(_12975_),
    .b(_12980_),
    .c(net911),
    .o1(_12981_));
 b15aoi022an1n04x5 _21759_ (.a(_12968_),
    .b(_12909_),
    .c(_12959_),
    .d(_12851_),
    .o1(_12982_));
 b15norp02an1n12x5 _21760_ (.a(net892),
    .b(net890),
    .o1(_12983_));
 b15nand02ar1n03x5 _21761_ (.a(net902),
    .b(_12983_),
    .o1(_12984_));
 b15bfn001ah1n64x5 load_slew623 (.a(net624),
    .o(net623));
 b15nonb02ar1n08x5 _21763_ (.a(net894),
    .b(net887),
    .out0(_12986_));
 b15nor002al1n32x5 _21764_ (.a(net905),
    .b(net897),
    .o1(_12987_));
 b15aoi022al1n02x5 _21765_ (.a(net908),
    .b(_12940_),
    .c(_12986_),
    .d(_12987_),
    .o1(_12988_));
 b15oai112ah1n06x5 _21766_ (.a(net911),
    .b(_12982_),
    .c(_12984_),
    .d(_12988_),
    .o1(_12989_));
 b15nonb02an1n04x5 _21767_ (.a(net897),
    .b(net908),
    .out0(_12990_));
 b15nano23as1n24x5 _21768_ (.a(\us10.a[5] ),
    .b(net895),
    .c(net888),
    .d(net891),
    .out0(_12991_));
 b15nand02ar1n02x5 _21769_ (.a(_12990_),
    .b(_12991_),
    .o1(_12992_));
 b15nand03al1n12x5 _21770_ (.a(_12851_),
    .b(_12881_),
    .c(_12883_),
    .o1(_12993_));
 b15oaoi13al1n03x5 _21771_ (.a(net902),
    .b(_12992_),
    .c(_12993_),
    .d(_12782_),
    .o1(_12994_));
 b15nand02ar1n32x5 _21772_ (.a(_12916_),
    .b(_12798_),
    .o1(_12995_));
 b15nand02al1n02x5 _21773_ (.a(_12832_),
    .b(_12782_),
    .o1(_12996_));
 b15nor002ah1n02x5 _21774_ (.a(net892),
    .b(net899),
    .o1(_12997_));
 b15nonb02aq1n08x5 _21775_ (.a(net902),
    .b(net890),
    .out0(_12998_));
 b15aoi022al1n08x5 _21776_ (.a(_12848_),
    .b(_12997_),
    .c(_12998_),
    .d(_12811_),
    .o1(_12999_));
 b15oai022ar1n06x5 _21777_ (.a(_12844_),
    .b(_12995_),
    .c(_12996_),
    .d(_12999_),
    .o1(_13000_));
 b15bfn001as1n64x5 load_slew622 (.a(\us03.a[7] ),
    .o(net622));
 b15bfn001ah1n64x5 max_length621 (.a(\us03.a[7] ),
    .o(net621));
 b15nand02an1n16x5 _21780_ (.a(_12916_),
    .b(_12874_),
    .o1(_13003_));
 b15oai012al1n06x5 _21781_ (.a(_12950_),
    .b(_12932_),
    .c(_13003_),
    .o1(_13004_));
 b15oai013ah1n04x5 _21782_ (.a(_12989_),
    .b(_12994_),
    .c(_13000_),
    .d(_13004_),
    .o1(_13005_));
 b15aoi013ar1n02x5 _21783_ (.a(net902),
    .b(_12881_),
    .c(_12879_),
    .d(_12822_),
    .o1(_13006_));
 b15nandp2aq1n32x5 _21784_ (.a(_12881_),
    .b(_12822_),
    .o1(_13007_));
 b15aoi112ar1n02x5 _21785_ (.a(_12851_),
    .b(_13006_),
    .c(_13007_),
    .d(_12800_),
    .o1(_13008_));
 b15nandp2al1n12x5 _21786_ (.a(_12950_),
    .b(net901),
    .o1(_13009_));
 b15aoai13aq1n04x5 _21787_ (.a(_13008_),
    .b(_13009_),
    .c(_12782_),
    .d(_12991_),
    .o1(_13010_));
 b15nanb02as1n24x5 _21788_ (.a(net896),
    .b(net893),
    .out0(_13011_));
 b15orn002aq1n08x5 _21789_ (.a(net886),
    .b(net889),
    .o(_13012_));
 b15nor002as1n24x5 _21790_ (.a(_13011_),
    .b(_13012_),
    .o1(_13013_));
 b15oaoi13al1n04x5 _21791_ (.a(net908),
    .b(_13009_),
    .c(_13013_),
    .d(net902),
    .o1(_13014_));
 b15nandp2an1n48x5 _21792_ (.a(net912),
    .b(net907),
    .o1(_13015_));
 b15bfn001ah1n64x5 load_slew620 (.a(\us13.a[0] ),
    .o(net620));
 b15aoai13as1n03x5 _21794_ (.a(_12851_),
    .b(_12909_),
    .c(_13015_),
    .d(_13013_),
    .o1(_13017_));
 b15oai112ar1n16x5 _21795_ (.a(_13005_),
    .b(_13010_),
    .c(_13014_),
    .d(_13017_),
    .o1(_13018_));
 b15nor004as1n12x5 _21796_ (.a(_12839_),
    .b(_12963_),
    .c(_12981_),
    .d(_13018_),
    .o1(_13019_));
 b15xor002as1n16x5 _21797_ (.a(_12776_),
    .b(_13019_),
    .out0(_13020_));
 b15bfn001as1n64x5 max_length619 (.a(\us13.a[0] ),
    .o(net619));
 b15inv040as1n40x5 _21799_ (.a(net782),
    .o1(_13022_));
 b15bfn001as1n64x5 max_length618 (.a(\us13.a[0] ),
    .o(net618));
 b15bfn001ah1n48x5 wire617 (.a(\us13.a[1] ),
    .o(net617));
 b15bfn001as1n48x5 load_slew616 (.a(net617),
    .o(net616));
 b15bfn001as1n64x5 max_length615 (.a(net616),
    .o(net615));
 b15bfn001ah1n48x5 max_length614 (.a(net617),
    .o(net614));
 b15bfn001ah1n64x5 max_length613 (.a(\us13.a[2] ),
    .o(net613));
 b15bfn001as1n48x5 load_slew612 (.a(\us13.a[2] ),
    .o(net612));
 b15orn002al1n08x5 _21807_ (.a(net776),
    .b(net777),
    .o(_13030_));
 b15bfn001ah1n64x5 load_slew611 (.a(\us13.a[2] ),
    .o(net611));
 b15bfn001ah1n64x5 max_length610 (.a(\us13.a[3] ),
    .o(net610));
 b15orn002ah1n16x5 _21810_ (.a(net795),
    .b(net787),
    .o(_13033_));
 b15bfn001ah1n64x5 max_length609 (.a(\us13.a[3] ),
    .o(net609));
 b15bfn001as1n48x5 load_slew608 (.a(net610),
    .o(net608));
 b15bfn001ah1n64x5 wire607 (.a(\us13.a[4] ),
    .o(net607));
 b15xor002ar1n02x5 _21814_ (.a(net769),
    .b(net791),
    .out0(_13037_));
 b15nor004as1n02x5 _21815_ (.a(net773),
    .b(_13030_),
    .c(_13033_),
    .d(_13037_),
    .o1(_13038_));
 b15bfn001as1n64x5 max_length606 (.a(net607),
    .o(net606));
 b15nanb02as1n24x5 _21817_ (.a(net794),
    .b(net793),
    .out0(_13040_));
 b15bfn001ah1n64x5 load_slew605 (.a(net606),
    .o(net605));
 b15bfn001as1n64x5 max_length604 (.a(\us13.a[5] ),
    .o(net604));
 b15bfn001as1n64x5 max_length603 (.a(\us13.a[5] ),
    .o(net603));
 b15bfn001ah1n64x5 load_slew602 (.a(net603),
    .o(net602));
 b15nanb02ah1n12x5 _21822_ (.a(net773),
    .b(net769),
    .out0(_13045_));
 b15nor002aq1n12x5 _21823_ (.a(_13030_),
    .b(_13045_),
    .o1(_13046_));
 b15aoi013aq1n04x5 _21824_ (.a(_13038_),
    .b(_13040_),
    .c(net786),
    .d(_13046_),
    .o1(_13047_));
 b15bfn001as1n48x5 wire601 (.a(\us13.a[6] ),
    .o(net601));
 b15bfn001ah1n64x5 wire600 (.a(net601),
    .o(net600));
 b15nonb02as1n16x5 _21827_ (.a(net788),
    .b(net792),
    .out0(_13050_));
 b15bfn001ah1n64x5 load_slew599 (.a(net601),
    .o(net599));
 b15nand02ar1n48x5 _21829_ (.a(net770),
    .b(net772),
    .o1(_13052_));
 b15nanb02aq1n24x5 _21830_ (.a(net777),
    .b(net774),
    .out0(_13053_));
 b15norp02as1n12x5 _21831_ (.a(_13052_),
    .b(_13053_),
    .o1(_13054_));
 b15nand02ar1n02x5 _21832_ (.a(_13050_),
    .b(_13054_),
    .o1(_13055_));
 b15bfn001as1n48x5 load_slew598 (.a(\us13.a[7] ),
    .o(net598));
 b15nonb02an1n12x5 _21834_ (.a(net771),
    .b(net789),
    .out0(_13057_));
 b15bfn001as1n48x5 load_slew597 (.a(\us13.a[7] ),
    .o(net597));
 b15bfn001as1n64x5 load_slew596 (.a(net598),
    .o(net596));
 b15bfn001as1n48x5 wire595 (.a(\us23.a[0] ),
    .o(net595));
 b15bfn001ah1n64x5 load_slew594 (.a(net595),
    .o(net594));
 b15nor004ar1n08x5 _21839_ (.a(net775),
    .b(net778),
    .c(net768),
    .d(net790),
    .o1(_13062_));
 b15inv020ah1n64x5 _21840_ (.a(net793),
    .o1(_13063_));
 b15bfn001as1n48x5 max_length593 (.a(net594),
    .o(net593));
 b15nand02ar1n32x5 _21842_ (.a(net774),
    .b(net768),
    .o1(_13065_));
 b15inv000an1n16x5 _21843_ (.a(\us21.a[4] ),
    .o1(_13066_));
 b15inv000an1n64x5 _21844_ (.a(net796),
    .o1(_13067_));
 b15aoi112al1n03x5 _21845_ (.a(_13063_),
    .b(_13065_),
    .c(_13066_),
    .d(_13067_),
    .o1(_13068_));
 b15oai012aq1n08x5 _21846_ (.a(_13057_),
    .b(_13062_),
    .c(_13068_),
    .o1(_13069_));
 b15bfn001as1n48x5 max_length592 (.a(net594),
    .o(net592));
 b15bfn001as1n64x5 max_length591 (.a(net593),
    .o(net591));
 b15nonb02as1n16x5 _21849_ (.a(net793),
    .b(net794),
    .out0(_13072_));
 b15bfn001as1n48x5 load_slew590 (.a(\us23.a[1] ),
    .o(net590));
 b15bfn001as1n64x5 max_length589 (.a(net590),
    .o(net589));
 b15nona23ah1n12x5 _21852_ (.a(net774),
    .b(net768),
    .c(net771),
    .d(net777),
    .out0(_13075_));
 b15norp03ar1n02x5 _21853_ (.a(net785),
    .b(_13072_),
    .c(_13075_),
    .o1(_13076_));
 b15bfn001ah1n64x5 max_length588 (.a(net590),
    .o(net588));
 b15nanb02as1n24x5 _21855_ (.a(net774),
    .b(net777),
    .out0(_13078_));
 b15orn002an1n12x5 _21856_ (.a(net768),
    .b(net771),
    .o(_13079_));
 b15nor002ar1n04x5 _21857_ (.a(_13078_),
    .b(_13079_),
    .o1(_13080_));
 b15aoi013aq1n03x5 _21858_ (.a(_13076_),
    .b(_13080_),
    .c(_13072_),
    .d(net785),
    .o1(_13081_));
 b15nand04ah1n02x5 _21859_ (.a(_13047_),
    .b(_13055_),
    .c(_13069_),
    .d(_13081_),
    .o1(_13082_));
 b15nand02ar1n08x5 _21860_ (.a(_13022_),
    .b(_13082_),
    .o1(_13083_));
 b15bfn001as1n64x5 max_length587 (.a(net588),
    .o(net587));
 b15bfn001ah1n64x5 load_slew586 (.a(\us23.a[2] ),
    .o(net586));
 b15nona23as1n32x5 _21863_ (.a(net777),
    .b(net769),
    .c(net773),
    .d(net774),
    .out0(_13086_));
 b15bfn001as1n48x5 load_slew585 (.a(net586),
    .o(net585));
 b15bfn001as1n48x5 load_slew584 (.a(\us23.a[2] ),
    .o(net584));
 b15nanb02as1n04x5 _21866_ (.a(net786),
    .b(net796),
    .out0(_13089_));
 b15nano23as1n24x5 _21867_ (.a(net775),
    .b(net771),
    .c(\us21.a[7] ),
    .d(net778),
    .out0(_13090_));
 b15nonb02as1n16x5 _21868_ (.a(net779),
    .b(\us21.a[5] ),
    .out0(_13091_));
 b15and002as1n32x5 _21869_ (.a(\us21.a[7] ),
    .b(\us21.a[6] ),
    .o(_13092_));
 b15bfn001ah1n64x5 wire583 (.a(\us23.a[3] ),
    .o(net583));
 b15aoi013ar1n03x5 _21871_ (.a(_13090_),
    .b(_13091_),
    .c(_13092_),
    .d(net781),
    .o1(_13094_));
 b15nandp2al1n08x5 _21872_ (.a(_13067_),
    .b(net786),
    .o1(_13095_));
 b15oai022as1n06x5 _21873_ (.a(_13086_),
    .b(_13089_),
    .c(_13094_),
    .d(_13095_),
    .o1(_13096_));
 b15bfn001as1n64x5 max_length582 (.a(net583),
    .o(net582));
 b15bfn001ah1n64x5 max_length581 (.a(net583),
    .o(net581));
 b15bfn001as1n48x5 max_length580 (.a(net583),
    .o(net580));
 b15nano23as1n24x5 _21877_ (.a(net768),
    .b(net771),
    .c(net775),
    .d(net778),
    .out0(_13100_));
 b15nandp2ar1n08x5 _21878_ (.a(\us21.a[0] ),
    .b(_13100_),
    .o1(_13101_));
 b15bfn001as1n64x5 wire579 (.a(\us23.a[4] ),
    .o(net579));
 b15bfn001as1n64x5 max_length578 (.a(net579),
    .o(net578));
 b15nonb02ah1n06x5 _21881_ (.a(net768),
    .b(net775),
    .out0(_13104_));
 b15bfn001ah1n48x5 max_length577 (.a(net579),
    .o(net577));
 b15norp02aq1n02x5 _21883_ (.a(net768),
    .b(net793),
    .o1(_13106_));
 b15bfn001as1n64x5 wire576 (.a(\us23.a[5] ),
    .o(net576));
 b15aoi022aq1n08x5 _21885_ (.a(net793),
    .b(_13104_),
    .c(_13106_),
    .d(net775),
    .o1(_13108_));
 b15bfn001as1n64x5 wire575 (.a(net576),
    .o(net575));
 b15bfn001ah1n64x5 max_length574 (.a(net575),
    .o(net574));
 b15bfn001as1n64x5 load_slew573 (.a(\us23.a[6] ),
    .o(net573));
 b15nonb02aq1n04x5 _21889_ (.a(net789),
    .b(net771),
    .out0(_13112_));
 b15nandp2ar1n05x5 _21890_ (.a(net778),
    .b(_13112_),
    .o1(_13113_));
 b15inv040as1n40x5 _21891_ (.a(net788),
    .o1(_13114_));
 b15aoi022ar1n12x5 _21892_ (.a(\us21.a[0] ),
    .b(_13100_),
    .c(_13090_),
    .d(_13114_),
    .o1(_13115_));
 b15oai222as1n16x5 _21893_ (.a(net789),
    .b(_13101_),
    .c(_13108_),
    .d(_13113_),
    .e(_13115_),
    .f(net793),
    .o1(_13116_));
 b15bfn001as1n48x5 max_length572 (.a(net573),
    .o(net572));
 b15bfn001ah1n64x5 max_length571 (.a(net573),
    .o(net571));
 b15bfn001ah1n64x5 load_slew570 (.a(\us23.a[7] ),
    .o(net570));
 b15aoi022ar1n02x5 _21897_ (.a(net791),
    .b(_13096_),
    .c(_13116_),
    .d(net781),
    .o1(_13120_));
 b15bfn001as1n64x5 max_length569 (.a(\us23.a[7] ),
    .o(net569));
 b15bfn001as1n64x5 max_length568 (.a(\us23.a[7] ),
    .o(net568));
 b15bfn001ah1n64x5 load_slew567 (.a(\us33.a[0] ),
    .o(net567));
 b15norp02as1n48x5 _21901_ (.a(net788),
    .b(net782),
    .o1(_13124_));
 b15nand03as1n12x5 _21902_ (.a(_13092_),
    .b(_13091_),
    .c(_13124_),
    .o1(_13125_));
 b15nand02ah1n02x5 _21903_ (.a(net793),
    .b(_13125_),
    .o1(_13126_));
 b15nand02an1n24x5 _21904_ (.a(net787),
    .b(net780),
    .o1(_13127_));
 b15nonb02as1n16x5 _21905_ (.a(net768),
    .b(net771),
    .out0(_13128_));
 b15and002as1n32x5 _21906_ (.a(net775),
    .b(\us21.a[4] ),
    .o(_13129_));
 b15nand02an1n48x5 _21907_ (.a(_13128_),
    .b(_13129_),
    .o1(_13130_));
 b15nonb02ah1n12x5 _21908_ (.a(net768),
    .b(net778),
    .out0(_13131_));
 b15nand02as1n03x5 _21909_ (.a(_13124_),
    .b(_13131_),
    .o1(_13132_));
 b15bfn001ah1n64x5 load_slew566 (.a(\us33.a[0] ),
    .o(net566));
 b15xor002ar1n03x5 _21911_ (.a(net774),
    .b(net771),
    .out0(_13134_));
 b15oai022an1n06x5 _21912_ (.a(_13127_),
    .b(_13130_),
    .c(_13132_),
    .d(_13134_),
    .o1(_13135_));
 b15bfn001ah1n64x5 load_slew565 (.a(net567),
    .o(net565));
 b15oai112al1n12x5 _21914_ (.a(_13067_),
    .b(_13126_),
    .c(_13135_),
    .d(net793),
    .o1(_13137_));
 b15bfn001ah1n48x5 max_length564 (.a(net565),
    .o(net564));
 b15bfn001as1n64x5 max_length563 (.a(\us33.a[1] ),
    .o(net563));
 b15orn002as1n12x5 _21917_ (.a(net785),
    .b(net780),
    .o(_13140_));
 b15nona23al1n32x5 _21918_ (.a(net776),
    .b(net772),
    .c(net769),
    .d(net779),
    .out0(_13141_));
 b15nona23aq1n32x5 _21919_ (.a(net774),
    .b(net777),
    .c(net769),
    .d(net773),
    .out0(_13142_));
 b15aoi112ar1n02x5 _21920_ (.a(_13063_),
    .b(_13140_),
    .c(_13141_),
    .d(_13142_),
    .o1(_13143_));
 b15bfn001as1n64x5 max_length562 (.a(\us33.a[1] ),
    .o(net562));
 b15bfn001as1n64x5 max_length561 (.a(net563),
    .o(net561));
 b15nonb02al1n08x5 _21923_ (.a(net781),
    .b(net791),
    .out0(_13146_));
 b15nano23aq1n16x5 _21924_ (.a(net776),
    .b(net779),
    .c(net770),
    .d(net772),
    .out0(_13147_));
 b15bfn001as1n48x5 max_length560 (.a(net563),
    .o(net560));
 b15norp03an1n08x5 _21926_ (.a(_13114_),
    .b(_13079_),
    .c(_13053_),
    .o1(_13149_));
 b15oaoi13al1n02x5 _21927_ (.a(_13143_),
    .b(_13146_),
    .c(_13147_),
    .d(_13149_),
    .o1(_13150_));
 b15bfn001as1n64x5 max_length559 (.a(\us33.a[2] ),
    .o(net559));
 b15bfn001ah1n64x5 load_slew558 (.a(\us33.a[2] ),
    .o(net558));
 b15bfn001as1n48x5 max_length557 (.a(\us33.a[2] ),
    .o(net557));
 b15nanb02al1n12x5 _21931_ (.a(net768),
    .b(net777),
    .out0(_13154_));
 b15nanb03ah1n02x5 _21932_ (.a(net790),
    .b(net771),
    .c(net774),
    .out0(_13155_));
 b15nanb02ah1n16x5 _21933_ (.a(net771),
    .b(net790),
    .out0(_13156_));
 b15aoi112as1n04x5 _21934_ (.a(net780),
    .b(_13154_),
    .c(_13155_),
    .d(_13156_),
    .o1(_13157_));
 b15bfn001ah1n64x5 load_slew556 (.a(\us33.a[3] ),
    .o(net556));
 b15nona23al1n32x5 _21936_ (.a(net770),
    .b(net772),
    .c(net776),
    .d(net779),
    .out0(_13159_));
 b15nor002ah1n02x5 _21937_ (.a(net781),
    .b(_13159_),
    .o1(_13160_));
 b15ornc04ah1n24x5 _21938_ (.a(net774),
    .b(net777),
    .c(net769),
    .d(net773),
    .o(_13161_));
 b15nor002aq1n08x5 _21939_ (.a(_13022_),
    .b(_13161_),
    .o1(_13162_));
 b15oaoi13ar1n02x5 _21940_ (.a(_13157_),
    .b(net795),
    .c(_13160_),
    .d(_13162_),
    .o1(_13163_));
 b15bfn001ah1n64x5 max_length555 (.a(net556),
    .o(net555));
 b15oai022ar1n02x5 _21942_ (.a(net795),
    .b(_13150_),
    .c(_13163_),
    .d(net785),
    .o1(_13165_));
 b15nano22aq1n05x5 _21943_ (.a(_13120_),
    .b(_13137_),
    .c(_13165_),
    .out0(_13166_));
 b15bfn001ah1n64x5 load_slew554 (.a(\us33.a[3] ),
    .o(net554));
 b15bfn001ah1n48x5 load_slew553 (.a(net554),
    .o(net553));
 b15bfn001ah1n64x5 load_slew552 (.a(\us33.a[4] ),
    .o(net552));
 b15bfn001ah1n64x5 wire551 (.a(\us33.a[4] ),
    .o(net551));
 b15nano23as1n24x5 _21948_ (.a(net776),
    .b(net770),
    .c(net772),
    .d(net779),
    .out0(_13171_));
 b15bfn001as1n48x5 max_length550 (.a(net552),
    .o(net550));
 b15nandp2ar1n04x5 _21950_ (.a(net784),
    .b(_13171_),
    .o1(_13173_));
 b15inv020an1n32x5 _21951_ (.a(net774),
    .o1(_13174_));
 b15bfn001as1n64x5 max_length549 (.a(\us33.a[5] ),
    .o(net549));
 b15norp02as1n48x5 _21953_ (.a(net770),
    .b(net772),
    .o1(_13176_));
 b15bfn001ah1n48x5 load_slew548 (.a(net549),
    .o(net548));
 b15oai112an1n04x5 _21955_ (.a(_13174_),
    .b(_13176_),
    .c(_13022_),
    .d(_13066_),
    .o1(_13178_));
 b15oai012aq1n06x5 _21956_ (.a(_13173_),
    .b(_13178_),
    .c(_13067_),
    .o1(_13179_));
 b15bfn001as1n48x5 max_length547 (.a(net549),
    .o(net547));
 b15andc04as1n16x5 _21958_ (.a(net776),
    .b(net779),
    .c(net770),
    .d(net772),
    .o(_13181_));
 b15aoi012ar1n02x5 _21959_ (.a(net795),
    .b(net790),
    .c(_13181_),
    .o1(_13182_));
 b15nand02al1n04x5 _21960_ (.a(net790),
    .b(_13171_),
    .o1(_13183_));
 b15norp02as1n48x5 _21961_ (.a(net774),
    .b(net777),
    .o1(_13184_));
 b15nandp2ah1n32x5 _21962_ (.a(_13184_),
    .b(_13128_),
    .o1(_13185_));
 b15aoi013an1n03x5 _21963_ (.a(_13182_),
    .b(_13183_),
    .c(_13185_),
    .d(net795),
    .o1(_13186_));
 b15bfn001as1n64x5 max_length546 (.a(\us33.a[6] ),
    .o(net546));
 b15bfn001ah1n64x5 max_length545 (.a(\us33.a[6] ),
    .o(net545));
 b15norp03ar1n03x5 _21966_ (.a(net769),
    .b(net794),
    .c(net783),
    .o1(_13189_));
 b15bfn001as1n48x5 load_slew544 (.a(\us33.a[7] ),
    .o(net544));
 b15aoai13ah1n04x5 _21968_ (.a(_13184_),
    .b(_13189_),
    .c(net769),
    .d(net783),
    .o1(_13191_));
 b15bfn001ah1n64x5 wire543 (.a(\us33.a[7] ),
    .o(net543));
 b15orn002aq1n12x5 _21970_ (.a(net794),
    .b(net783),
    .o(_13193_));
 b15nandp2ah1n08x5 _21971_ (.a(net774),
    .b(net777),
    .o1(_13194_));
 b15oai013as1n12x5 _21972_ (.a(_13191_),
    .b(_13193_),
    .c(_13194_),
    .d(net769),
    .o1(_13195_));
 b15nonb02aq1n06x5 _21973_ (.a(net793),
    .b(net771),
    .out0(_13196_));
 b15aoi222aq1n06x5 _21974_ (.a(_13063_),
    .b(_13179_),
    .c(_13186_),
    .d(net783),
    .e(_13195_),
    .f(_13196_),
    .o1(_13197_));
 b15bfn001ah1n48x5 max_length542 (.a(ld_r),
    .o(net542));
 b15bfn001as1n48x5 max_length541 (.a(ld_r),
    .o(net541));
 b15bfn001ah1n64x5 max_length540 (.a(net542),
    .o(net540));
 b15xor002ar1n02x5 _21978_ (.a(\us21.a[4] ),
    .b(net773),
    .out0(_13201_));
 b15nor004aq1n03x5 _21979_ (.a(_13174_),
    .b(net792),
    .c(net784),
    .d(_13201_),
    .o1(_13202_));
 b15and002aq1n12x5 _21980_ (.a(\us21.a[6] ),
    .b(net784),
    .o(_13203_));
 b15aoi012an1n06x5 _21981_ (.a(_13202_),
    .b(_13203_),
    .c(_13184_),
    .o1(_13204_));
 b15bfn001as1n48x5 max_length539 (.a(net540),
    .o(net539));
 b15nanb02an1n16x5 _21983_ (.a(\us21.a[0] ),
    .b(net768),
    .out0(_13206_));
 b15oaoi13as1n08x5 _21984_ (.a(_13114_),
    .b(_13197_),
    .c(_13204_),
    .d(_13206_),
    .o1(_13207_));
 b15nonb02as1n16x5 _21985_ (.a(net776),
    .b(net779),
    .out0(_13208_));
 b15nandp3al1n24x5 _21986_ (.a(net784),
    .b(_13092_),
    .c(_13208_),
    .o1(_13209_));
 b15nand02as1n16x5 _21987_ (.a(net794),
    .b(net787),
    .o1(_13210_));
 b15nanb02as1n24x5 _21988_ (.a(net782),
    .b(net788),
    .out0(_13211_));
 b15bfn001ah1n64x5 max_length538 (.a(ld_r),
    .o(net538));
 b15nano23as1n24x5 _21990_ (.a(net779),
    .b(net772),
    .c(net770),
    .d(net776),
    .out0(_13213_));
 b15nandp2al1n03x5 _21991_ (.a(net793),
    .b(_13213_),
    .o1(_13214_));
 b15nonb02as1n16x5 _21992_ (.a(net784),
    .b(net789),
    .out0(_13215_));
 b15bfn001as1n48x5 max_length537 (.a(net538),
    .o(net537));
 b15nonb02ah1n16x5 _21994_ (.a(net794),
    .b(net790),
    .out0(_13217_));
 b15aoi013al1n03x5 _21995_ (.a(_13215_),
    .b(_13217_),
    .c(_13174_),
    .d(net787),
    .o1(_13218_));
 b15and002aq1n12x5 _21996_ (.a(net778),
    .b(net768),
    .o(_13219_));
 b15nand02an1n02x5 _21997_ (.a(net773),
    .b(_13219_),
    .o1(_13220_));
 b15oai222aq1n08x5 _21998_ (.a(_13209_),
    .b(_13210_),
    .c(_13211_),
    .d(_13214_),
    .e(_13218_),
    .f(_13220_),
    .o1(_13221_));
 b15nonb02as1n16x5 _21999_ (.a(net773),
    .b(net769),
    .out0(_13222_));
 b15bfn001ah1n64x5 max_length536 (.a(net537),
    .o(net536));
 b15nandp3al1n04x5 _22001_ (.a(net795),
    .b(net791),
    .c(net786),
    .o1(_13224_));
 b15nand04aq1n08x5 _22002_ (.a(net781),
    .b(_13033_),
    .c(_13222_),
    .d(_13224_),
    .o1(_13225_));
 b15aoi012al1n04x5 _22003_ (.a(_13184_),
    .b(_13129_),
    .c(net786),
    .o1(_13226_));
 b15nandp2aq1n32x5 _22004_ (.a(_13184_),
    .b(_13222_),
    .o1(_13227_));
 b15norp02as1n12x5 _22005_ (.a(net795),
    .b(net791),
    .o1(_13228_));
 b15aoi112as1n08x5 _22006_ (.a(_13225_),
    .b(_13226_),
    .c(_13227_),
    .d(_13228_),
    .o1(_13229_));
 b15nandp2al1n02x5 _22007_ (.a(net795),
    .b(_13215_),
    .o1(_13230_));
 b15nonb02al1n12x5 _22008_ (.a(\us21.a[4] ),
    .b(\us21.a[7] ),
    .out0(_13231_));
 b15and002an1n02x5 _22009_ (.a(net773),
    .b(net792),
    .o(_13232_));
 b15nor002ar1n08x5 _22010_ (.a(net771),
    .b(net793),
    .o1(_13233_));
 b15nonb03ah1n02x5 _22011_ (.a(\us21.a[7] ),
    .b(\us21.a[4] ),
    .c(net775),
    .out0(_13234_));
 b15aoi022ar1n02x5 _22012_ (.a(_13231_),
    .b(_13232_),
    .c(_13233_),
    .d(_13234_),
    .o1(_13235_));
 b15norp02aq1n03x5 _22013_ (.a(_13230_),
    .b(_13235_),
    .o1(_13236_));
 b15nor002an1n12x5 _22014_ (.a(net778),
    .b(net768),
    .o1(_13237_));
 b15inv020as1n03x5 _22015_ (.a(_13237_),
    .o1(_13238_));
 b15nonb03ah1n12x5 _22016_ (.a(net787),
    .b(net780),
    .c(net794),
    .out0(_13239_));
 b15nor002ar1n06x5 _22017_ (.a(net774),
    .b(net790),
    .o1(_13240_));
 b15nand03ar1n04x5 _22018_ (.a(net771),
    .b(_13239_),
    .c(_13240_),
    .o1(_13241_));
 b15nor003ar1n02x5 _22019_ (.a(net774),
    .b(net787),
    .c(net780),
    .o1(_13242_));
 b15bfn001ah1n48x5 max_length535 (.a(net538),
    .o(net535));
 b15and002aq1n24x5 _22021_ (.a(net786),
    .b(net783),
    .o(_13244_));
 b15oaoi13as1n03x5 _22022_ (.a(_13242_),
    .b(net774),
    .c(_13244_),
    .d(_13239_),
    .o1(_13245_));
 b15oaoi13aq1n08x5 _22023_ (.a(_13238_),
    .b(_13241_),
    .c(_13245_),
    .d(_13156_),
    .o1(_13246_));
 b15nor004an1n04x5 _22024_ (.a(_13221_),
    .b(_13229_),
    .c(_13236_),
    .d(_13246_),
    .o1(_13247_));
 b15nandp3an1n04x5 _22025_ (.a(_13213_),
    .b(_13215_),
    .c(_13217_),
    .o1(_13248_));
 b15nor004as1n12x5 _22026_ (.a(net776),
    .b(net779),
    .c(net770),
    .d(net772),
    .o1(_13249_));
 b15bfn001as1n48x5 max_length534 (.a(ld_r),
    .o(net534));
 b15nonb02as1n16x5 _22028_ (.a(net786),
    .b(net783),
    .out0(_13251_));
 b15and002as1n16x5 _22029_ (.a(\us21.a[0] ),
    .b(net792),
    .o(_13252_));
 b15nand03an1n06x5 _22030_ (.a(_13249_),
    .b(_13251_),
    .c(_13252_),
    .o1(_13253_));
 b15orn002as1n04x5 _22031_ (.a(net792),
    .b(net785),
    .o(_13254_));
 b15nand03as1n24x5 _22032_ (.a(_13022_),
    .b(_13176_),
    .c(_13208_),
    .o1(_13255_));
 b15oai112al1n16x5 _22033_ (.a(_13248_),
    .b(_13253_),
    .c(_13254_),
    .d(_13255_),
    .o1(_13256_));
 b15norp03as1n02x5 _22034_ (.a(net771),
    .b(net793),
    .c(net783),
    .o1(_13257_));
 b15nonb03aq1n02x5 _22035_ (.a(\us21.a[0] ),
    .b(net789),
    .c(net775),
    .out0(_13258_));
 b15and002aq1n03x5 _22036_ (.a(net775),
    .b(net789),
    .o(_13259_));
 b15oai112ah1n06x5 _22037_ (.a(_13219_),
    .b(_13257_),
    .c(_13258_),
    .d(_13259_),
    .o1(_13260_));
 b15oai012ah1n06x5 _22038_ (.a(_13260_),
    .b(_13209_),
    .c(_13033_),
    .o1(_13261_));
 b15and002aq1n12x5 _22039_ (.a(net793),
    .b(net789),
    .o(_13262_));
 b15and002ar1n08x5 _22040_ (.a(net778),
    .b(net795),
    .o(_13263_));
 b15nano23ah1n02x5 _22041_ (.a(net771),
    .b(net783),
    .c(net775),
    .d(net768),
    .out0(_13264_));
 b15nano23ar1n03x5 _22042_ (.a(net775),
    .b(net768),
    .c(net771),
    .d(net783),
    .out0(_13265_));
 b15oai112aq1n08x5 _22043_ (.a(_13262_),
    .b(_13263_),
    .c(_13264_),
    .d(_13265_),
    .o1(_13266_));
 b15nano22as1n08x5 _22044_ (.a(net795),
    .b(net787),
    .c(net780),
    .out0(_13267_));
 b15nand02as1n03x5 _22045_ (.a(_13090_),
    .b(_13267_),
    .o1(_13268_));
 b15nandp3as1n08x5 _22046_ (.a(_13092_),
    .b(_13208_),
    .c(_13215_),
    .o1(_13269_));
 b15aoai13al1n08x5 _22047_ (.a(_13266_),
    .b(_13063_),
    .c(_13268_),
    .d(_13269_),
    .o1(_13270_));
 b15nand03al1n02x5 _22048_ (.a(_13124_),
    .b(_13176_),
    .c(_13208_),
    .o1(_13271_));
 b15nand02al1n24x5 _22049_ (.a(net792),
    .b(_13249_),
    .o1(_13272_));
 b15oaoi13aq1n04x5 _22050_ (.a(net795),
    .b(_13271_),
    .c(_13272_),
    .d(_13127_),
    .o1(_13273_));
 b15nor004as1n12x5 _22051_ (.a(_13256_),
    .b(_13261_),
    .c(_13270_),
    .d(_13273_),
    .o1(_13274_));
 b15nand02al1n02x5 _22052_ (.a(_13176_),
    .b(_13215_),
    .o1(_13275_));
 b15bfn001ah1n64x5 load_slew533 (.a(net534),
    .o(net533));
 b15nanb02as1n24x5 _22054_ (.a(net791),
    .b(net795),
    .out0(_13277_));
 b15bfn001ah1n24x5 wire532 (.a(\u0.w[0][1] ),
    .o(net532));
 b15nandp3an1n02x5 _22056_ (.a(_13091_),
    .b(_13040_),
    .c(_13277_),
    .o1(_13279_));
 b15oaoi13al1n04x5 _22057_ (.a(_13275_),
    .b(_13279_),
    .c(_13053_),
    .d(_13228_),
    .o1(_13280_));
 b15bfn001as1n24x5 wire531 (.a(\u0.w[2][1] ),
    .o(net531));
 b15nand04ah1n04x5 _22059_ (.a(net795),
    .b(_13129_),
    .c(_13222_),
    .d(_13254_),
    .o1(_13282_));
 b15nand02ah1n06x5 _22060_ (.a(_13114_),
    .b(_13277_),
    .o1(_13283_));
 b15bfn001ah1n32x5 wire530 (.a(\u0.w[2][3] ),
    .o(net530));
 b15oaoi13an1n03x5 _22062_ (.a(net781),
    .b(_13282_),
    .c(_13283_),
    .d(_13130_),
    .o1(_13285_));
 b15xor002aq1n08x5 _22063_ (.a(net771),
    .b(net789),
    .out0(_13286_));
 b15aoi022as1n06x5 _22064_ (.a(_13057_),
    .b(_13219_),
    .c(_13237_),
    .d(_13286_),
    .o1(_13287_));
 b15nor004an1n06x5 _22065_ (.a(_13174_),
    .b(net783),
    .c(_13277_),
    .d(_13287_),
    .o1(_13288_));
 b15nand04al1n06x5 _22066_ (.a(_13184_),
    .b(_13196_),
    .c(_13206_),
    .d(_13215_),
    .o1(_13289_));
 b15nand03aq1n03x5 _22067_ (.a(_13022_),
    .b(_13050_),
    .c(_13090_),
    .o1(_13290_));
 b15inv000ah1n16x5 _22068_ (.a(net771),
    .o1(_13291_));
 b15nand04as1n12x5 _22069_ (.a(net775),
    .b(_13291_),
    .c(net795),
    .d(net783),
    .o1(_13292_));
 b15aoi022ar1n02x5 _22070_ (.a(_13063_),
    .b(_13131_),
    .c(_13231_),
    .d(_13262_),
    .o1(_13293_));
 b15oai112ah1n06x5 _22071_ (.a(_13289_),
    .b(_13290_),
    .c(_13292_),
    .d(_13293_),
    .o1(_13294_));
 b15nor004ah1n04x5 _22072_ (.a(_13280_),
    .b(_13285_),
    .c(_13288_),
    .d(_13294_),
    .o1(_13295_));
 b15nandp3aq1n12x5 _22073_ (.o1(_13296_),
    .a(_13247_),
    .b(_13274_),
    .c(_13295_));
 b15nano23as1n24x5 _22074_ (.a(_13083_),
    .b(_13166_),
    .c(_13207_),
    .d(_13296_),
    .out0(_13297_));
 b15bfn001ah1n24x5 wire529 (.a(\u0.w[2][8] ),
    .o(net529));
 b15bfn001ah1n24x5 wire528 (.a(\u0.w[2][9] ),
    .o(net528));
 b15bfn001as1n24x5 wire527 (.a(\u0.w[2][16] ),
    .o(net527));
 b15bfn001as1n24x5 wire526 (.a(\u0.w[2][17] ),
    .o(net526));
 b15orn002ah1n32x5 _22079_ (.a(net643),
    .b(net647),
    .o(_13302_));
 b15bfn001as1n24x5 wire525 (.a(\u0.w[2][18] ),
    .o(net525));
 b15bfn001as1n24x5 wire524 (.a(\u0.w[2][19] ),
    .o(net524));
 b15bfn001as1n24x5 wire523 (.a(\u0.w[2][24] ),
    .o(net523));
 b15nanb02as1n24x5 _22083_ (.a(net654),
    .b(net650),
    .out0(_13306_));
 b15bfn001as1n24x5 wire522 (.a(\u0.w[2][25] ),
    .o(net522));
 b15bfn001as1n24x5 wire521 (.a(\u0.w[2][26] ),
    .o(net521));
 b15bfn001as1n48x5 load_slew520 (.a(\u0.tmp_w[0] ),
    .o(net520));
 b15nand02aq1n24x5 _22087_ (.a(net666),
    .b(net655),
    .o1(_13310_));
 b15norp03aq1n02x5 _22088_ (.a(_13302_),
    .b(_13306_),
    .c(_13310_),
    .o1(_13311_));
 b15bfn001as1n48x5 load_slew519 (.a(net520),
    .o(net519));
 b15inv020aq1n64x5 _22090_ (.a(net655),
    .o1(_13313_));
 b15bfn001as1n48x5 max_length518 (.a(net520),
    .o(net518));
 b15nanb02as1n24x5 _22092_ (.a(net646),
    .b(net643),
    .out0(_13315_));
 b15bfn001as1n48x5 load_slew517 (.a(\u0.tmp_w[1] ),
    .o(net517));
 b15bfn001ah1n64x5 max_length516 (.a(net517),
    .o(net516));
 b15nandp2ah1n48x5 _22095_ (.a(net649),
    .b(net652),
    .o1(_13318_));
 b15bfn001as1n48x5 max_length515 (.a(net517),
    .o(net515));
 b15norp02ar1n08x5 _22097_ (.a(_13315_),
    .b(_13318_),
    .o1(_13320_));
 b15bfn001as1n48x5 max_length514 (.a(\u0.tmp_w[1] ),
    .o(net514));
 b15bfn001as1n64x5 max_length513 (.a(\u0.tmp_w[2] ),
    .o(net513));
 b15bfn001as1n64x5 max_length512 (.a(\u0.tmp_w[2] ),
    .o(net512));
 b15nanb02as1n24x5 _22101_ (.a(net649),
    .b(net652),
    .out0(_13324_));
 b15norp03aq1n16x5 _22102_ (.a(net659),
    .b(_13324_),
    .c(_13302_),
    .o1(_13325_));
 b15oaoi13al1n04x5 _22103_ (.a(_13311_),
    .b(_13313_),
    .c(_13320_),
    .d(_13325_),
    .o1(_13326_));
 b15bfn001as1n64x5 max_length511 (.a(net512),
    .o(net511));
 b15bfn001as1n48x5 load_slew510 (.a(net511),
    .o(net510));
 b15bfn001ah1n64x5 load_slew509 (.a(\u0.tmp_w[3] ),
    .o(net509));
 b15nona23as1n32x5 _22107_ (.a(net645),
    .b(net648),
    .c(net651),
    .d(net653),
    .out0(_13330_));
 b15bfn001as1n48x5 wire508 (.a(net509),
    .o(net508));
 b15bfn001ah1n64x5 wire507 (.a(net509),
    .o(net507));
 b15bfn001ah1n64x5 load_slew506 (.a(\u0.tmp_w[4] ),
    .o(net506));
 b15bfn001as1n64x5 max_length505 (.a(\u0.tmp_w[4] ),
    .o(net505));
 b15bfn001as1n64x5 max_length504 (.a(\u0.tmp_w[4] ),
    .o(net504));
 b15nand04as1n16x5 _22113_ (.a(net651),
    .b(net653),
    .c(net645),
    .d(net648),
    .o1(_13336_));
 b15bfn001ah1n48x5 load_slew503 (.a(net506),
    .o(net503));
 b15nona22ah1n04x5 _22115_ (.a(net665),
    .b(net661),
    .c(net657),
    .out0(_13338_));
 b15oai022an1n12x5 _22116_ (.a(net657),
    .b(_13330_),
    .c(_13336_),
    .d(_13338_),
    .o1(_13339_));
 b15inv000as1n64x5 _22117_ (.a(\us32.a[1] ),
    .o1(_13340_));
 b15bfn001ah1n64x5 wire502 (.a(\u0.tmp_w[5] ),
    .o(net502));
 b15bfn001as1n64x5 load_slew501 (.a(net502),
    .o(net501));
 b15nandp2as1n48x5 _22120_ (.a(net643),
    .b(net647),
    .o1(_13343_));
 b15bfn001as1n64x5 max_length500 (.a(net501),
    .o(net500));
 b15nanb02as1n24x5 _22122_ (.a(net662),
    .b(net656),
    .out0(_13345_));
 b15nor004an1n04x5 _22123_ (.a(_13340_),
    .b(_13324_),
    .c(_13343_),
    .d(_13345_),
    .o1(_13346_));
 b15nanb02as1n24x5 _22124_ (.a(net655),
    .b(net660),
    .out0(_13347_));
 b15bfn001as1n48x5 max_length499 (.a(net502),
    .o(net499));
 b15nor003al1n04x5 _22126_ (.a(_13306_),
    .b(_13343_),
    .c(_13347_),
    .o1(_13349_));
 b15orn002al1n32x5 _22127_ (.a(net649),
    .b(net652),
    .o(_13350_));
 b15bfn001ah1n48x5 wire498 (.a(\u0.tmp_w[6] ),
    .o(net498));
 b15nor004ar1n06x5 _22129_ (.a(net663),
    .b(_13315_),
    .c(_13347_),
    .d(_13350_),
    .o1(_13352_));
 b15nor004ar1n08x5 _22130_ (.a(_13339_),
    .b(_13346_),
    .c(_13349_),
    .d(_13352_),
    .o1(_13353_));
 b15bfn001ah1n64x5 load_slew497 (.a(net498),
    .o(net497));
 b15inv000ah1n64x5 _22132_ (.a(net668),
    .o1(_13355_));
 b15bfn001ah1n64x5 load_slew496 (.a(net497),
    .o(net496));
 b15bfn001as1n48x5 wire495 (.a(net498),
    .o(net495));
 b15oai022al1n12x5 _22135_ (.a(net663),
    .b(_13326_),
    .c(_13353_),
    .d(_13355_),
    .o1(_13358_));
 b15bfn001ah1n64x5 wire494 (.a(\u0.tmp_w[7] ),
    .o(net494));
 b15bfn001ah1n64x5 load_slew493 (.a(net494),
    .o(net493));
 b15nano23as1n24x5 _22138_ (.a(net651),
    .b(net648),
    .c(net645),
    .d(net653),
    .out0(_13361_));
 b15norp02ah1n48x5 _22139_ (.a(net658),
    .b(net662),
    .o1(_13362_));
 b15bfn001ah1n64x5 load_slew492 (.a(net493),
    .o(net492));
 b15nand02ar1n02x5 _22141_ (.a(_13361_),
    .b(_13362_),
    .o1(_13364_));
 b15bfn001as1n48x5 load_slew491 (.a(net493),
    .o(net491));
 b15bfn001ah1n64x5 wire490 (.a(\u0.tmp_w[8] ),
    .o(net490));
 b15nanb02as1n24x5 _22144_ (.a(net666),
    .b(net659),
    .out0(_13367_));
 b15nor002an1n08x5 _22145_ (.a(net663),
    .b(_13367_),
    .o1(_13368_));
 b15bfn001ah1n64x5 load_slew489 (.a(net490),
    .o(net489));
 b15bfn001as1n48x5 max_length488 (.a(net490),
    .o(net488));
 b15nonb02as1n16x5 _22148_ (.a(net663),
    .b(net659),
    .out0(_13371_));
 b15bfn001as1n48x5 max_length487 (.a(net488),
    .o(net487));
 b15inv000aq1n06x5 _22150_ (.a(net649),
    .o1(_13373_));
 b15inv000al1n24x5 _22151_ (.a(net654),
    .o1(_13374_));
 b15and002aq1n32x5 _22152_ (.a(net645),
    .b(net648),
    .o(_13375_));
 b15bfn001ah1n48x5 max_length486 (.a(net488),
    .o(net486));
 b15nand04ah1n16x5 _22154_ (.a(net655),
    .b(_13373_),
    .c(_13374_),
    .d(_13375_),
    .o1(_13377_));
 b15oai013al1n03x5 _22155_ (.a(_13364_),
    .b(_13368_),
    .c(_13371_),
    .d(_13377_),
    .o1(_13378_));
 b15bfn001as1n64x5 max_length485 (.a(\u0.tmp_w[9] ),
    .o(net485));
 b15and002al1n32x5 _22157_ (.a(\us32.a[1] ),
    .b(net658),
    .o(_13380_));
 b15bfn001ah1n64x5 load_slew484 (.a(\u0.tmp_w[9] ),
    .o(net484));
 b15nonb02ah1n16x5 _22159_ (.a(net647),
    .b(net644),
    .out0(_13382_));
 b15nand02ar1n02x5 _22160_ (.a(_13380_),
    .b(_13382_),
    .o1(_13383_));
 b15bfn001as1n48x5 wire483 (.a(net485),
    .o(net483));
 b15nonb02as1n16x5 _22162_ (.a(net651),
    .b(net653),
    .out0(_13385_));
 b15bfn001ah1n64x5 max_length482 (.a(\u0.tmp_w[10] ),
    .o(net482));
 b15norp02as1n04x5 _22164_ (.a(net668),
    .b(net662),
    .o1(_13387_));
 b15nonb02as1n16x5 _22165_ (.a(net654),
    .b(net650),
    .out0(_13388_));
 b15aoi022ar1n02x5 _22166_ (.a(net660),
    .b(_13385_),
    .c(_13387_),
    .d(_13388_),
    .o1(_13389_));
 b15nona23as1n32x5 _22167_ (.a(net652),
    .b(net646),
    .c(net643),
    .d(net649),
    .out0(_13390_));
 b15bfn001as1n64x5 max_length481 (.a(net482),
    .o(net481));
 b15nanb02aq1n24x5 _22169_ (.a(net663),
    .b(net656),
    .out0(_13392_));
 b15oai022an1n04x5 _22170_ (.a(_13383_),
    .b(_13389_),
    .c(_13390_),
    .d(_13392_),
    .o1(_13393_));
 b15bfn001as1n48x5 load_slew480 (.a(net481),
    .o(net480));
 b15bfn001ah1n64x5 load_slew479 (.a(net481),
    .o(net479));
 b15norp02aq1n02x5 _22173_ (.a(net668),
    .b(net658),
    .o1(_13396_));
 b15and003al1n08x5 _22174_ (.a(net654),
    .b(net643),
    .c(net647),
    .o(_13397_));
 b15orn002an1n16x5 _22175_ (.a(\us32.a[1] ),
    .b(net650),
    .o(_13398_));
 b15nandp2aq1n32x5 _22176_ (.a(net662),
    .b(net650),
    .o1(_13399_));
 b15bfn001ah1n64x5 wire478 (.a(\u0.tmp_w[11] ),
    .o(net478));
 b15nand04aq1n04x5 _22178_ (.a(_13396_),
    .b(_13397_),
    .c(_13398_),
    .d(_13399_),
    .o1(_13401_));
 b15norp02ah1n32x5 _22179_ (.a(net645),
    .b(net648),
    .o1(_13402_));
 b15nor002ah1n24x5 _22180_ (.a(net663),
    .b(net655),
    .o1(_13403_));
 b15aoi022ar1n02x5 _22181_ (.a(_13402_),
    .b(_13380_),
    .c(_13403_),
    .d(_13375_),
    .o1(_13404_));
 b15bfn001ah1n48x5 wire477 (.a(net478),
    .o(net477));
 b15bfn001ah1n64x5 load_slew476 (.a(\u0.tmp_w[11] ),
    .o(net476));
 b15nonb02an1n12x5 _22184_ (.a(net650),
    .b(net662),
    .out0(_13407_));
 b15nand02an1n03x5 _22185_ (.a(net654),
    .b(_13407_),
    .o1(_13408_));
 b15oa0012al1n06x5 _22186_ (.a(_13401_),
    .b(_13404_),
    .c(_13408_),
    .o(_13409_));
 b15and002al1n32x5 _22187_ (.a(net658),
    .b(net662),
    .o(_13410_));
 b15bfn001as1n64x5 max_length475 (.a(\u0.tmp_w[12] ),
    .o(net475));
 b15nor002as1n08x5 _22189_ (.a(net667),
    .b(_13330_),
    .o1(_13412_));
 b15nandp2ar1n04x5 _22190_ (.a(_13410_),
    .b(_13412_),
    .o1(_13413_));
 b15nona23ar1n12x5 _22191_ (.a(_13378_),
    .b(_13393_),
    .c(_13409_),
    .d(_13413_),
    .out0(_13414_));
 b15nano23as1n24x5 _22192_ (.a(net653),
    .b(net645),
    .c(net648),
    .d(net651),
    .out0(_13415_));
 b15nand02aq1n24x5 _22193_ (.a(net657),
    .b(_13415_),
    .o1(_13416_));
 b15nonb02as1n16x5 _22194_ (.a(net668),
    .b(\us32.a[1] ),
    .out0(_13417_));
 b15nonb02as1n16x5 _22195_ (.a(net665),
    .b(net667),
    .out0(_13418_));
 b15bfn001as1n48x5 max_length474 (.a(\u0.tmp_w[12] ),
    .o(net474));
 b15norp03ar1n02x5 _22197_ (.a(net660),
    .b(_13417_),
    .c(_13418_),
    .o1(_13420_));
 b15inv000an1n64x5 _22198_ (.a(net659),
    .o1(_13421_));
 b15bfn001as1n48x5 load_slew473 (.a(\u0.tmp_w[12] ),
    .o(net473));
 b15nanb02as1n24x5 _22200_ (.a(net663),
    .b(net666),
    .out0(_13423_));
 b15bfn001ah1n64x5 max_length472 (.a(\u0.tmp_w[13] ),
    .o(net472));
 b15nanb02as1n24x5 _22202_ (.a(net666),
    .b(net663),
    .out0(_13425_));
 b15bfn001as1n48x5 max_length471 (.a(\u0.tmp_w[13] ),
    .o(net471));
 b15aoi012ar1n02x5 _22204_ (.a(_13421_),
    .b(_13423_),
    .c(_13425_),
    .o1(_13427_));
 b15orn003ah1n02x5 _22205_ (.a(_13416_),
    .b(_13420_),
    .c(_13427_),
    .o(_13428_));
 b15bfn001as1n48x5 load_slew470 (.a(net471),
    .o(net470));
 b15nonb02ar1n08x5 _22207_ (.a(net650),
    .b(net647),
    .out0(_13430_));
 b15nand02an1n32x5 _22208_ (.a(net654),
    .b(net644),
    .o1(_13431_));
 b15norp02ar1n08x5 _22209_ (.a(net668),
    .b(_13431_),
    .o1(_13432_));
 b15bfn001as1n64x5 max_length469 (.a(net470),
    .o(net469));
 b15nonb02ar1n06x5 _22211_ (.a(net654),
    .b(net644),
    .out0(_13434_));
 b15nonb02as1n04x5 _22212_ (.a(net644),
    .b(net654),
    .out0(_13435_));
 b15nor003ah1n04x5 _22213_ (.a(net662),
    .b(_13434_),
    .c(_13435_),
    .o1(_13436_));
 b15oai112ah1n12x5 _22214_ (.a(_13380_),
    .b(_13430_),
    .c(_13432_),
    .d(_13436_),
    .o1(_13437_));
 b15norp02aq1n16x5 _22215_ (.a(_13306_),
    .b(_13343_),
    .o1(_13438_));
 b15aoi012al1n04x5 _22216_ (.a(_13313_),
    .b(_13423_),
    .c(_13438_),
    .o1(_13439_));
 b15bfn001ah1n64x5 load_slew468 (.a(\u0.tmp_w[14] ),
    .o(net468));
 b15nanb02as1n24x5 _22218_ (.a(net645),
    .b(net648),
    .out0(_13441_));
 b15norp02ar1n48x5 _22219_ (.a(_13318_),
    .b(_13441_),
    .o1(_13442_));
 b15bfn001as1n64x5 max_length467 (.a(net468),
    .o(net467));
 b15oai112ah1n06x5 _22221_ (.a(net660),
    .b(_13425_),
    .c(_13442_),
    .d(net656),
    .o1(_13444_));
 b15oai112aq1n16x5 _22222_ (.a(_13428_),
    .b(_13437_),
    .c(_13439_),
    .d(_13444_),
    .o1(_13445_));
 b15bfn001ah1n64x5 load_slew466 (.a(net468),
    .o(net466));
 b15orn002an1n24x5 _22224_ (.a(net657),
    .b(net661),
    .o(_13447_));
 b15nor002an1n03x5 _22225_ (.a(_13423_),
    .b(_13447_),
    .o1(_13448_));
 b15bfn001as1n64x5 max_length465 (.a(\u0.tmp_w[15] ),
    .o(net465));
 b15nanb03an1n08x5 _22227_ (.a(net656),
    .b(net660),
    .c(net666),
    .out0(_13450_));
 b15aoi012al1n02x5 _22228_ (.a(_13340_),
    .b(_13345_),
    .c(_13450_),
    .o1(_13451_));
 b15oai112ar1n06x5 _22229_ (.a(_13373_),
    .b(_13382_),
    .c(_13448_),
    .d(_13451_),
    .o1(_13452_));
 b15bfn001as1n64x5 max_length464 (.a(\u0.tmp_w[15] ),
    .o(net464));
 b15nanb02aq1n12x5 _22231_ (.a(net666),
    .b(net655),
    .out0(_13454_));
 b15nor002as1n03x5 _22232_ (.a(net646),
    .b(_13454_),
    .o1(_13455_));
 b15bfn001ah1n64x5 load_slew463 (.a(net464),
    .o(net463));
 b15bfn001as1n48x5 load_slew462 (.a(net463),
    .o(net462));
 b15bfn001ah1n64x5 load_slew461 (.a(\u0.tmp_w[16] ),
    .o(net461));
 b15inv040as1n16x5 _22236_ (.a(net647),
    .o1(_13459_));
 b15rm6013en1n04x5 _22237_ (.a(net663),
    .b(net666),
    .c(_13459_),
    .carryb(_13460_));
 b15aoai13ah1n04x5 _22238_ (.a(net643),
    .b(_13455_),
    .c(_13460_),
    .d(_13362_),
    .o1(_13461_));
 b15oaoi13as1n04x5 _22239_ (.a(net652),
    .b(_13452_),
    .c(_13461_),
    .d(_13373_),
    .o1(_13462_));
 b15nor004as1n12x5 _22240_ (.a(_13358_),
    .b(_13414_),
    .c(_13445_),
    .d(_13462_),
    .o1(_13463_));
 b15bfn001ah1n64x5 max_length460 (.a(net461),
    .o(net460));
 b15bfn001ah1n64x5 wire459 (.a(\u0.tmp_w[16] ),
    .o(net459));
 b15oai012an1n02x5 _22243_ (.a(net663),
    .b(_13306_),
    .c(_13343_),
    .o1(_13466_));
 b15oai022an1n08x5 _22244_ (.a(_13315_),
    .b(_13350_),
    .c(_13441_),
    .d(_13318_),
    .o1(_13467_));
 b15bfn001as1n64x5 max_length458 (.a(\u0.tmp_w[17] ),
    .o(net458));
 b15oai112aq1n08x5 _22246_ (.a(net657),
    .b(_13466_),
    .c(_13467_),
    .d(net663),
    .o1(_13469_));
 b15bfn001as1n64x5 max_length457 (.a(\u0.tmp_w[17] ),
    .o(net457));
 b15bfn001ah1n64x5 max_length456 (.a(net457),
    .o(net456));
 b15norp02aq1n02x5 _22249_ (.a(_13355_),
    .b(net657),
    .o1(_13472_));
 b15aoi012al1n02x5 _22250_ (.a(net661),
    .b(_13442_),
    .c(_13472_),
    .o1(_13473_));
 b15bfn001ah1n48x5 max_length455 (.a(net457),
    .o(net455));
 b15bfn001as1n48x5 max_length454 (.a(\u0.tmp_w[18] ),
    .o(net454));
 b15bfn001ah1n64x5 wire453 (.a(\u0.tmp_w[18] ),
    .o(net453));
 b15norp02as1n03x5 _22254_ (.a(net653),
    .b(_13343_),
    .o1(_13477_));
 b15and002al1n16x5 _22255_ (.a(net658),
    .b(net651),
    .o(_13478_));
 b15nona22ah1n24x5 _22256_ (.a(net645),
    .b(net648),
    .c(\us32.a[4] ),
    .out0(_13479_));
 b15bfn001ah1n64x5 load_slew452 (.a(net453),
    .o(net452));
 b15nor002ar1n06x5 _22258_ (.a(net665),
    .b(net653),
    .o1(_13481_));
 b15aob012an1n04x5 _22259_ (.a(_13479_),
    .b(_13375_),
    .c(_13481_),
    .out0(_13482_));
 b15norp02ar1n12x5 _22260_ (.a(net657),
    .b(net651),
    .o1(_13483_));
 b15aoi022ah1n12x5 _22261_ (.a(_13477_),
    .b(_13478_),
    .c(_13482_),
    .d(_13483_),
    .o1(_13484_));
 b15oai112al1n06x5 _22262_ (.a(_13469_),
    .b(_13473_),
    .c(net667),
    .d(_13484_),
    .o1(_13485_));
 b15nor004as1n12x5 _22263_ (.a(net651),
    .b(net653),
    .c(net645),
    .d(net648),
    .o1(_13486_));
 b15nandp3as1n03x5 _22264_ (.a(_13355_),
    .b(net657),
    .c(_13486_),
    .o1(_13487_));
 b15nandp2an1n32x5 _22265_ (.a(net665),
    .b(net667),
    .o1(_13488_));
 b15nanb02aq1n16x5 _22266_ (.a(_13479_),
    .b(_13483_),
    .out0(_13489_));
 b15oai112ar1n06x5 _22267_ (.a(net661),
    .b(_13487_),
    .c(_13488_),
    .d(_13489_),
    .o1(_13490_));
 b15nand02al1n12x5 _22268_ (.a(net657),
    .b(_13486_),
    .o1(_13491_));
 b15oaoi13ar1n03x5 _22269_ (.a(net665),
    .b(_13491_),
    .c(_13489_),
    .d(net667),
    .o1(_13492_));
 b15oai012an1n06x5 _22270_ (.a(_13485_),
    .b(_13490_),
    .c(_13492_),
    .o1(_13493_));
 b15nona23as1n32x5 _22271_ (.a(net652),
    .b(net643),
    .c(net646),
    .d(net649),
    .out0(_13494_));
 b15bfn001ah1n64x5 wire451 (.a(\u0.tmp_w[19] ),
    .o(net451));
 b15nano23as1n24x5 _22273_ (.a(net652),
    .b(net646),
    .c(net643),
    .d(net649),
    .out0(_13496_));
 b15nandp2al1n03x5 _22274_ (.a(net657),
    .b(_13496_),
    .o1(_13497_));
 b15aoi112ar1n02x5 _22275_ (.a(net665),
    .b(net661),
    .c(_13494_),
    .d(_13497_),
    .o1(_13498_));
 b15nandp2ah1n16x5 _22276_ (.a(net657),
    .b(net661),
    .o1(_13499_));
 b15nona23as1n32x5 _22277_ (.a(net649),
    .b(net643),
    .c(net646),
    .d(net652),
    .out0(_13500_));
 b15bfn001as1n64x5 max_length450 (.a(net451),
    .o(net450));
 b15oai022al1n02x5 _22279_ (.a(net657),
    .b(_13494_),
    .c(_13499_),
    .d(_13500_),
    .o1(_13502_));
 b15aoai13an1n03x5 _22280_ (.a(net667),
    .b(_13498_),
    .c(_13502_),
    .d(net665),
    .o1(_13503_));
 b15nanb02aq1n16x5 _22281_ (.a(net657),
    .b(net667),
    .out0(_13504_));
 b15nonb02as1n16x5 _22282_ (.a(net644),
    .b(net647),
    .out0(_13505_));
 b15and002aq1n16x5 _22283_ (.a(net649),
    .b(net652),
    .o(_13506_));
 b15nand02aq1n06x5 _22284_ (.a(_13505_),
    .b(_13506_),
    .o1(_13507_));
 b15oai022al1n04x5 _22285_ (.a(_13336_),
    .b(_13454_),
    .c(_13504_),
    .d(_13507_),
    .o1(_13508_));
 b15nand02ar1n16x5 _22286_ (.a(_13388_),
    .b(_13375_),
    .o1(_13509_));
 b15nand02ah1n16x5 _22287_ (.a(_13385_),
    .b(_13375_),
    .o1(_13510_));
 b15nanb02as1n16x5 _22288_ (.a(net655),
    .b(net663),
    .out0(_13511_));
 b15oai022aq1n06x5 _22289_ (.a(_13392_),
    .b(_13509_),
    .c(_13510_),
    .d(_13511_),
    .o1(_13512_));
 b15nano22ar1n05x5 _22290_ (.a(net649),
    .b(net652),
    .c(net664),
    .out0(_13513_));
 b15orn002ah1n16x5 _22291_ (.a(net665),
    .b(net667),
    .o(_13514_));
 b15norp02an1n32x5 _22292_ (.a(net650),
    .b(net654),
    .o1(_13515_));
 b15aoai13ah1n03x5 _22293_ (.a(_13375_),
    .b(_13513_),
    .c(_13514_),
    .d(_13515_),
    .o1(_13516_));
 b15bfn001as1n64x5 max_length449 (.a(net451),
    .o(net449));
 b15nonb02aq1n06x5 _22295_ (.a(net647),
    .b(net650),
    .out0(_13518_));
 b15nona22as1n08x5 _22296_ (.a(_13434_),
    .b(_13435_),
    .c(_13518_),
    .out0(_13519_));
 b15oai022aq1n12x5 _22297_ (.a(net656),
    .b(_13516_),
    .c(_13519_),
    .d(_13310_),
    .o1(_13520_));
 b15oai013ar1n06x5 _22298_ (.a(net659),
    .b(_13508_),
    .c(_13512_),
    .d(_13520_),
    .o1(_13521_));
 b15nano22ah1n06x5 _22299_ (.a(net654),
    .b(net647),
    .c(net644),
    .out0(_13522_));
 b15and002ah1n16x5 _22300_ (.a(net668),
    .b(net661),
    .o(_13523_));
 b15oai112al1n12x5 _22301_ (.a(_13478_),
    .b(_13522_),
    .c(_13523_),
    .d(_13418_),
    .o1(_13524_));
 b15bfn001as1n48x5 load_slew448 (.a(net449),
    .o(net448));
 b15nand04al1n08x5 _22303_ (.a(_13313_),
    .b(_13421_),
    .c(_13505_),
    .d(_13515_),
    .o1(_13526_));
 b15aoai13ah1n08x5 _22304_ (.a(_13524_),
    .b(_13526_),
    .c(_13488_),
    .d(_13514_),
    .o1(_13527_));
 b15nonb02aq1n16x5 _22305_ (.a(net666),
    .b(net660),
    .out0(_13528_));
 b15oai012aq1n03x5 _22306_ (.a(_13528_),
    .b(_13496_),
    .c(_13415_),
    .o1(_13529_));
 b15nandp2an1n12x5 _22307_ (.a(net665),
    .b(net661),
    .o1(_13530_));
 b15nandp2al1n16x5 _22308_ (.a(_13505_),
    .b(_13388_),
    .o1(_13531_));
 b15oaoi13al1n08x5 _22309_ (.a(net655),
    .b(_13529_),
    .c(_13530_),
    .d(_13531_),
    .o1(_13532_));
 b15orn002ar1n16x5 _22310_ (.a(net651),
    .b(net645),
    .o(_13533_));
 b15and002ah1n12x5 _22311_ (.a(\us32.a[4] ),
    .b(net648),
    .o(_13534_));
 b15oai012as1n03x5 _22312_ (.a(_13534_),
    .b(_13418_),
    .c(_13417_),
    .o1(_13535_));
 b15norp02as1n08x5 _22313_ (.a(\us32.a[4] ),
    .b(net648),
    .o1(_13536_));
 b15nand03an1n06x5 _22314_ (.a(_13423_),
    .b(_13425_),
    .c(_13536_),
    .o1(_13537_));
 b15aoi112ah1n06x5 _22315_ (.a(_13347_),
    .b(_13533_),
    .c(_13535_),
    .d(_13537_),
    .o1(_13538_));
 b15nandp3ar1n02x5 _22316_ (.a(net657),
    .b(_13388_),
    .c(_13402_),
    .o1(_13539_));
 b15nanb02aq1n04x5 _22317_ (.a(net665),
    .b(net659),
    .out0(_13540_));
 b15nand04aq1n03x5 _22318_ (.a(_13313_),
    .b(_13402_),
    .c(_13385_),
    .d(_13540_),
    .o1(_13541_));
 b15oai022ar1n02x5 _22319_ (.a(net667),
    .b(_13499_),
    .c(_13504_),
    .d(net661),
    .o1(_13542_));
 b15aoi022an1n02x5 _22320_ (.a(_13539_),
    .b(_13541_),
    .c(_13542_),
    .d(net665),
    .o1(_13543_));
 b15nor004an1n06x5 _22321_ (.a(_13527_),
    .b(_13532_),
    .c(_13538_),
    .d(_13543_),
    .o1(_13544_));
 b15and003as1n03x5 _22322_ (.a(_13503_),
    .b(_13521_),
    .c(_13544_),
    .o(_13545_));
 b15and003as1n24x5 _22323_ (.a(_13463_),
    .b(_13493_),
    .c(_13545_),
    .o(_13546_));
 b15nanb02as1n24x5 _22324_ (.a(net635),
    .b(net639),
    .out0(_13547_));
 b15andc04as1n16x5 _22325_ (.a(\us03.a[5] ),
    .b(\us03.a[4] ),
    .c(\us03.a[7] ),
    .d(net625),
    .o(_13548_));
 b15nandp2aq1n03x5 _22326_ (.a(net633),
    .b(_13548_),
    .o1(_13549_));
 b15oai022aq1n02x5 _22327_ (.a(_12565_),
    .b(_13547_),
    .c(_13549_),
    .d(net642),
    .o1(_13550_));
 b15nandp2aq1n02x5 _22328_ (.a(net633),
    .b(_12752_),
    .o1(_13551_));
 b15aoi012al1n02x5 _22329_ (.a(_12615_),
    .b(_13551_),
    .c(_12565_),
    .o1(_13552_));
 b15nandp2aq1n03x5 _22330_ (.a(_12519_),
    .b(_12643_),
    .o1(_13553_));
 b15aoi012al1n02x5 _22331_ (.a(_12563_),
    .b(_12523_),
    .c(net638),
    .o1(_13554_));
 b15nona22an1n08x5 _22332_ (.a(net638),
    .b(net634),
    .c(net624),
    .out0(_13555_));
 b15nor002ah1n06x5 _22333_ (.a(net627),
    .b(_12671_),
    .o1(_13556_));
 b15aoi022aq1n08x5 _22334_ (.a(net627),
    .b(_12723_),
    .c(_13556_),
    .d(_12662_),
    .o1(_13557_));
 b15oai022ah1n06x5 _22335_ (.a(_13553_),
    .b(_13554_),
    .c(_13555_),
    .d(_13557_),
    .o1(_13558_));
 b15oai013ah1n04x5 _22336_ (.a(net632),
    .b(_13550_),
    .c(_13552_),
    .d(_13558_),
    .o1(_13559_));
 b15orn003ar1n16x5 _22337_ (.a(net638),
    .b(net631),
    .c(net634),
    .o(_13560_));
 b15aoi112ar1n02x5 _22338_ (.a(_12550_),
    .b(_12718_),
    .c(_12697_),
    .d(net641),
    .o1(_13561_));
 b15oaoi13aq1n03x5 _22339_ (.a(_13560_),
    .b(_13561_),
    .c(net641),
    .d(_12771_),
    .o1(_13562_));
 b15xor002ah1n12x5 _22340_ (.a(net638),
    .b(net641),
    .out0(_13563_));
 b15and002ah1n04x5 _22341_ (.a(_12646_),
    .b(_13563_),
    .o(_13564_));
 b15nonb02as1n16x5 _22342_ (.a(net640),
    .b(net637),
    .out0(_13565_));
 b15aoi012an1n02x5 _22343_ (.a(_12697_),
    .b(_13565_),
    .c(_13548_),
    .o1(_13566_));
 b15and002ah1n16x5 _22344_ (.a(net630),
    .b(net633),
    .o(_13567_));
 b15nand02an1n04x5 _22345_ (.a(_13567_),
    .b(_13565_),
    .o1(_13568_));
 b15obai22aq1n08x5 _22346_ (.a(_13564_),
    .b(_13566_),
    .c(_12594_),
    .d(_13568_),
    .out0(_13569_));
 b15nandp2ah1n24x5 _22347_ (.a(\us03.a[1] ),
    .b(\us03.a[0] ),
    .o1(_13570_));
 b15aoi013an1n02x5 _22348_ (.a(net632),
    .b(_12586_),
    .c(_12593_),
    .d(_13570_),
    .o1(_13571_));
 b15oai112aq1n02x5 _22349_ (.a(_12586_),
    .b(_12593_),
    .c(_12654_),
    .d(net638),
    .o1(_13572_));
 b15aoi112ah1n03x5 _22350_ (.a(net633),
    .b(_13571_),
    .c(_13572_),
    .d(_12684_),
    .o1(_13573_));
 b15bfn001as1n48x5 load_slew447 (.a(\u0.tmp_w[20] ),
    .o(net447));
 b15nor003ah1n02x5 _22352_ (.a(net637),
    .b(net633),
    .c(_12613_),
    .o1(_13575_));
 b15aoai13al1n06x5 _22353_ (.a(net640),
    .b(_13575_),
    .c(_12718_),
    .d(_12598_),
    .o1(_13576_));
 b15norp03ar1n03x5 _22354_ (.a(net637),
    .b(_12601_),
    .c(_12677_),
    .o1(_13577_));
 b15oai012ar1n06x5 _22355_ (.a(_12511_),
    .b(_12599_),
    .c(_13577_),
    .o1(_13578_));
 b15nona23ar1n12x5 _22356_ (.a(_13569_),
    .b(_13573_),
    .c(_13576_),
    .d(_13578_),
    .out0(_13579_));
 b15nanb02as1n24x5 _22357_ (.a(net630),
    .b(net636),
    .out0(_13580_));
 b15bfn001ah1n64x5 load_slew446 (.a(\u0.tmp_w[20] ),
    .o(net446));
 b15nor003ah1n02x5 _22359_ (.a(net639),
    .b(_13580_),
    .c(_12760_),
    .o1(_13582_));
 b15nor002an1n03x5 _22360_ (.a(_12566_),
    .b(_12654_),
    .o1(_13583_));
 b15bfn001as1n48x5 max_length445 (.a(net447),
    .o(net445));
 b15nor003as1n03x5 _22362_ (.a(_12766_),
    .b(_12552_),
    .c(_13580_),
    .o1(_13585_));
 b15oaoi13an1n08x5 _22363_ (.a(_13582_),
    .b(net639),
    .c(_13583_),
    .d(_13585_),
    .o1(_13586_));
 b15oai012aq1n03x5 _22364_ (.a(_12648_),
    .b(_12753_),
    .c(_13580_),
    .o1(_13587_));
 b15aob012aq1n04x5 _22365_ (.a(_13586_),
    .b(_13587_),
    .c(net638),
    .out0(_13588_));
 b15norp02al1n12x5 _22366_ (.a(net640),
    .b(_12591_),
    .o1(_13589_));
 b15nand03an1n03x5 _22367_ (.a(net637),
    .b(_13548_),
    .c(_13589_),
    .o1(_13590_));
 b15oai022ar1n04x5 _22368_ (.a(_12553_),
    .b(_12601_),
    .c(_12591_),
    .d(_12766_),
    .o1(_13591_));
 b15aoi022al1n06x5 _22369_ (.a(_12523_),
    .b(_12646_),
    .c(_13591_),
    .d(_12511_),
    .o1(_13592_));
 b15oai013ah1n06x5 _22370_ (.a(_13590_),
    .b(_13592_),
    .c(_12549_),
    .d(net637),
    .o1(_13593_));
 b15nor004ar1n08x5 _22371_ (.a(_13562_),
    .b(_13579_),
    .c(_13588_),
    .d(_13593_),
    .o1(_13594_));
 b15nano22ar1n24x5 _22372_ (.a(\us03.a[4] ),
    .b(net621),
    .c(net624),
    .out0(_13595_));
 b15aoai13as1n02x5 _22373_ (.a(net631),
    .b(_12610_),
    .c(_13595_),
    .d(net634),
    .o1(_13596_));
 b15nandp2ar1n03x5 _22374_ (.a(net634),
    .b(_12610_),
    .o1(_13597_));
 b15aoi112ah1n04x5 _22375_ (.a(net627),
    .b(_13570_),
    .c(_13596_),
    .d(_13597_),
    .o1(_13598_));
 b15nanb02as1n24x5 _22376_ (.a(net641),
    .b(net634),
    .out0(_13599_));
 b15norp03ar1n02x5 _22377_ (.a(net638),
    .b(net631),
    .c(net627),
    .o1(_13600_));
 b15aoi012ar1n02x5 _22378_ (.a(_13600_),
    .b(_12722_),
    .c(net638),
    .o1(_13601_));
 b15inv020aq1n12x5 _22379_ (.a(net623),
    .o1(_13602_));
 b15nona23as1n05x5 _22380_ (.a(_13599_),
    .b(_13601_),
    .c(_12723_),
    .d(_13602_),
    .out0(_13603_));
 b15nor003aq1n02x5 _22381_ (.a(_12545_),
    .b(_12683_),
    .c(_12771_),
    .o1(_13604_));
 b15nor002aq1n06x5 _22382_ (.a(_12707_),
    .b(_12646_),
    .o1(_13605_));
 b15orn002as1n24x5 _22383_ (.a(net626),
    .b(net628),
    .o(_13606_));
 b15norp02al1n16x5 _22384_ (.a(_12569_),
    .b(_13606_),
    .o1(_13607_));
 b15aoi013al1n06x5 _22385_ (.a(_13604_),
    .b(_13605_),
    .c(_13565_),
    .d(_13607_),
    .o1(_13608_));
 b15bfn001as1n48x5 load_slew444 (.a(net447),
    .o(net444));
 b15oai022ar1n04x5 _22387_ (.a(_12553_),
    .b(_13570_),
    .c(_13563_),
    .d(_12766_),
    .o1(_13610_));
 b15nand03ar1n08x5 _22388_ (.a(_12587_),
    .b(_13567_),
    .c(_13610_),
    .o1(_13611_));
 b15norp03ar1n04x5 _22389_ (.a(_12511_),
    .b(net621),
    .c(_12547_),
    .o1(_13612_));
 b15nor002ar1n03x5 _22390_ (.a(net624),
    .b(_13580_),
    .o1(_13613_));
 b15aoai13al1n08x5 _22391_ (.a(_13612_),
    .b(_13613_),
    .c(net624),
    .d(_13605_),
    .o1(_13614_));
 b15nand04as1n16x5 _22392_ (.a(_13603_),
    .b(_13608_),
    .c(_13611_),
    .d(_13614_),
    .o1(_13615_));
 b15nor002ar1n08x5 _22393_ (.a(net639),
    .b(_12545_),
    .o1(_13616_));
 b15aoi012ar1n02x5 _22394_ (.a(_12766_),
    .b(_12580_),
    .c(net624),
    .o1(_13617_));
 b15nanb02an1n02x5 _22395_ (.a(net627),
    .b(net635),
    .out0(_13618_));
 b15nandp2al1n03x5 _22396_ (.a(\us03.a[4] ),
    .b(net624),
    .o1(_13619_));
 b15nor002al1n02x5 _22397_ (.a(_13618_),
    .b(_13619_),
    .o1(_13620_));
 b15oai112aq1n06x5 _22398_ (.a(net621),
    .b(_13616_),
    .c(_13617_),
    .d(_13620_),
    .o1(_13621_));
 b15norp02ar1n02x5 _22399_ (.a(_12683_),
    .b(_12771_),
    .o1(_13622_));
 b15aoai13aq1n03x5 _22400_ (.a(_12545_),
    .b(_13622_),
    .c(_12700_),
    .d(_12554_),
    .o1(_13623_));
 b15nor002aq1n06x5 _22401_ (.a(_12581_),
    .b(_12750_),
    .o1(_13624_));
 b15aoai13al1n04x5 _22402_ (.a(_12707_),
    .b(_13624_),
    .c(_12581_),
    .d(_12550_),
    .o1(_13625_));
 b15nor003al1n06x5 _22403_ (.a(_12511_),
    .b(_12591_),
    .c(_12677_),
    .o1(_13626_));
 b15nor004an1n08x5 _22404_ (.a(_12549_),
    .b(_13606_),
    .c(_12591_),
    .d(_13563_),
    .o1(_13627_));
 b15norp02ar1n24x5 _22405_ (.a(_12766_),
    .b(_12717_),
    .o1(_13628_));
 b15aoi112as1n08x5 _22406_ (.a(_13626_),
    .b(_13627_),
    .c(_13628_),
    .d(_12598_),
    .o1(_13629_));
 b15nand04aq1n12x5 _22407_ (.a(_13621_),
    .b(_13623_),
    .c(_13625_),
    .d(_13629_),
    .o1(_13630_));
 b15aoi112ah1n04x5 _22408_ (.a(_12591_),
    .b(_13570_),
    .c(_12750_),
    .d(_12714_),
    .o1(_13631_));
 b15nor004ah1n02x5 _22409_ (.a(net628),
    .b(_12552_),
    .c(_12722_),
    .d(_12725_),
    .o1(_13632_));
 b15and003ar1n02x5 _22410_ (.a(net628),
    .b(_12595_),
    .c(_12651_),
    .o(_13633_));
 b15oai012ar1n03x5 _22411_ (.a(_12717_),
    .b(_12552_),
    .c(net634),
    .o1(_13634_));
 b15aoi112al1n03x5 _22412_ (.a(_13631_),
    .b(_13632_),
    .c(_13633_),
    .d(_13634_),
    .o1(_13635_));
 b15norp03ar1n02x5 _22413_ (.a(net631),
    .b(net634),
    .c(_12613_),
    .o1(_13636_));
 b15and003ar1n02x5 _22414_ (.a(net627),
    .b(_12595_),
    .c(_12707_),
    .o(_13637_));
 b15oaoi13ah1n02x5 _22415_ (.a(_13636_),
    .b(_13637_),
    .c(_13595_),
    .d(_12610_),
    .o1(_13638_));
 b15nano23al1n02x5 _22416_ (.a(_12587_),
    .b(_12722_),
    .c(_13547_),
    .d(net628),
    .out0(_13639_));
 b15nanb02aq1n02x5 _22417_ (.a(net635),
    .b(net627),
    .out0(_13640_));
 b15norp03ah1n03x5 _22418_ (.a(_12552_),
    .b(_13640_),
    .c(_12754_),
    .o1(_13641_));
 b15nor002an1n03x5 _22419_ (.a(_13639_),
    .b(_13641_),
    .o1(_13642_));
 b15nor004al1n02x5 _22420_ (.a(_12766_),
    .b(_12552_),
    .c(_12580_),
    .d(_12629_),
    .o1(_13643_));
 b15and002al1n16x5 _22421_ (.a(net639),
    .b(net635),
    .o(_13644_));
 b15aoi013al1n03x5 _22422_ (.a(_13643_),
    .b(_13644_),
    .c(_12611_),
    .d(net631),
    .o1(_13645_));
 b15nand04an1n08x5 _22423_ (.a(_13635_),
    .b(_13638_),
    .c(_13642_),
    .d(_13645_),
    .o1(_13646_));
 b15nor004ah1n08x5 _22424_ (.a(_13598_),
    .b(_13615_),
    .c(_13630_),
    .d(_13646_),
    .o1(_13647_));
 b15bfn001as1n48x5 load_slew443 (.a(\u0.tmp_w[21] ),
    .o(net443));
 b15aoi022ar1n04x5 _22426_ (.a(_12570_),
    .b(_13567_),
    .c(_12718_),
    .d(_13589_),
    .o1(_13649_));
 b15mdn022ah1n04x5 _22427_ (.a(_12689_),
    .b(_12726_),
    .o1(_13650_),
    .sa(_12581_));
 b15aoi022aq1n02x5 _22428_ (.a(_12707_),
    .b(_13565_),
    .c(_13650_),
    .d(net630),
    .o1(_13651_));
 b15oai022aq1n08x5 _22429_ (.a(_12581_),
    .b(_13649_),
    .c(_13651_),
    .d(_12714_),
    .o1(_13652_));
 b15aoai13ah1n03x5 _22430_ (.a(net642),
    .b(_12570_),
    .c(_12538_),
    .d(_12606_),
    .o1(_13653_));
 b15orn002as1n04x5 _22431_ (.a(\us03.a[5] ),
    .b(net624),
    .o(_13654_));
 b15norp03as1n02x5 _22432_ (.a(net642),
    .b(\us03.a[4] ),
    .c(_13654_),
    .o1(_13655_));
 b15and002as1n04x5 _22433_ (.a(net628),
    .b(net623),
    .o(_13656_));
 b15aoi012an1n06x5 _22434_ (.a(_13655_),
    .b(_13656_),
    .c(\us03.a[5] ),
    .o1(_13657_));
 b15oai013ar1n12x5 _22435_ (.a(_13653_),
    .b(_13657_),
    .c(\us03.a[7] ),
    .d(net639),
    .o1(_13658_));
 b15nandp3ar1n02x5 _22436_ (.a(net641),
    .b(_12597_),
    .c(_12720_),
    .o1(_13659_));
 b15orn002ar1n08x5 _22437_ (.a(net627),
    .b(net621),
    .o(_13660_));
 b15oai013al1n04x5 _22438_ (.a(_13659_),
    .b(_13660_),
    .c(net624),
    .d(_12601_),
    .o1(_13661_));
 b15aoi122an1n04x5 _22439_ (.a(_13652_),
    .b(_13658_),
    .c(_12707_),
    .d(_12581_),
    .e(_13661_),
    .o1(_13662_));
 b15andc04as1n16x5 _22440_ (.a(_13559_),
    .b(_13594_),
    .c(_13647_),
    .d(_13662_),
    .o(_13663_));
 b15xnr002as1n16x5 _22441_ (.a(_13546_),
    .b(_13663_),
    .out0(_13664_));
 b15xor002aq1n12x5 _22442_ (.a(_13297_),
    .b(_13664_),
    .out0(_13665_));
 b15xor002as1n16x5 _22443_ (.a(_13020_),
    .b(_13665_),
    .out0(_13666_));
 b15bfn001as1n64x5 max_length442 (.a(net443),
    .o(net442));
 b15bfn001as1n64x5 max_length441 (.a(net443),
    .o(net441));
 b15bfn001as1n48x5 load_slew440 (.a(net441),
    .o(net440));
 b15mdn022ar1n02x5 _22447_ (.a(_12505_),
    .b(_13666_),
    .o1(_13670_),
    .sa(net537));
 b15xor002ar1n02x5 _22448_ (.a(net520),
    .b(_13670_),
    .out0(_00121_));
 b15bfn001ah1n64x5 load_slew439 (.a(\u0.tmp_w[22] ),
    .o(net439));
 b15nanb02aq1n06x5 _22450_ (.a(\text_in_r[1] ),
    .b(net533),
    .out0(_13672_));
 b15nandp2as1n08x5 _22451_ (.a(_12636_),
    .b(_13595_),
    .o1(_13673_));
 b15oai122an1n02x5 _22452_ (.a(net640),
    .b(_12566_),
    .c(_12709_),
    .d(_12751_),
    .e(_13673_),
    .o1(_13674_));
 b15nor004al1n02x5 _22453_ (.a(_12581_),
    .b(_12569_),
    .c(_13606_),
    .d(_12601_),
    .o1(_13675_));
 b15norp02ah1n04x5 _22454_ (.a(net639),
    .b(net635),
    .o1(_13676_));
 b15ao0022ar1n02x5 _22455_ (.a(\us03.a[5] ),
    .b(_13644_),
    .c(_13676_),
    .d(_12523_),
    .o(_13677_));
 b15aoi013al1n03x5 _22456_ (.a(_13675_),
    .b(_13677_),
    .c(_12587_),
    .d(_12545_),
    .o1(_13678_));
 b15nor004an1n03x5 _22457_ (.a(net631),
    .b(net628),
    .c(_12717_),
    .d(_13640_),
    .o1(_13679_));
 b15aoi013aq1n06x5 _22458_ (.a(_13679_),
    .b(_12554_),
    .c(net635),
    .d(net631),
    .o1(_13680_));
 b15oai112aq1n12x5 _22459_ (.a(_12511_),
    .b(_13678_),
    .c(_13680_),
    .d(net639),
    .o1(_13681_));
 b15and002al1n04x5 _22460_ (.a(_13674_),
    .b(_13681_),
    .o(_13682_));
 b15norp02al1n48x5 _22461_ (.a(_12549_),
    .b(_13606_),
    .o1(_13683_));
 b15aoai13as1n02x5 _22462_ (.a(_12643_),
    .b(_12550_),
    .c(net638),
    .d(_13683_),
    .o1(_13684_));
 b15oai022ar1n12x5 _22463_ (.a(_13599_),
    .b(_12524_),
    .c(_12600_),
    .d(_12738_),
    .o1(_13685_));
 b15nanb02as1n24x5 _22464_ (.a(net639),
    .b(\us03.a[2] ),
    .out0(_13686_));
 b15nano22ah1n03x5 _22465_ (.a(_12610_),
    .b(_12675_),
    .c(_13686_),
    .out0(_13687_));
 b15nano23aq1n24x5 _22466_ (.a(net622),
    .b(net625),
    .c(net626),
    .d(net629),
    .out0(_13688_));
 b15aoi012ar1n02x5 _22467_ (.a(net632),
    .b(_12579_),
    .c(_13688_),
    .o1(_13689_));
 b15oai013al1n03x5 _22468_ (.a(_13689_),
    .b(_12643_),
    .c(_12619_),
    .d(_12581_),
    .o1(_13690_));
 b15nor003aq1n06x5 _22469_ (.a(_13685_),
    .b(_13687_),
    .c(_13690_),
    .o1(_13691_));
 b15bfn001ah1n64x5 load_slew438 (.a(\u0.tmp_w[22] ),
    .o(net438));
 b15nandp3ar1n02x5 _22471_ (.a(_12511_),
    .b(\us03.a[2] ),
    .c(_12597_),
    .o1(_13693_));
 b15oaoi13ah1n02x5 _22472_ (.a(net639),
    .b(_13693_),
    .c(_13673_),
    .d(_12511_),
    .o1(_13694_));
 b15nandp2ah1n05x5 _22473_ (.a(net635),
    .b(_12597_),
    .o1(_13695_));
 b15oab012al1n02x5 _22474_ (.a(_13694_),
    .b(_13695_),
    .c(_13570_),
    .out0(_13696_));
 b15aoi022ah1n06x5 _22475_ (.a(_13684_),
    .b(_13691_),
    .c(_13696_),
    .d(net632),
    .o1(_13697_));
 b15bfn001as1n48x5 load_slew437 (.a(net439),
    .o(net437));
 b15aoai13an1n02x5 _22477_ (.a(net630),
    .b(_12752_),
    .c(_12645_),
    .d(_12581_),
    .o1(_13699_));
 b15norp02an1n24x5 _22478_ (.a(net641),
    .b(net631),
    .o1(_13700_));
 b15nor003ah1n08x5 _22479_ (.a(net627),
    .b(net621),
    .c(net623),
    .o1(_13701_));
 b15aoi022ar1n24x5 _22480_ (.a(_12587_),
    .b(_12722_),
    .c(_13700_),
    .d(_13701_),
    .o1(_13702_));
 b15oaoi13aq1n04x5 _22481_ (.a(_12515_),
    .b(_13699_),
    .c(_13702_),
    .d(_12745_),
    .o1(_13703_));
 b15aoi012ar1n02x5 _22482_ (.a(_12591_),
    .b(_12603_),
    .c(_12762_),
    .o1(_13704_));
 b15aoai13ar1n02x5 _22483_ (.a(_12677_),
    .b(net640),
    .c(net637),
    .d(_12750_),
    .o1(_13705_));
 b15aoi012aq1n02x5 _22484_ (.a(_13703_),
    .b(_13704_),
    .c(_13705_),
    .o1(_13706_));
 b15nand02an1n08x5 _22485_ (.a(\us03.a[5] ),
    .b(net624),
    .o1(_13707_));
 b15aoi012al1n04x5 _22486_ (.a(_12632_),
    .b(_12637_),
    .c(net642),
    .o1(_13708_));
 b15nor003ah1n03x5 _22487_ (.a(_13547_),
    .b(_13707_),
    .c(_13708_),
    .o1(_13709_));
 b15nandp2ah1n03x5 _22488_ (.a(net635),
    .b(_12697_),
    .o1(_13710_));
 b15nor002ar1n08x5 _22489_ (.a(net634),
    .b(_12700_),
    .o1(_13711_));
 b15nano23an1n24x5 _22490_ (.a(\us03.a[5] ),
    .b(net622),
    .c(net625),
    .d(\us03.a[4] ),
    .out0(_13712_));
 b15aob012al1n02x5 _22491_ (.a(_13710_),
    .b(_13711_),
    .c(_13712_),
    .out0(_13713_));
 b15oai012ar1n06x5 _22492_ (.a(net632),
    .b(_13709_),
    .c(_13713_),
    .o1(_13714_));
 b15nandp2aq1n03x5 _22493_ (.a(\us03.a[1] ),
    .b(_12657_),
    .o1(_13715_));
 b15aoi012ar1n02x5 _22494_ (.a(_13715_),
    .b(_12684_),
    .c(\us03.a[3] ),
    .o1(_13716_));
 b15nonb02an1n08x5 _22495_ (.a(net627),
    .b(net624),
    .out0(_13717_));
 b15norp03ar1n02x5 _22496_ (.a(\us03.a[2] ),
    .b(\us03.a[4] ),
    .c(\us03.a[7] ),
    .o1(_13718_));
 b15aoai13as1n03x5 _22497_ (.a(_13717_),
    .b(_13718_),
    .c(\us03.a[2] ),
    .d(_12637_),
    .o1(_13719_));
 b15aob012ar1n06x5 _22498_ (.a(_13716_),
    .b(_13719_),
    .c(_12545_),
    .out0(_13720_));
 b15and003as1n04x5 _22499_ (.a(_13706_),
    .b(_13714_),
    .c(_13720_),
    .o(_13721_));
 b15nanb02al1n12x5 _22500_ (.a(net637),
    .b(net630),
    .out0(_13722_));
 b15norp02ah1n04x5 _22501_ (.a(_12515_),
    .b(_13722_),
    .o1(_13723_));
 b15norp02ar1n02x5 _22502_ (.a(net641),
    .b(_12771_),
    .o1(_13724_));
 b15aoai13an1n03x5 _22503_ (.a(_13723_),
    .b(_13724_),
    .c(_12550_),
    .d(net641),
    .o1(_13725_));
 b15norp02al1n02x5 _22504_ (.a(_13606_),
    .b(_13547_),
    .o1(_13726_));
 b15nanb02al1n24x5 _22505_ (.a(net630),
    .b(net641),
    .out0(_13727_));
 b15oai012al1n02x5 _22506_ (.a(_12717_),
    .b(_13727_),
    .c(_13602_),
    .o1(_13728_));
 b15oai012an1n02x5 _22507_ (.a(_12747_),
    .b(_13580_),
    .c(net641),
    .o1(_13729_));
 b15nor003ar1n02x5 _22508_ (.a(net638),
    .b(_12569_),
    .c(_12547_),
    .o1(_13730_));
 b15aoi022as1n04x5 _22509_ (.a(_13726_),
    .b(_13728_),
    .c(_13729_),
    .d(_13730_),
    .o1(_13731_));
 b15norp03ah1n03x5 _22510_ (.a(_12553_),
    .b(_12717_),
    .c(_13560_),
    .o1(_13732_));
 b15nanb02aq1n04x5 _22511_ (.a(net638),
    .b(net642),
    .out0(_13733_));
 b15nor004as1n04x5 _22512_ (.a(net631),
    .b(_12552_),
    .c(_12553_),
    .d(_13733_),
    .o1(_13734_));
 b15nanb02ar1n12x5 _22513_ (.a(\us03.a[7] ),
    .b(net627),
    .out0(_13735_));
 b15norp02an1n08x5 _22514_ (.a(_12751_),
    .b(_13735_),
    .o1(_13736_));
 b15oai022ar1n08x5 _22515_ (.a(_13599_),
    .b(_12669_),
    .c(_12689_),
    .d(_12692_),
    .o1(_13737_));
 b15aoi112an1n08x5 _22516_ (.a(_13732_),
    .b(_13734_),
    .c(_13736_),
    .d(_13737_),
    .o1(_13738_));
 b15nona22an1n02x5 _22517_ (.a(net637),
    .b(net636),
    .c(net629),
    .out0(_13739_));
 b15oaoi13aq1n08x5 _22518_ (.a(_13739_),
    .b(_12743_),
    .c(_12710_),
    .d(net626),
    .o1(_13740_));
 b15aoai13ah1n08x5 _22519_ (.a(net630),
    .b(_13740_),
    .c(_13650_),
    .d(_13683_),
    .o1(_13741_));
 b15nand04an1n12x5 _22520_ (.a(_13725_),
    .b(_13731_),
    .c(_13738_),
    .d(_13741_),
    .o1(_13742_));
 b15nand03al1n03x5 _22521_ (.a(_13712_),
    .b(_12720_),
    .c(_13565_),
    .o1(_13743_));
 b15nand04al1n02x5 _22522_ (.a(_12586_),
    .b(_12593_),
    .c(_13570_),
    .d(_12707_),
    .o1(_13744_));
 b15norp02ar1n04x5 _22523_ (.a(net627),
    .b(net621),
    .o1(_13745_));
 b15nano22al1n03x5 _22524_ (.a(net627),
    .b(net621),
    .c(net639),
    .out0(_13746_));
 b15oai112al1n12x5 _22525_ (.a(_12687_),
    .b(_12646_),
    .c(_13745_),
    .d(_13746_),
    .o1(_13747_));
 b15nandp3as1n04x5 _22526_ (.a(_13743_),
    .b(_13744_),
    .c(_13747_),
    .o1(_13748_));
 b15nonb03ar1n02x5 _22527_ (.a(net630),
    .b(net633),
    .c(net641),
    .out0(_13749_));
 b15aoai13ah1n02x5 _22528_ (.a(net637),
    .b(_13749_),
    .c(_12707_),
    .d(net641),
    .o1(_13750_));
 b15oaoi13al1n04x5 _22529_ (.a(_12714_),
    .b(_13750_),
    .c(_12649_),
    .d(_12591_),
    .o1(_13751_));
 b15nor002an1n03x5 _22530_ (.a(_12566_),
    .b(_12591_),
    .o1(_13752_));
 b15nanb02al1n08x5 _22531_ (.a(net633),
    .b(net632),
    .out0(_13753_));
 b15aoi112al1n02x5 _22532_ (.a(net641),
    .b(_13753_),
    .c(_12553_),
    .d(_12766_),
    .o1(_13754_));
 b15aoai13ar1n02x5 _22533_ (.a(net638),
    .b(_13752_),
    .c(_13754_),
    .d(_12587_),
    .o1(_13755_));
 b15nanb03ar1n02x5 _22534_ (.a(net624),
    .b(net621),
    .c(net633),
    .out0(_13756_));
 b15aoi112aq1n02x5 _22535_ (.a(net641),
    .b(_12547_),
    .c(_13756_),
    .d(_12569_),
    .o1(_13757_));
 b15nor002ar1n08x5 _22536_ (.a(_12689_),
    .b(_12771_),
    .o1(_13758_));
 b15oai112as1n06x5 _22537_ (.a(net637),
    .b(net630),
    .c(_13757_),
    .d(_13758_),
    .o1(_13759_));
 b15nona23aq1n05x5 _22538_ (.a(_13748_),
    .b(_13751_),
    .c(_13755_),
    .d(_13759_),
    .out0(_13760_));
 b15norp02as1n04x5 _22539_ (.a(net642),
    .b(_12762_),
    .o1(_13761_));
 b15qgbxo2an1n05x5 _22540_ (.a(\us03.a[4] ),
    .b(\us03.a[7] ),
    .out0(_13762_));
 b15oaoi13ah1n03x5 _22541_ (.a(net639),
    .b(_12760_),
    .c(_13762_),
    .d(_13654_),
    .o1(_13763_));
 b15oai012aq1n12x5 _22542_ (.a(_12707_),
    .b(_13761_),
    .c(_13763_),
    .o1(_13764_));
 b15nand04ah1n08x5 _22543_ (.a(_12657_),
    .b(_12649_),
    .c(_12610_),
    .d(_12641_),
    .o1(_13765_));
 b15nandp2ah1n03x5 _22544_ (.a(_13764_),
    .b(_13765_),
    .o1(_13766_));
 b15nor004as1n12x5 _22545_ (.a(_13615_),
    .b(_13742_),
    .c(_13760_),
    .d(_13766_),
    .o1(_13767_));
 b15nona23as1n32x5 _22546_ (.a(_13682_),
    .b(_13697_),
    .c(_13721_),
    .d(_13767_),
    .out0(_13768_));
 b15nandp2ah1n24x5 _22547_ (.a(_12822_),
    .b(_12798_),
    .o1(_13769_));
 b15nanb02as1n24x5 _22548_ (.a(net893),
    .b(net896),
    .out0(_13770_));
 b15nand02ah1n04x5 _22549_ (.a(net893),
    .b(net889),
    .o1(_13771_));
 b15oai022ar1n02x5 _22550_ (.a(net889),
    .b(_13770_),
    .c(_13771_),
    .d(net896),
    .o1(_13772_));
 b15norp02ar1n02x5 _22551_ (.a(net886),
    .b(net912),
    .o1(_13773_));
 b15aoi022ar1n02x5 _22552_ (.a(_12789_),
    .b(_12971_),
    .c(_13772_),
    .d(_13773_),
    .o1(_13774_));
 b15oai022ar1n04x5 _22553_ (.a(_12932_),
    .b(_13769_),
    .c(_13774_),
    .d(_12851_),
    .o1(_13775_));
 b15bfn001ah1n64x5 load_slew436 (.a(\u0.tmp_w[23] ),
    .o(net436));
 b15bfn001as1n48x5 load_slew435 (.a(\u0.tmp_w[23] ),
    .o(net435));
 b15bfn001as1n48x5 max_length434 (.a(net435),
    .o(net434));
 b15bfn001as1n48x5 max_length433 (.a(net435),
    .o(net433));
 b15norp02ar1n02x5 _22558_ (.a(net896),
    .b(_12931_),
    .o1(_13780_));
 b15norp02ar1n02x5 _22559_ (.a(net889),
    .b(net898),
    .o1(_13781_));
 b15aoai13ar1n02x5 _22560_ (.a(net893),
    .b(_13780_),
    .c(_13781_),
    .d(net896),
    .o1(_13782_));
 b15nand02ah1n04x5 _22561_ (.a(net898),
    .b(_12883_),
    .o1(_13783_));
 b15oaoi13an1n03x5 _22562_ (.a(_12867_),
    .b(_13782_),
    .c(_13783_),
    .d(net889),
    .o1(_13784_));
 b15oai012an1n06x5 _22563_ (.a(net906),
    .b(_13775_),
    .c(_13784_),
    .o1(_13785_));
 b15nor002an1n12x5 _22564_ (.a(net912),
    .b(net903),
    .o1(_13786_));
 b15inv000al1n05x5 _22565_ (.a(_13786_),
    .o1(_13787_));
 b15nandp3al1n02x5 _22566_ (.a(net905),
    .b(net897),
    .c(_12825_),
    .o1(_13788_));
 b15and003an1n02x5 _22567_ (.a(net910),
    .b(net905),
    .c(net901),
    .o(_13789_));
 b15oai013as1n03x5 _22568_ (.a(_13788_),
    .b(_13789_),
    .c(_12917_),
    .d(net897),
    .o1(_13790_));
 b15oai012ar1n04x5 _22569_ (.a(_12971_),
    .b(_12995_),
    .c(net905),
    .o1(_13791_));
 b15oai012aq1n02x5 _22570_ (.a(_12851_),
    .b(_12909_),
    .c(_12959_),
    .o1(_13792_));
 b15nandp2aq1n04x5 _22571_ (.a(net912),
    .b(_12959_),
    .o1(_13793_));
 b15norp02as1n48x5 _22572_ (.a(net907),
    .b(net903),
    .o1(_13794_));
 b15aoi012ar1n06x5 _22573_ (.a(_13792_),
    .b(_13793_),
    .c(_13794_),
    .o1(_13795_));
 b15aoi022ar1n08x5 _22574_ (.a(_13787_),
    .b(_13790_),
    .c(_13791_),
    .d(_13795_),
    .o1(_13796_));
 b15nonb02as1n16x5 _22575_ (.a(net905),
    .b(net901),
    .out0(_13797_));
 b15nano23as1n24x5 _22576_ (.a(net886),
    .b(net889),
    .c(net893),
    .d(net896),
    .out0(_13798_));
 b15nandp3ar1n02x5 _22577_ (.a(net910),
    .b(_12851_),
    .c(_13798_),
    .o1(_13799_));
 b15oai012aq1n02x5 _22578_ (.a(_13799_),
    .b(_12790_),
    .c(net910),
    .o1(_13800_));
 b15and002as1n24x5 _22579_ (.a(net913),
    .b(net908),
    .o(_13801_));
 b15bfn001as1n64x5 max_length432 (.a(\u0.tmp_w[24] ),
    .o(net432));
 b15nandp2al1n24x5 _22581_ (.a(_12796_),
    .b(_12848_),
    .o1(_13803_));
 b15aoai13ar1n02x5 _22582_ (.a(net901),
    .b(_12910_),
    .c(_13801_),
    .d(_13803_),
    .o1(_13804_));
 b15nand03ah1n16x5 _22583_ (.a(net901),
    .b(_12796_),
    .c(_12848_),
    .o1(_13805_));
 b15aoi012ar1n02x5 _22584_ (.a(_12851_),
    .b(_12917_),
    .c(_13805_),
    .o1(_13806_));
 b15aoi022aq1n04x5 _22585_ (.a(_13797_),
    .b(_13800_),
    .c(_13804_),
    .d(_13806_),
    .o1(_13807_));
 b15and003ar1n02x5 _22586_ (.a(_12851_),
    .b(_13798_),
    .c(_13786_),
    .o(_13808_));
 b15nano23as1n24x5 _22587_ (.a(net896),
    .b(net886),
    .c(\us10.a[6] ),
    .d(\us10.a[5] ),
    .out0(_13809_));
 b15bfn001as1n64x5 max_length431 (.a(\u0.tmp_w[24] ),
    .o(net431));
 b15aoi112as1n02x5 _22589_ (.a(net907),
    .b(_13808_),
    .c(_13809_),
    .d(net898),
    .o1(_13811_));
 b15nona23aq1n08x5 _22590_ (.a(net893),
    .b(net886),
    .c(net889),
    .d(net896),
    .out0(_13812_));
 b15qgbno2an1n10x5 _22591_ (.a(net898),
    .b(_13812_),
    .o1(_13813_));
 b15aoi022as1n02x5 _22592_ (.a(net898),
    .b(_12909_),
    .c(_12971_),
    .d(_13813_),
    .o1(_13814_));
 b15bfn001as1n48x5 load_slew430 (.a(net432),
    .o(net430));
 b15aoi012an1n08x5 _22594_ (.a(_13811_),
    .b(_13814_),
    .c(net907),
    .o1(_13816_));
 b15nano23as1n24x5 _22595_ (.a(net892),
    .b(net887),
    .c(net891),
    .d(net894),
    .out0(_13817_));
 b15nandp3as1n03x5 _22596_ (.a(_12968_),
    .b(_12904_),
    .c(_13817_),
    .o1(_13818_));
 b15oai112as1n16x5 _22597_ (.a(_12911_),
    .b(_13818_),
    .c(_12790_),
    .d(_12827_),
    .o1(_13819_));
 b15oai012aq1n08x5 _22598_ (.a(_13011_),
    .b(_13770_),
    .c(_13794_),
    .o1(_13820_));
 b15aoi012ar1n02x5 _22599_ (.a(net910),
    .b(net905),
    .c(net901),
    .o1(_13821_));
 b15orn003aq1n04x5 _22600_ (.a(_13794_),
    .b(_13789_),
    .c(_13821_),
    .o(_13822_));
 b15nand04ar1n06x5 _22601_ (.a(net897),
    .b(_12881_),
    .c(_13820_),
    .d(_13822_),
    .o1(_13823_));
 b15bfn001as1n48x5 max_length429 (.a(net432),
    .o(net429));
 b15bfn001as1n64x5 max_length428 (.a(\u0.tmp_w[25] ),
    .o(net428));
 b15and002ar1n04x5 _22604_ (.a(net910),
    .b(net899),
    .o(_13826_));
 b15norp02aq1n12x5 _22605_ (.a(net891),
    .b(net904),
    .o1(_13827_));
 b15xor002an1n12x5 _22606_ (.a(net908),
    .b(_13827_),
    .out0(_13828_));
 b15nand04aq1n12x5 _22607_ (.a(net886),
    .b(_12916_),
    .c(_13826_),
    .d(_13828_),
    .o1(_13829_));
 b15nanb03as1n06x5 _22608_ (.a(_13819_),
    .b(_13823_),
    .c(_13829_),
    .out0(_13830_));
 b15nano23aq1n16x5 _22609_ (.a(_13796_),
    .b(_13807_),
    .c(_13816_),
    .d(_13830_),
    .out0(_13831_));
 b15nonb03as1n04x5 _22610_ (.a(net909),
    .b(net904),
    .c(net891),
    .out0(_13832_));
 b15and002ah1n03x5 _22611_ (.a(net891),
    .b(net904),
    .o(_13833_));
 b15oai112an1n12x5 _22612_ (.a(net888),
    .b(_12916_),
    .c(_13832_),
    .d(_13833_),
    .o1(_13834_));
 b15nanb02as1n24x5 _22613_ (.a(net907),
    .b(net903),
    .out0(_13835_));
 b15oai112an1n04x5 _22614_ (.a(net898),
    .b(_13834_),
    .c(_13835_),
    .d(_13812_),
    .o1(_13836_));
 b15oai112an1n06x5 _22615_ (.a(_12950_),
    .b(_13836_),
    .c(_13013_),
    .d(net898),
    .o1(_13837_));
 b15nandp3as1n12x5 _22616_ (.o1(_13838_),
    .a(_12820_),
    .b(_12796_),
    .c(_12874_));
 b15aoai13ar1n04x5 _22617_ (.a(_12874_),
    .b(_12796_),
    .c(_12916_),
    .d(_12820_),
    .o1(_13839_));
 b15oaoi13aq1n04x5 _22618_ (.a(net912),
    .b(_13838_),
    .c(_13839_),
    .d(_12782_),
    .o1(_13840_));
 b15aoi013as1n03x5 _22619_ (.a(_13840_),
    .b(_12957_),
    .c(net903),
    .d(net912),
    .o1(_13841_));
 b15oai012an1n12x5 _22620_ (.a(_13837_),
    .b(_13841_),
    .c(net898),
    .o1(_13842_));
 b15orn002as1n16x5 _22621_ (.a(net910),
    .b(net908),
    .o(_13843_));
 b15nonb03ar1n06x5 _22622_ (.a(net890),
    .b(net904),
    .c(net887),
    .out0(_13844_));
 b15nand03al1n03x5 _22623_ (.a(_12796_),
    .b(_13843_),
    .c(_13844_),
    .o1(_13845_));
 b15nandp2as1n12x5 _22624_ (.a(net904),
    .b(_12991_),
    .o1(_13846_));
 b15aoai13an1n03x5 _22625_ (.a(net900),
    .b(_13801_),
    .c(_13845_),
    .d(_13846_),
    .o1(_13847_));
 b15and002aq1n02x5 _22626_ (.a(net892),
    .b(net890),
    .o(_13848_));
 b15nandp3ar1n02x5 _22627_ (.a(net894),
    .b(_13848_),
    .c(_13015_),
    .o1(_13849_));
 b15norp02ar1n08x5 _22628_ (.a(\us10.a[6] ),
    .b(net909),
    .o1(_13850_));
 b15nand02ar1n02x5 _22629_ (.a(_12916_),
    .b(_13850_),
    .o1(_13851_));
 b15aoi012ar1n02x5 _22630_ (.a(_12869_),
    .b(_13849_),
    .c(_13851_),
    .o1(_13852_));
 b15oai112aq1n02x5 _22631_ (.a(_12883_),
    .b(_12798_),
    .c(_12912_),
    .d(_13794_),
    .o1(_13853_));
 b15nonb02as1n04x5 _22632_ (.a(net888),
    .b(\us10.a[5] ),
    .out0(_13854_));
 b15xor002ar1n02x5 _22633_ (.a(net895),
    .b(net904),
    .out0(_13855_));
 b15aoi013an1n03x5 _22634_ (.a(_12991_),
    .b(_13854_),
    .c(_13855_),
    .d(net891),
    .o1(_13856_));
 b15oai112al1n06x5 _22635_ (.a(_12851_),
    .b(_13853_),
    .c(_13856_),
    .d(_12950_),
    .o1(_13857_));
 b15oai012as1n04x5 _22636_ (.a(_13847_),
    .b(_13852_),
    .c(_13857_),
    .o1(_13858_));
 b15qgbno2an1n10x5 _22637_ (.a(net887),
    .b(net904),
    .o1(_13859_));
 b15nonb02as1n16x5 _22638_ (.a(net904),
    .b(net909),
    .out0(_13860_));
 b15bfn001as1n64x5 max_length427 (.a(\u0.tmp_w[25] ),
    .o(net427));
 b15aoi012ar1n02x5 _22640_ (.a(_13859_),
    .b(_13860_),
    .c(net887),
    .o1(_13862_));
 b15nor003ah1n03x5 _22641_ (.a(_12865_),
    .b(_12938_),
    .c(_13862_),
    .o1(_13863_));
 b15bfn001as1n64x5 max_length426 (.a(net428),
    .o(net426));
 b15aoi013ar1n02x5 _22643_ (.a(_12851_),
    .b(_12796_),
    .c(_13794_),
    .d(_12798_),
    .o1(_13865_));
 b15nand03ar1n08x5 _22644_ (.a(_12796_),
    .b(_12874_),
    .c(_12877_),
    .o1(_13866_));
 b15oai012ar1n04x5 _22645_ (.a(_13865_),
    .b(_13866_),
    .c(_12820_),
    .o1(_13867_));
 b15aoi012aq1n02x5 _22646_ (.a(net900),
    .b(_13809_),
    .c(_13860_),
    .o1(_13868_));
 b15nano22ar1n02x5 _22647_ (.a(\us10.a[5] ),
    .b(net891),
    .c(net888),
    .out0(_13869_));
 b15aoi022ah1n02x5 _22648_ (.a(_13832_),
    .b(_13854_),
    .c(_13869_),
    .d(_13860_),
    .o1(_13870_));
 b15nandp2as1n12x5 _22649_ (.a(net894),
    .b(_12950_),
    .o1(_13871_));
 b15nandp2as1n04x5 _22650_ (.a(net888),
    .b(net909),
    .o1(_13872_));
 b15aoi022an1n04x5 _22651_ (.a(_12822_),
    .b(_13827_),
    .c(_13833_),
    .d(_12883_),
    .o1(_13873_));
 b15oai122ar1n12x5 _22652_ (.a(_13868_),
    .b(_13870_),
    .c(_13871_),
    .d(_13872_),
    .e(_13873_),
    .o1(_13874_));
 b15nano23ar1n02x5 _22653_ (.a(net894),
    .b(\us10.a[6] ),
    .c(net904),
    .d(net888),
    .out0(_13875_));
 b15aoai13ar1n02x5 _22654_ (.a(net892),
    .b(_13875_),
    .c(_13850_),
    .d(_12940_),
    .o1(_13876_));
 b15nanb02ar1n02x5 _22655_ (.a(_12929_),
    .b(_13833_),
    .out0(_13877_));
 b15aoi012ar1n02x5 _22656_ (.a(_12950_),
    .b(_13876_),
    .c(_13877_),
    .o1(_13878_));
 b15oai022ah1n04x5 _22657_ (.a(_13863_),
    .b(_13867_),
    .c(_13874_),
    .d(_13878_),
    .o1(_13879_));
 b15nor003al1n03x5 _22658_ (.a(net899),
    .b(_13812_),
    .c(_13843_),
    .o1(_13880_));
 b15oai012ar1n04x5 _22659_ (.a(_12820_),
    .b(_12875_),
    .c(_12900_),
    .o1(_13881_));
 b15inv000al1n10x5 _22660_ (.a(net893),
    .o1(_13882_));
 b15and002ar1n24x5 _22661_ (.a(net894),
    .b(net887),
    .o(_13883_));
 b15norp02al1n32x5 _22662_ (.a(net895),
    .b(net888),
    .o1(_13884_));
 b15oai112al1n08x5 _22663_ (.a(_13882_),
    .b(net899),
    .c(_13883_),
    .d(_13884_),
    .o1(_13885_));
 b15nandp2ar1n03x5 _22664_ (.a(_12822_),
    .b(_12987_),
    .o1(_13886_));
 b15oaoi13aq1n04x5 _22665_ (.a(net889),
    .b(_13885_),
    .c(_13886_),
    .d(net886),
    .o1(_13887_));
 b15oai013ah1n03x5 _22666_ (.a(net902),
    .b(net899),
    .c(_12904_),
    .d(_13007_),
    .o1(_13888_));
 b15oai022aq1n08x5 _22667_ (.a(_13880_),
    .b(_13881_),
    .c(_13887_),
    .d(_13888_),
    .o1(_13889_));
 b15nandp3aq1n12x5 _22668_ (.o1(_13890_),
    .a(_13858_),
    .b(_13879_),
    .c(_13889_));
 b15nano23as1n24x5 _22669_ (.a(_13785_),
    .b(_13831_),
    .c(_13842_),
    .d(_13890_),
    .out0(_13891_));
 b15xor002as1n12x5 _22670_ (.a(_13768_),
    .b(_13891_),
    .out0(_13892_));
 b15xor002al1n12x5 _22671_ (.a(_13664_),
    .b(_13892_),
    .out0(_13893_));
 b15norp02ar1n03x5 _22672_ (.a(_13390_),
    .b(_13499_),
    .o1(_13894_));
 b15bfn001as1n48x5 max_length425 (.a(net427),
    .o(net425));
 b15nandp2an1n08x5 _22674_ (.a(net661),
    .b(_13486_),
    .o1(_13896_));
 b15nonb03al1n12x5 _22675_ (.a(net644),
    .b(net647),
    .c(net654),
    .out0(_13897_));
 b15aoai13ar1n08x5 _22676_ (.a(_13478_),
    .b(_13897_),
    .c(_13522_),
    .d(net661),
    .o1(_13898_));
 b15aoi012ar1n02x5 _22677_ (.a(_13355_),
    .b(_13896_),
    .c(_13898_),
    .o1(_13899_));
 b15oab012ar1n02x5 _22678_ (.a(net665),
    .b(_13894_),
    .c(_13899_),
    .out0(_13900_));
 b15nor003as1n06x5 _22679_ (.a(_13318_),
    .b(_13441_),
    .c(_13450_),
    .o1(_13901_));
 b15orn003ah1n02x5 _22680_ (.a(net657),
    .b(net653),
    .c(net648),
    .o(_13902_));
 b15nand04as1n06x5 _22681_ (.a(net667),
    .b(net657),
    .c(net653),
    .d(net648),
    .o1(_13903_));
 b15aoi112ar1n08x5 _22682_ (.a(_13530_),
    .b(_13533_),
    .c(_13902_),
    .d(_13903_),
    .o1(_13904_));
 b15nonb03as1n12x5 _22683_ (.a(net656),
    .b(net660),
    .c(net664),
    .out0(_13905_));
 b15aoi112ar1n06x5 _22684_ (.a(_13901_),
    .b(_13904_),
    .c(_13905_),
    .d(_13412_),
    .o1(_13906_));
 b15norp02as1n02x5 _22685_ (.a(_13423_),
    .b(_13494_),
    .o1(_13907_));
 b15aoai13al1n08x5 _22686_ (.a(_13362_),
    .b(_13907_),
    .c(_13423_),
    .d(_13320_),
    .o1(_13908_));
 b15bfn001ah1n64x5 max_length424 (.a(\u0.tmp_w[26] ),
    .o(net424));
 b15nona23al1n05x5 _22688_ (.a(net649),
    .b(net643),
    .c(net652),
    .d(net666),
    .out0(_13910_));
 b15oaoi13aq1n08x5 _22689_ (.a(_13340_),
    .b(_13910_),
    .c(_13343_),
    .d(_13306_),
    .o1(_13911_));
 b15nor002ah1n02x5 _22690_ (.a(_13355_),
    .b(_13500_),
    .o1(_13912_));
 b15oai022ar1n02x5 _22691_ (.a(_13306_),
    .b(_13343_),
    .c(_13398_),
    .d(_13479_),
    .o1(_13913_));
 b15aoi112ar1n02x5 _22692_ (.a(_13911_),
    .b(_13912_),
    .c(_13355_),
    .d(_13913_),
    .o1(_13914_));
 b15oai112as1n04x5 _22693_ (.a(_13906_),
    .b(_13908_),
    .c(_13345_),
    .d(_13914_),
    .o1(_13915_));
 b15norp02ar1n48x5 _22694_ (.a(_13340_),
    .b(net658),
    .o1(_13916_));
 b15nonb02ar1n16x5 _22695_ (.a(net648),
    .b(\us32.a[4] ),
    .out0(_13917_));
 b15nand03ar1n04x5 _22696_ (.a(_13407_),
    .b(_13916_),
    .c(_13917_),
    .o1(_13918_));
 b15nor003al1n02x5 _22697_ (.a(_13318_),
    .b(_13441_),
    .c(_13447_),
    .o1(_13919_));
 b15nonb02ah1n12x5 _22698_ (.a(net662),
    .b(net650),
    .out0(_13920_));
 b15aoi013aq1n02x5 _22699_ (.a(_13919_),
    .b(_13897_),
    .c(_13920_),
    .d(net656),
    .o1(_13921_));
 b15nand02an1n02x5 _22700_ (.a(_13438_),
    .b(_13410_),
    .o1(_13922_));
 b15aoi013aq1n04x5 _22701_ (.a(_13355_),
    .b(_13918_),
    .c(_13921_),
    .d(_13922_),
    .o1(_13923_));
 b15nor002al1n16x5 _22702_ (.a(_13324_),
    .b(_13302_),
    .o1(_13924_));
 b15nor002aq1n03x5 _22703_ (.a(_13313_),
    .b(_13418_),
    .o1(_13925_));
 b15aoi022ah1n04x5 _22704_ (.a(_13924_),
    .b(_13916_),
    .c(_13925_),
    .d(_13361_),
    .o1(_13926_));
 b15nand03as1n06x5 _22705_ (.a(net655),
    .b(_13402_),
    .c(_13385_),
    .o1(_13927_));
 b15andc04as1n16x5 _22706_ (.a(net650),
    .b(net654),
    .c(net643),
    .d(net647),
    .o(_13928_));
 b15nand02ar1n02x5 _22707_ (.a(_13313_),
    .b(_13928_),
    .o1(_13929_));
 b15aob012ar1n02x5 _22708_ (.a(net664),
    .b(_13927_),
    .c(_13929_),
    .out0(_13930_));
 b15aoi012al1n02x5 _22709_ (.a(net659),
    .b(_13926_),
    .c(_13930_),
    .o1(_13931_));
 b15ornc04aq1n03x5 _22710_ (.a(_13900_),
    .b(_13915_),
    .c(_13923_),
    .d(_13931_),
    .o(_13932_));
 b15bfn001as1n64x5 max_length423 (.a(\u0.tmp_w[26] ),
    .o(net423));
 b15nonb03as1n12x5 _22712_ (.a(net647),
    .b(net645),
    .c(net653),
    .out0(_13934_));
 b15aoi022ar1n02x5 _22713_ (.a(_13505_),
    .b(_13418_),
    .c(_13934_),
    .d(_13417_),
    .o1(_13935_));
 b15orn003ar1n02x5 _22714_ (.a(net651),
    .b(_13447_),
    .c(_13935_),
    .o(_13936_));
 b15norp03al1n02x5 _22715_ (.a(_13479_),
    .b(_13392_),
    .c(_13399_),
    .o1(_13937_));
 b15nano23as1n24x5 _22716_ (.a(net645),
    .b(net648),
    .c(net651),
    .d(\us32.a[4] ),
    .out0(_13938_));
 b15nor002al1n24x5 _22717_ (.a(net665),
    .b(net667),
    .o1(_13939_));
 b15aoi013an1n02x5 _22718_ (.a(_13937_),
    .b(_13938_),
    .c(_13939_),
    .d(_13410_),
    .o1(_13940_));
 b15nanb02aq1n08x5 _22719_ (.a(net660),
    .b(net663),
    .out0(_13941_));
 b15ornc04al1n12x5 _22720_ (.a(net649),
    .b(net652),
    .c(net643),
    .d(net646),
    .o(_13942_));
 b15nor002ah1n04x5 _22721_ (.a(_13941_),
    .b(_13942_),
    .o1(_13943_));
 b15norp02aq1n04x5 _22722_ (.a(_13315_),
    .b(_13350_),
    .o1(_13944_));
 b15nonb02as1n16x5 _22723_ (.a(net662),
    .b(net656),
    .out0(_13945_));
 b15aoi013ah1n06x5 _22724_ (.a(_13943_),
    .b(_13944_),
    .c(_13945_),
    .d(_13425_),
    .o1(_13946_));
 b15nand03as1n04x5 _22725_ (.a(_13936_),
    .b(_13940_),
    .c(_13946_),
    .o1(_13947_));
 b15bfn001as1n64x5 max_length422 (.a(\u0.tmp_w[26] ),
    .o(net422));
 b15orn002aq1n12x5 _22727_ (.a(net667),
    .b(net661),
    .o(_13949_));
 b15and002ah1n08x5 _22728_ (.a(net665),
    .b(net667),
    .o(_13950_));
 b15nand02an1n02x5 _22729_ (.a(net659),
    .b(_13950_),
    .o1(_13951_));
 b15nand04an1n02x5 _22730_ (.a(net657),
    .b(_13949_),
    .c(_13934_),
    .d(_13951_),
    .o1(_13952_));
 b15nandp3aq1n08x5 _22731_ (.a(net663),
    .b(net657),
    .c(net659),
    .o1(_13953_));
 b15aoi112al1n02x5 _22732_ (.a(_13431_),
    .b(_13953_),
    .c(net666),
    .d(net646),
    .o1(_13954_));
 b15norp03ah1n24x5 _22733_ (.a(net654),
    .b(net643),
    .c(net647),
    .o1(_13955_));
 b15aoi013ah1n03x5 _22734_ (.a(_13954_),
    .b(_13955_),
    .c(_13410_),
    .d(_13418_),
    .o1(_13956_));
 b15aoi012ar1n02x5 _22735_ (.a(net651),
    .b(_13952_),
    .c(_13956_),
    .o1(_13957_));
 b15nonb02as1n06x5 _22736_ (.a(net656),
    .b(net660),
    .out0(_13958_));
 b15bfn001ah1n64x5 max_length421 (.a(net422),
    .o(net421));
 b15nand02aq1n16x5 _22738_ (.a(net663),
    .b(net655),
    .o1(_13960_));
 b15oaoi13an1n03x5 _22739_ (.a(net666),
    .b(_13960_),
    .c(_13347_),
    .d(net663),
    .o1(_13961_));
 b15oai012an1n08x5 _22740_ (.a(_13928_),
    .b(_13958_),
    .c(_13961_),
    .o1(_13962_));
 b15aoi012ar1n06x5 _22741_ (.a(_13534_),
    .b(_13536_),
    .c(_13355_),
    .o1(_13963_));
 b15nor004al1n12x5 _22742_ (.a(_13418_),
    .b(_13447_),
    .c(_13533_),
    .d(_13963_),
    .o1(_13964_));
 b15nonb02as1n16x5 _22743_ (.a(net660),
    .b(net663),
    .out0(_13965_));
 b15nand04al1n03x5 _22744_ (.a(_13355_),
    .b(_13505_),
    .c(_13506_),
    .d(_13965_),
    .o1(_13966_));
 b15orn002aq1n12x5 _22745_ (.a(net660),
    .b(net649),
    .o(_13967_));
 b15inv020ar1n08x5 _22746_ (.a(_13435_),
    .o1(_13968_));
 b15oai013al1n04x5 _22747_ (.a(_13966_),
    .b(_13967_),
    .c(_13968_),
    .d(_13355_),
    .o1(_13969_));
 b15bfn001ah1n64x5 wire420 (.a(\u0.tmp_w[27] ),
    .o(net420));
 b15bfn001as1n64x5 max_length419 (.a(net420),
    .o(net419));
 b15aoi012aq1n02x5 _22750_ (.a(_13964_),
    .b(_13969_),
    .c(net657),
    .o1(_13972_));
 b15nona23an1n04x5 _22751_ (.a(_13947_),
    .b(_13957_),
    .c(_13962_),
    .d(_13972_),
    .out0(_13973_));
 b15oai012ar1n02x5 _22752_ (.a(_13402_),
    .b(net653),
    .c(net651),
    .o1(_13974_));
 b15oaoi13ar1n02x5 _22753_ (.a(net665),
    .b(net667),
    .c(_13374_),
    .d(_13924_),
    .o1(_13975_));
 b15nor004an1n02x5 _22754_ (.a(_13347_),
    .b(_13950_),
    .c(_13974_),
    .d(_13975_),
    .o1(_13976_));
 b15xor002as1n16x5 _22755_ (.a(net668),
    .b(net662),
    .out0(_13977_));
 b15nand03ar1n02x5 _22756_ (.a(_13380_),
    .b(_13442_),
    .c(_13977_),
    .o1(_13978_));
 b15norp02al1n03x5 _22757_ (.a(_13315_),
    .b(_13306_),
    .o1(_13979_));
 b15norp02al1n08x5 _22758_ (.a(_13350_),
    .b(_13441_),
    .o1(_13980_));
 b15oai112al1n06x5 _22759_ (.a(_13945_),
    .b(_13939_),
    .c(_13979_),
    .d(_13980_),
    .o1(_13981_));
 b15norp02an1n03x5 _22760_ (.a(_13514_),
    .b(_13447_),
    .o1(_13982_));
 b15nand02ar1n02x5 _22761_ (.a(_13467_),
    .b(_13982_),
    .o1(_13983_));
 b15nandp3aq1n02x5 _22762_ (.a(_13978_),
    .b(_13981_),
    .c(_13983_),
    .o1(_13984_));
 b15xnr002ah1n16x5 _22763_ (.a(net650),
    .b(\us32.a[7] ),
    .out0(_13985_));
 b15norp03ar1n02x5 _22764_ (.a(net648),
    .b(_13953_),
    .c(_13985_),
    .o1(_13986_));
 b15bfn001as1n64x5 max_length418 (.a(net419),
    .o(net418));
 b15aoi013ar1n02x5 _22766_ (.a(_13986_),
    .b(_13985_),
    .c(_13982_),
    .d(net648),
    .o1(_13988_));
 b15orn002ar1n02x5 _22767_ (.a(net653),
    .b(_13988_),
    .o(_13989_));
 b15norp02aq1n03x5 _22768_ (.a(net657),
    .b(_13330_),
    .o1(_13990_));
 b15bfn001ah1n48x5 max_length417 (.a(net420),
    .o(net417));
 b15aoai13ar1n04x5 _22770_ (.a(net667),
    .b(_13894_),
    .c(_13990_),
    .d(_13421_),
    .o1(_13992_));
 b15nona23ar1n05x5 _22771_ (.a(_13976_),
    .b(_13984_),
    .c(_13989_),
    .d(_13992_),
    .out0(_13993_));
 b15norp02ar1n02x5 _22772_ (.a(_13340_),
    .b(_13500_),
    .o1(_13994_));
 b15aoai13ar1n02x5 _22773_ (.a(_13945_),
    .b(_13994_),
    .c(_13340_),
    .d(_13438_),
    .o1(_13995_));
 b15norp02al1n32x5 _22774_ (.a(_13324_),
    .b(_13343_),
    .o1(_13996_));
 b15aoai13ah1n03x5 _22775_ (.a(_13371_),
    .b(_13990_),
    .c(_13355_),
    .d(_13996_),
    .o1(_13997_));
 b15aoi012al1n06x5 _22776_ (.a(net656),
    .b(_13977_),
    .c(net664),
    .o1(_13998_));
 b15norp03an1n24x5 _22777_ (.a(net646),
    .b(_13431_),
    .c(_13399_),
    .o1(_13999_));
 b15nor002ar1n24x5 _22778_ (.a(_13302_),
    .b(_13306_),
    .o1(_14000_));
 b15aoai13ah1n02x5 _22779_ (.a(_13998_),
    .b(_13999_),
    .c(_13421_),
    .d(_14000_),
    .o1(_14001_));
 b15nor002aq1n06x5 _22780_ (.a(net655),
    .b(_13494_),
    .o1(_14002_));
 b15nonb03ar1n08x5 _22781_ (.a(net666),
    .b(net649),
    .c(net664),
    .out0(_14003_));
 b15and003ar1n02x5 _22782_ (.a(net655),
    .b(_13375_),
    .c(_14003_),
    .o(_14004_));
 b15oai012ah1n03x5 _22783_ (.a(net660),
    .b(_14002_),
    .c(_14004_),
    .o1(_14005_));
 b15nand04al1n03x5 _22784_ (.a(_13995_),
    .b(_13997_),
    .c(_14001_),
    .d(_14005_),
    .o1(_14006_));
 b15aoi022aq1n02x5 _22785_ (.a(_13945_),
    .b(_13397_),
    .c(_13955_),
    .d(_13958_),
    .o1(_14007_));
 b15nanb02an1n02x5 _22786_ (.a(_14007_),
    .b(_14003_),
    .out0(_14008_));
 b15oai012as1n02x5 _22787_ (.a(_13448_),
    .b(_13928_),
    .c(_13415_),
    .o1(_14009_));
 b15nor002al1n02x5 _22788_ (.a(_13368_),
    .b(_13528_),
    .o1(_14010_));
 b15oai112as1n06x5 _22789_ (.a(_14008_),
    .b(_14009_),
    .c(_14010_),
    .d(_13927_),
    .o1(_14011_));
 b15nanb02al1n08x5 _22790_ (.a(net651),
    .b(net645),
    .out0(_14012_));
 b15oai022ar1n02x5 _22791_ (.a(_13447_),
    .b(_14012_),
    .c(_13985_),
    .d(_13499_),
    .o1(_14013_));
 b15nandp3ar1n02x5 _22792_ (.a(_13418_),
    .b(_13917_),
    .c(_14013_),
    .o1(_14014_));
 b15bfn001as1n64x5 max_length416 (.a(\u0.tmp_w[28] ),
    .o(net416));
 b15oai022ar1n02x5 _22794_ (.a(net659),
    .b(_13509_),
    .c(_13951_),
    .d(_13330_),
    .o1(_14016_));
 b15aob012an1n02x5 _22795_ (.a(_14014_),
    .b(_14016_),
    .c(net657),
    .out0(_14017_));
 b15orn003as1n02x5 _22796_ (.a(_14006_),
    .b(_14011_),
    .c(_14017_),
    .o(_14018_));
 b15nor004an1n08x5 _22797_ (.a(_13932_),
    .b(_13973_),
    .c(_13993_),
    .d(_14018_),
    .o1(_14019_));
 b15nonb02al1n12x5 _22798_ (.a(net788),
    .b(net796),
    .out0(_14020_));
 b15aoi012ar1n02x5 _22799_ (.a(_13022_),
    .b(_13147_),
    .c(_14020_),
    .o1(_14021_));
 b15nandp2ar1n05x5 _22800_ (.a(net788),
    .b(_13147_),
    .o1(_14022_));
 b15nandp2ah1n05x5 _22801_ (.a(_13114_),
    .b(_13171_),
    .o1(_14023_));
 b15aoai13as1n02x5 _22802_ (.a(_14021_),
    .b(net791),
    .c(_14022_),
    .d(_14023_),
    .o1(_14024_));
 b15nanb02as1n24x5 _22803_ (.a(net769),
    .b(net773),
    .out0(_14025_));
 b15nor004ah1n04x5 _22804_ (.a(net795),
    .b(_13063_),
    .c(_13194_),
    .d(_14025_),
    .o1(_14026_));
 b15oaoi13al1n04x5 _22805_ (.a(_13194_),
    .b(_13045_),
    .c(net793),
    .d(_14025_),
    .o1(_14027_));
 b15aoai13as1n08x5 _22806_ (.a(_13114_),
    .b(_14026_),
    .c(_14027_),
    .d(net795),
    .o1(_14028_));
 b15nanb02as1n24x5 _22807_ (.a(net789),
    .b(net792),
    .out0(_14029_));
 b15nano23as1n24x5 _22808_ (.a(net779),
    .b(net770),
    .c(net772),
    .d(net776),
    .out0(_14030_));
 b15aoai13ar1n03x5 _22809_ (.a(_14029_),
    .b(_14030_),
    .c(net791),
    .d(_13181_),
    .o1(_14031_));
 b15aoi022ar1n02x5 _22810_ (.a(_13114_),
    .b(_13171_),
    .c(_13181_),
    .d(net791),
    .o1(_14032_));
 b15oai112al1n06x5 _22811_ (.a(_14028_),
    .b(_14031_),
    .c(_14032_),
    .d(_13067_),
    .o1(_14033_));
 b15nandp2ah1n24x5 _22812_ (.a(_13176_),
    .b(_13208_),
    .o1(_14034_));
 b15nonb02as1n16x5 _22813_ (.a(net790),
    .b(net785),
    .out0(_14035_));
 b15nandp2ah1n04x5 _22814_ (.a(net796),
    .b(_14035_),
    .o1(_14036_));
 b15oai022ah1n02x5 _22815_ (.a(net796),
    .b(_14034_),
    .c(_14036_),
    .d(_13142_),
    .o1(_14037_));
 b15oai022as1n06x5 _22816_ (.a(_14024_),
    .b(_14033_),
    .c(_14037_),
    .d(net782),
    .o1(_14038_));
 b15aoi022ar1n04x5 _22817_ (.a(_13128_),
    .b(_13129_),
    .c(_13213_),
    .d(_13063_),
    .o1(_14039_));
 b15oai112aq1n08x5 _22818_ (.a(_13022_),
    .b(_13272_),
    .c(_14039_),
    .d(net788),
    .o1(_14040_));
 b15bfn001as1n64x5 max_length415 (.a(net416),
    .o(net415));
 b15nand03an1n03x5 _22820_ (.a(_13066_),
    .b(net789),
    .c(_13092_),
    .o1(_14042_));
 b15oai012al1n08x5 _22821_ (.a(_13231_),
    .b(_13196_),
    .c(_13057_),
    .o1(_14043_));
 b15aoi012aq1n06x5 _22822_ (.a(net775),
    .b(_14042_),
    .c(_14043_),
    .o1(_14044_));
 b15oai112ah1n16x5 _22823_ (.a(_13067_),
    .b(_14040_),
    .c(_14044_),
    .d(_13022_),
    .o1(_14045_));
 b15oai012an1n02x5 _22824_ (.a(net788),
    .b(_13252_),
    .c(_13227_),
    .o1(_14046_));
 b15bfn001as1n48x5 max_length414 (.a(net416),
    .o(net414));
 b15nonb02aq1n02x5 _22826_ (.a(net792),
    .b(net770),
    .out0(_14048_));
 b15norp02ar1n02x5 _22827_ (.a(net772),
    .b(net784),
    .o1(_14049_));
 b15oai112al1n02x5 _22828_ (.a(_13208_),
    .b(_14048_),
    .c(_14049_),
    .d(_13203_),
    .o1(_14050_));
 b15nor003al1n08x5 _22829_ (.a(net796),
    .b(net788),
    .c(net784),
    .o1(_14051_));
 b15oai012an1n02x5 _22830_ (.a(_14050_),
    .b(_14051_),
    .c(_13227_),
    .o1(_14052_));
 b15nandp2al1n12x5 _22831_ (.a(net782),
    .b(_13050_),
    .o1(_14053_));
 b15oai112aq1n08x5 _22832_ (.a(_14046_),
    .b(_14052_),
    .c(net796),
    .d(_14053_),
    .o1(_14054_));
 b15nonb02as1n03x5 _22833_ (.a(net796),
    .b(net779),
    .out0(_14055_));
 b15nand02al1n02x5 _22834_ (.a(_13092_),
    .b(_14055_),
    .o1(_14056_));
 b15bfn001as1n64x5 max_length413 (.a(\u0.tmp_w[29] ),
    .o(net413));
 b15nonb03as1n12x5 _22836_ (.a(net779),
    .b(net770),
    .c(net772),
    .out0(_14058_));
 b15nand02ar1n02x5 _22837_ (.a(_13067_),
    .b(_14058_),
    .o1(_14059_));
 b15aoi112an1n03x5 _22838_ (.a(net776),
    .b(net784),
    .c(_14056_),
    .d(_14059_),
    .o1(_14060_));
 b15norp02aq1n04x5 _22839_ (.a(net791),
    .b(_13255_),
    .o1(_14061_));
 b15bfn001ah1n64x5 wire412 (.a(net413),
    .o(net412));
 b15nandp2aq1n16x5 _22841_ (.a(net790),
    .b(net780),
    .o1(_14063_));
 b15nor003al1n02x5 _22842_ (.a(net796),
    .b(_13086_),
    .c(_14063_),
    .o1(_14064_));
 b15oai013as1n04x5 _22843_ (.a(net788),
    .b(_14060_),
    .c(_14061_),
    .d(_14064_),
    .o1(_14065_));
 b15nand03ah1n08x5 _22844_ (.a(net782),
    .b(_13092_),
    .c(_13091_),
    .o1(_14066_));
 b15nanb02as1n24x5 _22845_ (.a(net792),
    .b(net789),
    .out0(_14067_));
 b15aoi012al1n02x5 _22846_ (.a(_14066_),
    .b(_14067_),
    .c(_14029_),
    .o1(_14068_));
 b15bfn001ah1n64x5 max_length411 (.a(net413),
    .o(net411));
 b15aoi013an1n06x5 _22848_ (.a(_14068_),
    .b(_13124_),
    .c(_14030_),
    .d(net791),
    .o1(_14070_));
 b15oai112as1n16x5 _22849_ (.a(_14054_),
    .b(_14065_),
    .c(_14070_),
    .d(net796),
    .o1(_14071_));
 b15nand03ah1n02x5 _22850_ (.a(_13114_),
    .b(net782),
    .c(_13213_),
    .o1(_14072_));
 b15nandp2an1n04x5 _22851_ (.a(net796),
    .b(_13171_),
    .o1(_14073_));
 b15oaoi13as1n08x5 _22852_ (.a(net792),
    .b(_14072_),
    .c(_14073_),
    .d(net782),
    .o1(_14074_));
 b15and002al1n12x5 _22853_ (.a(net775),
    .b(net771),
    .o(_14075_));
 b15nonb03an1n04x5 _22854_ (.a(net778),
    .b(net768),
    .c(net790),
    .out0(_14076_));
 b15nano22ah1n05x5 _22855_ (.a(net768),
    .b(net790),
    .c(net778),
    .out0(_14077_));
 b15oai112aq1n16x5 _22856_ (.a(_13239_),
    .b(_14075_),
    .c(_14076_),
    .d(_14077_),
    .o1(_14078_));
 b15xor002ar1n02x5 _22857_ (.a(net794),
    .b(net785),
    .out0(_14079_));
 b15nona23an1n04x5 _22858_ (.a(_14079_),
    .b(_14063_),
    .c(_13128_),
    .d(_13184_),
    .out0(_14080_));
 b15nandp3ah1n04x5 _22859_ (.a(net790),
    .b(_13124_),
    .c(_13171_),
    .o1(_14081_));
 b15nano22an1n02x5 _22860_ (.a(net774),
    .b(net777),
    .c(net783),
    .out0(_14082_));
 b15oai112as1n06x5 _22861_ (.a(_14035_),
    .b(_13176_),
    .c(_14082_),
    .d(_13184_),
    .o1(_14083_));
 b15nand04al1n12x5 _22862_ (.a(_14078_),
    .b(_14080_),
    .c(_14081_),
    .d(_14083_),
    .o1(_14084_));
 b15nanb02as1n24x5 _22863_ (.a(net787),
    .b(net780),
    .out0(_14085_));
 b15orn002ar1n02x5 _22864_ (.a(net774),
    .b(net793),
    .o(_14086_));
 b15oai112aq1n02x5 _22865_ (.a(_14086_),
    .b(_14058_),
    .c(_13174_),
    .d(_13040_),
    .o1(_14087_));
 b15oaoi13aq1n04x5 _22866_ (.a(_14085_),
    .b(_14087_),
    .c(_13277_),
    .d(_13185_),
    .o1(_14088_));
 b15norp02al1n08x5 _22867_ (.a(net791),
    .b(net786),
    .o1(_14089_));
 b15aoi012ar1n06x5 _22868_ (.a(net794),
    .b(net793),
    .c(net786),
    .o1(_14090_));
 b15oai112ar1n04x5 _22869_ (.a(_13092_),
    .b(_13208_),
    .c(_14089_),
    .d(_14090_),
    .o1(_14091_));
 b15orn003ar1n02x5 _22870_ (.a(_13052_),
    .b(_13078_),
    .c(_13224_),
    .o(_14092_));
 b15aoi012aq1n02x5 _22871_ (.a(_13022_),
    .b(_14091_),
    .c(_14092_),
    .o1(_14093_));
 b15nor004aq1n06x5 _22872_ (.a(_14074_),
    .b(_14084_),
    .c(_14088_),
    .d(_14093_),
    .o1(_14094_));
 b15nanb02aq1n12x5 _22873_ (.a(net781),
    .b(net791),
    .out0(_14095_));
 b15nor003al1n08x5 _22874_ (.a(_13052_),
    .b(_13078_),
    .c(_14095_),
    .o1(_14096_));
 b15oai012ah1n02x5 _22875_ (.a(net785),
    .b(_13162_),
    .c(_14096_),
    .o1(_14097_));
 b15norp02as1n08x5 _22876_ (.a(_13141_),
    .b(_14067_),
    .o1(_14098_));
 b15nor002ah1n04x5 _22877_ (.a(_13052_),
    .b(_13078_),
    .o1(_14099_));
 b15aoai13al1n02x5 _22878_ (.a(_13022_),
    .b(_14098_),
    .c(_14099_),
    .d(net795),
    .o1(_14100_));
 b15nand03an1n06x5 _22879_ (.a(net777),
    .b(net785),
    .c(net783),
    .o1(_14101_));
 b15oai012ar1n02x5 _22880_ (.a(_14101_),
    .b(_13140_),
    .c(net777),
    .o1(_14102_));
 b15orn002ah1n12x5 _22881_ (.a(net794),
    .b(net790),
    .o(_14103_));
 b15nonb02aq1n06x5 _22882_ (.a(net775),
    .b(net768),
    .out0(_14104_));
 b15and003ar1n02x5 _22883_ (.a(net773),
    .b(_14103_),
    .c(_14104_),
    .o(_14105_));
 b15ao0022an1n04x5 _22884_ (.a(_13090_),
    .b(_13239_),
    .c(_14102_),
    .d(_14105_),
    .o(_14106_));
 b15and002ah1n16x5 _22885_ (.a(net775),
    .b(net768),
    .o(_14107_));
 b15oai112ah1n06x5 _22886_ (.a(_13291_),
    .b(_14107_),
    .c(_13217_),
    .d(_13072_),
    .o1(_14108_));
 b15nand04aq1n04x5 _22887_ (.a(_13174_),
    .b(_13040_),
    .c(_13222_),
    .d(_13277_),
    .o1(_14109_));
 b15aoi012al1n06x5 _22888_ (.a(_14101_),
    .b(_14108_),
    .c(_14109_),
    .o1(_14110_));
 b15nano23al1n06x5 _22889_ (.a(_14097_),
    .b(_14100_),
    .c(_14106_),
    .d(_14110_),
    .out0(_14111_));
 b15aoi022ar1n02x5 _22890_ (.a(net795),
    .b(_13147_),
    .c(_13050_),
    .d(_13249_),
    .o1(_14112_));
 b15aob012al1n06x5 _22891_ (.a(_13022_),
    .b(_13047_),
    .c(_14112_),
    .out0(_14113_));
 b15nandp2aq1n24x5 _22892_ (.a(_13129_),
    .b(_13222_),
    .o1(_14114_));
 b15nona22ar1n32x5 _22893_ (.a(net789),
    .b(net780),
    .c(net795),
    .out0(_14115_));
 b15nand02an1n08x5 _22894_ (.a(_13124_),
    .b(_13240_),
    .o1(_14116_));
 b15nonb02ah1n06x5 _22895_ (.a(net773),
    .b(net794),
    .out0(_14117_));
 b15aoi012ar1n06x5 _22896_ (.a(_14058_),
    .b(_14117_),
    .c(_13131_),
    .o1(_14118_));
 b15nand02ah1n08x5 _22897_ (.a(_13244_),
    .b(_13252_),
    .o1(_14119_));
 b15nandp2as1n05x5 _22898_ (.a(_13092_),
    .b(_13208_),
    .o1(_14120_));
 b15oai222as1n16x5 _22899_ (.a(_14114_),
    .b(_14115_),
    .c(_14116_),
    .d(_14118_),
    .e(_14119_),
    .f(_14120_),
    .o1(_14121_));
 b15bfn001as1n64x5 wire410 (.a(\u0.tmp_w[30] ),
    .o(net410));
 b15nandp2ah1n05x5 _22901_ (.a(net769),
    .b(net791),
    .o1(_14123_));
 b15nano22ar1n16x5 _22902_ (.a(net774),
    .b(net778),
    .c(net771),
    .out0(_14124_));
 b15nanb02ar1n02x5 _22903_ (.a(_13193_),
    .b(_14124_),
    .out0(_14125_));
 b15nand04al1n02x5 _22904_ (.a(net773),
    .b(net794),
    .c(net783),
    .d(_13184_),
    .o1(_14126_));
 b15aoi012ah1n02x5 _22905_ (.a(_14123_),
    .b(_14125_),
    .c(_14126_),
    .o1(_14127_));
 b15nonb02aq1n04x5 _22906_ (.a(net778),
    .b(net780),
    .out0(_14128_));
 b15and002aq1n12x5 _22907_ (.a(net771),
    .b(net789),
    .o(_14129_));
 b15nand02ah1n06x5 _22908_ (.a(_14128_),
    .b(_14129_),
    .o1(_14130_));
 b15norp02aq1n12x5 _22909_ (.a(net776),
    .b(net769),
    .o1(_14131_));
 b15nandp2ar1n02x5 _22910_ (.a(_13252_),
    .b(_14131_),
    .o1(_14132_));
 b15oaoi13aq1n04x5 _22911_ (.a(_14130_),
    .b(_14132_),
    .c(_13065_),
    .d(_13252_),
    .o1(_14133_));
 b15norp03al1n08x5 _22912_ (.a(_14121_),
    .b(_14127_),
    .c(_14133_),
    .o1(_14134_));
 b15nand04as1n16x5 _22913_ (.a(_14094_),
    .b(_14111_),
    .c(_14113_),
    .d(_14134_),
    .o1(_14135_));
 b15nano23as1n24x5 _22914_ (.a(_14038_),
    .b(_14045_),
    .c(_14071_),
    .d(_14135_),
    .out0(_14136_));
 b15xor002as1n06x5 _22915_ (.a(net402),
    .b(_14136_),
    .out0(_14137_));
 b15xor002ar1n16x5 _22916_ (.a(_12776_),
    .b(_14137_),
    .out0(_14138_));
 b15xor002as1n12x5 _22917_ (.a(_13893_),
    .b(_14138_),
    .out0(_14139_));
 b15bfn001as1n64x5 max_length409 (.a(net410),
    .o(net409));
 b15oai012an1n24x5 _22919_ (.a(_13672_),
    .b(_14139_),
    .c(net533),
    .o1(_14141_));
 b15xor002al1n04x5 _22920_ (.a(_09932_),
    .b(_14141_),
    .out0(_00122_));
 b15nanb02ah1n04x5 _22921_ (.a(\text_in_r[2] ),
    .b(net533),
    .out0(_14142_));
 b15nanb02aq1n24x5 _22922_ (.a(net903),
    .b(net907),
    .out0(_14143_));
 b15nand02an1n08x5 _22923_ (.a(net901),
    .b(_12922_),
    .o1(_14144_));
 b15oai012ar1n02x5 _22924_ (.a(_12848_),
    .b(_12883_),
    .c(_12822_),
    .o1(_14145_));
 b15oai022ah1n04x5 _22925_ (.a(_12857_),
    .b(_14143_),
    .c(_14144_),
    .d(_14145_),
    .o1(_14146_));
 b15orn002aq1n08x5 _22926_ (.a(net889),
    .b(net912),
    .o(_14147_));
 b15oai012aq1n02x5 _22927_ (.a(_12811_),
    .b(net901),
    .c(_12832_),
    .o1(_14148_));
 b15oai012ar1n06x5 _22928_ (.a(net905),
    .b(_14147_),
    .c(_14148_),
    .o1(_14149_));
 b15oai112al1n08x5 _22929_ (.a(_12782_),
    .b(_13003_),
    .c(_12912_),
    .d(_13803_),
    .o1(_14150_));
 b15aoai13as1n06x5 _22930_ (.a(net897),
    .b(_14146_),
    .c(_14149_),
    .d(_14150_),
    .o1(_14151_));
 b15nandp2an1n16x5 _22931_ (.a(net886),
    .b(net889),
    .o1(_14152_));
 b15nor002ah1n04x5 _22932_ (.a(_14152_),
    .b(_13770_),
    .o1(_14153_));
 b15nor002as1n08x5 _22933_ (.a(net903),
    .b(_12877_),
    .o1(_14154_));
 b15aoi022an1n08x5 _22934_ (.a(net905),
    .b(_14153_),
    .c(_13013_),
    .d(_14154_),
    .o1(_14155_));
 b15oai012ar1n16x5 _22935_ (.a(_14151_),
    .b(_14155_),
    .c(net898),
    .o1(_14156_));
 b15and003aq1n03x5 _22936_ (.a(\us10.a[5] ),
    .b(net895),
    .c(net891),
    .o(_14157_));
 b15ao0022ar1n06x5 _22937_ (.a(_12864_),
    .b(_12916_),
    .c(_14157_),
    .d(net909),
    .o(_14158_));
 b15nand03al1n12x5 _22938_ (.a(net886),
    .b(_14154_),
    .c(_14158_),
    .o1(_14159_));
 b15oai013ar1n02x5 _22939_ (.a(_12851_),
    .b(_14152_),
    .c(_13011_),
    .d(_12913_),
    .o1(_14160_));
 b15aoi013al1n02x5 _22940_ (.a(_14160_),
    .b(_12909_),
    .c(_13794_),
    .d(net912),
    .o1(_14161_));
 b15nor002an1n03x5 _22941_ (.a(net901),
    .b(_13015_),
    .o1(_14162_));
 b15norp03ar1n02x5 _22942_ (.a(net911),
    .b(_13797_),
    .c(_13860_),
    .o1(_14163_));
 b15oai012al1n02x5 _22943_ (.a(_12959_),
    .b(_14162_),
    .c(_14163_),
    .o1(_14164_));
 b15nona23an1n16x5 _22944_ (.a(net893),
    .b(net889),
    .c(net886),
    .d(net896),
    .out0(_14165_));
 b15oai013al1n08x5 _22945_ (.a(net898),
    .b(_13015_),
    .c(_14165_),
    .d(net903),
    .o1(_14166_));
 b15oai022ar1n06x5 _22946_ (.a(net907),
    .b(_13012_),
    .c(_12913_),
    .d(_14152_),
    .o1(_14167_));
 b15aoi122ar1n04x5 _22947_ (.a(_14166_),
    .b(_14167_),
    .c(_12883_),
    .d(_13794_),
    .e(_13013_),
    .o1(_14168_));
 b15aoi022an1n02x5 _22948_ (.a(_14159_),
    .b(_14161_),
    .c(_14164_),
    .d(_14168_),
    .o1(_14169_));
 b15nor004al1n03x5 _22949_ (.a(net893),
    .b(net886),
    .c(_14147_),
    .d(_12960_),
    .o1(_14170_));
 b15aoi012ar1n02x5 _22950_ (.a(_12832_),
    .b(net901),
    .c(_14170_),
    .o1(_14171_));
 b15nand02ar1n02x5 _22951_ (.a(_12820_),
    .b(_14170_),
    .o1(_14172_));
 b15nanb02ar1n06x5 _22952_ (.a(net886),
    .b(net889),
    .out0(_14173_));
 b15mdn022aq1n03x5 _22953_ (.a(_14173_),
    .b(_12956_),
    .o1(_14174_),
    .sa(_13882_));
 b15nand04ar1n06x5 _22954_ (.a(net901),
    .b(_12851_),
    .c(_12922_),
    .d(_14174_),
    .o1(_14175_));
 b15aoi013an1n03x5 _22955_ (.a(_14171_),
    .b(_14172_),
    .c(_14175_),
    .d(_12832_),
    .o1(_14176_));
 b15nand02al1n24x5 _22956_ (.a(net903),
    .b(net898),
    .o1(_14177_));
 b15oai022al1n02x5 _22957_ (.a(_12857_),
    .b(_12954_),
    .c(_12800_),
    .d(_14177_),
    .o1(_14178_));
 b15oai013al1n04x5 _22958_ (.a(_12924_),
    .b(_12973_),
    .c(net901),
    .d(net897),
    .o1(_14179_));
 b15aoai13ah1n04x5 _22959_ (.a(net911),
    .b(_14178_),
    .c(_14179_),
    .d(net906),
    .o1(_14180_));
 b15aoi022as1n04x5 _22960_ (.a(_12968_),
    .b(_12825_),
    .c(_12909_),
    .d(_12863_),
    .o1(_14181_));
 b15nandp2ah1n03x5 _22961_ (.a(net905),
    .b(_14181_),
    .o1(_14182_));
 b15aoi013al1n02x5 _22962_ (.a(net905),
    .b(_12968_),
    .c(_12991_),
    .d(_12950_),
    .o1(_14183_));
 b15nanb02ah1n12x5 _22963_ (.a(net897),
    .b(net910),
    .out0(_14184_));
 b15nand02ar1n08x5 _22964_ (.a(net901),
    .b(_12789_),
    .o1(_14185_));
 b15aoai13ah1n03x5 _22965_ (.a(_14183_),
    .b(_14184_),
    .c(_12800_),
    .d(_14185_),
    .o1(_14186_));
 b15nandp3as1n04x5 _22966_ (.a(net897),
    .b(_12796_),
    .c(_12874_),
    .o1(_14187_));
 b15nandp2as1n04x5 _22967_ (.a(_12950_),
    .b(_12991_),
    .o1(_14188_));
 b15oai012ar1n08x5 _22968_ (.a(_14187_),
    .b(_14188_),
    .c(net897),
    .o1(_14189_));
 b15aoai13as1n08x5 _22969_ (.a(_14182_),
    .b(_14186_),
    .c(_12820_),
    .d(_14189_),
    .o1(_14190_));
 b15nona23ar1n16x5 _22970_ (.a(_14169_),
    .b(_14176_),
    .c(_14180_),
    .d(_14190_),
    .out0(_14191_));
 b15nand02ar1n24x5 _22971_ (.a(net907),
    .b(net900),
    .o1(_14192_));
 b15oai022ar1n02x5 _22972_ (.a(net899),
    .b(_13011_),
    .c(_14192_),
    .d(_13770_),
    .o1(_14193_));
 b15and003ar1n02x5 _22973_ (.a(_12848_),
    .b(_12971_),
    .c(_14193_),
    .o(_14194_));
 b15nand03ar1n16x5 _22974_ (.a(net898),
    .b(_12916_),
    .c(_12874_),
    .o1(_14195_));
 b15nandp3ar1n12x5 _22975_ (.o1(_14196_),
    .a(_12851_),
    .b(_12916_),
    .c(_12848_));
 b15oaoi13ah1n08x5 _22976_ (.a(net901),
    .b(_14195_),
    .c(_14196_),
    .d(_12904_),
    .o1(_14197_));
 b15nanb02ar1n06x5 _22977_ (.a(net900),
    .b(net887),
    .out0(_14198_));
 b15nand03ah1n02x5 _22978_ (.a(net890),
    .b(_12916_),
    .c(_13797_),
    .o1(_14199_));
 b15oaoi13al1n08x5 _22979_ (.a(_14198_),
    .b(_14199_),
    .c(_12949_),
    .d(_13835_),
    .o1(_14200_));
 b15nor003as1n04x5 _22980_ (.a(_14194_),
    .b(_14197_),
    .c(_14200_),
    .o1(_14201_));
 b15oai112as1n02x5 _22981_ (.a(_12851_),
    .b(_13794_),
    .c(_12825_),
    .d(net913),
    .o1(_14202_));
 b15aoi022an1n06x5 _22982_ (.a(net888),
    .b(_12883_),
    .c(_13884_),
    .d(\us10.a[5] ),
    .o1(_14203_));
 b15oaoi13an1n08x5 _22983_ (.a(_14202_),
    .b(net913),
    .c(_12864_),
    .d(_14203_),
    .o1(_14204_));
 b15nanb02al1n16x5 _22984_ (.a(net904),
    .b(net900),
    .out0(_14205_));
 b15nonb02al1n03x5 _22985_ (.a(net891),
    .b(net909),
    .out0(_14206_));
 b15aoi022ah1n06x5 _22986_ (.a(net909),
    .b(_12798_),
    .c(_14206_),
    .d(net888),
    .o1(_14207_));
 b15nandp2aq1n03x5 _22987_ (.a(net912),
    .b(_12883_),
    .o1(_14208_));
 b15oaoi13as1n08x5 _22988_ (.a(_14205_),
    .b(_13866_),
    .c(_14207_),
    .d(_14208_),
    .o1(_14209_));
 b15and002aq1n04x5 _22989_ (.a(net909),
    .b(net900),
    .o(_14210_));
 b15nonb02aq1n06x5 _22990_ (.a(net891),
    .b(\us10.a[5] ),
    .out0(_14211_));
 b15nonb03al1n02x5 _22991_ (.a(net904),
    .b(net888),
    .c(net895),
    .out0(_14212_));
 b15nano23ar1n03x5 _22992_ (.a(net895),
    .b(net888),
    .c(net913),
    .d(net904),
    .out0(_14213_));
 b15oai112ar1n08x5 _22993_ (.a(_14210_),
    .b(_14211_),
    .c(_14212_),
    .d(_14213_),
    .o1(_14214_));
 b15orn002al1n02x5 _22994_ (.a(net888),
    .b(net913),
    .o(_14215_));
 b15nand04ar1n12x5 _22995_ (.a(_12863_),
    .b(_13872_),
    .c(_14215_),
    .d(_14157_),
    .o1(_14216_));
 b15nano22an1n03x5 _22996_ (.a(net904),
    .b(net900),
    .c(net909),
    .out0(_14217_));
 b15oai112an1n04x5 _22997_ (.a(_12874_),
    .b(_14217_),
    .c(_12893_),
    .d(_12883_),
    .o1(_14218_));
 b15nand04al1n08x5 _22998_ (.a(net894),
    .b(_12848_),
    .c(_12908_),
    .d(_13801_),
    .o1(_14219_));
 b15nand04aq1n08x5 _22999_ (.a(_14214_),
    .b(_14216_),
    .c(_14218_),
    .d(_14219_),
    .o1(_14220_));
 b15aoi012aq1n04x5 _23000_ (.a(_12789_),
    .b(_12798_),
    .c(_12822_),
    .o1(_14221_));
 b15nand02al1n06x5 _23001_ (.a(_12968_),
    .b(_12877_),
    .o1(_14222_));
 b15nonb02al1n12x5 _23002_ (.a(net900),
    .b(net913),
    .out0(_14223_));
 b15nand02as1n04x5 _23003_ (.a(_14211_),
    .b(_14223_),
    .o1(_14224_));
 b15aoi022as1n08x5 _23004_ (.a(_13797_),
    .b(_13884_),
    .c(_13860_),
    .d(_13883_),
    .o1(_14225_));
 b15aoi012ah1n06x5 _23005_ (.a(_13854_),
    .b(_12798_),
    .c(\us10.a[5] ),
    .o1(_14226_));
 b15nand02al1n06x5 _23006_ (.a(_12832_),
    .b(_12863_),
    .o1(_14227_));
 b15oai222as1n16x5 _23007_ (.a(_14221_),
    .b(_14222_),
    .c(_14224_),
    .d(_14225_),
    .e(_14226_),
    .f(_14227_),
    .o1(_14228_));
 b15nor004as1n12x5 _23008_ (.a(_14204_),
    .b(_14209_),
    .c(_14220_),
    .d(_14228_),
    .o1(_14229_));
 b15nandp2al1n08x5 _23009_ (.a(net905),
    .b(_13817_),
    .o1(_14230_));
 b15oai022ar1n06x5 _23010_ (.a(_12950_),
    .b(_12902_),
    .c(_14230_),
    .d(net899),
    .o1(_14231_));
 b15oai013al1n04x5 _23011_ (.a(net902),
    .b(_12949_),
    .c(_12978_),
    .d(net911),
    .o1(_14232_));
 b15and003aq1n04x5 _23012_ (.a(net892),
    .b(net890),
    .c(net900),
    .o(_14233_));
 b15nandp2an1n08x5 _23013_ (.a(_12940_),
    .b(_14233_),
    .o1(_14234_));
 b15oai122as1n04x5 _23014_ (.a(_12820_),
    .b(_12875_),
    .c(_12960_),
    .d(_14234_),
    .e(_12879_),
    .o1(_14235_));
 b15nand03ah1n12x5 _23015_ (.a(_12851_),
    .b(_12796_),
    .c(_12874_),
    .o1(_14236_));
 b15oaoi13aq1n03x5 _23016_ (.a(net911),
    .b(_14236_),
    .c(_14234_),
    .d(_12782_),
    .o1(_14237_));
 b15oai022an1n08x5 _23017_ (.a(_14231_),
    .b(_14232_),
    .c(_14235_),
    .d(_14237_),
    .o1(_14238_));
 b15aoai13ar1n06x5 _23018_ (.a(_12904_),
    .b(_12909_),
    .c(_12822_),
    .d(_12881_),
    .o1(_14239_));
 b15oai122an1n12x5 _23019_ (.a(net902),
    .b(_12904_),
    .c(_14236_),
    .d(_14239_),
    .e(_12851_),
    .o1(_14240_));
 b15nonb02an1n08x5 _23020_ (.a(net887),
    .b(net900),
    .out0(_14241_));
 b15aoi022ah1n02x5 _23021_ (.a(net894),
    .b(_14241_),
    .c(_14223_),
    .d(_13884_),
    .o1(_14242_));
 b15nandp2aq1n02x5 _23022_ (.a(net906),
    .b(_12983_),
    .o1(_14243_));
 b15oai022al1n08x5 _23023_ (.a(_12954_),
    .b(_14165_),
    .c(_14242_),
    .d(_14243_),
    .o1(_14244_));
 b15oai012ah1n08x5 _23024_ (.a(_14240_),
    .b(_14244_),
    .c(net902),
    .o1(_14245_));
 b15nand04as1n16x5 _23025_ (.a(_14201_),
    .b(_14229_),
    .c(_14238_),
    .d(_14245_),
    .o1(_14246_));
 b15norp03as1n24x5 _23026_ (.a(_14156_),
    .b(_14191_),
    .c(_14246_),
    .o1(_14247_));
 b15norp02ar1n02x5 _23027_ (.a(_13086_),
    .b(_13089_),
    .o1(_14248_));
 b15nor002aq1n16x5 _23028_ (.a(_13030_),
    .b(_14025_),
    .o1(_14249_));
 b15aoai13an1n02x5 _23029_ (.a(net782),
    .b(_14248_),
    .c(_14249_),
    .d(net788),
    .o1(_14250_));
 b15nandp2al1n02x5 _23030_ (.a(_13244_),
    .b(_13090_),
    .o1(_14251_));
 b15nand03al1n02x5 _23031_ (.a(_13184_),
    .b(_13124_),
    .c(_13222_),
    .o1(_14252_));
 b15aoai13aq1n03x5 _23032_ (.a(net791),
    .b(net796),
    .c(_14251_),
    .d(_14252_),
    .o1(_14253_));
 b15nor002an1n24x5 _23033_ (.a(net779),
    .b(\us21.a[6] ),
    .o1(_14254_));
 b15aoi022an1n08x5 _23034_ (.a(_13174_),
    .b(_14254_),
    .c(_14129_),
    .d(_13129_),
    .o1(_14255_));
 b15qgbin1an1n15x5 _23035_ (.a(net768),
    .o1(_14256_));
 b15oai013ah1n12x5 _23036_ (.a(_13063_),
    .b(net784),
    .c(_14255_),
    .d(_14256_),
    .o1(_14257_));
 b15nand02ar1n02x5 _23037_ (.a(net788),
    .b(_14030_),
    .o1(_14258_));
 b15oaoi13an1n03x5 _23038_ (.a(_13022_),
    .b(_14258_),
    .c(_14034_),
    .d(net788),
    .o1(_14259_));
 b15obai22ah1n06x5 _23039_ (.a(_14250_),
    .b(_14253_),
    .c(_14257_),
    .d(_14259_),
    .out0(_14260_));
 b15aoai13al1n02x5 _23040_ (.a(net792),
    .b(_13171_),
    .c(_13091_),
    .d(_13092_),
    .o1(_14261_));
 b15aoi012an1n02x5 _23041_ (.a(_13211_),
    .b(_14073_),
    .c(_14261_),
    .o1(_14262_));
 b15nand03ar1n03x5 _23042_ (.a(net792),
    .b(net788),
    .c(_13249_),
    .o1(_14263_));
 b15oai013as1n03x5 _23043_ (.a(_14263_),
    .b(_14020_),
    .c(_13159_),
    .d(net792),
    .o1(_14264_));
 b15aoi012al1n06x5 _23044_ (.a(_14262_),
    .b(_14264_),
    .c(_13022_),
    .o1(_14265_));
 b15nanb03an1n12x5 _23045_ (.a(net771),
    .b(net768),
    .c(net778),
    .out0(_14266_));
 b15nand02al1n04x5 _23046_ (.a(_13174_),
    .b(net794),
    .o1(_14267_));
 b15aoi112as1n06x5 _23047_ (.a(_14085_),
    .b(_14266_),
    .c(_14267_),
    .d(net790),
    .o1(_14268_));
 b15xor002aq1n08x5 _23048_ (.a(net777),
    .b(net785),
    .out0(_14269_));
 b15nanb02al1n08x5 _23049_ (.a(net780),
    .b(net771),
    .out0(_14270_));
 b15nano23an1n02x5 _23050_ (.a(_13252_),
    .b(_14269_),
    .c(_14270_),
    .d(_13065_),
    .out0(_14271_));
 b15norp03ar1n02x5 _23051_ (.a(_13086_),
    .b(_14085_),
    .c(_14103_),
    .o1(_14272_));
 b15nor002aq1n06x5 _23052_ (.a(_13142_),
    .b(_14095_),
    .o1(_14273_));
 b15orn003as1n02x5 _23053_ (.a(_14271_),
    .b(_14272_),
    .c(_14273_),
    .o(_14274_));
 b15nand03ah1n06x5 _23054_ (.a(_13146_),
    .b(_13129_),
    .c(_13222_),
    .o1(_14275_));
 b15nand03ar1n08x5 _23055_ (.a(net794),
    .b(_13125_),
    .c(_14275_),
    .o1(_14276_));
 b15oai112ah1n04x5 _23056_ (.a(_13128_),
    .b(_13129_),
    .c(_13251_),
    .d(_13215_),
    .o1(_14277_));
 b15oai112an1n12x5 _23057_ (.a(_13067_),
    .b(_14277_),
    .c(_13272_),
    .d(_14085_),
    .o1(_14278_));
 b15aoi112as1n08x5 _23058_ (.a(_14268_),
    .b(_14274_),
    .c(_14276_),
    .d(_14278_),
    .o1(_14279_));
 b15norp03ar1n03x5 _23059_ (.a(net769),
    .b(_13078_),
    .c(_14036_),
    .o1(_14280_));
 b15and002ar1n24x5 _23060_ (.a(net794),
    .b(net785),
    .o(_14281_));
 b15oai112al1n12x5 _23061_ (.a(_13131_),
    .b(_13233_),
    .c(_14281_),
    .d(_13174_),
    .o1(_14282_));
 b15aoi012ar1n06x5 _23062_ (.a(_13022_),
    .b(_13072_),
    .c(_13171_),
    .o1(_14283_));
 b15nor004ah1n06x5 _23063_ (.a(net776),
    .b(net779),
    .c(net772),
    .d(net788),
    .o1(_14284_));
 b15and002ah1n12x5 _23064_ (.a(net773),
    .b(\us21.a[0] ),
    .o(_14285_));
 b15aoi013ah1n04x5 _23065_ (.a(_14284_),
    .b(_14285_),
    .c(net787),
    .d(_13129_),
    .o1(_14286_));
 b15oai112as1n16x5 _23066_ (.a(_14282_),
    .b(_14283_),
    .c(_14286_),
    .d(_14256_),
    .o1(_14287_));
 b15nand04as1n16x5 _23067_ (.a(net776),
    .b(net779),
    .c(net770),
    .d(net772),
    .o1(_14288_));
 b15oai022as1n06x5 _23068_ (.a(_13063_),
    .b(_14288_),
    .c(_14103_),
    .d(_13159_),
    .o1(_14289_));
 b15aoai13an1n06x5 _23069_ (.a(_14280_),
    .b(_14287_),
    .c(_13114_),
    .d(_14289_),
    .o1(_14290_));
 b15nand04an1n16x5 _23070_ (.a(_14260_),
    .b(_14265_),
    .c(_14279_),
    .d(_14290_),
    .o1(_14291_));
 b15nand03ar1n03x5 _23071_ (.a(net796),
    .b(net784),
    .c(_13249_),
    .o1(_14292_));
 b15nandp2al1n04x5 _23072_ (.a(net784),
    .b(_13249_),
    .o1(_14293_));
 b15nandp3an1n08x5 _23073_ (.a(_13022_),
    .b(_13128_),
    .c(_13129_),
    .o1(_14294_));
 b15aoai13ah1n03x5 _23074_ (.a(_14292_),
    .b(net791),
    .c(_14293_),
    .d(_14294_),
    .o1(_14295_));
 b15nand02as1n32x5 _23075_ (.a(_13091_),
    .b(_13176_),
    .o1(_14296_));
 b15oai022ah1n04x5 _23076_ (.a(_13040_),
    .b(_14296_),
    .c(_13075_),
    .d(_13277_),
    .o1(_14297_));
 b15aoai13an1n04x5 _23077_ (.a(net786),
    .b(_14295_),
    .c(_14297_),
    .d(_14287_),
    .o1(_14298_));
 b15nand04aq1n04x5 _23078_ (.a(_13114_),
    .b(_13091_),
    .c(_13176_),
    .d(_13040_),
    .o1(_14299_));
 b15oai112al1n12x5 _23079_ (.a(net781),
    .b(_14299_),
    .c(_13095_),
    .d(_13130_),
    .o1(_14300_));
 b15nor002ar1n08x5 _23080_ (.a(net794),
    .b(net785),
    .o1(_14301_));
 b15oai022an1n06x5 _23081_ (.a(_13141_),
    .b(_14029_),
    .c(_14301_),
    .d(_13185_),
    .o1(_14302_));
 b15oai012al1n06x5 _23082_ (.a(_13282_),
    .b(_13283_),
    .c(_13130_),
    .o1(_14303_));
 b15oai013al1n08x5 _23083_ (.a(_14300_),
    .b(_14302_),
    .c(net781),
    .d(_14303_),
    .o1(_14304_));
 b15nanb02ah1n02x5 _23084_ (.a(_14096_),
    .b(_14275_),
    .out0(_14305_));
 b15oai022aq1n06x5 _23085_ (.a(net781),
    .b(_13142_),
    .c(_13154_),
    .d(_13292_),
    .o1(_14306_));
 b15nand02as1n03x5 _23086_ (.a(net785),
    .b(_13255_),
    .o1(_14307_));
 b15oai022ah1n08x5 _23087_ (.a(net785),
    .b(_14305_),
    .c(_14306_),
    .d(_14307_),
    .o1(_14308_));
 b15nand04as1n02x5 _23088_ (.a(_13092_),
    .b(_13208_),
    .c(_13072_),
    .d(_13251_),
    .o1(_14309_));
 b15oai012aq1n08x5 _23089_ (.a(_14309_),
    .b(_14296_),
    .c(_14053_),
    .o1(_14310_));
 b15oaoi13al1n04x5 _23090_ (.a(_14034_),
    .b(_14119_),
    .c(_13072_),
    .d(net781),
    .o1(_14311_));
 b15oai012as1n04x5 _23091_ (.a(_14066_),
    .b(_13161_),
    .c(net781),
    .o1(_14312_));
 b15nonb03as1n12x5 _23092_ (.a(net794),
    .b(net793),
    .c(net785),
    .out0(_14313_));
 b15aoi112ar1n08x5 _23093_ (.a(_14310_),
    .b(_14311_),
    .c(_14312_),
    .d(_14313_),
    .o1(_14314_));
 b15nand04aq1n16x5 _23094_ (.a(_14298_),
    .b(_14304_),
    .c(_14308_),
    .d(_14314_),
    .o1(_14315_));
 b15nand04as1n16x5 _23095_ (.a(_13063_),
    .b(_13092_),
    .c(_13091_),
    .d(_13244_),
    .o1(_14316_));
 b15nor002aq1n06x5 _23096_ (.a(net791),
    .b(net784),
    .o1(_14317_));
 b15nandp2ar1n03x5 _23097_ (.a(_13181_),
    .b(_14317_),
    .o1(_14318_));
 b15aoi013ar1n02x5 _23098_ (.a(net796),
    .b(_13176_),
    .c(_13208_),
    .d(_13215_),
    .o1(_14319_));
 b15nano22ar1n02x5 _23099_ (.a(net792),
    .b(net782),
    .c(net788),
    .out0(_14320_));
 b15oai112al1n02x5 _23100_ (.a(_13092_),
    .b(_14320_),
    .c(_13208_),
    .d(_13091_),
    .o1(_14321_));
 b15nand04aq1n04x5 _23101_ (.a(_14316_),
    .b(_14318_),
    .c(_14319_),
    .d(_14321_),
    .o1(_14322_));
 b15nand03al1n03x5 _23102_ (.a(net782),
    .b(_13184_),
    .c(_13222_),
    .o1(_14323_));
 b15nandp2ar1n02x5 _23103_ (.a(_13124_),
    .b(_13249_),
    .o1(_14324_));
 b15nandp2ar1n02x5 _23104_ (.a(_13147_),
    .b(_13251_),
    .o1(_14325_));
 b15aoi013an1n03x5 _23105_ (.a(_13063_),
    .b(_14323_),
    .c(_14324_),
    .d(_14325_),
    .o1(_14326_));
 b15oai013aq1n03x5 _23106_ (.a(net796),
    .b(net792),
    .c(_13211_),
    .d(_13227_),
    .o1(_14327_));
 b15oaoi13as1n02x5 _23107_ (.a(_13086_),
    .b(_13211_),
    .c(_13215_),
    .d(net792),
    .o1(_14328_));
 b15oai022an1n08x5 _23108_ (.a(_14322_),
    .b(_14326_),
    .c(_14327_),
    .d(_14328_),
    .o1(_14329_));
 b15aoi012ar1n04x5 _23109_ (.a(_14287_),
    .b(_14289_),
    .c(_13114_),
    .o1(_14330_));
 b15oaoi13an1n04x5 _23110_ (.a(_13075_),
    .b(_13210_),
    .c(net795),
    .d(_14029_),
    .o1(_14331_));
 b15nandp3as1n03x5 _23111_ (.a(_13174_),
    .b(net793),
    .c(_13092_),
    .o1(_14332_));
 b15oai022ah1n12x5 _23112_ (.a(_13142_),
    .b(_13277_),
    .c(_14269_),
    .d(_14332_),
    .o1(_14333_));
 b15oai012ar1n08x5 _23113_ (.a(_14067_),
    .b(_14035_),
    .c(_13067_),
    .o1(_14334_));
 b15aoi112al1n08x5 _23114_ (.a(_14331_),
    .b(_14333_),
    .c(_14334_),
    .d(_13054_),
    .o1(_14335_));
 b15aoai13aq1n08x5 _23115_ (.a(_14329_),
    .b(_13022_),
    .c(_14330_),
    .d(_14335_),
    .o1(_14336_));
 b15norp03as1n24x5 _23116_ (.a(_14291_),
    .b(_14315_),
    .c(_14336_),
    .o1(_14337_));
 b15xnr002an1n16x5 _23117_ (.a(_14247_),
    .b(_14337_),
    .out0(_14338_));
 b15aoai13ar1n02x5 _23118_ (.a(_13380_),
    .b(_13412_),
    .c(_13996_),
    .d(net667),
    .o1(_14339_));
 b15oab012ar1n02x5 _23119_ (.a(_13421_),
    .b(_13330_),
    .c(_13504_),
    .out0(_14340_));
 b15norp03ar1n02x5 _23120_ (.a(_13315_),
    .b(_13423_),
    .c(_13350_),
    .o1(_14341_));
 b15oai022ar1n04x5 _23121_ (.a(_13324_),
    .b(_13343_),
    .c(_13350_),
    .d(_13315_),
    .o1(_14342_));
 b15aoai13an1n03x5 _23122_ (.a(net657),
    .b(_14341_),
    .c(_14342_),
    .d(_13418_),
    .o1(_14343_));
 b15aoi012ar1n02x5 _23123_ (.a(net661),
    .b(_13996_),
    .c(_13472_),
    .o1(_14344_));
 b15aoi022as1n02x5 _23124_ (.a(_14339_),
    .b(_14340_),
    .c(_14343_),
    .d(_14344_),
    .o1(_14345_));
 b15aoi022ar1n02x5 _23125_ (.a(_14000_),
    .b(_13371_),
    .c(_13368_),
    .d(_13924_),
    .o1(_14346_));
 b15norp02aq1n03x5 _23126_ (.a(net657),
    .b(_14346_),
    .o1(_14347_));
 b15aoai13al1n02x5 _23127_ (.a(_13340_),
    .b(_13897_),
    .c(_13522_),
    .d(net668),
    .o1(_14348_));
 b15and002ar1n02x5 _23128_ (.a(net668),
    .b(net645),
    .o(_14349_));
 b15aoai13aq1n02x5 _23129_ (.a(_14349_),
    .b(_13536_),
    .c(_13534_),
    .d(\us32.a[1] ),
    .o1(_14350_));
 b15aob012an1n12x5 _23130_ (.a(_13407_),
    .b(_14348_),
    .c(_14350_),
    .out0(_14351_));
 b15norp03ar1n02x5 _23131_ (.a(net667),
    .b(_13315_),
    .c(_13318_),
    .o1(_14352_));
 b15oai112an1n02x5 _23132_ (.a(net663),
    .b(net661),
    .c(_13912_),
    .d(_14352_),
    .o1(_14353_));
 b15nor003ah1n02x5 _23133_ (.a(_13355_),
    .b(_13315_),
    .c(_13318_),
    .o1(_14354_));
 b15norp02ar1n02x5 _23134_ (.a(net667),
    .b(_13500_),
    .o1(_14355_));
 b15oai022an1n02x5 _23135_ (.a(_13371_),
    .b(_13965_),
    .c(_14354_),
    .d(_14355_),
    .o1(_14356_));
 b15nand04aq1n04x5 _23136_ (.a(_13896_),
    .b(_14351_),
    .c(_14353_),
    .d(_14356_),
    .o1(_14357_));
 b15aoi112ah1n04x5 _23137_ (.a(_14345_),
    .b(_14347_),
    .c(_14357_),
    .d(net657),
    .o1(_14358_));
 b15aoai13ah1n03x5 _23138_ (.a(_13380_),
    .b(_13325_),
    .c(_13523_),
    .d(_13438_),
    .o1(_14359_));
 b15aoai13al1n04x5 _23139_ (.a(_13368_),
    .b(_14002_),
    .c(net655),
    .d(_13996_),
    .o1(_14360_));
 b15nanb02al1n12x5 _23140_ (.a(net657),
    .b(net651),
    .out0(_14361_));
 b15norp02as1n03x5 _23141_ (.a(_13431_),
    .b(_14361_),
    .o1(_14362_));
 b15orn002ar1n08x5 _23142_ (.a(net654),
    .b(net643),
    .o(_14363_));
 b15nor003ah1n04x5 _23143_ (.a(net649),
    .b(_13310_),
    .c(_14363_),
    .o1(_14364_));
 b15oai112al1n16x5 _23144_ (.a(net646),
    .b(_13965_),
    .c(_14362_),
    .d(_14364_),
    .o1(_14365_));
 b15qgbno3an1n05x5 _23145_ (.o1(_14366_),
    .a(net667),
    .b(net655),
    .c(net659));
 b15nand02al1n02x5 _23146_ (.a(_13496_),
    .b(_14366_),
    .o1(_14367_));
 b15aob012al1n12x5 _23147_ (.a(_13340_),
    .b(_13416_),
    .c(_14367_),
    .out0(_14368_));
 b15nand04ah1n12x5 _23148_ (.a(_14359_),
    .b(_14360_),
    .c(_14365_),
    .d(_14368_),
    .o1(_14369_));
 b15aoi112ar1n02x5 _23149_ (.a(net655),
    .b(_13528_),
    .c(_13367_),
    .d(net663),
    .o1(_14370_));
 b15aoai13ah1n02x5 _23150_ (.a(_14370_),
    .b(_14000_),
    .c(net659),
    .d(_13980_),
    .o1(_14371_));
 b15nor003al1n02x5 _23151_ (.a(net659),
    .b(_13330_),
    .c(_13939_),
    .o1(_14372_));
 b15aoi012ar1n04x5 _23152_ (.a(_14372_),
    .b(_13965_),
    .c(_13415_),
    .o1(_14373_));
 b15oai012ar1n08x5 _23153_ (.a(_14371_),
    .b(_14373_),
    .c(net655),
    .o1(_14374_));
 b15aoi012ar1n02x5 _23154_ (.a(_13355_),
    .b(_13447_),
    .c(_13499_),
    .o1(_14375_));
 b15aoai13ar1n02x5 _23155_ (.a(_13442_),
    .b(_14375_),
    .c(net655),
    .d(_13418_),
    .o1(_14376_));
 b15inv000ah1n16x5 _23156_ (.a(net644),
    .o1(_14377_));
 b15nand02ah1n04x5 _23157_ (.a(net654),
    .b(_14377_),
    .o1(_14378_));
 b15orn002aq1n04x5 _23158_ (.a(net668),
    .b(net658),
    .o(_14379_));
 b15orn003ah1n03x5 _23159_ (.a(_13459_),
    .b(_14379_),
    .c(_13399_),
    .o(_14380_));
 b15orn003ar1n08x5 _23160_ (.a(net664),
    .b(_14378_),
    .c(_14380_),
    .o(_14381_));
 b15nand04aq1n04x5 _23161_ (.a(_13313_),
    .b(_13514_),
    .c(_13530_),
    .d(_13979_),
    .o1(_14382_));
 b15nandp3al1n04x5 _23162_ (.a(_14376_),
    .b(_14381_),
    .c(_14382_),
    .o1(_14383_));
 b15norp02ar1n02x5 _23163_ (.a(_13318_),
    .b(_13960_),
    .o1(_14384_));
 b15aoi012ar1n02x5 _23164_ (.a(_13350_),
    .b(_13504_),
    .c(_13960_),
    .o1(_14385_));
 b15oai112an1n04x5 _23165_ (.a(net659),
    .b(_13375_),
    .c(_14384_),
    .d(_14385_),
    .o1(_14386_));
 b15oaoi13ah1n03x5 _23166_ (.a(_13942_),
    .b(_13367_),
    .c(net663),
    .d(_13528_),
    .o1(_14387_));
 b15nanb02as1n24x5 _23167_ (.a(net659),
    .b(net666),
    .out0(_14388_));
 b15aoi012as1n02x5 _23168_ (.a(_13494_),
    .b(_14388_),
    .c(_13425_),
    .o1(_14389_));
 b15oai012ar1n08x5 _23169_ (.a(_13313_),
    .b(_14387_),
    .c(_14389_),
    .o1(_14390_));
 b15nor004al1n02x5 _23170_ (.a(net667),
    .b(net659),
    .c(_13315_),
    .d(_13318_),
    .o1(_14391_));
 b15aoi013as1n02x5 _23171_ (.a(_14391_),
    .b(_13514_),
    .c(_13996_),
    .d(net659),
    .o1(_14392_));
 b15oai112aq1n08x5 _23172_ (.a(_14386_),
    .b(_14390_),
    .c(net655),
    .d(_14392_),
    .o1(_14393_));
 b15nor004as1n08x5 _23173_ (.a(_14369_),
    .b(_14374_),
    .c(_14383_),
    .d(_14393_),
    .o1(_14394_));
 b15and003as1n04x5 _23174_ (.a(_13421_),
    .b(_13403_),
    .c(_13938_),
    .o(_14395_));
 b15nor003as1n02x5 _23175_ (.a(_13340_),
    .b(net651),
    .c(_13479_),
    .o1(_14396_));
 b15nor004as1n03x5 _23176_ (.a(net664),
    .b(net653),
    .c(_13343_),
    .d(_13399_),
    .o1(_14397_));
 b15oaoi13ar1n04x5 _23177_ (.a(_14395_),
    .b(net656),
    .c(_14396_),
    .d(_14397_),
    .o1(_14398_));
 b15norp02ar1n02x5 _23178_ (.a(_13425_),
    .b(_13347_),
    .o1(_14399_));
 b15nand02as1n08x5 _23179_ (.a(net651),
    .b(net645),
    .o1(_14400_));
 b15oai012ar1n02x5 _23180_ (.a(_14400_),
    .b(_13302_),
    .c(net651),
    .o1(_14401_));
 b15nand03as1n03x5 _23181_ (.a(net668),
    .b(net651),
    .c(net644),
    .o1(_14402_));
 b15oai022ar1n02x5 _23182_ (.a(net651),
    .b(_13441_),
    .c(_14402_),
    .d(net647),
    .o1(_14403_));
 b15aoi022al1n02x5 _23183_ (.a(_14399_),
    .b(_14401_),
    .c(_14403_),
    .d(_13905_),
    .o1(_14404_));
 b15oai022an1n06x5 _23184_ (.a(net668),
    .b(_14398_),
    .c(_14404_),
    .d(_13374_),
    .o1(_14405_));
 b15nanb02as1n06x5 _23185_ (.a(net645),
    .b(net651),
    .out0(_14406_));
 b15oai112ar1n02x5 _23186_ (.a(net657),
    .b(_13917_),
    .c(_14406_),
    .d(net665),
    .o1(_14407_));
 b15aoi012ar1n02x5 _23187_ (.a(_14377_),
    .b(_13488_),
    .c(net651),
    .o1(_14408_));
 b15oai012an1n04x5 _23188_ (.a(_13340_),
    .b(_13483_),
    .c(_13478_),
    .o1(_14409_));
 b15oa0022an1n02x5 _23189_ (.a(_14407_),
    .b(_14408_),
    .c(_14409_),
    .d(_13479_),
    .o(_14410_));
 b15aoi013ar1n02x5 _23190_ (.a(_13421_),
    .b(_13950_),
    .c(_13496_),
    .d(_13313_),
    .o1(_14411_));
 b15aoi022ar1n04x5 _23191_ (.a(_13421_),
    .b(_14410_),
    .c(_14411_),
    .d(_13416_),
    .o1(_14412_));
 b15orn002ar1n12x5 _23192_ (.a(_14405_),
    .b(_14412_),
    .o(_14413_));
 b15nano23an1n03x5 _23193_ (.a(net657),
    .b(net661),
    .c(net645),
    .d(net667),
    .out0(_14414_));
 b15oab012ah1n06x5 _23194_ (.a(_14414_),
    .b(_14012_),
    .c(_14388_),
    .out0(_14415_));
 b15nanb02as1n16x5 _23195_ (.a(net654),
    .b(net647),
    .out0(_14416_));
 b15oai022ah1n06x5 _23196_ (.a(_13968_),
    .b(_14380_),
    .c(_14415_),
    .d(_14416_),
    .o1(_14417_));
 b15nandp3al1n04x5 _23197_ (.a(_13515_),
    .b(_13382_),
    .c(_13362_),
    .o1(_14418_));
 b15aoi022ah1n04x5 _23198_ (.a(_13434_),
    .b(_13407_),
    .c(_13920_),
    .d(_13435_),
    .o1(_14419_));
 b15nanb02aq1n06x5 _23199_ (.a(net647),
    .b(net658),
    .out0(_14420_));
 b15oaoi13an1n08x5 _23200_ (.a(_13355_),
    .b(_14418_),
    .c(_14419_),
    .d(_14420_),
    .o1(_14421_));
 b15oai012ar1n16x5 _23201_ (.a(net664),
    .b(_14417_),
    .c(_14421_),
    .o1(_14422_));
 b15nanb02ah1n12x5 _23202_ (.a(_13947_),
    .b(_14422_),
    .out0(_14423_));
 b15nano23as1n24x5 _23203_ (.a(_14358_),
    .b(_14394_),
    .c(_14413_),
    .d(_14423_),
    .out0(_14424_));
 b15aob012ar1n02x5 _23204_ (.a(_13656_),
    .b(net627),
    .c(net639),
    .out0(_14425_));
 b15oai013al1n02x5 _23205_ (.a(net631),
    .b(_12657_),
    .c(_13556_),
    .d(_14425_),
    .o1(_14426_));
 b15xor002al1n02x5 _23206_ (.a(net642),
    .b(\us03.a[7] ),
    .out0(_14427_));
 b15aoi013an1n03x5 _23207_ (.a(_12515_),
    .b(net628),
    .c(_13717_),
    .d(_14427_),
    .o1(_14428_));
 b15aoi012ah1n04x5 _23208_ (.a(_13701_),
    .b(_12587_),
    .c(net627),
    .o1(_14429_));
 b15oai013ar1n02x5 _23209_ (.a(_14428_),
    .b(_14429_),
    .c(_12700_),
    .d(net628),
    .o1(_14430_));
 b15oai012as1n04x5 _23210_ (.a(_12515_),
    .b(_12714_),
    .c(_12615_),
    .o1(_14431_));
 b15aoi012aq1n02x5 _23211_ (.a(_14426_),
    .b(_14430_),
    .c(_14431_),
    .o1(_14432_));
 b15nor002as1n03x5 _23212_ (.a(net641),
    .b(_12760_),
    .o1(_14433_));
 b15aoai13an1n06x5 _23213_ (.a(_13676_),
    .b(_14433_),
    .c(net641),
    .d(_12752_),
    .o1(_14434_));
 b15nanb03ah1n03x5 _23214_ (.a(net627),
    .b(net621),
    .c(net623),
    .out0(_14435_));
 b15aoai13ar1n03x5 _23215_ (.a(_14435_),
    .b(_12581_),
    .c(_12552_),
    .d(_13660_),
    .o1(_14436_));
 b15nand04al1n03x5 _23216_ (.a(net642),
    .b(_12515_),
    .c(net628),
    .d(_14436_),
    .o1(_14437_));
 b15norp02ar1n02x5 _23217_ (.a(_12511_),
    .b(_12569_),
    .o1(_14438_));
 b15aoi012ar1n02x5 _23218_ (.a(net639),
    .b(_12766_),
    .c(_13618_),
    .o1(_14439_));
 b15aoai13ar1n02x5 _23219_ (.a(_14438_),
    .b(_14439_),
    .c(net635),
    .d(_12586_),
    .o1(_14440_));
 b15aoi012ar1n08x5 _23220_ (.a(net632),
    .b(net635),
    .c(_13688_),
    .o1(_14441_));
 b15nand04al1n04x5 _23221_ (.a(_14434_),
    .b(_14437_),
    .c(_14440_),
    .d(_14441_),
    .o1(_14442_));
 b15nanb02ar1n02x5 _23222_ (.a(net627),
    .b(net639),
    .out0(_14443_));
 b15norp02ar1n02x5 _23223_ (.a(net642),
    .b(\us03.a[7] ),
    .o1(_14444_));
 b15norp02ar1n02x5 _23224_ (.a(\us03.a[2] ),
    .b(net628),
    .o1(_14445_));
 b15aoai13al1n02x5 _23225_ (.a(_14444_),
    .b(_14445_),
    .c(\us03.a[2] ),
    .d(_12666_),
    .o1(_14446_));
 b15oaoi13an1n03x5 _23226_ (.a(_14443_),
    .b(_14446_),
    .c(net628),
    .d(_12552_),
    .o1(_14447_));
 b15oab012ah1n06x5 _23227_ (.a(_14432_),
    .b(_14442_),
    .c(_14447_),
    .out0(_14448_));
 b15nand02an1n08x5 _23228_ (.a(net635),
    .b(_12671_),
    .o1(_14449_));
 b15aoi012ar1n02x5 _23229_ (.a(net631),
    .b(_12515_),
    .c(net621),
    .o1(_14450_));
 b15and003aq1n02x5 _23230_ (.a(_12563_),
    .b(_14449_),
    .c(_14450_),
    .o(_14451_));
 b15nand02an1n02x5 _23231_ (.a(_12632_),
    .b(_12636_),
    .o1(_14452_));
 b15nandp2ar1n05x5 _23232_ (.a(\us03.a[4] ),
    .b(\us03.a[7] ),
    .o1(_14453_));
 b15oaoi13an1n08x5 _23233_ (.a(_12545_),
    .b(_14452_),
    .c(_14453_),
    .d(\us03.a[5] ),
    .o1(_14454_));
 b15oai112an1n12x5 _23234_ (.a(_12581_),
    .b(_13602_),
    .c(_14451_),
    .d(_14454_),
    .o1(_14455_));
 b15nona23al1n12x5 _23235_ (.a(_12639_),
    .b(_12650_),
    .c(_13586_),
    .d(_14455_),
    .out0(_14456_));
 b15aoi012ar1n02x5 _23236_ (.a(net639),
    .b(net641),
    .c(_13712_),
    .o1(_14457_));
 b15aoi112al1n02x5 _23237_ (.a(_13580_),
    .b(_14457_),
    .c(_12566_),
    .d(_12619_),
    .o1(_14458_));
 b15aoi122ar1n02x5 _23238_ (.a(net631),
    .b(_12550_),
    .c(_12551_),
    .d(_13624_),
    .e(_12515_),
    .o1(_14459_));
 b15and002ar1n02x5 _23239_ (.a(net639),
    .b(_12689_),
    .o(_14460_));
 b15aoi022ar1n02x5 _23240_ (.a(_12570_),
    .b(_13676_),
    .c(_14460_),
    .d(_13607_),
    .o1(_14461_));
 b15aoi012ar1n02x5 _23241_ (.a(_14459_),
    .b(_14461_),
    .c(net631),
    .o1(_14462_));
 b15norp02ar1n02x5 _23242_ (.a(_12551_),
    .b(_12751_),
    .o1(_14463_));
 b15oai012al1n03x5 _23243_ (.a(_14463_),
    .b(_13761_),
    .c(_13548_),
    .o1(_14464_));
 b15oai112al1n02x5 _23244_ (.a(net641),
    .b(_13628_),
    .c(_13644_),
    .d(_12545_),
    .o1(_14465_));
 b15nona23aq1n05x5 _23245_ (.a(_14458_),
    .b(_14462_),
    .c(_14464_),
    .d(_14465_),
    .out0(_14466_));
 b15norp02ar1n02x5 _23246_ (.a(_12545_),
    .b(_13644_),
    .o1(_14467_));
 b15aoai13al1n03x5 _23247_ (.a(_14467_),
    .b(_13683_),
    .c(_12718_),
    .d(_13711_),
    .o1(_14468_));
 b15norp03ar1n02x5 _23248_ (.a(_13580_),
    .b(_12615_),
    .c(_12677_),
    .o1(_14469_));
 b15aoi012aq1n02x5 _23249_ (.a(_14469_),
    .b(_13723_),
    .c(_12718_),
    .o1(_14470_));
 b15oa0022ar1n04x5 _23250_ (.a(_12566_),
    .b(_13568_),
    .c(_13560_),
    .d(_12594_),
    .o(_14471_));
 b15norp02an1n24x5 _23251_ (.a(_12766_),
    .b(_12552_),
    .o1(_14472_));
 b15norp02ar1n08x5 _23252_ (.a(_12545_),
    .b(_12771_),
    .o1(_14473_));
 b15nandp2ar1n08x5 _23253_ (.a(_13733_),
    .b(_13547_),
    .o1(_14474_));
 b15and003aq1n04x5 _23254_ (.a(_12662_),
    .b(_12593_),
    .c(_12641_),
    .o(_14475_));
 b15aoi222ah1n06x5 _23255_ (.a(_14472_),
    .b(_13564_),
    .c(_14473_),
    .d(_14474_),
    .e(_14475_),
    .f(net633),
    .o1(_14476_));
 b15nand04ah1n08x5 _23256_ (.a(_14468_),
    .b(_14470_),
    .c(_14471_),
    .d(_14476_),
    .o1(_14477_));
 b15aoai13ar1n02x5 _23257_ (.a(_12685_),
    .b(net642),
    .c(net632),
    .d(_12554_),
    .o1(_14478_));
 b15nor002ah1n04x5 _23258_ (.a(net635),
    .b(_13570_),
    .o1(_14479_));
 b15nano23ar1n02x5 _23259_ (.a(net632),
    .b(_12725_),
    .c(_14479_),
    .d(_12619_),
    .out0(_14480_));
 b15oai022ar1n02x5 _23260_ (.a(_13753_),
    .b(_12750_),
    .c(_12754_),
    .d(_12677_),
    .o1(_14481_));
 b15oab012ar1n02x5 _23261_ (.a(_14478_),
    .b(_14480_),
    .c(_14481_),
    .out0(_14482_));
 b15aoai13aq1n06x5 _23262_ (.a(net637),
    .b(_12643_),
    .c(_13567_),
    .d(net641),
    .o1(_14483_));
 b15aoai13ah1n04x5 _23263_ (.a(net630),
    .b(_12613_),
    .c(_12726_),
    .d(_12581_),
    .o1(_14484_));
 b15oai112ah1n16x5 _23264_ (.a(_14483_),
    .b(_14484_),
    .c(net630),
    .d(_13683_),
    .o1(_14485_));
 b15oai022ar1n02x5 _23265_ (.a(net639),
    .b(_14453_),
    .c(_13762_),
    .d(net642),
    .o1(_14486_));
 b15and003an1n02x5 _23266_ (.a(\us03.a[3] ),
    .b(_13717_),
    .c(_14486_),
    .o(_14487_));
 b15norp02al1n04x5 _23267_ (.a(_12629_),
    .b(_13619_),
    .o1(_14488_));
 b15nanb02ar1n06x5 _23268_ (.a(net627),
    .b(\us03.a[7] ),
    .out0(_14489_));
 b15oai012as1n06x5 _23269_ (.a(_14489_),
    .b(_13735_),
    .c(_12511_),
    .o1(_14490_));
 b15aoai13al1n08x5 _23270_ (.a(_12515_),
    .b(_14487_),
    .c(_14488_),
    .d(_14490_),
    .o1(_14491_));
 b15nona23an1n05x5 _23271_ (.a(_14477_),
    .b(_14482_),
    .c(_14485_),
    .d(_14491_),
    .out0(_14492_));
 b15nor004as1n12x5 _23272_ (.a(_14448_),
    .b(_14456_),
    .c(_14466_),
    .d(_14492_),
    .o1(_14493_));
 b15qgbxo2an1n05x5 _23273_ (.a(_13768_),
    .b(_14493_),
    .out0(_14494_));
 b15xor002as1n06x5 _23274_ (.a(_14424_),
    .b(_14494_),
    .out0(_14495_));
 b15xnr002as1n12x5 _23275_ (.a(_14338_),
    .b(_14495_),
    .out0(_14496_));
 b15oai012ah1n16x5 _23276_ (.a(_14142_),
    .b(_14496_),
    .c(net533),
    .o1(_14497_));
 b15xor002ar1n03x5 _23277_ (.a(_09892_),
    .b(_14497_),
    .out0(_00123_));
 b15nanb02ar1n02x5 _23278_ (.a(\text_in_r[3] ),
    .b(net537),
    .out0(_14498_));
 b15nonb02an1n08x5 _23279_ (.a(net653),
    .b(net647),
    .out0(_14499_));
 b15nandp3ar1n02x5 _23280_ (.a(_13945_),
    .b(_13985_),
    .c(_14499_),
    .o1(_14500_));
 b15oaoi13as1n02x5 _23281_ (.a(net666),
    .b(_14500_),
    .c(_13390_),
    .d(_13313_),
    .o1(_14501_));
 b15nand04ar1n03x5 _23282_ (.a(net666),
    .b(_13506_),
    .c(_13382_),
    .d(_13362_),
    .o1(_14502_));
 b15oai112ah1n02x5 _23283_ (.a(net664),
    .b(_14502_),
    .c(_13977_),
    .d(_13927_),
    .o1(_14503_));
 b15oaoi13al1n02x5 _23284_ (.a(_13315_),
    .b(_13350_),
    .c(_13347_),
    .d(_13318_),
    .o1(_14504_));
 b15oai022ah1n04x5 _23285_ (.a(_14501_),
    .b(_14503_),
    .c(_14504_),
    .d(net664),
    .o1(_14505_));
 b15nor003al1n12x5 _23286_ (.a(net655),
    .b(_13315_),
    .c(_13350_),
    .o1(_14506_));
 b15norp03al1n02x5 _23287_ (.a(_13355_),
    .b(_13313_),
    .c(_13336_),
    .o1(_14507_));
 b15oai012al1n03x5 _23288_ (.a(net659),
    .b(_14506_),
    .c(_14507_),
    .o1(_14508_));
 b15nanb02as1n16x5 _23289_ (.a(net647),
    .b(net654),
    .out0(_14509_));
 b15mdn022an1n06x5 _23290_ (.a(_14416_),
    .b(_14509_),
    .o1(_14510_),
    .sa(_13355_));
 b15nor002ar1n12x5 _23291_ (.a(net650),
    .b(net644),
    .o1(_14511_));
 b15aoai13as1n03x5 _23292_ (.a(_13380_),
    .b(_13928_),
    .c(_14510_),
    .d(_14511_),
    .o1(_14512_));
 b15oai012ah1n03x5 _23293_ (.a(_13479_),
    .b(_13343_),
    .c(net653),
    .o1(_14513_));
 b15aoi022ar1n12x5 _23294_ (.a(_13375_),
    .b(_13481_),
    .c(_14513_),
    .d(net668),
    .o1(_14514_));
 b15nand02al1n04x5 _23295_ (.a(net649),
    .b(_13410_),
    .o1(_14515_));
 b15oai022an1n12x5 _23296_ (.a(net660),
    .b(_14512_),
    .c(_14514_),
    .d(_14515_),
    .o1(_14516_));
 b15nor003ah1n04x5 _23297_ (.a(net659),
    .b(_13315_),
    .c(_13350_),
    .o1(_14517_));
 b15aoai13aq1n02x5 _23298_ (.a(net655),
    .b(_14517_),
    .c(_13999_),
    .d(_13418_),
    .o1(_14518_));
 b15nor002ar1n02x5 _23299_ (.a(_13431_),
    .b(_13967_),
    .o1(_14519_));
 b15nand02ar1n02x5 _23300_ (.a(net656),
    .b(net652),
    .o1(_14520_));
 b15oai012ar1n04x5 _23301_ (.a(_14520_),
    .b(_13350_),
    .c(net656),
    .o1(_14521_));
 b15nor002as1n03x5 _23302_ (.a(_13421_),
    .b(net643),
    .o1(_14522_));
 b15aoi012aq1n04x5 _23303_ (.a(_14519_),
    .b(_14521_),
    .c(_14522_),
    .o1(_14523_));
 b15oai013as1n06x5 _23304_ (.a(_14518_),
    .b(_14523_),
    .c(_13459_),
    .d(_13423_),
    .o1(_14524_));
 b15nano23aq1n08x5 _23305_ (.a(_14505_),
    .b(_14508_),
    .c(_14516_),
    .d(_14524_),
    .out0(_14525_));
 b15nand02ar1n02x5 _23306_ (.a(_13313_),
    .b(_13415_),
    .o1(_14526_));
 b15aob012ah1n04x5 _23307_ (.a(_13371_),
    .b(_13487_),
    .c(_14526_),
    .out0(_14527_));
 b15nand03an1n06x5 _23308_ (.a(_13425_),
    .b(_13410_),
    .c(_13486_),
    .o1(_14528_));
 b15nand04aq1n08x5 _23309_ (.a(_13906_),
    .b(_13908_),
    .c(_14527_),
    .d(_14528_),
    .o1(_14529_));
 b15norp03aq1n02x5 _23310_ (.a(net652),
    .b(net646),
    .c(_13399_),
    .o1(_14530_));
 b15aobi12ar1n02x5 _23311_ (.a(net649),
    .b(net652),
    .c(net666),
    .out0(_14531_));
 b15oaoi13an1n02x5 _23312_ (.a(_13459_),
    .b(_13324_),
    .c(_14531_),
    .d(net660),
    .o1(_14532_));
 b15oai112an1n06x5 _23313_ (.a(net643),
    .b(_13916_),
    .c(_14530_),
    .d(_14532_),
    .o1(_14533_));
 b15norp03an1n02x5 _23314_ (.a(_13313_),
    .b(_13425_),
    .c(_13494_),
    .o1(_14534_));
 b15aoi012an1n04x5 _23315_ (.a(_14534_),
    .b(_13403_),
    .c(_13928_),
    .o1(_14535_));
 b15norp03as1n02x5 _23316_ (.a(_13459_),
    .b(_13306_),
    .c(_13511_),
    .o1(_14536_));
 b15nor003ah1n02x5 _23317_ (.a(net649),
    .b(_13392_),
    .c(_14509_),
    .o1(_14537_));
 b15oai012al1n06x5 _23318_ (.a(net643),
    .b(_14536_),
    .c(_14537_),
    .o1(_14538_));
 b15aoai13as1n08x5 _23319_ (.a(_14533_),
    .b(_13421_),
    .c(_14535_),
    .d(_14538_),
    .o1(_14539_));
 b15nor002ah1n02x5 _23320_ (.a(_13425_),
    .b(_13942_),
    .o1(_14540_));
 b15bfn001as1n48x5 load_slew408 (.a(net409),
    .o(net408));
 b15aoai13aq1n08x5 _23322_ (.a(_13362_),
    .b(_14540_),
    .c(_13340_),
    .d(_14000_),
    .o1(_14542_));
 b15nano22ah1n06x5 _23323_ (.a(net649),
    .b(net644),
    .c(net646),
    .out0(_14543_));
 b15nano23al1n02x5 _23324_ (.a(net659),
    .b(_14543_),
    .c(net653),
    .d(_13392_),
    .out0(_14544_));
 b15norp03ar1n02x5 _23325_ (.a(_13302_),
    .b(_13306_),
    .c(_13447_),
    .o1(_14545_));
 b15oai013as1n02x5 _23326_ (.a(net666),
    .b(_14506_),
    .c(_14544_),
    .d(_14545_),
    .o1(_14546_));
 b15norp03aq1n02x5 _23327_ (.a(net648),
    .b(_13338_),
    .c(_14406_),
    .o1(_14547_));
 b15oai022aq1n02x5 _23328_ (.a(net651),
    .b(_13343_),
    .c(_14406_),
    .d(net648),
    .o1(_14548_));
 b15aoai13as1n04x5 _23329_ (.a(_13374_),
    .b(_14547_),
    .c(_14548_),
    .d(_13945_),
    .o1(_14549_));
 b15aoi022aq1n02x5 _23330_ (.a(_13924_),
    .b(_13905_),
    .c(_13982_),
    .d(_13928_),
    .o1(_14550_));
 b15nand04an1n08x5 _23331_ (.a(_14542_),
    .b(_14546_),
    .c(_14549_),
    .d(_14550_),
    .o1(_14551_));
 b15nandp3ar1n02x5 _23332_ (.a(net653),
    .b(_13905_),
    .c(_14543_),
    .o1(_14552_));
 b15oai012aq1n04x5 _23333_ (.a(_14552_),
    .b(_13953_),
    .c(_13519_),
    .o1(_14553_));
 b15nandp3ar1n02x5 _23334_ (.a(_13421_),
    .b(_13415_),
    .c(_13380_),
    .o1(_14554_));
 b15oaoi13an1n02x5 _23335_ (.a(_13355_),
    .b(_14554_),
    .c(_13494_),
    .d(_13347_),
    .o1(_14555_));
 b15xor002an1n03x5 _23336_ (.a(net657),
    .b(net653),
    .out0(_14556_));
 b15nor004al1n08x5 _23337_ (.a(net651),
    .b(_13441_),
    .c(_13949_),
    .d(_14556_),
    .o1(_14557_));
 b15norp03ar1n02x5 _23338_ (.a(_13479_),
    .b(_13504_),
    .c(_13967_),
    .o1(_14558_));
 b15oai012aq1n02x5 _23339_ (.a(net663),
    .b(_14557_),
    .c(_14558_),
    .o1(_14559_));
 b15nona23as1n24x5 _23340_ (.a(net649),
    .b(net652),
    .c(net643),
    .d(net646),
    .out0(_14560_));
 b15aoi012aq1n04x5 _23341_ (.a(_14560_),
    .b(_13941_),
    .c(_13423_),
    .o1(_14561_));
 b15nor004an1n06x5 _23342_ (.a(net663),
    .b(net660),
    .c(_13318_),
    .d(_13441_),
    .o1(_14562_));
 b15oai012ar1n16x5 _23343_ (.a(net655),
    .b(_14561_),
    .c(_14562_),
    .o1(_14563_));
 b15nona23al1n05x5 _23344_ (.a(_14553_),
    .b(_14555_),
    .c(_14559_),
    .d(_14563_),
    .out0(_14564_));
 b15nor004as1n08x5 _23345_ (.a(_14529_),
    .b(_14539_),
    .c(_14551_),
    .d(_14564_),
    .o1(_14565_));
 b15obai22ar1n02x5 _23346_ (.a(_13367_),
    .b(_13330_),
    .c(_14388_),
    .d(_13942_),
    .out0(_14566_));
 b15aoi012al1n02x5 _23347_ (.a(net655),
    .b(_14566_),
    .c(_13340_),
    .o1(_14567_));
 b15xnr002as1n04x5 _23348_ (.a(net662),
    .b(net643),
    .out0(_14568_));
 b15oai013as1n08x5 _23349_ (.a(net658),
    .b(_13398_),
    .c(_14509_),
    .d(_14568_),
    .o1(_14569_));
 b15nor004an1n06x5 _23350_ (.a(net660),
    .b(_13423_),
    .c(_13306_),
    .d(_13343_),
    .o1(_14570_));
 b15mdn022an1n06x5 _23351_ (.a(_14388_),
    .b(_13977_),
    .o1(_14571_),
    .sa(net664));
 b15aoi112ah1n08x5 _23352_ (.a(_14569_),
    .b(_14570_),
    .c(_14571_),
    .d(_13361_),
    .o1(_14572_));
 b15nor002al1n06x5 _23353_ (.a(net666),
    .b(_13343_),
    .o1(_14573_));
 b15aoi012ar1n02x5 _23354_ (.a(_13941_),
    .b(_13306_),
    .c(_13324_),
    .o1(_14574_));
 b15aoai13aq1n02x5 _23355_ (.a(_14573_),
    .b(_14574_),
    .c(_13388_),
    .d(_13965_),
    .o1(_14575_));
 b15aoi012al1n04x5 _23356_ (.a(_14567_),
    .b(_14572_),
    .c(_14575_),
    .o1(_14576_));
 b15nor004ah1n04x5 _23357_ (.a(net646),
    .b(_13431_),
    .c(_13392_),
    .d(_13399_),
    .o1(_14577_));
 b15nand04as1n12x5 _23358_ (.a(net656),
    .b(_13421_),
    .c(_13505_),
    .d(_13506_),
    .o1(_14578_));
 b15oaoi13as1n02x5 _23359_ (.a(_13340_),
    .b(_14578_),
    .c(_13347_),
    .d(_13330_),
    .o1(_14579_));
 b15nor003ah1n06x5 _23360_ (.a(net666),
    .b(_14577_),
    .c(_14579_),
    .o1(_14580_));
 b15oai012ar1n02x5 _23361_ (.a(_13390_),
    .b(_13500_),
    .c(net663),
    .o1(_14581_));
 b15aoi022ar1n02x5 _23362_ (.a(_13371_),
    .b(_13496_),
    .c(_14581_),
    .d(net659),
    .o1(_14582_));
 b15oab012al1n02x5 _23363_ (.a(_13355_),
    .b(_14572_),
    .c(_14582_),
    .out0(_14583_));
 b15oab012as1n08x5 _23364_ (.c(_14583_),
    .a(_14576_),
    .b(_14580_),
    .out0(_14584_));
 b15nandp3as1n24x5 _23365_ (.a(_14525_),
    .b(_14565_),
    .c(_14584_),
    .o1(_14585_));
 b15xor002as1n12x5 _23366_ (.a(_14493_),
    .b(_14585_),
    .out0(_14586_));
 b15nonb02ah1n04x5 _23367_ (.a(net907),
    .b(net898),
    .out0(_14587_));
 b15oai012al1n02x5 _23368_ (.a(_14587_),
    .b(_12973_),
    .c(net901),
    .o1(_14588_));
 b15nandp2aq1n05x5 _23369_ (.a(_12874_),
    .b(_12822_),
    .o1(_14589_));
 b15oai012ar1n03x5 _23370_ (.a(_12987_),
    .b(_14589_),
    .c(_13009_),
    .o1(_14590_));
 b15nonb02ah1n12x5 _23371_ (.a(net910),
    .b(net901),
    .out0(_14591_));
 b15norp02an1n12x5 _23372_ (.a(net892),
    .b(net887),
    .o1(_14592_));
 b15nona23aq1n02x5 _23373_ (.a(net890),
    .b(_14591_),
    .c(_14592_),
    .d(net894),
    .out0(_14593_));
 b15nand02an1n02x5 _23374_ (.a(net890),
    .b(_12940_),
    .o1(_14594_));
 b15oai013ah1n04x5 _23375_ (.a(_14593_),
    .b(_14594_),
    .c(_13009_),
    .d(net892),
    .o1(_14595_));
 b15oai012as1n04x5 _23376_ (.a(_14588_),
    .b(_14590_),
    .c(_14595_),
    .o1(_14596_));
 b15nandp2ah1n02x5 _23377_ (.a(net910),
    .b(_13798_),
    .o1(_14597_));
 b15oai012ar1n02x5 _23378_ (.a(_14597_),
    .b(_14144_),
    .c(_13803_),
    .o1(_14598_));
 b15oai022ar1n02x5 _23379_ (.a(_12857_),
    .b(_13797_),
    .c(_13787_),
    .d(_13803_),
    .o1(_14599_));
 b15norp02ar1n04x5 _23380_ (.a(_14598_),
    .b(_14599_),
    .o1(_14600_));
 b15aoi012ah1n06x5 _23381_ (.a(_14596_),
    .b(_14600_),
    .c(net897),
    .o1(_14601_));
 b15nandp3al1n04x5 _23382_ (.a(net898),
    .b(_12883_),
    .c(_12798_),
    .o1(_14602_));
 b15oai112aq1n04x5 _23383_ (.a(_14196_),
    .b(_14602_),
    .c(_12910_),
    .d(_14195_),
    .o1(_14603_));
 b15aoi012aq1n02x5 _23384_ (.a(_13835_),
    .b(_14195_),
    .c(_14196_),
    .o1(_14604_));
 b15aoi013as1n02x5 _23385_ (.a(net911),
    .b(net905),
    .c(_14195_),
    .d(_14196_),
    .o1(_14605_));
 b15oai013as1n06x5 _23386_ (.a(_14603_),
    .b(_14604_),
    .c(_14605_),
    .d(_14162_),
    .o1(_14606_));
 b15oai012ar1n02x5 _23387_ (.a(_13797_),
    .b(_12959_),
    .c(_13809_),
    .o1(_14607_));
 b15oaoi13ar1n02x5 _23388_ (.a(net899),
    .b(_14607_),
    .c(_13769_),
    .d(_12879_),
    .o1(_14608_));
 b15aoai13ah1n08x5 _23389_ (.a(_14211_),
    .b(_12912_),
    .c(_13794_),
    .d(net913),
    .o1(_14609_));
 b15nanb02aq1n12x5 _23390_ (.a(net890),
    .b(net892),
    .out0(_14610_));
 b15oai012an1n02x5 _23391_ (.a(_14609_),
    .b(_14144_),
    .c(_14610_),
    .o1(_14611_));
 b15aoi013al1n03x5 _23392_ (.a(_14608_),
    .b(_14611_),
    .c(net899),
    .d(_13884_),
    .o1(_14612_));
 b15aoi012as1n02x5 _23393_ (.a(_12883_),
    .b(_13848_),
    .c(_12832_),
    .o1(_14613_));
 b15norp03aq1n12x5 _23394_ (.a(_12851_),
    .b(_12869_),
    .c(_14613_),
    .o1(_14614_));
 b15aoi012an1n02x5 _23395_ (.a(net905),
    .b(_13809_),
    .c(_14614_),
    .o1(_14615_));
 b15orn002an1n12x5 _23396_ (.a(net894),
    .b(net890),
    .o(_14616_));
 b15norp02ar1n02x5 _23397_ (.a(_12912_),
    .b(_14616_),
    .o1(_14617_));
 b15nanb02aq1n03x5 _23398_ (.a(net902),
    .b(net890),
    .out0(_14618_));
 b15obai22aq1n02x5 _23399_ (.a(_14617_),
    .b(_14591_),
    .c(_14618_),
    .d(_12832_),
    .out0(_14619_));
 b15aoi013ar1n03x5 _23400_ (.a(_14614_),
    .b(_14619_),
    .c(net899),
    .d(_12811_),
    .o1(_14620_));
 b15oai112as1n08x5 _23401_ (.a(_14606_),
    .b(_14612_),
    .c(_14615_),
    .d(_14620_),
    .o1(_14621_));
 b15nandp3ar1n02x5 _23402_ (.a(net908),
    .b(net900),
    .c(_13809_),
    .o1(_14622_));
 b15oai112al1n02x5 _23403_ (.a(_12950_),
    .b(_14622_),
    .c(_13846_),
    .d(net908),
    .o1(_14623_));
 b15oai022an1n02x5 _23404_ (.a(_12960_),
    .b(_13846_),
    .c(_14165_),
    .d(_12954_),
    .o1(_14624_));
 b15oai012as1n04x5 _23405_ (.a(_14623_),
    .b(_14624_),
    .c(_12950_),
    .o1(_14625_));
 b15nonb02ah1n02x5 _23406_ (.a(net913),
    .b(net900),
    .out0(_14626_));
 b15oai012an1n04x5 _23407_ (.a(_14626_),
    .b(_12789_),
    .c(_12825_),
    .o1(_14627_));
 b15nand02ar1n32x5 _23408_ (.a(net904),
    .b(_12851_),
    .o1(_14628_));
 b15oai012al1n04x5 _23409_ (.a(_14627_),
    .b(_12875_),
    .c(_14628_),
    .o1(_14629_));
 b15aoai13al1n08x5 _23410_ (.a(_14233_),
    .b(_13884_),
    .c(_13883_),
    .d(_12950_),
    .o1(_14630_));
 b15qgbna2an1n05x5 _23411_ (.o1(_14631_),
    .a(_12851_),
    .b(_13794_));
 b15oai012ah1n02x5 _23412_ (.a(_14630_),
    .b(_14631_),
    .c(_12885_),
    .o1(_14632_));
 b15aoi022as1n06x5 _23413_ (.a(_12879_),
    .b(_14629_),
    .c(_14632_),
    .d(net911),
    .o1(_14633_));
 b15norp02ah1n02x5 _23414_ (.a(net886),
    .b(_13770_),
    .o1(_14634_));
 b15aoi013ar1n02x5 _23415_ (.a(_14634_),
    .b(_12912_),
    .c(_12822_),
    .d(net886),
    .o1(_14635_));
 b15orn002al1n04x5 _23416_ (.a(_12931_),
    .b(_14635_),
    .o(_14636_));
 b15aoi022an1n06x5 _23417_ (.a(_13826_),
    .b(_14592_),
    .c(_14241_),
    .d(net892),
    .o1(_14637_));
 b15nor003al1n08x5 _23418_ (.a(_14143_),
    .b(_14616_),
    .c(_14637_),
    .o1(_14638_));
 b15nandp2as1n04x5 _23419_ (.a(net892),
    .b(_13883_),
    .o1(_14639_));
 b15aoi112an1n03x5 _23420_ (.a(_12932_),
    .b(_12938_),
    .c(_14639_),
    .d(_12870_),
    .o1(_14640_));
 b15norp03aq1n02x5 _23421_ (.a(_13794_),
    .b(_12875_),
    .c(_12900_),
    .o1(_14641_));
 b15nor003ah1n04x5 _23422_ (.a(_14638_),
    .b(_14640_),
    .c(_14641_),
    .o1(_14642_));
 b15nand04an1n16x5 _23423_ (.a(_14625_),
    .b(_14633_),
    .c(_14636_),
    .d(_14642_),
    .o1(_14643_));
 b15nand03ar1n03x5 _23424_ (.a(_12950_),
    .b(_12825_),
    .c(_12818_),
    .o1(_14644_));
 b15oai022ar1n02x5 _23425_ (.a(_12913_),
    .b(_14610_),
    .c(_14618_),
    .d(net892),
    .o1(_14645_));
 b15aoi022ar1n02x5 _23426_ (.a(_12913_),
    .b(_12959_),
    .c(_12940_),
    .d(_14645_),
    .o1(_14646_));
 b15oai012al1n03x5 _23427_ (.a(_14644_),
    .b(_14646_),
    .c(_14184_),
    .o1(_14647_));
 b15nandp2aq1n02x5 _23428_ (.a(net911),
    .b(_13809_),
    .o1(_14648_));
 b15nor002aq1n06x5 _23429_ (.a(net890),
    .b(_12904_),
    .o1(_14649_));
 b15nor002as1n04x5 _23430_ (.a(_13771_),
    .b(_13801_),
    .o1(_14650_));
 b15aoi022as1n06x5 _23431_ (.a(_14592_),
    .b(_14649_),
    .c(_14650_),
    .d(net887),
    .o1(_14651_));
 b15oaoi13ah1n08x5 _23432_ (.a(_14628_),
    .b(_14648_),
    .c(_14651_),
    .d(net894),
    .o1(_14652_));
 b15nand02ah1n04x5 _23433_ (.a(_12820_),
    .b(_12877_),
    .o1(_14653_));
 b15oai022as1n06x5 _23434_ (.a(_14653_),
    .b(_13007_),
    .c(_13822_),
    .d(_13803_),
    .o1(_14654_));
 b15nandp3al1n03x5 _23435_ (.a(net901),
    .b(_12796_),
    .c(_12874_),
    .o1(_14655_));
 b15nand03an1n03x5 _23436_ (.a(_12881_),
    .b(_12883_),
    .c(_14591_),
    .o1(_14656_));
 b15aoai13as1n04x5 _23437_ (.a(net905),
    .b(_12851_),
    .c(_14655_),
    .d(_14656_),
    .o1(_14657_));
 b15aoi012aq1n08x5 _23438_ (.a(net905),
    .b(_13798_),
    .c(_12908_),
    .o1(_14658_));
 b15nand04ar1n12x5 _23439_ (.a(_12950_),
    .b(_12851_),
    .c(_12916_),
    .d(_12874_),
    .o1(_14659_));
 b15oai112an1n12x5 _23440_ (.a(_14658_),
    .b(_14659_),
    .c(_12950_),
    .d(_14181_),
    .o1(_14660_));
 b15aoi022ar1n16x5 _23441_ (.a(_12851_),
    .b(_14654_),
    .c(_14657_),
    .d(_14660_),
    .o1(_14661_));
 b15aoi012aq1n02x5 _23442_ (.a(_12990_),
    .b(_12960_),
    .c(net910),
    .o1(_14662_));
 b15oai122ah1n08x5 _23443_ (.a(_12820_),
    .b(_13843_),
    .c(_14187_),
    .d(_14662_),
    .e(_13007_),
    .o1(_14663_));
 b15oai012al1n02x5 _23444_ (.a(net902),
    .b(_13843_),
    .c(_12993_),
    .o1(_14664_));
 b15nand03al1n08x5 _23445_ (.a(_12864_),
    .b(_12822_),
    .c(_14626_),
    .o1(_14665_));
 b15nanb02ar1n02x5 _23446_ (.a(net911),
    .b(net899),
    .out0(_14666_));
 b15nand02al1n06x5 _23447_ (.a(net894),
    .b(net890),
    .o1(_14667_));
 b15oa0022ar1n02x5 _23448_ (.a(_14616_),
    .b(_14666_),
    .c(_14667_),
    .d(_14184_),
    .o(_14668_));
 b15oaoi13al1n03x5 _23449_ (.a(net887),
    .b(_14665_),
    .c(_14668_),
    .d(net892),
    .o1(_14669_));
 b15oaoi13ar1n03x5 _23450_ (.a(_12782_),
    .b(_14630_),
    .c(_12993_),
    .d(_12950_),
    .o1(_14670_));
 b15oai013aq1n04x5 _23451_ (.a(_14663_),
    .b(_14664_),
    .c(_14669_),
    .d(_14670_),
    .o1(_14671_));
 b15nona23al1n12x5 _23452_ (.a(_14647_),
    .b(_14652_),
    .c(_14661_),
    .d(_14671_),
    .out0(_14672_));
 b15nor004as1n12x5 _23453_ (.a(_14601_),
    .b(_14621_),
    .c(_14643_),
    .d(_14672_),
    .o1(_14673_));
 b15aoai13al1n02x5 _23454_ (.a(_13067_),
    .b(net785),
    .c(_13129_),
    .d(_13222_),
    .o1(_14674_));
 b15qgbao4an1n05x5 _23455_ (.o1(_14675_),
    .a(_14674_),
    .b(_13227_),
    .c(_14120_),
    .d(net785));
 b15aoi012ar1n02x5 _23456_ (.a(_14077_),
    .b(_13217_),
    .c(_13231_),
    .o1(_14676_));
 b15nand02al1n03x5 _23457_ (.a(net787),
    .b(_14075_),
    .o1(_14677_));
 b15nanb02al1n06x5 _23458_ (.a(net790),
    .b(net778),
    .out0(_14678_));
 b15aoai13an1n02x5 _23459_ (.a(_14285_),
    .b(_13062_),
    .c(_14107_),
    .d(_14678_),
    .o1(_14679_));
 b15oai022ar1n02x5 _23460_ (.a(_14676_),
    .b(_14677_),
    .c(_14679_),
    .d(net787),
    .o1(_14680_));
 b15oai012aq1n02x5 _23461_ (.a(net787),
    .b(_13100_),
    .c(_14030_),
    .o1(_14681_));
 b15nand04ar1n02x5 _23462_ (.a(net790),
    .b(_13092_),
    .c(_13091_),
    .d(_13033_),
    .o1(_14682_));
 b15nanb02al1n02x5 _23463_ (.a(net778),
    .b(net790),
    .out0(_14683_));
 b15nand04aq1n03x5 _23464_ (.a(_13057_),
    .b(_14107_),
    .c(_14678_),
    .d(_14683_),
    .o1(_14684_));
 b15nandp3ar1n02x5 _23465_ (.a(_14681_),
    .b(_14682_),
    .c(_14684_),
    .o1(_14685_));
 b15oai013aq1n02x5 _23466_ (.a(net780),
    .b(_14675_),
    .c(_14680_),
    .d(_14685_),
    .o1(_14686_));
 b15nandp2an1n04x5 _23467_ (.a(net778),
    .b(net768),
    .o1(_14687_));
 b15oai013ah1n02x5 _23468_ (.a(net774),
    .b(_13156_),
    .c(_13211_),
    .d(_14687_),
    .o1(_14688_));
 b15nand04ar1n03x5 _23469_ (.a(net771),
    .b(net790),
    .c(_13219_),
    .d(_13267_),
    .o1(_14689_));
 b15nano22ar1n02x5 _23470_ (.a(net778),
    .b(net768),
    .c(net780),
    .out0(_14690_));
 b15nonb02an1n02x5 _23471_ (.a(net780),
    .b(net778),
    .out0(_14691_));
 b15oaoi13aq1n02x5 _23472_ (.a(_14690_),
    .b(_14691_),
    .c(net768),
    .d(net795),
    .o1(_14692_));
 b15oai013as1n02x5 _23473_ (.a(_14689_),
    .b(_14692_),
    .c(_14029_),
    .d(net771),
    .o1(_14693_));
 b15oai012ar1n03x5 _23474_ (.a(_14688_),
    .b(_14693_),
    .c(net774),
    .o1(_14694_));
 b15nano22ah1n05x5 _23475_ (.a(net775),
    .b(net787),
    .c(net768),
    .out0(_14695_));
 b15aoi022an1n04x5 _23476_ (.a(_13114_),
    .b(_13104_),
    .c(_14695_),
    .d(net780),
    .o1(_14696_));
 b15nor003aq1n02x5 _23477_ (.a(net778),
    .b(_13291_),
    .c(_14696_),
    .o1(_14697_));
 b15nanb02al1n02x5 _23478_ (.a(net768),
    .b(net787),
    .out0(_14698_));
 b15oa0022ar1n02x5 _23479_ (.a(_14256_),
    .b(_14085_),
    .c(_14698_),
    .d(net780),
    .o(_14699_));
 b15nand02ar1n02x5 _23480_ (.a(net790),
    .b(_14124_),
    .o1(_14700_));
 b15oai022ar1n02x5 _23481_ (.a(net790),
    .b(_13125_),
    .c(_14699_),
    .d(_14700_),
    .o1(_14701_));
 b15nona23al1n24x5 _23482_ (.a(net777),
    .b(net773),
    .c(net769),
    .d(net776),
    .out0(_14702_));
 b15oai022as1n08x5 _23483_ (.a(_14053_),
    .b(_13185_),
    .c(_14702_),
    .d(_14095_),
    .o1(_14703_));
 b15oai013ar1n02x5 _23484_ (.a(net794),
    .b(_14697_),
    .c(_14701_),
    .d(_14703_),
    .o1(_14704_));
 b15and003ah1n03x5 _23485_ (.a(_14686_),
    .b(_14694_),
    .c(_14704_),
    .o(_14705_));
 b15aoi012ah1n02x5 _23486_ (.a(_14115_),
    .b(_13161_),
    .c(_13130_),
    .o1(_14706_));
 b15oai013an1n04x5 _23487_ (.a(_14081_),
    .b(_13211_),
    .c(_14296_),
    .d(net790),
    .o1(_14707_));
 b15nand02aq1n08x5 _23488_ (.a(net774),
    .b(net783),
    .o1(_14708_));
 b15oai022ar1n02x5 _23489_ (.a(net774),
    .b(_14025_),
    .c(_14708_),
    .d(_13045_),
    .o1(_14709_));
 b15and003an1n02x5 _23490_ (.a(net777),
    .b(_14281_),
    .c(_14709_),
    .o(_14710_));
 b15xor002as1n08x5 _23491_ (.a(net793),
    .b(net786),
    .out0(_14711_));
 b15nor002aq1n03x5 _23492_ (.a(_13067_),
    .b(_14711_),
    .o1(_14712_));
 b15oab012ar1n03x5 _23493_ (.a(_13184_),
    .b(_13194_),
    .c(_14090_),
    .out0(_14713_));
 b15nor004ar1n08x5 _23494_ (.a(net783),
    .b(_14025_),
    .c(_14712_),
    .d(_14713_),
    .o1(_14714_));
 b15nor004an1n08x5 _23495_ (.a(_14706_),
    .b(_14707_),
    .c(_14710_),
    .d(_14714_),
    .o1(_14715_));
 b15nandp3ar1n02x5 _23496_ (.a(net774),
    .b(net790),
    .c(_13244_),
    .o1(_14716_));
 b15oaoi13as1n02x5 _23497_ (.a(_14716_),
    .b(_14266_),
    .c(_13238_),
    .d(_13291_),
    .o1(_14717_));
 b15nandp2ah1n03x5 _23498_ (.a(_14254_),
    .b(_14020_),
    .o1(_14718_));
 b15oai012an1n06x5 _23499_ (.a(_14718_),
    .b(_13291_),
    .c(_13066_),
    .o1(_14719_));
 b15aoi013an1n02x5 _23500_ (.a(_14717_),
    .b(_14719_),
    .c(_14131_),
    .d(net783),
    .o1(_14720_));
 b15norp02as1n03x5 _23501_ (.a(net774),
    .b(net771),
    .o1(_14721_));
 b15norp03aq1n02x5 _23502_ (.a(net778),
    .b(net768),
    .c(net790),
    .o1(_14722_));
 b15oai112an1n06x5 _23503_ (.a(_13267_),
    .b(_14721_),
    .c(_14722_),
    .d(_13219_),
    .o1(_14723_));
 b15oai013ah1n02x5 _23504_ (.a(_14723_),
    .b(_13277_),
    .c(_13127_),
    .d(_14034_),
    .o1(_14724_));
 b15norp02an1n12x5 _23505_ (.a(_13022_),
    .b(_13141_),
    .o1(_14725_));
 b15oai012aq1n06x5 _23506_ (.a(_13053_),
    .b(_13078_),
    .c(_13063_),
    .o1(_14726_));
 b15nor002aq1n03x5 _23507_ (.a(_14025_),
    .b(_14115_),
    .o1(_14727_));
 b15nona22an1n02x5 _23508_ (.a(net774),
    .b(net794),
    .c(net780),
    .out0(_14728_));
 b15oai022an1n08x5 _23509_ (.a(net780),
    .b(_13086_),
    .c(_14266_),
    .d(_14728_),
    .o1(_14729_));
 b15aoi222as1n12x5 _23510_ (.a(_14313_),
    .b(_14725_),
    .c(_14726_),
    .d(_14727_),
    .e(_14729_),
    .f(_14035_),
    .o1(_14730_));
 b15nor002an1n04x5 _23511_ (.a(_13065_),
    .b(_14270_),
    .o1(_14731_));
 b15nor003al1n08x5 _23512_ (.a(net775),
    .b(net789),
    .c(_13079_),
    .o1(_14732_));
 b15oai112al1n12x5 _23513_ (.a(net790),
    .b(_13263_),
    .c(_14731_),
    .d(_14732_),
    .o1(_14733_));
 b15norp02ah1n02x5 _23514_ (.a(_13063_),
    .b(_13161_),
    .o1(_14734_));
 b15nand02ar1n02x5 _23515_ (.a(net778),
    .b(_13211_),
    .o1(_14735_));
 b15and003ar1n03x5 _23516_ (.a(_13063_),
    .b(_13104_),
    .c(_14117_),
    .o(_14736_));
 b15aoi022ar1n02x5 _23517_ (.a(_13239_),
    .b(_14734_),
    .c(_14735_),
    .d(_14736_),
    .o1(_14737_));
 b15nand03ah1n03x5 _23518_ (.a(_14730_),
    .b(_14733_),
    .c(_14737_),
    .o1(_14738_));
 b15nano23al1n06x5 _23519_ (.a(_14715_),
    .b(_14720_),
    .c(_14724_),
    .d(_14738_),
    .out0(_14739_));
 b15oai012al1n02x5 _23520_ (.a(net794),
    .b(_14035_),
    .c(_13255_),
    .o1(_14740_));
 b15oai012aq1n02x5 _23521_ (.a(_14085_),
    .b(_13211_),
    .c(net790),
    .o1(_14741_));
 b15aoi012an1n04x5 _23522_ (.a(_14740_),
    .b(_14741_),
    .c(_13090_),
    .o1(_14742_));
 b15aoai13as1n06x5 _23523_ (.a(_14128_),
    .b(_14732_),
    .c(_14107_),
    .d(_13286_),
    .o1(_14743_));
 b15norp02ar1n02x5 _23524_ (.a(net775),
    .b(_13079_),
    .o1(_14744_));
 b15oab012ar1n02x5 _23525_ (.a(_14678_),
    .b(_14744_),
    .c(_14731_),
    .out0(_14745_));
 b15oai012aq1n03x5 _23526_ (.a(_14698_),
    .b(_14085_),
    .c(_14256_),
    .o1(_14746_));
 b15aoi013an1n04x5 _23527_ (.a(_14745_),
    .b(_14746_),
    .c(_14124_),
    .d(_13063_),
    .o1(_14747_));
 b15aoi013as1n08x5 _23528_ (.a(_14742_),
    .b(_14743_),
    .c(_14747_),
    .d(_13067_),
    .o1(_14748_));
 b15nanb02ar1n12x5 _23529_ (.a(net790),
    .b(net771),
    .out0(_14749_));
 b15nor002aq1n03x5 _23530_ (.a(net779),
    .b(net784),
    .o1(_14750_));
 b15aoi012ar1n08x5 _23531_ (.a(_14750_),
    .b(_13215_),
    .c(net779),
    .o1(_14751_));
 b15orn003ah1n02x5 _23532_ (.a(_13065_),
    .b(_14749_),
    .c(_14751_),
    .o(_14752_));
 b15norp02aq1n03x5 _23533_ (.a(_13127_),
    .b(_13183_),
    .o1(_14753_));
 b15aoi112ah1n04x5 _23534_ (.a(_13067_),
    .b(_14753_),
    .c(_13046_),
    .d(_13124_),
    .o1(_14754_));
 b15nandp2al1n05x5 _23535_ (.a(net787),
    .b(_13181_),
    .o1(_14755_));
 b15nand04an1n12x5 _23536_ (.a(net782),
    .b(_13185_),
    .c(_14023_),
    .d(_14755_),
    .o1(_14756_));
 b15nonb02aq1n08x5 _23537_ (.a(net790),
    .b(net780),
    .out0(_14757_));
 b15aoi012al1n02x5 _23538_ (.a(_13146_),
    .b(_14120_),
    .c(_14757_),
    .o1(_14758_));
 b15oai012as1n02x5 _23539_ (.a(_13185_),
    .b(_14702_),
    .c(_13114_),
    .o1(_14759_));
 b15oai112as1n06x5 _23540_ (.a(_14756_),
    .b(_14758_),
    .c(net793),
    .d(_14759_),
    .o1(_14760_));
 b15aoi012ar1n04x5 _23541_ (.a(net794),
    .b(_13054_),
    .c(_13251_),
    .o1(_14761_));
 b15aoi022as1n12x5 _23542_ (.a(_14752_),
    .b(_14754_),
    .c(_14760_),
    .d(_14761_),
    .o1(_14762_));
 b15nano23as1n24x5 _23543_ (.a(_14705_),
    .b(_14739_),
    .c(_14748_),
    .d(_14762_),
    .out0(_14763_));
 b15xor002as1n12x5 _23544_ (.a(_14673_),
    .b(_14763_),
    .out0(_14764_));
 b15xor002ah1n08x5 _23545_ (.a(_14586_),
    .b(_14764_),
    .out0(_14765_));
 b15oaoi13ar1n02x5 _23546_ (.a(net640),
    .b(_12589_),
    .c(_12684_),
    .d(net637),
    .o1(_14766_));
 b15norp03aq1n08x5 _23547_ (.a(net633),
    .b(_12553_),
    .c(_12717_),
    .o1(_14767_));
 b15aob012ar1n02x5 _23548_ (.a(_12589_),
    .b(_14767_),
    .c(net640),
    .out0(_14768_));
 b15aoai13ar1n02x5 _23549_ (.a(net632),
    .b(_14766_),
    .c(_14768_),
    .d(net637),
    .o1(_14769_));
 b15inv040aq1n03x5 _23550_ (.a(_14769_),
    .o1(_14770_));
 b15oai022al1n04x5 _23551_ (.a(_12511_),
    .b(_12714_),
    .c(_12684_),
    .d(net632),
    .o1(_14771_));
 b15aoi122ar1n04x5 _23552_ (.a(net636),
    .b(_12736_),
    .c(net632),
    .d(_14771_),
    .e(net637),
    .o1(_14772_));
 b15nand04ar1n03x5 _23553_ (.a(net632),
    .b(_12563_),
    .c(_12564_),
    .d(_12649_),
    .o1(_14773_));
 b15oai013al1n02x5 _23554_ (.a(_14773_),
    .b(_12595_),
    .c(_12623_),
    .d(net632),
    .o1(_14774_));
 b15oai012ah1n02x5 _23555_ (.a(_12704_),
    .b(_12600_),
    .c(_12545_),
    .o1(_14775_));
 b15aoi012ar1n04x5 _23556_ (.a(_14774_),
    .b(_14775_),
    .c(_13565_),
    .o1(_14776_));
 b15oaoi13ah1n02x5 _23557_ (.a(net640),
    .b(_12565_),
    .c(_12760_),
    .d(net637),
    .o1(_14777_));
 b15oai122al1n08x5 _23558_ (.a(_12545_),
    .b(_12524_),
    .c(_12595_),
    .d(_12750_),
    .e(_12511_),
    .o1(_14778_));
 b15oai022al1n06x5 _23559_ (.a(_12545_),
    .b(_13688_),
    .c(_14777_),
    .d(_14778_),
    .o1(_14779_));
 b15aoi013ar1n06x5 _23560_ (.a(_14772_),
    .b(_14776_),
    .c(_14779_),
    .d(net636),
    .o1(_14780_));
 b15norp02ar1n02x5 _23561_ (.a(_12545_),
    .b(_13688_),
    .o1(_14781_));
 b15aoi122ar1n02x5 _23562_ (.a(_13570_),
    .b(_13673_),
    .c(_14781_),
    .d(_13549_),
    .e(_12545_),
    .o1(_14782_));
 b15nand04ar1n02x5 _23563_ (.a(_12545_),
    .b(_12519_),
    .c(_12563_),
    .d(_12657_),
    .o1(_14783_));
 b15oaoi13ar1n03x5 _23564_ (.a(_12643_),
    .b(_14783_),
    .c(_12545_),
    .d(_12619_),
    .o1(_14784_));
 b15oai022ar1n02x5 _23565_ (.a(_12565_),
    .b(_13580_),
    .c(_12760_),
    .d(net633),
    .o1(_14785_));
 b15oaoi13aq1n03x5 _23566_ (.a(_14782_),
    .b(net637),
    .c(_14784_),
    .d(_14785_),
    .o1(_14786_));
 b15oai022al1n02x5 _23567_ (.a(_12600_),
    .b(_12658_),
    .c(_12747_),
    .d(_12524_),
    .o1(_14787_));
 b15aob012ar1n03x5 _23568_ (.a(net637),
    .b(_14472_),
    .c(_13589_),
    .out0(_14788_));
 b15nand02ar1n02x5 _23569_ (.a(net640),
    .b(_12707_),
    .o1(_14789_));
 b15oai022ar1n04x5 _23570_ (.a(_12747_),
    .b(_12762_),
    .c(_14789_),
    .d(_12677_),
    .o1(_14790_));
 b15oai022aq1n06x5 _23571_ (.a(net637),
    .b(_14787_),
    .c(_14788_),
    .d(_14790_),
    .o1(_14791_));
 b15nand03an1n02x5 _23572_ (.a(net633),
    .b(_12554_),
    .c(_12603_),
    .o1(_14792_));
 b15aoai13an1n04x5 _23573_ (.a(_13547_),
    .b(_13628_),
    .c(_12554_),
    .d(_13686_),
    .o1(_14793_));
 b15oaoi13al1n04x5 _23574_ (.a(net630),
    .b(_14792_),
    .c(_14793_),
    .d(_12511_),
    .o1(_14794_));
 b15nano23as1n08x5 _23575_ (.a(_14786_),
    .b(_14791_),
    .c(_14794_),
    .d(_13569_),
    .out0(_14795_));
 b15nandp2al1n08x5 _23576_ (.a(_12720_),
    .b(_13624_),
    .o1(_14796_));
 b15oai112an1n08x5 _23577_ (.a(_13567_),
    .b(_12700_),
    .c(_13548_),
    .d(_13683_),
    .o1(_14797_));
 b15nand02ah1n03x5 _23578_ (.a(_12580_),
    .b(_12725_),
    .o1(_14798_));
 b15oai012as1n03x5 _23579_ (.a(net634),
    .b(net621),
    .c(net638),
    .o1(_14799_));
 b15nor003al1n04x5 _23580_ (.a(net624),
    .b(_13606_),
    .c(_13727_),
    .o1(_14800_));
 b15aoi022an1n12x5 _23581_ (.a(_12724_),
    .b(_14798_),
    .c(_14799_),
    .d(_14800_),
    .o1(_14801_));
 b15nor002ar1n03x5 _23582_ (.a(_12581_),
    .b(_12726_),
    .o1(_14802_));
 b15nand02ar1n02x5 _23583_ (.a(net633),
    .b(net626),
    .o1(_14803_));
 b15oai012an1n04x5 _23584_ (.a(_14803_),
    .b(net626),
    .c(net630),
    .o1(_14804_));
 b15nor003ah1n02x5 _23585_ (.a(_12662_),
    .b(_12717_),
    .c(_12649_),
    .o1(_14805_));
 b15aoi022as1n06x5 _23586_ (.a(_12577_),
    .b(_14802_),
    .c(_14804_),
    .d(_14805_),
    .o1(_14806_));
 b15nand04aq1n16x5 _23587_ (.a(_14796_),
    .b(_14797_),
    .c(_14801_),
    .d(_14806_),
    .o1(_14807_));
 b15aoi012ar1n02x5 _23588_ (.a(_13727_),
    .b(_13673_),
    .c(_13695_),
    .o1(_14808_));
 b15nor004an1n02x5 _23589_ (.a(_12598_),
    .b(_12603_),
    .c(_12613_),
    .d(_12646_),
    .o1(_14809_));
 b15oai222aq1n12x5 _23590_ (.a(_12613_),
    .b(_12747_),
    .c(_12771_),
    .d(_13560_),
    .e(_12751_),
    .f(_12542_),
    .o1(_14810_));
 b15nonb02al1n06x5 _23591_ (.a(\us03.a[3] ),
    .b(net642),
    .out0(_14811_));
 b15nand03ah1n08x5 _23592_ (.a(_12632_),
    .b(_12635_),
    .c(_14811_),
    .o1(_14812_));
 b15nand03an1n02x5 _23593_ (.a(_12707_),
    .b(_12603_),
    .c(_13688_),
    .o1(_14813_));
 b15oai112al1n08x5 _23594_ (.a(_14812_),
    .b(_14813_),
    .c(_12684_),
    .d(_12709_),
    .o1(_14814_));
 b15ornc04aq1n06x5 _23595_ (.a(_14808_),
    .b(_14809_),
    .c(_14810_),
    .d(_14814_),
    .o(_14815_));
 b15oab012al1n02x5 _23596_ (.a(_13758_),
    .b(_13551_),
    .c(net642),
    .out0(_14816_));
 b15oai012ar1n02x5 _23597_ (.a(_12584_),
    .b(_13700_),
    .c(net637),
    .o1(_14817_));
 b15aoi022al1n04x5 _23598_ (.a(_13700_),
    .b(_13548_),
    .c(_14817_),
    .d(_14472_),
    .o1(_14818_));
 b15oai022aq1n08x5 _23599_ (.a(_12629_),
    .b(_14816_),
    .c(_14818_),
    .d(net633),
    .o1(_14819_));
 b15aoai13ar1n02x5 _23600_ (.a(_12581_),
    .b(net640),
    .c(_12515_),
    .d(_12524_),
    .o1(_14820_));
 b15aoi012ar1n02x5 _23601_ (.a(_12515_),
    .b(_13712_),
    .c(_12615_),
    .o1(_14821_));
 b15aoi112al1n02x5 _23602_ (.a(net632),
    .b(_14821_),
    .c(_12524_),
    .d(_12566_),
    .o1(_14822_));
 b15oai112an1n08x5 _23603_ (.a(_12714_),
    .b(_13710_),
    .c(_12685_),
    .d(_12565_),
    .o1(_14823_));
 b15ao0022aq1n06x5 _23604_ (.a(_14820_),
    .b(_14822_),
    .c(_14823_),
    .d(net632),
    .o(_14824_));
 b15nor004as1n12x5 _23605_ (.a(_14807_),
    .b(_14815_),
    .c(_14819_),
    .d(_14824_),
    .o1(_14825_));
 b15nona23as1n32x5 _23606_ (.a(_14770_),
    .b(_14780_),
    .c(_14795_),
    .d(_14825_),
    .out0(_14826_));
 b15xor002aq1n12x5 _23607_ (.a(_13664_),
    .b(_14826_),
    .out0(_14827_));
 b15xor002as1n16x5 _23608_ (.a(_14765_),
    .b(_14827_),
    .out0(_14828_));
 b15oai012ar1n02x5 _23609_ (.a(_14498_),
    .b(_14828_),
    .c(net537),
    .o1(_14829_));
 b15xor002ar1n02x5 _23610_ (.a(_10038_),
    .b(_14829_),
    .out0(_00124_));
 b15nanb02al1n12x5 _23611_ (.a(\text_in_r[4] ),
    .b(net533),
    .out0(_14830_));
 b15obai22aq1n04x5 _23612_ (.a(_14254_),
    .b(_13228_),
    .c(_14749_),
    .d(_13066_),
    .out0(_14831_));
 b15nand03ah1n08x5 _23613_ (.a(_13124_),
    .b(_14131_),
    .c(_14831_),
    .o1(_14832_));
 b15aob012aq1n04x5 _23614_ (.a(_14832_),
    .b(_14306_),
    .c(_14089_),
    .out0(_14833_));
 b15oai022ar1n02x5 _23615_ (.a(_13209_),
    .b(_13210_),
    .c(_13211_),
    .d(_13214_),
    .o1(_14834_));
 b15oaoi13ar1n02x5 _23616_ (.a(net795),
    .b(_13255_),
    .c(_14288_),
    .d(_14067_),
    .o1(_14835_));
 b15aoai13ar1n02x5 _23617_ (.a(_14030_),
    .b(_13244_),
    .c(_13210_),
    .d(net793),
    .o1(_14836_));
 b15aob012ar1n02x5 _23618_ (.a(_13140_),
    .b(_13262_),
    .c(net783),
    .out0(_14837_));
 b15aoi012ar1n02x5 _23619_ (.a(_14836_),
    .b(_14837_),
    .c(_13067_),
    .o1(_14838_));
 b15orn003an1n03x5 _23620_ (.a(_14834_),
    .b(_14835_),
    .c(_14838_),
    .o(_14839_));
 b15nandp3aq1n03x5 _23621_ (.a(_13092_),
    .b(_13208_),
    .c(_13267_),
    .o1(_14840_));
 b15oai013an1n12x5 _23622_ (.a(_14840_),
    .b(_14114_),
    .c(_13252_),
    .d(_14085_),
    .o1(_14841_));
 b15aoi012ar1n02x5 _23623_ (.a(_14085_),
    .b(_13067_),
    .c(net774),
    .o1(_14842_));
 b15nand03ah1n03x5 _23624_ (.a(net773),
    .b(_13237_),
    .c(_14842_),
    .o1(_14843_));
 b15norp02an1n02x5 _23625_ (.a(net795),
    .b(_13022_),
    .o1(_14844_));
 b15oai112al1n08x5 _23626_ (.a(_14104_),
    .b(_14129_),
    .c(_14844_),
    .d(net777),
    .o1(_14845_));
 b15nanb03al1n08x5 _23627_ (.a(_14841_),
    .b(_14843_),
    .c(_14845_),
    .out0(_14846_));
 b15nand03aq1n03x5 _23628_ (.a(_13046_),
    .b(_13040_),
    .c(_13251_),
    .o1(_14847_));
 b15oai013aq1n08x5 _23629_ (.a(_14847_),
    .b(_14711_),
    .c(_13193_),
    .d(_13086_),
    .o1(_14848_));
 b15nor004as1n06x5 _23630_ (.a(_14833_),
    .b(_14839_),
    .c(_14846_),
    .d(_14848_),
    .o1(_14849_));
 b15nandp2as1n03x5 _23631_ (.a(net781),
    .b(_14333_),
    .o1(_14850_));
 b15nor003as1n03x5 _23632_ (.a(\us21.a[4] ),
    .b(net773),
    .c(net792),
    .o1(_14851_));
 b15and003ar1n03x5 _23633_ (.a(_13124_),
    .b(_14107_),
    .c(_14851_),
    .o(_14852_));
 b15nano23an1n08x5 _23634_ (.a(\us21.a[7] ),
    .b(net771),
    .c(net789),
    .d(net775),
    .out0(_14853_));
 b15aoai13ar1n03x5 _23635_ (.a(net778),
    .b(_14853_),
    .c(_13233_),
    .d(_14107_),
    .o1(_14854_));
 b15oai012al1n06x5 _23636_ (.a(_14854_),
    .b(_13185_),
    .c(_13114_),
    .o1(_14855_));
 b15aoai13ah1n08x5 _23637_ (.a(\us21.a[0] ),
    .b(_14852_),
    .c(_14855_),
    .d(net783),
    .o1(_14856_));
 b15ao0022ah1n03x5 _23638_ (.a(_13128_),
    .b(_14281_),
    .c(_14117_),
    .d(_14256_),
    .o(_14857_));
 b15aoi013aq1n06x5 _23639_ (.a(_14061_),
    .b(_14857_),
    .c(_13129_),
    .d(_14317_),
    .o1(_14858_));
 b15mdn022as1n02x5 _23640_ (.a(_14301_),
    .b(_14281_),
    .o1(_14859_),
    .sa(net777));
 b15nor004ah1n04x5 _23641_ (.a(net780),
    .b(_13065_),
    .c(_13156_),
    .d(_14859_),
    .o1(_14860_));
 b15aoi022an1n04x5 _23642_ (.a(_14103_),
    .b(_14075_),
    .c(_14721_),
    .d(_13072_),
    .o1(_14861_));
 b15oab012ah1n06x5 _23643_ (.a(_14860_),
    .b(_14861_),
    .c(_13132_),
    .out0(_14862_));
 b15nandp3ar1n02x5 _23644_ (.a(_13067_),
    .b(_14035_),
    .c(_13171_),
    .o1(_14863_));
 b15aoai13as1n03x5 _23645_ (.a(_14863_),
    .b(_13227_),
    .c(_13095_),
    .d(_14036_),
    .o1(_14864_));
 b15oai022ah1n02x5 _23646_ (.a(_13142_),
    .b(_13193_),
    .c(_14063_),
    .d(_13159_),
    .o1(_14865_));
 b15aoi022as1n08x5 _23647_ (.a(_13022_),
    .b(_14864_),
    .c(_14865_),
    .d(net786),
    .o1(_14866_));
 b15nand04an1n16x5 _23648_ (.a(_14856_),
    .b(_14858_),
    .c(_14862_),
    .d(_14866_),
    .o1(_14867_));
 b15nano22al1n02x5 _23649_ (.a(net770),
    .b(net772),
    .c(\us21.a[0] ),
    .out0(_14868_));
 b15nonb03an1n02x5 _23650_ (.a(net796),
    .b(net772),
    .c(net770),
    .out0(_14869_));
 b15oai112ah1n06x5 _23651_ (.a(net792),
    .b(_13091_),
    .c(_14868_),
    .d(_14869_),
    .o1(_14870_));
 b15oai112ar1n08x5 _23652_ (.a(_13022_),
    .b(_14870_),
    .c(_14296_),
    .d(_14067_),
    .o1(_14871_));
 b15norp02ar1n08x5 _23653_ (.a(net773),
    .b(\us21.a[0] ),
    .o1(_14872_));
 b15nand04an1n06x5 _23654_ (.a(\us21.a[4] ),
    .b(_14035_),
    .c(_14107_),
    .d(_14872_),
    .o1(_14873_));
 b15nor002ah1n12x5 _23655_ (.a(net768),
    .b(net794),
    .o1(_14874_));
 b15aoai13aq1n04x5 _23656_ (.a(_14874_),
    .b(_14851_),
    .c(_13091_),
    .d(_13232_),
    .o1(_14875_));
 b15oai112ar1n16x5 _23657_ (.a(_13091_),
    .b(_13176_),
    .c(_14020_),
    .d(_14313_),
    .o1(_14876_));
 b15aoai13ah1n03x5 _23658_ (.a(_13171_),
    .b(_13050_),
    .c(_14029_),
    .d(\us21.a[0] ),
    .o1(_14877_));
 b15nand04al1n12x5 _23659_ (.a(_14873_),
    .b(_14875_),
    .c(_14876_),
    .d(_14877_),
    .o1(_14878_));
 b15aoi012ar1n02x5 _23660_ (.a(_13022_),
    .b(_14035_),
    .c(_13213_),
    .o1(_14879_));
 b15nor002ar1n02x5 _23661_ (.a(net787),
    .b(_13252_),
    .o1(_14880_));
 b15oai112aq1n08x5 _23662_ (.a(_14755_),
    .b(_14879_),
    .c(_14880_),
    .d(_14034_),
    .o1(_14881_));
 b15aoi022ar1n02x5 _23663_ (.a(net787),
    .b(_13249_),
    .c(_13181_),
    .d(_13063_),
    .o1(_14882_));
 b15nor002aq1n03x5 _23664_ (.a(_13067_),
    .b(_14882_),
    .o1(_14883_));
 b15oai013ar1n12x5 _23665_ (.a(_14871_),
    .b(_14878_),
    .c(_14881_),
    .d(_14883_),
    .o1(_14884_));
 b15xor002ar1n03x5 _23666_ (.a(net768),
    .b(net789),
    .out0(_14885_));
 b15nand03an1n06x5 _23667_ (.a(_14075_),
    .b(_14691_),
    .c(_14885_),
    .o1(_14886_));
 b15aoai13ar1n02x5 _23668_ (.a(_14128_),
    .b(_14853_),
    .c(_14104_),
    .d(_13112_),
    .o1(_14887_));
 b15nandp3ah1n03x5 _23669_ (.a(_13063_),
    .b(_14886_),
    .c(_14887_),
    .o1(_14888_));
 b15nand02ar1n02x5 _23670_ (.a(net780),
    .b(_13104_),
    .o1(_14889_));
 b15aoi012ar1n02x5 _23671_ (.a(_14254_),
    .b(_13057_),
    .c(net778),
    .o1(_14890_));
 b15oai022ah1n04x5 _23672_ (.a(_13086_),
    .b(_14115_),
    .c(_14889_),
    .d(_14890_),
    .o1(_14891_));
 b15oai012an1n12x5 _23673_ (.a(_14888_),
    .b(_14891_),
    .c(_13063_),
    .o1(_14892_));
 b15nand02an1n03x5 _23674_ (.a(net794),
    .b(_14124_),
    .o1(_14893_));
 b15norp03ar1n02x5 _23675_ (.a(net778),
    .b(net771),
    .c(net794),
    .o1(_14894_));
 b15aoai13aq1n03x5 _23676_ (.a(_13240_),
    .b(_14894_),
    .c(_14285_),
    .d(net778),
    .o1(_14895_));
 b15aob012al1n24x5 _23677_ (.a(_13251_),
    .b(_14893_),
    .c(_14895_),
    .out0(_14896_));
 b15oai112as1n16x5 _23678_ (.a(_14884_),
    .b(_14892_),
    .c(_14896_),
    .d(\us21.a[7] ),
    .o1(_14897_));
 b15nano23as1n24x5 _23679_ (.a(_14849_),
    .b(_14850_),
    .c(_14867_),
    .d(_14897_),
    .out0(_14898_));
 b15nona22an1n08x5 _23680_ (.a(net894),
    .b(net887),
    .c(net890),
    .out0(_14899_));
 b15nanb02ar1n12x5 _23681_ (.a(net890),
    .b(net908),
    .out0(_14900_));
 b15nandp2al1n08x5 _23682_ (.a(net894),
    .b(net887),
    .o1(_14901_));
 b15oaoi13an1n04x5 _23683_ (.a(net892),
    .b(_14899_),
    .c(_14900_),
    .d(_14901_),
    .o1(_14902_));
 b15aoai13ah1n08x5 _23684_ (.a(net900),
    .b(_14902_),
    .c(_14649_),
    .d(_13883_),
    .o1(_14903_));
 b15nand02ar1n02x5 _23685_ (.a(net897),
    .b(_13798_),
    .o1(_14904_));
 b15aob012as1n03x5 _23686_ (.a(net905),
    .b(_14659_),
    .c(_14904_),
    .out0(_14905_));
 b15and002ar1n02x5 _23687_ (.a(_14903_),
    .b(_14905_),
    .o(_14906_));
 b15nand03ar1n03x5 _23688_ (.a(net890),
    .b(_12883_),
    .c(_13843_),
    .o1(_14907_));
 b15oai013ah1n03x5 _23689_ (.a(_14907_),
    .b(_12938_),
    .c(_13011_),
    .d(net908),
    .o1(_14908_));
 b15nandp2aq1n08x5 _23690_ (.a(net887),
    .b(_14908_),
    .o1(_14909_));
 b15nandp2ah1n05x5 _23691_ (.a(net910),
    .b(net901),
    .o1(_14910_));
 b15oai112aq1n06x5 _23692_ (.a(_12782_),
    .b(_13769_),
    .c(_14910_),
    .d(_12875_),
    .o1(_14911_));
 b15aoi013ar1n04x5 _23693_ (.a(_13801_),
    .b(_13838_),
    .c(net905),
    .d(_13769_),
    .o1(_14912_));
 b15aoi012aq1n08x5 _23694_ (.a(net897),
    .b(_14911_),
    .c(_14912_),
    .o1(_14913_));
 b15oaoi13ah1n04x5 _23695_ (.a(net901),
    .b(_14906_),
    .c(_14909_),
    .d(_14913_),
    .o1(_14914_));
 b15aoi022an1n02x5 _23696_ (.a(net908),
    .b(_12957_),
    .c(_13809_),
    .d(_13860_),
    .o1(_14915_));
 b15and003ar1n02x5 _23697_ (.a(_12782_),
    .b(_12822_),
    .c(_12998_),
    .o(_14916_));
 b15nonb03ar1n02x5 _23698_ (.a(net890),
    .b(net908),
    .c(net894),
    .out0(_14917_));
 b15oab012ar1n02x5 _23699_ (.a(net892),
    .b(_12998_),
    .c(_14917_),
    .out0(_14918_));
 b15and002ar1n02x5 _23700_ (.a(_12832_),
    .b(_12998_),
    .o(_14919_));
 b15oai122as1n04x5 _23701_ (.a(net887),
    .b(net911),
    .c(_14916_),
    .d(_14918_),
    .e(_14919_),
    .o1(_14920_));
 b15and003aq1n04x5 _23702_ (.a(net899),
    .b(_14915_),
    .c(_14920_),
    .o(_14921_));
 b15nona23as1n12x5 _23703_ (.a(net887),
    .b(_12820_),
    .c(_12796_),
    .d(_14900_),
    .out0(_14922_));
 b15aoi013ar1n02x5 _23704_ (.a(net897),
    .b(_12796_),
    .c(_12848_),
    .d(_12910_),
    .o1(_14923_));
 b15oai112ah1n02x5 _23705_ (.a(_14922_),
    .b(_14923_),
    .c(_14653_),
    .d(_14589_),
    .o1(_14924_));
 b15nand02ar1n02x5 _23706_ (.a(net902),
    .b(_13817_),
    .o1(_14925_));
 b15oaoi13al1n02x5 _23707_ (.a(_13015_),
    .b(_14925_),
    .c(net902),
    .d(_12917_),
    .o1(_14926_));
 b15aoi013al1n04x5 _23708_ (.a(net913),
    .b(net904),
    .c(_12916_),
    .d(_12848_),
    .o1(_14927_));
 b15nandp2al1n04x5 _23709_ (.a(_13794_),
    .b(_13817_),
    .o1(_14928_));
 b15aoi013ah1n08x5 _23710_ (.a(_14927_),
    .b(_14928_),
    .c(net913),
    .d(_13846_),
    .o1(_14929_));
 b15norp03as1n04x5 _23711_ (.a(_14924_),
    .b(_14926_),
    .c(_14929_),
    .o1(_14930_));
 b15aoi022an1n02x5 _23712_ (.a(net902),
    .b(_12916_),
    .c(_12796_),
    .d(_13794_),
    .o1(_14931_));
 b15nand02an1n02x5 _23713_ (.a(net910),
    .b(_12798_),
    .o1(_14932_));
 b15oai222al1n08x5 _23714_ (.a(_12995_),
    .b(_13843_),
    .c(_12913_),
    .d(_12800_),
    .e(_14931_),
    .f(_14932_),
    .o1(_14933_));
 b15norp02al1n04x5 _23715_ (.a(_12851_),
    .b(_14933_),
    .o1(_14934_));
 b15oai022al1n12x5 _23716_ (.a(_14913_),
    .b(_14921_),
    .c(_14930_),
    .d(_14934_),
    .o1(_14935_));
 b15nona23al1n12x5 _23717_ (.a(net896),
    .b(net886),
    .c(net889),
    .d(net893),
    .out0(_14936_));
 b15aoi013al1n02x5 _23718_ (.a(_14936_),
    .b(_14143_),
    .c(_12954_),
    .d(net912),
    .o1(_14937_));
 b15xor002ar1n03x5 _23719_ (.a(net903),
    .b(_12987_),
    .out0(_14938_));
 b15oai012an1n04x5 _23720_ (.a(_14937_),
    .b(_14938_),
    .c(net912),
    .o1(_14939_));
 b15nand03al1n02x5 _23721_ (.a(_12820_),
    .b(_12954_),
    .c(_12960_),
    .o1(_14940_));
 b15oai012al1n03x5 _23722_ (.a(_12950_),
    .b(_12820_),
    .c(_14587_),
    .o1(_14941_));
 b15norp02aq1n08x5 _23723_ (.a(_13770_),
    .b(_13012_),
    .o1(_14942_));
 b15oai112an1n08x5 _23724_ (.a(_14940_),
    .b(_14941_),
    .c(_14942_),
    .d(_12825_),
    .o1(_14943_));
 b15oai022an1n06x5 _23725_ (.a(net898),
    .b(_14942_),
    .c(_12825_),
    .d(_14177_),
    .o1(_14944_));
 b15aoai13as1n08x5 _23726_ (.a(_14939_),
    .b(_14943_),
    .c(_14944_),
    .d(net912),
    .o1(_14945_));
 b15nor002al1n02x5 _23727_ (.a(_14143_),
    .b(_14223_),
    .o1(_14946_));
 b15oai112ah1n02x5 _23728_ (.a(_12851_),
    .b(_12789_),
    .c(_13835_),
    .d(net910),
    .o1(_14947_));
 b15oaoi13al1n04x5 _23729_ (.a(_14946_),
    .b(_14947_),
    .c(_12851_),
    .d(_13803_),
    .o1(_14948_));
 b15oai022ah1n06x5 _23730_ (.a(net910),
    .b(_12857_),
    .c(_12995_),
    .d(_13843_),
    .o1(_14949_));
 b15aoi112as1n08x5 _23731_ (.a(_14945_),
    .b(_14948_),
    .c(_14949_),
    .d(_12863_),
    .o1(_14950_));
 b15nand03ar1n02x5 _23732_ (.a(_12782_),
    .b(_12993_),
    .c(_14234_),
    .o1(_14951_));
 b15oai012al1n02x5 _23733_ (.a(net908),
    .b(net899),
    .c(_13007_),
    .o1(_14952_));
 b15and003ah1n04x5 _23734_ (.a(_12820_),
    .b(_14951_),
    .c(_14952_),
    .o(_14953_));
 b15norp03aq1n03x5 _23735_ (.a(_14152_),
    .b(_13011_),
    .c(_13797_),
    .o1(_14954_));
 b15aoai13al1n06x5 _23736_ (.a(net911),
    .b(_14954_),
    .c(_12957_),
    .d(_12863_),
    .o1(_14955_));
 b15and002an1n02x5 _23737_ (.a(net893),
    .b(net899),
    .o(_14956_));
 b15nona23an1n04x5 _23738_ (.a(_14147_),
    .b(net906),
    .c(_13884_),
    .d(_14956_),
    .out0(_14957_));
 b15norp02al1n02x5 _23739_ (.a(net906),
    .b(_12857_),
    .o1(_14958_));
 b15aoi012al1n04x5 _23740_ (.a(_14958_),
    .b(_12909_),
    .c(net906),
    .o1(_14959_));
 b15oai112ah1n12x5 _23741_ (.a(_14955_),
    .b(_14957_),
    .c(_14959_),
    .d(_12932_),
    .o1(_14960_));
 b15mdn022ar1n02x5 _23742_ (.a(_13883_),
    .b(_13884_),
    .o1(_14961_),
    .sa(_12782_));
 b15oai013ar1n02x5 _23743_ (.a(_12924_),
    .b(_14610_),
    .c(_14961_),
    .d(_12950_),
    .o1(_14962_));
 b15nand03as1n12x5 _23744_ (.a(_12881_),
    .b(_12883_),
    .c(_12877_),
    .o1(_14963_));
 b15aoi012ar1n02x5 _23745_ (.a(_13884_),
    .b(_13883_),
    .c(net906),
    .o1(_14964_));
 b15nand02ar1n02x5 _23746_ (.a(_12983_),
    .b(_14591_),
    .o1(_14965_));
 b15oai122as1n02x5 _23747_ (.a(_14963_),
    .b(_14964_),
    .c(_14965_),
    .d(_13003_),
    .e(_13835_),
    .o1(_14966_));
 b15cmbn22al1n04x5 _23748_ (.clk1(_14962_),
    .clk2(_14966_),
    .clkout(_14967_),
    .s(net899));
 b15norp03ar1n02x5 _23749_ (.a(net886),
    .b(_12931_),
    .c(_12971_),
    .o1(_14968_));
 b15oai012al1n02x5 _23750_ (.a(_12931_),
    .b(_14147_),
    .c(net898),
    .o1(_14969_));
 b15aoi013aq1n03x5 _23751_ (.a(_14968_),
    .b(_14969_),
    .c(net903),
    .d(net886),
    .o1(_14970_));
 b15nor003as1n08x5 _23752_ (.a(_12782_),
    .b(_13770_),
    .c(_14970_),
    .o1(_14971_));
 b15nor004as1n12x5 _23753_ (.a(_14953_),
    .b(_14960_),
    .c(_14967_),
    .d(_14971_),
    .o1(_14972_));
 b15nona23as1n32x5 _23754_ (.a(_14914_),
    .b(_14935_),
    .c(_14950_),
    .d(_14972_),
    .out0(_14973_));
 b15xor002an1n16x5 _23755_ (.a(_14898_),
    .b(_14973_),
    .out0(_14974_));
 b15xnr002ah1n08x5 _23756_ (.a(_13663_),
    .b(_14826_),
    .out0(_14975_));
 b15xor002al1n16x5 _23757_ (.a(_14974_),
    .b(_14975_),
    .out0(_14976_));
 b15and003an1n02x5 _23758_ (.a(_12538_),
    .b(_12595_),
    .c(_12641_),
    .o(_14977_));
 b15oai022as1n02x5 _23759_ (.a(_12684_),
    .b(_12654_),
    .c(_12750_),
    .d(_13722_),
    .o1(_14978_));
 b15nanb02an1n03x5 _23760_ (.a(net629),
    .b(net621),
    .out0(_14979_));
 b15oab012aq1n04x5 _23761_ (.a(_12723_),
    .b(_13727_),
    .c(_14979_),
    .out0(_14980_));
 b15nor002ar1n06x5 _23762_ (.a(_13707_),
    .b(_14980_),
    .o1(_14981_));
 b15oai013ar1n08x5 _23763_ (.a(net635),
    .b(_14977_),
    .c(_14978_),
    .d(_14981_),
    .o1(_14982_));
 b15nand03ar1n04x5 _23764_ (.a(\us03.a[2] ),
    .b(_13570_),
    .c(_12611_),
    .o1(_14983_));
 b15oai112ar1n08x5 _23765_ (.a(\us03.a[3] ),
    .b(_14983_),
    .c(_13715_),
    .d(_12714_),
    .o1(_14984_));
 b15nor003an1n04x5 _23766_ (.a(\us03.a[1] ),
    .b(_12551_),
    .c(_12714_),
    .o1(_14985_));
 b15nor003al1n04x5 _23767_ (.a(\us03.a[2] ),
    .b(_12603_),
    .c(_12762_),
    .o1(_14986_));
 b15oai013as1n08x5 _23768_ (.a(_14984_),
    .b(_14985_),
    .c(_14986_),
    .d(\us03.a[3] ),
    .o1(_14987_));
 b15aoai13aq1n03x5 _23769_ (.a(_12601_),
    .b(net637),
    .c(_13599_),
    .d(_12584_),
    .o1(_14988_));
 b15aoi012aq1n06x5 _23770_ (.a(_14810_),
    .b(_14988_),
    .c(_13548_),
    .o1(_14989_));
 b15aoi012al1n02x5 _23771_ (.a(_12601_),
    .b(_12594_),
    .c(_12753_),
    .o1(_14990_));
 b15oai022ar1n06x5 _23772_ (.a(_13580_),
    .b(_12684_),
    .c(_12654_),
    .d(_12762_),
    .o1(_14991_));
 b15aoi012al1n06x5 _23773_ (.a(_14990_),
    .b(_14991_),
    .c(_12581_),
    .o1(_14992_));
 b15nand04as1n16x5 _23774_ (.a(_14982_),
    .b(_14987_),
    .c(_14989_),
    .d(_14992_),
    .o1(_14993_));
 b15nonb03ar1n03x5 _23775_ (.a(net628),
    .b(net623),
    .c(net627),
    .out0(_14994_));
 b15aoai13ar1n02x5 _23776_ (.a(net642),
    .b(_14994_),
    .c(_12636_),
    .d(_12687_),
    .o1(_14995_));
 b15aoai13ar1n02x5 _23777_ (.a(net639),
    .b(\us03.a[7] ),
    .c(_12688_),
    .d(_14995_),
    .o1(_14996_));
 b15oai022ar1n06x5 _23778_ (.a(net642),
    .b(_13735_),
    .c(_14489_),
    .d(\us03.a[2] ),
    .o1(_14997_));
 b15aoai13ah1n03x5 _23779_ (.a(_14996_),
    .b(net639),
    .c(_13656_),
    .d(_14997_),
    .o1(_14998_));
 b15aoi012as1n02x5 _23780_ (.a(_12554_),
    .b(_12611_),
    .c(_12581_),
    .o1(_14999_));
 b15oaoi13ah1n04x5 _23781_ (.a(net631),
    .b(_14998_),
    .c(_14999_),
    .d(_12580_),
    .o1(_15000_));
 b15oaoi13ah1n03x5 _23782_ (.a(_13688_),
    .b(_12615_),
    .c(_12645_),
    .d(_12752_),
    .o1(_15001_));
 b15aoi112ar1n08x5 _23783_ (.a(_13580_),
    .b(_15001_),
    .c(_12677_),
    .d(net640),
    .o1(_15002_));
 b15aoi012al1n02x5 _23784_ (.a(_13688_),
    .b(_12564_),
    .c(_12563_),
    .o1(_15003_));
 b15oai022as1n06x5 _23785_ (.a(_12600_),
    .b(_13580_),
    .c(_13722_),
    .d(_15003_),
    .o1(_15004_));
 b15xor002ar1n02x5 _23786_ (.a(net630),
    .b(net629),
    .out0(_15005_));
 b15nano23ar1n02x5 _23787_ (.a(net626),
    .b(_12564_),
    .c(_12580_),
    .d(_15005_),
    .out0(_15006_));
 b15orn003an1n03x5 _23788_ (.a(_12581_),
    .b(_12769_),
    .c(_15006_),
    .o(_15007_));
 b15oai122al1n16x5 _23789_ (.a(_12581_),
    .b(_12600_),
    .c(_13580_),
    .d(_12677_),
    .e(_12747_),
    .o1(_15008_));
 b15aoi122as1n08x5 _23790_ (.a(_15002_),
    .b(_15004_),
    .c(net640),
    .d(_15007_),
    .e(_15008_),
    .o1(_15009_));
 b15norp02ah1n02x5 _23791_ (.a(_12601_),
    .b(_12677_),
    .o1(_15010_));
 b15aoai13aq1n08x5 _23792_ (.a(net637),
    .b(_15010_),
    .c(_13589_),
    .d(_13683_),
    .o1(_15011_));
 b15aoai13ar1n02x5 _23793_ (.a(_12747_),
    .b(_12581_),
    .c(_12545_),
    .d(_13599_),
    .o1(_15012_));
 b15nand02ah1n02x5 _23794_ (.a(_12554_),
    .b(_15012_),
    .o1(_15013_));
 b15and003al1n02x5 _23795_ (.a(net638),
    .b(_12641_),
    .c(_13595_),
    .o(_15014_));
 b15oai112al1n08x5 _23796_ (.a(_12515_),
    .b(_13570_),
    .c(_12724_),
    .d(_15014_),
    .o1(_15015_));
 b15nor003aq1n02x5 _23797_ (.a(_12569_),
    .b(_13606_),
    .c(_13727_),
    .o1(_15016_));
 b15oai112ah1n06x5 _23798_ (.a(net638),
    .b(_12515_),
    .c(_14473_),
    .d(_15016_),
    .o1(_15017_));
 b15nand04an1n12x5 _23799_ (.a(_15011_),
    .b(_15013_),
    .c(_15015_),
    .d(_15017_),
    .o1(_15018_));
 b15nandp3ar1n02x5 _23800_ (.a(_12707_),
    .b(_12700_),
    .c(_12697_),
    .o1(_15019_));
 b15aoi022ar1n02x5 _23801_ (.a(_12687_),
    .b(_12641_),
    .c(_12651_),
    .d(_12666_),
    .o1(_15020_));
 b15oai013aq1n02x5 _23802_ (.a(_15019_),
    .b(_15020_),
    .c(_13547_),
    .d(_12671_),
    .o1(_15021_));
 b15nor002ar1n06x5 _23803_ (.a(net642),
    .b(_12766_),
    .o1(_15022_));
 b15norp02ar1n02x5 _23804_ (.a(_12553_),
    .b(_12689_),
    .o1(_15023_));
 b15oai112an1n04x5 _23805_ (.a(_12593_),
    .b(_13616_),
    .c(_15022_),
    .d(_15023_),
    .o1(_15024_));
 b15nand03al1n02x5 _23806_ (.a(net634),
    .b(_13607_),
    .c(_13700_),
    .o1(_15025_));
 b15nona23al1n05x5 _23807_ (.a(_13748_),
    .b(_15021_),
    .c(_15024_),
    .d(_15025_),
    .out0(_15026_));
 b15nano23aq1n12x5 _23808_ (.a(_12605_),
    .b(_15009_),
    .c(_15018_),
    .d(_15026_),
    .out0(_15027_));
 b15norp02aq1n03x5 _23809_ (.a(_12750_),
    .b(_12751_),
    .o1(_15028_));
 b15nandp2aq1n02x5 _23810_ (.a(net627),
    .b(_12666_),
    .o1(_15029_));
 b15aoi022aq1n02x5 _23811_ (.a(net627),
    .b(_12687_),
    .c(_14994_),
    .d(net639),
    .o1(_15030_));
 b15oai022as1n06x5 _23812_ (.a(_15029_),
    .b(_13686_),
    .c(_15030_),
    .d(net635),
    .o1(_15031_));
 b15nor002aq1n03x5 _23813_ (.a(net631),
    .b(_12671_),
    .o1(_15032_));
 b15aoai13as1n08x5 _23814_ (.a(net642),
    .b(_15028_),
    .c(_15031_),
    .d(_15032_),
    .o1(_15033_));
 b15nona23as1n32x5 _23815_ (.a(_14993_),
    .b(_15000_),
    .c(_15027_),
    .d(_15033_),
    .out0(_15034_));
 b15aoi112ah1n04x5 _23816_ (.a(_13313_),
    .b(_13496_),
    .c(_13999_),
    .d(_13514_),
    .o1(_15035_));
 b15nor004al1n02x5 _23817_ (.a(_14377_),
    .b(_13417_),
    .c(_13399_),
    .d(_13917_),
    .o1(_15036_));
 b15nanb02ar1n02x5 _23818_ (.a(net668),
    .b(net647),
    .out0(_15037_));
 b15aob012al1n04x5 _23819_ (.a(\us32.a[1] ),
    .b(net654),
    .c(_15037_),
    .out0(_15038_));
 b15aoi022ar1n02x5 _23820_ (.a(net664),
    .b(_13325_),
    .c(_15036_),
    .d(_15038_),
    .o1(_15039_));
 b15aoi022an1n08x5 _23821_ (.a(_13924_),
    .b(_14388_),
    .c(_13977_),
    .d(_13996_),
    .o1(_15040_));
 b15oai012ar1n02x5 _23822_ (.a(_15039_),
    .b(_15040_),
    .c(net664),
    .o1(_15041_));
 b15oab012ar1n06x5 _23823_ (.a(_15035_),
    .b(_15041_),
    .c(net656),
    .out0(_15042_));
 b15aoi013aq1n02x5 _23824_ (.a(net668),
    .b(_13410_),
    .c(_13917_),
    .d(_13985_),
    .o1(_15043_));
 b15nand02al1n03x5 _23825_ (.a(_14418_),
    .b(_15043_),
    .o1(_15044_));
 b15nand03aq1n02x5 _23826_ (.a(_13459_),
    .b(_13515_),
    .c(_13362_),
    .o1(_15045_));
 b15nanb02ar1n02x5 _23827_ (.a(\us32.a[1] ),
    .b(net647),
    .out0(_15046_));
 b15nand04as1n02x5 _23828_ (.a(net644),
    .b(_13388_),
    .c(_14420_),
    .d(_15046_),
    .o1(_15047_));
 b15oai112an1n06x5 _23829_ (.a(_13377_),
    .b(_15045_),
    .c(_15047_),
    .d(_13362_),
    .o1(_15048_));
 b15nanb02as1n02x5 _23830_ (.a(net662),
    .b(net650),
    .out0(_15049_));
 b15nandp3ar1n02x5 _23831_ (.a(net658),
    .b(_13374_),
    .c(_13382_),
    .o1(_15050_));
 b15nand02ar1n02x5 _23832_ (.a(_13313_),
    .b(net644),
    .o1(_15051_));
 b15oaoi13as1n02x5 _23833_ (.a(_15049_),
    .b(_15050_),
    .c(_14509_),
    .d(_15051_),
    .o1(_15052_));
 b15oai013al1n06x5 _23834_ (.a(_15044_),
    .b(_15048_),
    .c(_15052_),
    .d(_13355_),
    .o1(_15053_));
 b15nandp3al1n03x5 _23835_ (.a(net647),
    .b(_13515_),
    .c(_13362_),
    .o1(_15054_));
 b15nand02al1n12x5 _23836_ (.a(net668),
    .b(net644),
    .o1(_15055_));
 b15oaoi13ah1n04x5 _23837_ (.a(_15054_),
    .b(_15055_),
    .c(net644),
    .d(_13340_),
    .o1(_15056_));
 b15aoi022aq1n04x5 _23838_ (.a(_13506_),
    .b(_13945_),
    .c(_13515_),
    .d(_13958_),
    .o1(_15057_));
 b15aoi012al1n02x5 _23839_ (.a(_13513_),
    .b(_13515_),
    .c(net656),
    .o1(_15058_));
 b15oai022an1n08x5 _23840_ (.a(_13488_),
    .b(_15057_),
    .c(_15058_),
    .d(_13367_),
    .o1(_15059_));
 b15nandp2aq1n16x5 _23841_ (.a(_13515_),
    .b(_13382_),
    .o1(_15060_));
 b15oai122as1n08x5 _23842_ (.a(_13377_),
    .b(_14379_),
    .c(_14560_),
    .d(_15060_),
    .e(_13347_),
    .o1(_15061_));
 b15aoi122an1n06x5 _23843_ (.a(_15056_),
    .b(_15059_),
    .c(_13402_),
    .d(_15061_),
    .e(_13340_),
    .o1(_15062_));
 b15aoi122ah1n06x5 _23844_ (.a(net656),
    .b(_13496_),
    .c(_13523_),
    .d(_13955_),
    .e(_14003_),
    .o1(_15063_));
 b15nandp3ar1n02x5 _23845_ (.a(net649),
    .b(_13523_),
    .c(_13934_),
    .o1(_15064_));
 b15nanb02al1n08x5 _23846_ (.a(net668),
    .b(net653),
    .out0(_15065_));
 b15orn003ar1n02x5 _23847_ (.a(_13302_),
    .b(_13398_),
    .c(_15065_),
    .o(_15066_));
 b15aoi013aq1n02x5 _23848_ (.a(_15063_),
    .b(_15064_),
    .c(_15066_),
    .d(net658),
    .o1(_15067_));
 b15nano23an1n08x5 _23849_ (.a(net658),
    .b(net645),
    .c(net648),
    .d(\us32.a[5] ),
    .out0(_15068_));
 b15qgbno2an1n05x5 _23850_ (.o1(_15069_),
    .a(_13421_),
    .b(_13374_));
 b15oai012al1n02x5 _23851_ (.a(net668),
    .b(net662),
    .c(net654),
    .o1(_15070_));
 b15xor002as1n02x5 _23852_ (.a(_13340_),
    .b(_15070_),
    .out0(_15071_));
 b15oaoi13aq1n04x5 _23853_ (.a(_15067_),
    .b(_15068_),
    .c(_15069_),
    .d(_15071_),
    .o1(_15072_));
 b15nand03al1n12x5 _23854_ (.a(_15053_),
    .b(_15062_),
    .c(_15072_),
    .o1(_15073_));
 b15nandp2al1n03x5 _23855_ (.a(net668),
    .b(net662),
    .o1(_15074_));
 b15oai022ar1n06x5 _23856_ (.a(net668),
    .b(_13345_),
    .c(_15074_),
    .d(net664),
    .o1(_15075_));
 b15aoai13an1n06x5 _23857_ (.a(_13442_),
    .b(_15075_),
    .c(_13977_),
    .d(_13916_),
    .o1(_15076_));
 b15nandp3ah1n04x5 _23858_ (.a(_13380_),
    .b(_13397_),
    .c(_13920_),
    .o1(_15077_));
 b15oai112as1n06x5 _23859_ (.a(net664),
    .b(_13367_),
    .c(_13345_),
    .d(_13355_),
    .o1(_15078_));
 b15oai112ar1n16x5 _23860_ (.a(_15076_),
    .b(_15077_),
    .c(_15078_),
    .d(_13390_),
    .o1(_15079_));
 b15oai012ar1n02x5 _23861_ (.a(net658),
    .b(net646),
    .c(_13418_),
    .o1(_15080_));
 b15nand02ah1n16x5 _23862_ (.a(_13313_),
    .b(_13459_),
    .o1(_15081_));
 b15norp03ar1n02x5 _23863_ (.a(_14377_),
    .b(_13417_),
    .c(_13408_),
    .o1(_15082_));
 b15and003ar1n02x5 _23864_ (.a(_15080_),
    .b(_15081_),
    .c(_15082_),
    .o(_15083_));
 b15nor004ar1n02x5 _23865_ (.a(net653),
    .b(_13505_),
    .c(_14361_),
    .d(_13382_),
    .o1(_15084_));
 b15aoai13ar1n02x5 _23866_ (.a(_13340_),
    .b(net666),
    .c(net660),
    .d(_13438_),
    .o1(_15085_));
 b15aoi022ar1n02x5 _23867_ (.a(_13418_),
    .b(_13438_),
    .c(_13523_),
    .d(_14000_),
    .o1(_15086_));
 b15aob012al1n02x5 _23868_ (.a(_15084_),
    .b(_15085_),
    .c(_15086_),
    .out0(_15087_));
 b15aoi022ar1n08x5 _23869_ (.a(_13415_),
    .b(_13371_),
    .c(_13361_),
    .d(_13417_),
    .o1(_15088_));
 b15norp02al1n02x5 _23870_ (.a(net657),
    .b(_15088_),
    .o1(_15089_));
 b15norp02ar1n02x5 _23871_ (.a(net667),
    .b(_13481_),
    .o1(_15090_));
 b15oai022al1n02x5 _23872_ (.a(_13374_),
    .b(_13425_),
    .c(_15090_),
    .d(net661),
    .o1(_15091_));
 b15aoi013an1n04x5 _23873_ (.a(_15089_),
    .b(_15091_),
    .c(_13478_),
    .d(_13375_),
    .o1(_15092_));
 b15nona23aq1n05x5 _23874_ (.a(_15079_),
    .b(_15083_),
    .c(_15087_),
    .d(_15092_),
    .out0(_15093_));
 b15nor004al1n02x5 _23875_ (.a(net649),
    .b(net643),
    .c(_14379_),
    .d(_14416_),
    .o1(_15094_));
 b15nor004al1n02x5 _23876_ (.a(net643),
    .b(net646),
    .c(_13423_),
    .d(_13306_),
    .o1(_15095_));
 b15oaoi13ah1n02x5 _23877_ (.a(_15094_),
    .b(net658),
    .c(_13938_),
    .d(_15095_),
    .o1(_15096_));
 b15aoi013al1n02x5 _23878_ (.a(_13340_),
    .b(_13396_),
    .c(_13920_),
    .d(_13955_),
    .o1(_15097_));
 b15aoi012ar1n02x5 _23879_ (.a(_13410_),
    .b(_13362_),
    .c(_14377_),
    .o1(_15098_));
 b15oai013ar1n03x5 _23880_ (.a(_15097_),
    .b(_15098_),
    .c(_13306_),
    .d(_13459_),
    .o1(_15099_));
 b15nandp2al1n12x5 _23881_ (.a(_13388_),
    .b(_13402_),
    .o1(_15100_));
 b15oai022ar1n06x5 _23882_ (.a(_15100_),
    .b(_13345_),
    .c(_13500_),
    .d(net656),
    .o1(_15101_));
 b15aoi012aq1n02x5 _23883_ (.a(_15099_),
    .b(_15101_),
    .c(net668),
    .o1(_15102_));
 b15oai013aq1n02x5 _23884_ (.a(_13340_),
    .b(net660),
    .c(_13310_),
    .d(_15060_),
    .o1(_15103_));
 b15aoi012ar1n06x5 _23885_ (.a(_15103_),
    .b(_14506_),
    .c(_13355_),
    .o1(_15104_));
 b15oai022aq1n08x5 _23886_ (.a(_13421_),
    .b(_15096_),
    .c(_15102_),
    .d(_15104_),
    .o1(_15105_));
 b15nor004as1n12x5 _23887_ (.a(_15042_),
    .b(_15073_),
    .c(_15093_),
    .d(_15105_),
    .o1(_15106_));
 b15xnr002an1n16x5 _23888_ (.a(_13546_),
    .b(_15106_),
    .out0(_15107_));
 b15xor002as1n06x5 _23889_ (.a(_15034_),
    .b(_15107_),
    .out0(_15108_));
 b15xor002an1n16x5 _23890_ (.a(_14976_),
    .b(_15108_),
    .out0(_15109_));
 b15bfn001as1n64x5 max_length407 (.a(net410),
    .o(net407));
 b15oai012as1n24x5 _23892_ (.a(_14830_),
    .b(_15109_),
    .c(net533),
    .o1(_15111_));
 b15xor002an1n02x5 _23893_ (.a(_09901_),
    .b(_15111_),
    .out0(_00125_));
 b15inv000ah1n10x5 _23894_ (.a(\text_in_r[5] ),
    .o1(_15112_));
 b15oai022ar1n02x5 _23895_ (.a(_14152_),
    .b(_13770_),
    .c(_14936_),
    .d(net898),
    .o1(_15113_));
 b15oai022ar1n02x5 _23896_ (.a(net907),
    .b(_14152_),
    .c(_14192_),
    .d(net886),
    .o1(_15114_));
 b15ao0022aq1n02x5 _23897_ (.a(net912),
    .b(_15113_),
    .c(_15114_),
    .d(_12883_),
    .o(_15115_));
 b15aoi022an1n08x5 _23898_ (.a(net899),
    .b(_12811_),
    .c(_14592_),
    .d(_12987_),
    .o1(_15116_));
 b15nor003ar1n06x5 _23899_ (.a(net889),
    .b(_13871_),
    .c(_15116_),
    .o1(_15117_));
 b15oai012ah1n02x5 _23900_ (.a(net901),
    .b(_12954_),
    .c(_12875_),
    .o1(_15118_));
 b15oai022aq1n08x5 _23901_ (.a(net901),
    .b(_15115_),
    .c(_15117_),
    .d(_15118_),
    .o1(_15119_));
 b15nand04ar1n02x5 _23902_ (.a(_12851_),
    .b(_12883_),
    .c(_12798_),
    .d(_13801_),
    .o1(_15120_));
 b15oai012al1n02x5 _23903_ (.a(_15120_),
    .b(_13793_),
    .c(_12851_),
    .o1(_15121_));
 b15aoi012an1n02x5 _23904_ (.a(_12863_),
    .b(_12968_),
    .c(net911),
    .o1(_15122_));
 b15aoi012an1n02x5 _23905_ (.a(_12987_),
    .b(_12968_),
    .c(net905),
    .o1(_15123_));
 b15oai022ar1n08x5 _23906_ (.a(net905),
    .b(_15122_),
    .c(_15123_),
    .d(net911),
    .o1(_15124_));
 b15aoi012al1n04x5 _23907_ (.a(_15121_),
    .b(_15124_),
    .c(_13809_),
    .o1(_15125_));
 b15nand04ar1n02x5 _23908_ (.a(net911),
    .b(_12964_),
    .c(_12883_),
    .d(_12798_),
    .o1(_15126_));
 b15oaoi13al1n02x5 _23909_ (.a(net905),
    .b(_15126_),
    .c(_13007_),
    .d(_12932_),
    .o1(_15127_));
 b15nand02ar1n02x5 _23910_ (.a(_12851_),
    .b(_12909_),
    .o1(_15128_));
 b15oai013ar1n02x5 _23911_ (.a(_15128_),
    .b(_12910_),
    .c(_13803_),
    .d(_12851_),
    .o1(_15129_));
 b15aoi013as1n02x5 _23912_ (.a(_15127_),
    .b(_15129_),
    .c(net901),
    .d(_13015_),
    .o1(_15130_));
 b15norp02ar1n03x5 _23913_ (.a(net898),
    .b(_14143_),
    .o1(_15131_));
 b15oai012ah1n04x5 _23914_ (.a(_14188_),
    .b(_13003_),
    .c(_12950_),
    .o1(_15132_));
 b15nand02ah1n04x5 _23915_ (.a(_12881_),
    .b(_12796_),
    .o1(_15133_));
 b15oai013ar1n04x5 _23916_ (.a(_14230_),
    .b(_15133_),
    .c(_13794_),
    .d(net911),
    .o1(_15134_));
 b15aoi122an1n04x5 _23917_ (.a(_12919_),
    .b(_15131_),
    .c(_15132_),
    .d(_15134_),
    .e(net898),
    .o1(_15135_));
 b15nand04as1n08x5 _23918_ (.a(_15119_),
    .b(_15125_),
    .c(_15130_),
    .d(_15135_),
    .o1(_15136_));
 b15oai022al1n02x5 _23919_ (.a(_13803_),
    .b(_12827_),
    .c(_12917_),
    .d(_12820_),
    .o1(_15137_));
 b15oai012ar1n03x5 _23920_ (.a(_13805_),
    .b(_13787_),
    .c(_12917_),
    .o1(_15138_));
 b15aoi022aq1n06x5 _23921_ (.a(net911),
    .b(_15137_),
    .c(_15138_),
    .d(net905),
    .o1(_15139_));
 b15aoi022al1n02x5 _23922_ (.a(net905),
    .b(_12991_),
    .c(_13860_),
    .d(_13798_),
    .o1(_15140_));
 b15nor002ar1n02x5 _23923_ (.a(_12950_),
    .b(_15140_),
    .o1(_15141_));
 b15aoi013ar1n04x5 _23924_ (.a(_15141_),
    .b(_13798_),
    .c(_12820_),
    .d(_12950_),
    .o1(_15142_));
 b15oai112aq1n02x5 _23925_ (.a(net901),
    .b(_12800_),
    .c(_13007_),
    .d(_12904_),
    .o1(_15143_));
 b15oaoi13an1n03x5 _23926_ (.a(_12877_),
    .b(_13803_),
    .c(_12782_),
    .d(_13007_),
    .o1(_15144_));
 b15oaoi13ar1n04x5 _23927_ (.a(_12851_),
    .b(_15143_),
    .c(_15144_),
    .d(net901),
    .o1(_15145_));
 b15aoi022aq1n12x5 _23928_ (.a(_12851_),
    .b(_15139_),
    .c(_15142_),
    .d(_15145_),
    .o1(_15146_));
 b15aoai13ar1n02x5 _23929_ (.a(net907),
    .b(_12851_),
    .c(_12796_),
    .d(_12874_),
    .o1(_15147_));
 b15aoai13ar1n02x5 _23930_ (.a(net912),
    .b(_12789_),
    .c(_12798_),
    .d(_12822_),
    .o1(_15148_));
 b15aoi022ar1n02x5 _23931_ (.a(_13769_),
    .b(_15147_),
    .c(_15148_),
    .d(_12851_),
    .o1(_15149_));
 b15nor003aq1n06x5 _23932_ (.a(net897),
    .b(_13801_),
    .c(_14589_),
    .o1(_15150_));
 b15oai012aq1n03x5 _23933_ (.a(_12820_),
    .b(_15149_),
    .c(_15150_),
    .o1(_15151_));
 b15norp03an1n16x5 _23934_ (.a(net903),
    .b(_12870_),
    .c(_12956_),
    .o1(_15152_));
 b15xor002aq1n06x5 _23935_ (.a(net902),
    .b(_12990_),
    .out0(_15153_));
 b15aoi022as1n06x5 _23936_ (.a(_14195_),
    .b(_14236_),
    .c(_15153_),
    .d(_12950_),
    .o1(_15154_));
 b15oai022an1n06x5 _23937_ (.a(_12879_),
    .b(_15152_),
    .c(_15154_),
    .d(_12909_),
    .o1(_15155_));
 b15nandp2ah1n03x5 _23938_ (.a(_12879_),
    .b(_15154_),
    .o1(_15156_));
 b15aoai13ar1n08x5 _23939_ (.a(_15151_),
    .b(_15155_),
    .c(_15156_),
    .d(_12851_),
    .o1(_15157_));
 b15aoi013ah1n03x5 _23940_ (.a(net905),
    .b(_13769_),
    .c(_14185_),
    .d(_14597_),
    .o1(_15158_));
 b15aoi022an1n06x5 _23941_ (.a(_13882_),
    .b(_13859_),
    .c(_12912_),
    .d(_12811_),
    .o1(_15159_));
 b15nor003ah1n06x5 _23942_ (.a(_12782_),
    .b(_14616_),
    .c(_15159_),
    .o1(_15160_));
 b15aoi012an1n02x5 _23943_ (.a(_13860_),
    .b(_14143_),
    .c(net911),
    .o1(_15161_));
 b15aoi012aq1n02x5 _23944_ (.a(_13798_),
    .b(_12909_),
    .c(net911),
    .o1(_15162_));
 b15oai222as1n08x5 _23945_ (.a(_12857_),
    .b(_12904_),
    .c(_15133_),
    .d(_15161_),
    .e(_15162_),
    .f(net901),
    .o1(_15163_));
 b15oai013ar1n08x5 _23946_ (.a(_12851_),
    .b(_15158_),
    .c(_15160_),
    .d(_15163_),
    .o1(_15164_));
 b15nor004ar1n02x5 _23947_ (.a(net905),
    .b(net898),
    .c(_14152_),
    .d(_13011_),
    .o1(_15165_));
 b15oai022al1n04x5 _23948_ (.a(net886),
    .b(_14205_),
    .c(_12960_),
    .d(_14152_),
    .o1(_15166_));
 b15aoi012ar1n02x5 _23949_ (.a(_15165_),
    .b(_15166_),
    .c(_12883_),
    .o1(_15167_));
 b15oai012ar1n02x5 _23950_ (.a(net903),
    .b(_13013_),
    .c(_13813_),
    .o1(_15168_));
 b15oaoi13al1n02x5 _23951_ (.a(_12782_),
    .b(_14602_),
    .c(_14936_),
    .d(net898),
    .o1(_15169_));
 b15aoi012al1n02x5 _23952_ (.a(_12851_),
    .b(_13769_),
    .c(_13838_),
    .o1(_15170_));
 b15nano23al1n05x5 _23953_ (.a(_15167_),
    .b(_15168_),
    .c(_15169_),
    .d(_15170_),
    .out0(_15171_));
 b15oai012an1n06x5 _23954_ (.a(_15164_),
    .b(_15171_),
    .c(net912),
    .o1(_15172_));
 b15nor004as1n12x5 _23955_ (.a(_15136_),
    .b(_15146_),
    .c(_15157_),
    .d(_15172_),
    .o1(_15173_));
 b15nor004ah1n03x5 _23956_ (.a(net641),
    .b(_12766_),
    .c(_12552_),
    .d(_12683_),
    .o1(_15174_));
 b15oai013ar1n06x5 _23957_ (.a(_12613_),
    .b(_12683_),
    .c(_12549_),
    .d(_13606_),
    .o1(_15175_));
 b15aoai13aq1n08x5 _23958_ (.a(net630),
    .b(_15174_),
    .c(_15175_),
    .d(net641),
    .o1(_15176_));
 b15nandp3an1n08x5 _23959_ (.a(_12519_),
    .b(_12563_),
    .c(_12598_),
    .o1(_15177_));
 b15nand04al1n16x5 _23960_ (.a(_13764_),
    .b(_13765_),
    .c(_15176_),
    .d(_15177_),
    .o1(_15178_));
 b15norp02ar1n02x5 _23961_ (.a(_12591_),
    .b(_12762_),
    .o1(_15179_));
 b15norp03al1n02x5 _23962_ (.a(_12552_),
    .b(_12553_),
    .c(_12658_),
    .o1(_15180_));
 b15oai013aq1n04x5 _23963_ (.a(net637),
    .b(_12577_),
    .c(_15179_),
    .d(_15180_),
    .o1(_15181_));
 b15and003al1n02x5 _23964_ (.a(_12646_),
    .b(_12697_),
    .c(_13563_),
    .o(_15182_));
 b15nanb03aq1n03x5 _23965_ (.a(net631),
    .b(net621),
    .c(net641),
    .out0(_15183_));
 b15aoi112ah1n04x5 _23966_ (.a(_12547_),
    .b(_15183_),
    .c(_13555_),
    .d(_12683_),
    .o1(_15184_));
 b15oai022as1n08x5 _23967_ (.a(_12601_),
    .b(_13654_),
    .c(_13707_),
    .d(net631),
    .o1(_15185_));
 b15nor002ah1n02x5 _23968_ (.a(_14979_),
    .b(_12649_),
    .o1(_15186_));
 b15aoi112an1n06x5 _23969_ (.a(_15182_),
    .b(_15184_),
    .c(_15185_),
    .d(_15186_),
    .o1(_15187_));
 b15nand03an1n16x5 _23970_ (.a(_12545_),
    .b(_12636_),
    .c(_13595_),
    .o1(_15188_));
 b15nand02ar1n02x5 _23971_ (.a(_13567_),
    .b(_13548_),
    .o1(_15189_));
 b15aob012al1n04x5 _23972_ (.a(_12511_),
    .b(_15188_),
    .c(_15189_),
    .out0(_15190_));
 b15oaoi13al1n03x5 _23973_ (.a(_12581_),
    .b(_12584_),
    .c(_12591_),
    .d(net640),
    .o1(_15191_));
 b15oai012as1n06x5 _23974_ (.a(_12645_),
    .b(_15191_),
    .c(_13567_),
    .o1(_15192_));
 b15nand04ah1n12x5 _23975_ (.a(_15181_),
    .b(_15187_),
    .c(_15190_),
    .d(_15192_),
    .o1(_15193_));
 b15nand02aq1n06x5 _23976_ (.a(_12657_),
    .b(_12724_),
    .o1(_15194_));
 b15norp03ar1n12x5 _23977_ (.a(_12545_),
    .b(_12547_),
    .c(_12549_),
    .o1(_15195_));
 b15oai012aq1n06x5 _23978_ (.a(_13547_),
    .b(_13686_),
    .c(_15195_),
    .o1(_15196_));
 b15nand03ah1n06x5 _23979_ (.a(net623),
    .b(_12722_),
    .c(_12723_),
    .o1(_15197_));
 b15aoi012as1n04x5 _23980_ (.a(_13752_),
    .b(_13567_),
    .c(_12550_),
    .o1(_15198_));
 b15aoi222as1n12x5 _23981_ (.a(net638),
    .b(_15194_),
    .c(_15196_),
    .d(_12511_),
    .e(_15197_),
    .f(_15198_),
    .o1(_15199_));
 b15aoai13ah1n03x5 _23982_ (.a(_13711_),
    .b(_14475_),
    .c(net632),
    .d(_12554_),
    .o1(_15200_));
 b15aoi022an1n04x5 _23983_ (.a(_12550_),
    .b(_12646_),
    .c(_13700_),
    .d(_13712_),
    .o1(_15201_));
 b15aoi022an1n04x5 _23984_ (.a(_12603_),
    .b(_12697_),
    .c(_12752_),
    .d(net642),
    .o1(_15202_));
 b15oai122aq1n12x5 _23985_ (.a(_15200_),
    .b(_15201_),
    .c(_12581_),
    .d(_12591_),
    .e(_15202_),
    .o1(_15203_));
 b15nor004as1n12x5 _23986_ (.a(_15178_),
    .b(_15193_),
    .c(_15199_),
    .d(_15203_),
    .o1(_15204_));
 b15nand03al1n03x5 _23987_ (.a(net632),
    .b(_14472_),
    .c(_12595_),
    .o1(_15205_));
 b15aoi012aq1n02x5 _23988_ (.a(_14472_),
    .b(_12570_),
    .c(net640),
    .o1(_15206_));
 b15oaoi13an1n04x5 _23989_ (.a(net635),
    .b(_15205_),
    .c(_15206_),
    .d(_12754_),
    .o1(_15207_));
 b15oai012as1n02x5 _23990_ (.a(_12597_),
    .b(_14479_),
    .c(_12551_),
    .o1(_15208_));
 b15aoi022ah1n02x5 _23991_ (.a(net635),
    .b(_12597_),
    .c(_12643_),
    .d(_12752_),
    .o1(_15209_));
 b15oaoi13al1n04x5 _23992_ (.a(net632),
    .b(_15208_),
    .c(_15209_),
    .d(\us03.a[1] ),
    .o1(_15210_));
 b15aoai13aq1n04x5 _23993_ (.a(net631),
    .b(_14433_),
    .c(_13683_),
    .d(_12515_),
    .o1(_15211_));
 b15oai112ah1n12x5 _23994_ (.a(_15188_),
    .b(_15211_),
    .c(_12511_),
    .d(_12542_),
    .o1(_15212_));
 b15aoi112ar1n08x5 _23995_ (.a(_15207_),
    .b(_15210_),
    .c(\us03.a[1] ),
    .d(_15212_),
    .o1(_15213_));
 b15oaoi13an1n03x5 _23996_ (.a(net633),
    .b(net630),
    .c(_12553_),
    .d(net622),
    .o1(_15214_));
 b15oai122as1n08x5 _23997_ (.a(net637),
    .b(_12601_),
    .c(_12718_),
    .d(_15214_),
    .e(_12511_),
    .o1(_15215_));
 b15nandp2aq1n04x5 _23998_ (.a(_13599_),
    .b(_12747_),
    .o1(_15216_));
 b15oai012al1n16x5 _23999_ (.a(_15215_),
    .b(_15216_),
    .c(net637),
    .o1(_15217_));
 b15aoi012ar1n02x5 _24000_ (.a(_12718_),
    .b(_12597_),
    .c(_12515_),
    .o1(_15218_));
 b15oai012ar1n06x5 _24001_ (.a(_12771_),
    .b(_15218_),
    .c(_12545_),
    .o1(_15219_));
 b15nor004aq1n03x5 _24002_ (.a(net642),
    .b(net635),
    .c(_12569_),
    .d(_13606_),
    .o1(_15220_));
 b15aoai13aq1n06x5 _24003_ (.a(net639),
    .b(_15220_),
    .c(_12718_),
    .d(net642),
    .o1(_15221_));
 b15aoi012al1n04x5 _24004_ (.a(net631),
    .b(_12515_),
    .c(_12554_),
    .o1(_15222_));
 b15nor003an1n03x5 _24005_ (.a(_12511_),
    .b(net627),
    .c(_12669_),
    .o1(_15223_));
 b15oaoi13ah1n03x5 _24006_ (.a(net639),
    .b(_12766_),
    .c(_12553_),
    .d(net642),
    .o1(_15224_));
 b15oaoi13ah1n04x5 _24007_ (.a(_15223_),
    .b(_13602_),
    .c(_15022_),
    .d(_15224_),
    .o1(_15225_));
 b15oai112as1n16x5 _24008_ (.a(_15221_),
    .b(_15222_),
    .c(_14449_),
    .d(_15225_),
    .o1(_15226_));
 b15aoi022ar1n02x5 _24009_ (.a(_12657_),
    .b(_13628_),
    .c(_12752_),
    .d(net639),
    .o1(_15227_));
 b15nor002ah1n03x5 _24010_ (.a(_12550_),
    .b(_12752_),
    .o1(_15228_));
 b15oai112an1n08x5 _24011_ (.a(\us03.a[3] ),
    .b(_15227_),
    .c(_15228_),
    .d(net642),
    .o1(_15229_));
 b15aoi022as1n08x5 _24012_ (.a(_15217_),
    .b(_15219_),
    .c(_15226_),
    .d(_15229_),
    .o1(_15230_));
 b15nand04as1n16x5 _24013_ (.a(_12544_),
    .b(_15204_),
    .c(_15213_),
    .d(_15230_),
    .o1(_15231_));
 b15xor002as1n12x5 _24014_ (.a(_15173_),
    .b(_15231_),
    .out0(_15232_));
 b15aoi022al1n02x5 _24015_ (.a(_13184_),
    .b(_13057_),
    .c(_13112_),
    .d(_13129_),
    .o1(_15233_));
 b15oai012aq1n06x5 _24016_ (.a(net783),
    .b(_13206_),
    .c(_15233_),
    .o1(_15234_));
 b15aoi012al1n04x5 _24017_ (.a(_14067_),
    .b(_13130_),
    .c(_13101_),
    .o1(_15235_));
 b15nona23ah1n02x5 _24018_ (.a(_13196_),
    .b(_13206_),
    .c(_14749_),
    .d(_13091_),
    .out0(_15236_));
 b15aoi022aq1n02x5 _24019_ (.a(_13063_),
    .b(_13100_),
    .c(_14029_),
    .d(_13181_),
    .o1(_15237_));
 b15oai012al1n08x5 _24020_ (.a(_15236_),
    .b(_15237_),
    .c(_13067_),
    .o1(_15238_));
 b15orn003ar1n04x5 _24021_ (.a(net780),
    .b(_14098_),
    .c(_14853_),
    .o(_15239_));
 b15oai022ah1n12x5 _24022_ (.a(_15234_),
    .b(_15235_),
    .c(_15238_),
    .d(_15239_),
    .o1(_15240_));
 b15nand04ar1n02x5 _24023_ (.a(_13063_),
    .b(_13124_),
    .c(_13129_),
    .d(_13222_),
    .o1(_15241_));
 b15oai112aq1n02x5 _24024_ (.a(net796),
    .b(_15241_),
    .c(_14063_),
    .d(_13159_),
    .o1(_15242_));
 b15aoi012ar1n02x5 _24025_ (.a(_14288_),
    .b(_14063_),
    .c(_14067_),
    .o1(_15243_));
 b15oai013aq1n04x5 _24026_ (.a(_15242_),
    .b(_15243_),
    .c(net796),
    .d(_14273_),
    .o1(_15244_));
 b15nandp2al1n05x5 _24027_ (.a(net796),
    .b(net791),
    .o1(_15245_));
 b15nandp2ah1n03x5 _24028_ (.a(_13067_),
    .b(_13050_),
    .o1(_15246_));
 b15aoi012an1n02x5 _24029_ (.a(_14296_),
    .b(_15245_),
    .c(_15246_),
    .o1(_15247_));
 b15aoi013ar1n06x5 _24030_ (.a(_15247_),
    .b(_14249_),
    .c(_14035_),
    .d(_13067_),
    .o1(_15248_));
 b15oai112ah1n12x5 _24031_ (.a(_15240_),
    .b(_15244_),
    .c(_15248_),
    .d(net781),
    .o1(_15249_));
 b15oai012ar1n03x5 _24032_ (.a(_13022_),
    .b(_14284_),
    .c(_15245_),
    .o1(_15250_));
 b15oai012an1n02x5 _24033_ (.a(net788),
    .b(_13249_),
    .c(_13213_),
    .o1(_15251_));
 b15oai012ar1n04x5 _24034_ (.a(net796),
    .b(net792),
    .c(_13249_),
    .o1(_15252_));
 b15aoi013ah1n03x5 _24035_ (.a(_15250_),
    .b(_15251_),
    .c(_15252_),
    .d(_13272_),
    .o1(_15253_));
 b15aoi022ar1n04x5 _24036_ (.a(net784),
    .b(_13091_),
    .c(_14750_),
    .d(net776),
    .o1(_15254_));
 b15nor003ah1n04x5 _24037_ (.a(net792),
    .b(_13052_),
    .c(_15254_),
    .o1(_15255_));
 b15and002ar1n02x5 _24038_ (.a(net770),
    .b(net796),
    .o(_15256_));
 b15oai112al1n06x5 _24039_ (.a(_13091_),
    .b(_13203_),
    .c(_14048_),
    .d(_15256_),
    .o1(_15257_));
 b15nand02an1n02x5 _24040_ (.a(_13067_),
    .b(_14131_),
    .o1(_15258_));
 b15aoi022ar1n04x5 _24041_ (.a(net779),
    .b(_13203_),
    .c(_14317_),
    .d(_14254_),
    .o1(_15259_));
 b15oai012al1n06x5 _24042_ (.a(_15257_),
    .b(_15258_),
    .c(_15259_),
    .o1(_15260_));
 b15oaoi13as1n08x5 _24043_ (.a(_15253_),
    .b(_13114_),
    .c(_15255_),
    .d(_15260_),
    .o1(_15261_));
 b15nandp3ar1n02x5 _24044_ (.a(net785),
    .b(_13040_),
    .c(_13277_),
    .o1(_15262_));
 b15aoi012ar1n02x5 _24045_ (.a(_13249_),
    .b(_13080_),
    .c(_15262_),
    .o1(_15263_));
 b15aoai13ar1n02x5 _24046_ (.a(net780),
    .b(_13277_),
    .c(_13080_),
    .d(net785),
    .o1(_15264_));
 b15oa0012ah1n03x5 _24047_ (.a(_14730_),
    .b(_15263_),
    .c(_15264_),
    .o(_15265_));
 b15aoi112ar1n02x5 _24048_ (.a(net789),
    .b(net780),
    .c(net778),
    .d(net795),
    .o1(_15266_));
 b15nand04as1n03x5 _24049_ (.a(_13291_),
    .b(_14107_),
    .c(_14683_),
    .d(_15266_),
    .o1(_15267_));
 b15aoi012ar1n08x5 _24050_ (.a(_14129_),
    .b(_14872_),
    .c(_13114_),
    .o1(_15268_));
 b15nand03ar1n06x5 _24051_ (.a(_14256_),
    .b(_14757_),
    .c(_13129_),
    .o1(_15269_));
 b15oai012ah1n06x5 _24052_ (.a(_15267_),
    .b(_15268_),
    .c(_15269_),
    .o1(_15270_));
 b15oai012aq1n06x5 _24053_ (.a(_14708_),
    .b(_13211_),
    .c(net774),
    .o1(_15271_));
 b15aoi013al1n08x5 _24054_ (.a(_15270_),
    .b(_15271_),
    .c(_14285_),
    .d(_13237_),
    .o1(_15272_));
 b15oai022ar1n08x5 _24055_ (.a(_13072_),
    .b(_14025_),
    .c(_13217_),
    .d(_13045_),
    .o1(_15273_));
 b15aoi013al1n06x5 _24056_ (.a(_13229_),
    .b(_15273_),
    .c(_13129_),
    .d(_13215_),
    .o1(_15274_));
 b15nand04an1n16x5 _24057_ (.a(_15261_),
    .b(_15265_),
    .c(_15272_),
    .d(_15274_),
    .o1(_15275_));
 b15norp03as1n04x5 _24058_ (.a(net791),
    .b(_13052_),
    .c(_13053_),
    .o1(_15276_));
 b15oai012al1n08x5 _24059_ (.a(_13067_),
    .b(_13149_),
    .c(_15276_),
    .o1(_15277_));
 b15and002ar1n02x5 _24060_ (.a(net791),
    .b(_13089_),
    .o(_15278_));
 b15oai112as1n06x5 _24061_ (.a(_13022_),
    .b(_15277_),
    .c(_15278_),
    .d(_14034_),
    .o1(_15279_));
 b15oai012al1n08x5 _24062_ (.a(_14022_),
    .b(_14281_),
    .c(_14034_),
    .o1(_15280_));
 b15nor002ah1n02x5 _24063_ (.a(net796),
    .b(_14711_),
    .o1(_15281_));
 b15aoi112an1n06x5 _24064_ (.a(_13185_),
    .b(_15281_),
    .c(net796),
    .d(_13050_),
    .o1(_15282_));
 b15oai013ah1n12x5 _24065_ (.a(_15279_),
    .b(_15280_),
    .c(_15282_),
    .d(_13022_),
    .o1(_15283_));
 b15nand03ar1n03x5 _24066_ (.a(\us21.a[0] ),
    .b(_13269_),
    .c(_14294_),
    .o1(_15284_));
 b15oaoi13al1n02x5 _24067_ (.a(_13114_),
    .b(_13209_),
    .c(_13086_),
    .d(net784),
    .o1(_15285_));
 b15oai013ah1n03x5 _24068_ (.a(_15284_),
    .b(_15285_),
    .c(\us21.a[0] ),
    .d(_13171_),
    .o1(_15286_));
 b15aob012an1n16x5 _24069_ (.a(net792),
    .b(_13173_),
    .c(_15286_),
    .out0(_15287_));
 b15nona23as1n32x5 _24070_ (.a(_15249_),
    .b(_15275_),
    .c(_15283_),
    .d(_15287_),
    .out0(_15288_));
 b15nor004ar1n02x5 _24071_ (.a(net662),
    .b(_13315_),
    .c(_13425_),
    .d(_13318_),
    .o1(_15289_));
 b15oaoi13ar1n02x5 _24072_ (.a(_13390_),
    .b(_15074_),
    .c(net664),
    .d(_13387_),
    .o1(_15290_));
 b15orn003ar1n02x5 _24073_ (.a(_13313_),
    .b(_15289_),
    .c(_15290_),
    .o(_15291_));
 b15nand02aq1n02x5 _24074_ (.a(net662),
    .b(net647),
    .o1(_15292_));
 b15nandp3ar1n03x5 _24075_ (.a(\us32.a[1] ),
    .b(_13388_),
    .c(_15055_),
    .o1(_15293_));
 b15oaoi13an1n08x5 _24076_ (.a(_15292_),
    .b(_15293_),
    .c(_13306_),
    .d(_15055_),
    .o1(_15294_));
 b15oai012ar1n02x5 _24077_ (.a(_13367_),
    .b(_13496_),
    .c(net664),
    .o1(_15295_));
 b15oaoi13ar1n03x5 _24078_ (.a(_15295_),
    .b(net664),
    .c(_13390_),
    .d(_13528_),
    .o1(_15296_));
 b15oai013ar1n06x5 _24079_ (.a(_15291_),
    .b(_15294_),
    .c(_15296_),
    .d(net656),
    .o1(_15297_));
 b15and002an1n04x5 _24080_ (.a(net667),
    .b(net655),
    .o(_15298_));
 b15aoi022an1n16x5 _24081_ (.a(_13928_),
    .b(_13939_),
    .c(_13486_),
    .d(_15298_),
    .o1(_15299_));
 b15oaoi13ar1n02x5 _24082_ (.a(net656),
    .b(_13318_),
    .c(_13350_),
    .d(net666),
    .o1(_15300_));
 b15aoai13an1n03x5 _24083_ (.a(_13382_),
    .b(_15300_),
    .c(_13425_),
    .d(_13506_),
    .o1(_15301_));
 b15aoai13as1n06x5 _24084_ (.a(_15297_),
    .b(_13421_),
    .c(_15299_),
    .d(_15301_),
    .o1(_15302_));
 b15nand02ar1n02x5 _24085_ (.a(net656),
    .b(_13397_),
    .o1(_15303_));
 b15oaoi13as1n02x5 _24086_ (.a(_13967_),
    .b(_15303_),
    .c(_15081_),
    .d(_14363_),
    .o1(_15304_));
 b15nand03ah1n02x5 _24087_ (.a(net656),
    .b(net650),
    .c(net654),
    .o1(_15305_));
 b15oaoi13aq1n08x5 _24088_ (.a(_15305_),
    .b(_13343_),
    .c(_13302_),
    .d(_13965_),
    .o1(_15306_));
 b15aoai13an1n08x5 _24089_ (.a(net668),
    .b(_15304_),
    .c(_15306_),
    .d(_13340_),
    .o1(_15307_));
 b15oai012as1n03x5 _24090_ (.a(_13450_),
    .b(_13410_),
    .c(net663),
    .o1(_15308_));
 b15oab012al1n02x5 _24091_ (.a(_13362_),
    .b(_13496_),
    .c(_13953_),
    .out0(_15309_));
 b15oai013ah1n03x5 _24092_ (.a(_13531_),
    .b(_13960_),
    .c(_13500_),
    .d(_13523_),
    .o1(_15310_));
 b15oai022ah1n06x5 _24093_ (.a(net666),
    .b(_15309_),
    .c(_15310_),
    .d(_14002_),
    .o1(_15311_));
 b15oai112aq1n12x5 _24094_ (.a(_14563_),
    .b(_15307_),
    .c(_15308_),
    .d(_15311_),
    .o1(_15312_));
 b15oai012ar1n02x5 _24095_ (.a(_13347_),
    .b(_13345_),
    .c(_13355_),
    .o1(_15313_));
 b15aoi022ar1n02x5 _24096_ (.a(_13355_),
    .b(_13410_),
    .c(_15313_),
    .d(_13340_),
    .o1(_15314_));
 b15norp03an1n02x5 _24097_ (.a(net664),
    .b(net656),
    .c(_14363_),
    .o1(_15315_));
 b15orn002ar1n02x5 _24098_ (.a(net650),
    .b(net647),
    .o(_15316_));
 b15oai022as1n04x5 _24099_ (.a(_13459_),
    .b(_15049_),
    .c(_15316_),
    .d(_13421_),
    .o1(_15317_));
 b15aoi222ar1n04x5 _24100_ (.a(_13380_),
    .b(_13442_),
    .c(_15315_),
    .d(_15317_),
    .e(_13938_),
    .f(_13945_),
    .o1(_15318_));
 b15oa0022al1n02x5 _24101_ (.a(_15100_),
    .b(_15314_),
    .c(_15318_),
    .d(net668),
    .o(_15319_));
 b15and002as1n02x5 _24102_ (.a(net650),
    .b(net644),
    .o(_15320_));
 b15aoai13aq1n04x5 _24103_ (.a(\us32.a[1] ),
    .b(_15320_),
    .c(_14511_),
    .d(net668),
    .o1(_15321_));
 b15aoi112ah1n03x5 _24104_ (.a(_13447_),
    .b(_14416_),
    .c(_14402_),
    .d(_15321_),
    .o1(_15322_));
 b15oai022as1n02x5 _24105_ (.a(_13302_),
    .b(_13399_),
    .c(_13967_),
    .d(_13343_),
    .o1(_15323_));
 b15aoi013al1n06x5 _24106_ (.a(_15322_),
    .b(_15323_),
    .c(net653),
    .d(_13998_),
    .o1(_15324_));
 b15nand02ar1n02x5 _24107_ (.a(net651),
    .b(_13536_),
    .o1(_15325_));
 b15aboi22ar1n02x5 _24108_ (.a(_14361_),
    .b(_13534_),
    .c(_13536_),
    .d(net657),
    .out0(_15326_));
 b15oai012as1n04x5 _24109_ (.a(_15325_),
    .b(_15326_),
    .c(net667),
    .o1(_15327_));
 b15oai012ar1n02x5 _24110_ (.a(net666),
    .b(_13905_),
    .c(_13916_),
    .o1(_15328_));
 b15oai112al1n02x5 _24111_ (.a(_13402_),
    .b(_13385_),
    .c(_13345_),
    .d(net666),
    .o1(_15329_));
 b15aoi012ar1n02x5 _24112_ (.a(net644),
    .b(_15329_),
    .c(net664),
    .o1(_15330_));
 b15and003aq1n04x5 _24113_ (.a(_15327_),
    .b(_15328_),
    .c(_15330_),
    .o(_15331_));
 b15aoi012al1n02x5 _24114_ (.a(_13345_),
    .b(net650),
    .c(_13355_),
    .o1(_15332_));
 b15aoi122al1n04x5 _24115_ (.a(_14395_),
    .b(_15306_),
    .c(net660),
    .d(_15332_),
    .e(_13934_),
    .o1(_15333_));
 b15oai012ar1n02x5 _24116_ (.a(net662),
    .b(_13403_),
    .c(net668),
    .o1(_15334_));
 b15oai012ar1n02x5 _24117_ (.a(net664),
    .b(net656),
    .c(_13387_),
    .o1(_15335_));
 b15aob012aq1n04x5 _24118_ (.a(_13944_),
    .b(_15334_),
    .c(_15335_),
    .out0(_15336_));
 b15aoi022ar1n02x5 _24119_ (.a(net656),
    .b(_13397_),
    .c(_13955_),
    .d(_13362_),
    .o1(_15337_));
 b15orn003al1n02x5 _24120_ (.a(_13340_),
    .b(net650),
    .c(_15337_),
    .o(_15338_));
 b15nand03aq1n08x5 _24121_ (.a(_15333_),
    .b(_15336_),
    .c(_15338_),
    .o1(_15339_));
 b15nano23ah1n08x5 _24122_ (.a(_15319_),
    .b(_15324_),
    .c(_15331_),
    .d(_15339_),
    .out0(_15340_));
 b15nand02ar1n02x5 _24123_ (.a(_13355_),
    .b(_14377_),
    .o1(_15341_));
 b15aoi112al1n02x5 _24124_ (.a(_13399_),
    .b(_14416_),
    .c(_15055_),
    .d(_15341_),
    .o1(_15342_));
 b15nand02ar1n02x5 _24125_ (.a(net668),
    .b(net654),
    .o1(_15343_));
 b15oai022ah1n02x5 _24126_ (.a(_13315_),
    .b(_15343_),
    .c(_14568_),
    .d(_14416_),
    .o1(_15344_));
 b15aoi013ah1n03x5 _24127_ (.a(_15342_),
    .b(_15344_),
    .c(net650),
    .d(_13340_),
    .o1(_15345_));
 b15nor002ar1n04x5 _24128_ (.a(net662),
    .b(net654),
    .o1(_15346_));
 b15oai112as1n06x5 _24129_ (.a(_13417_),
    .b(_14543_),
    .c(_15069_),
    .d(_15346_),
    .o1(_15347_));
 b15oai022al1n12x5 _24130_ (.a(_13355_),
    .b(_13533_),
    .c(_14400_),
    .d(_13949_),
    .o1(_15348_));
 b15aoi013ar1n08x5 _24131_ (.a(net658),
    .b(_14499_),
    .c(_15348_),
    .d(net664),
    .o1(_15349_));
 b15ao0022ar1n12x5 _24132_ (.a(net658),
    .b(_15345_),
    .c(_15347_),
    .d(_15349_),
    .o(_15350_));
 b15nona23as1n32x5 _24133_ (.a(_15302_),
    .b(_15312_),
    .c(_15340_),
    .d(_15350_),
    .out0(_15351_));
 b15xor002as1n16x5 _24134_ (.a(_15034_),
    .b(_15351_),
    .out0(_15352_));
 b15xor002ar1n12x5 _24135_ (.a(_15288_),
    .b(_15352_),
    .out0(_15353_));
 b15xor002an1n12x5 _24136_ (.a(_15232_),
    .b(_15353_),
    .out0(_15354_));
 b15mdn022as1n16x5 _24137_ (.a(_15112_),
    .b(_15354_),
    .o1(_15355_),
    .sa(net533));
 b15xor002ar1n02x5 _24138_ (.a(net500),
    .b(_15355_),
    .out0(_00126_));
 b15inv040ar1n06x5 _24139_ (.a(\text_in_r[6] ),
    .o1(_15356_));
 b15oai022ar1n02x5 _24140_ (.a(net894),
    .b(_12867_),
    .c(_14901_),
    .d(_13835_),
    .o1(_15357_));
 b15nandp3ar1n02x5 _24141_ (.a(net911),
    .b(_13848_),
    .c(_15357_),
    .o1(_15358_));
 b15nandp3ar1n02x5 _24142_ (.a(net909),
    .b(_12822_),
    .c(_12798_),
    .o1(_15359_));
 b15nand02ar1n02x5 _24143_ (.a(net890),
    .b(_12950_),
    .o1(_15360_));
 b15oaoi13ah1n02x5 _24144_ (.a(net903),
    .b(_15359_),
    .c(_15360_),
    .d(_12929_),
    .o1(_15361_));
 b15qgbxo2an1n10x5 _24145_ (.a(_12864_),
    .b(net904),
    .out0(_15362_));
 b15nor004an1n03x5 _24146_ (.a(net887),
    .b(net908),
    .c(_13011_),
    .d(_15362_),
    .o1(_15363_));
 b15nano23aq1n03x5 _24147_ (.a(_15358_),
    .b(net899),
    .c(_15361_),
    .d(_15363_),
    .out0(_15364_));
 b15aoai13ar1n02x5 _24148_ (.a(_12910_),
    .b(_15152_),
    .c(_13817_),
    .d(net903),
    .o1(_15365_));
 b15oai013aq1n06x5 _24149_ (.a(_14899_),
    .b(_13015_),
    .c(_14901_),
    .d(net890),
    .o1(_15366_));
 b15nandp3ar1n02x5 _24150_ (.a(net893),
    .b(_14154_),
    .c(_15366_),
    .o1(_15367_));
 b15nand02al1n04x5 _24151_ (.a(net896),
    .b(net903),
    .o1(_15368_));
 b15orn003ar1n02x5 _24152_ (.a(net893),
    .b(net886),
    .c(net889),
    .o(_15369_));
 b15oaoi13al1n02x5 _24153_ (.a(_15368_),
    .b(_15369_),
    .c(_13771_),
    .d(_13015_),
    .o1(_15370_));
 b15aoi112ar1n02x5 _24154_ (.a(net899),
    .b(_15370_),
    .c(_15152_),
    .d(_13801_),
    .o1(_15371_));
 b15and003ah1n02x5 _24155_ (.a(_15365_),
    .b(_15367_),
    .c(_15371_),
    .o(_15372_));
 b15nand02an1n03x5 _24156_ (.a(_12864_),
    .b(_12922_),
    .o1(_15373_));
 b15nanb02ar1n02x5 _24157_ (.a(\us10.a[5] ),
    .b(net909),
    .out0(_15374_));
 b15xor002ar1n03x5 _24158_ (.a(net888),
    .b(net913),
    .out0(_15375_));
 b15oai022ar1n06x5 _24159_ (.a(net888),
    .b(_12879_),
    .c(_15374_),
    .d(_15375_),
    .o1(_15376_));
 b15ao0012an1n02x5 _24160_ (.a(_14206_),
    .b(_12798_),
    .c(net909),
    .o(_15377_));
 b15aoi022aq1n08x5 _24161_ (.a(net891),
    .b(_15376_),
    .c(_15377_),
    .d(\us10.a[5] ),
    .o1(_15378_));
 b15oa0022aq1n02x5 _24162_ (.a(_15373_),
    .b(_14639_),
    .c(_15378_),
    .d(net894),
    .o(_15379_));
 b15oai022ah1n08x5 _24163_ (.a(_15364_),
    .b(_15372_),
    .c(_15379_),
    .d(_14628_),
    .o1(_15380_));
 b15nand02an1n02x5 _24164_ (.a(net899),
    .b(_13860_),
    .o1(_15381_));
 b15aoi012ar1n02x5 _24165_ (.a(_12909_),
    .b(_13860_),
    .c(_12825_),
    .o1(_15382_));
 b15oai022an1n02x5 _24166_ (.a(_12917_),
    .b(_15381_),
    .c(_15382_),
    .d(net899),
    .o1(_15383_));
 b15oai022aq1n02x5 _24167_ (.a(_12885_),
    .b(_12932_),
    .c(_12800_),
    .d(_14177_),
    .o1(_15384_));
 b15aoi112al1n04x5 _24168_ (.a(_12950_),
    .b(_15383_),
    .c(_15384_),
    .d(net906),
    .o1(_15385_));
 b15nor004al1n06x5 _24169_ (.a(net892),
    .b(_12832_),
    .c(net908),
    .d(_12998_),
    .o1(_15386_));
 b15oai022al1n12x5 _24170_ (.a(_12827_),
    .b(_14616_),
    .c(_14667_),
    .d(_12913_),
    .o1(_15387_));
 b15aoai13ah1n08x5 _24171_ (.a(_14241_),
    .b(_15386_),
    .c(_15387_),
    .d(net892),
    .o1(_15388_));
 b15nand02an1n04x5 _24172_ (.a(net899),
    .b(_15152_),
    .o1(_15389_));
 b15aoi013ah1n04x5 _24173_ (.a(_15385_),
    .b(_15388_),
    .c(_15389_),
    .d(_12950_),
    .o1(_15390_));
 b15oaoi13ar1n02x5 _24174_ (.a(_12950_),
    .b(_12800_),
    .c(_13769_),
    .d(net906),
    .o1(_15391_));
 b15nand02ar1n02x5 _24175_ (.a(net889),
    .b(_12877_),
    .o1(_15392_));
 b15aoi013as1n02x5 _24176_ (.a(_15391_),
    .b(_15392_),
    .c(_15373_),
    .d(_14634_),
    .o1(_15393_));
 b15oai012al1n08x5 _24177_ (.a(_12995_),
    .b(_13003_),
    .c(net911),
    .o1(_15394_));
 b15aoi022ar1n16x5 _24178_ (.a(net905),
    .b(_12909_),
    .c(_15394_),
    .d(net901),
    .o1(_15395_));
 b15oai022as1n06x5 _24179_ (.a(_12932_),
    .b(_15393_),
    .c(_15395_),
    .d(net899),
    .o1(_15396_));
 b15oai012an1n02x5 _24180_ (.a(net911),
    .b(_12885_),
    .c(_15381_),
    .o1(_15397_));
 b15xor002al1n02x5 _24181_ (.a(\us10.a[5] ),
    .b(net888),
    .out0(_15398_));
 b15nand04an1n06x5 _24182_ (.a(_12832_),
    .b(net891),
    .c(_14217_),
    .d(_15398_),
    .o1(_15399_));
 b15oai022ar1n02x5 _24183_ (.a(net899),
    .b(_12865_),
    .c(_14192_),
    .d(_12870_),
    .o1(_15400_));
 b15aob012ar1n04x5 _24184_ (.a(_15399_),
    .b(_15400_),
    .c(_13844_),
    .out0(_15401_));
 b15oai012ar1n06x5 _24185_ (.a(_15397_),
    .b(_15401_),
    .c(net911),
    .o1(_15402_));
 b15aoi012ar1n06x5 _24186_ (.a(_12789_),
    .b(_13817_),
    .c(net908),
    .o1(_15403_));
 b15nand02al1n04x5 _24187_ (.a(_12851_),
    .b(_12971_),
    .o1(_15404_));
 b15aoi022an1n06x5 _24188_ (.a(_12796_),
    .b(_12874_),
    .c(_12822_),
    .d(_12881_),
    .o1(_15405_));
 b15nand02ah1n03x5 _24189_ (.a(_12968_),
    .b(_12910_),
    .o1(_15406_));
 b15oai222ah1n12x5 _24190_ (.a(_15403_),
    .b(_15404_),
    .c(_15405_),
    .d(_14631_),
    .e(_12917_),
    .f(_15406_),
    .o1(_15407_));
 b15nand02ar1n02x5 _24191_ (.a(net892),
    .b(_12968_),
    .o1(_15408_));
 b15nandp3ar1n02x5 _24192_ (.a(net890),
    .b(_12940_),
    .c(_13801_),
    .o1(_15409_));
 b15aoi022ar1n02x5 _24193_ (.a(_12881_),
    .b(_12910_),
    .c(_13801_),
    .d(_12798_),
    .o1(_15410_));
 b15oaoi13as1n02x5 _24194_ (.a(_15408_),
    .b(_15409_),
    .c(_15410_),
    .d(_12832_),
    .o1(_15411_));
 b15norp02al1n02x5 _24195_ (.a(net892),
    .b(net902),
    .o1(_15412_));
 b15nano23ah1n02x5 _24196_ (.a(net887),
    .b(net890),
    .c(net900),
    .d(net894),
    .out0(_15413_));
 b15nano23ah1n02x5 _24197_ (.a(net894),
    .b(net900),
    .c(net890),
    .d(net887),
    .out0(_15414_));
 b15oai112al1n08x5 _24198_ (.a(_12922_),
    .b(_15412_),
    .c(_15413_),
    .d(_15414_),
    .o1(_15415_));
 b15nand04an1n06x5 _24199_ (.a(net908),
    .b(net902),
    .c(net900),
    .d(_12983_),
    .o1(_15416_));
 b15aoi012ah1n02x5 _24200_ (.a(_12986_),
    .b(_12940_),
    .c(net911),
    .o1(_15417_));
 b15oai122ar1n12x5 _24201_ (.a(_15415_),
    .b(_15416_),
    .c(_15417_),
    .d(_14628_),
    .e(_14963_),
    .o1(_15418_));
 b15nor004as1n06x5 _24202_ (.a(_13819_),
    .b(_15407_),
    .c(_15411_),
    .d(_15418_),
    .o1(_15419_));
 b15aoi022al1n08x5 _24203_ (.a(_12820_),
    .b(_13798_),
    .c(_12796_),
    .d(_12848_),
    .o1(_15420_));
 b15oai122ah1n12x5 _24204_ (.a(_13838_),
    .b(_15420_),
    .c(_12904_),
    .d(_13805_),
    .e(_12950_),
    .o1(_15421_));
 b15oaoi13al1n02x5 _24205_ (.a(_12977_),
    .b(_12949_),
    .c(_12870_),
    .d(_15362_),
    .o1(_15422_));
 b15aoi013ar1n02x5 _24206_ (.a(_12789_),
    .b(_12983_),
    .c(_12904_),
    .d(_13883_),
    .o1(_15423_));
 b15aoi022ar1n02x5 _24207_ (.a(net908),
    .b(_12940_),
    .c(_12986_),
    .d(_12910_),
    .o1(_15424_));
 b15oaoi13ah1n03x5 _24208_ (.a(_12820_),
    .b(_15423_),
    .c(_15424_),
    .d(_14610_),
    .o1(_15425_));
 b15oai013as1n03x5 _24209_ (.a(net899),
    .b(_15421_),
    .c(_15422_),
    .d(_15425_),
    .o1(_15426_));
 b15nand04ah1n08x5 _24210_ (.a(_14245_),
    .b(_15402_),
    .c(_15419_),
    .d(_15426_),
    .o1(_15427_));
 b15nor004as1n12x5 _24211_ (.a(_15380_),
    .b(_15390_),
    .c(_15396_),
    .d(_15427_),
    .o1(_15428_));
 b15aoi012ar1n02x5 _24212_ (.a(_13548_),
    .b(_13712_),
    .c(\us03.a[0] ),
    .o1(_15429_));
 b15oai022ah1n02x5 _24213_ (.a(_12511_),
    .b(_12760_),
    .c(_15429_),
    .d(_12581_),
    .o1(_15430_));
 b15oaoi13an1n03x5 _24214_ (.a(_12511_),
    .b(_12714_),
    .c(_12524_),
    .d(\us03.a[1] ),
    .o1(_15431_));
 b15oai013an1n08x5 _24215_ (.a(_12707_),
    .b(_12718_),
    .c(_15430_),
    .d(_15431_),
    .o1(_15432_));
 b15oai112aq1n02x5 _24216_ (.a(net632),
    .b(net636),
    .c(_12570_),
    .d(_13683_),
    .o1(_15433_));
 b15oai112ah1n06x5 _24217_ (.a(_12515_),
    .b(_12519_),
    .c(_12586_),
    .d(_12617_),
    .o1(_15434_));
 b15oaoi13aq1n04x5 _24218_ (.a(_12511_),
    .b(_15433_),
    .c(_15434_),
    .d(net632),
    .o1(_15435_));
 b15oai022an1n02x5 _24219_ (.a(_12662_),
    .b(_12601_),
    .c(_12591_),
    .d(_13606_),
    .o1(_15436_));
 b15nandp3aq1n02x5 _24220_ (.a(net642),
    .b(_12587_),
    .c(_15436_),
    .o1(_15437_));
 b15aoi022al1n06x5 _24221_ (.a(_12538_),
    .b(_12641_),
    .c(_12646_),
    .d(_13548_),
    .o1(_15438_));
 b15oaoi13an1n04x5 _24222_ (.a(net638),
    .b(_15437_),
    .c(_15438_),
    .d(net642),
    .o1(_15439_));
 b15nor004aq1n02x5 _24223_ (.a(net638),
    .b(_12766_),
    .c(_12717_),
    .d(_12689_),
    .o1(_15440_));
 b15aoi112ar1n02x5 _24224_ (.a(net632),
    .b(_15440_),
    .c(_12551_),
    .d(_12554_),
    .o1(_15441_));
 b15nand02ar1n02x5 _24225_ (.a(_14472_),
    .b(_14479_),
    .o1(_15442_));
 b15aoi013ah1n02x5 _24226_ (.a(_15441_),
    .b(_15442_),
    .c(net632),
    .d(_13695_),
    .o1(_15443_));
 b15oaoi13al1n03x5 _24227_ (.a(_12581_),
    .b(_12580_),
    .c(_12752_),
    .d(_12657_),
    .o1(_15444_));
 b15nanb02ar1n02x5 _24228_ (.a(_13686_),
    .b(_12762_),
    .out0(_15445_));
 b15oaoi13an1n02x5 _24229_ (.a(\us03.a[0] ),
    .b(_15445_),
    .c(_12550_),
    .d(\us03.a[2] ),
    .o1(_15446_));
 b15nor004ah1n04x5 _24230_ (.a(\us03.a[3] ),
    .b(_15228_),
    .c(_15444_),
    .d(_15446_),
    .o1(_15447_));
 b15nor004aq1n06x5 _24231_ (.a(_15435_),
    .b(_15439_),
    .c(_15443_),
    .d(_15447_),
    .o1(_15448_));
 b15aoai13as1n02x5 _24232_ (.a(_12581_),
    .b(_12577_),
    .c(_12597_),
    .d(_12545_),
    .o1(_15449_));
 b15aoi022aq1n02x5 _24233_ (.a(net641),
    .b(_12577_),
    .c(_13700_),
    .d(_12697_),
    .o1(_15450_));
 b15oai022al1n04x5 _24234_ (.a(net631),
    .b(_12692_),
    .c(_12669_),
    .d(_12654_),
    .o1(_15451_));
 b15nandp3al1n08x5 _24235_ (.a(net639),
    .b(_13556_),
    .c(_15451_),
    .o1(_15452_));
 b15aoi013ah1n04x5 _24236_ (.a(net634),
    .b(_15449_),
    .c(_15450_),
    .d(_15452_),
    .o1(_15453_));
 b15oai112ah1n06x5 _24237_ (.a(_13567_),
    .b(_12615_),
    .c(_12752_),
    .d(_14472_),
    .o1(_15454_));
 b15norp02an1n02x5 _24238_ (.a(_13727_),
    .b(_12771_),
    .o1(_15455_));
 b15oai012al1n06x5 _24239_ (.a(_13644_),
    .b(_15455_),
    .c(_12577_),
    .o1(_15456_));
 b15aoai13as1n04x5 _24240_ (.a(_13700_),
    .b(_14767_),
    .c(net633),
    .d(_13683_),
    .o1(_15457_));
 b15aoai13an1n06x5 _24241_ (.a(_12646_),
    .b(_12736_),
    .c(_12752_),
    .d(_12700_),
    .o1(_15458_));
 b15nand04an1n16x5 _24242_ (.a(_15454_),
    .b(_15456_),
    .c(_15457_),
    .d(_15458_),
    .o1(_15459_));
 b15nand02ar1n02x5 _24243_ (.a(_12545_),
    .b(_12611_),
    .o1(_15460_));
 b15oaoi13ar1n02x5 _24244_ (.a(net638),
    .b(_15460_),
    .c(_12601_),
    .d(_12600_),
    .o1(_15461_));
 b15nonb02ar1n02x5 _24245_ (.a(net623),
    .b(net639),
    .out0(_15462_));
 b15nano23an1n02x5 _24246_ (.a(net627),
    .b(net621),
    .c(net628),
    .d(net631),
    .out0(_15463_));
 b15aoai13al1n04x5 _24247_ (.a(_15462_),
    .b(_15463_),
    .c(_12723_),
    .d(_12651_),
    .o1(_15464_));
 b15aoi022as1n06x5 _24248_ (.a(_12515_),
    .b(_12666_),
    .c(_12687_),
    .d(_12551_),
    .o1(_15465_));
 b15oai013ar1n06x5 _24249_ (.a(_15464_),
    .b(_15465_),
    .c(_13660_),
    .d(_12629_),
    .o1(_15466_));
 b15nanb02ar1n02x5 _24250_ (.a(net634),
    .b(net628),
    .out0(_15467_));
 b15oai012an1n04x5 _24251_ (.a(_15467_),
    .b(_13686_),
    .c(net628),
    .o1(_15468_));
 b15nor002al1n04x5 _24252_ (.a(_12654_),
    .b(_14435_),
    .o1(_15469_));
 b15aoi022an1n08x5 _24253_ (.a(_12683_),
    .b(_15195_),
    .c(_15468_),
    .d(_15469_),
    .o1(_15470_));
 b15norp03as1n02x5 _24254_ (.a(_12552_),
    .b(_12553_),
    .c(_13563_),
    .o1(_15471_));
 b15oai012ar1n08x5 _24255_ (.a(_12720_),
    .b(_12763_),
    .c(_15471_),
    .o1(_15472_));
 b15nona23ah1n05x5 _24256_ (.a(_15461_),
    .b(_15466_),
    .c(_15470_),
    .d(_15472_),
    .out0(_15473_));
 b15nand02ar1n02x5 _24257_ (.a(_12611_),
    .b(_12646_),
    .o1(_15474_));
 b15and003an1n02x5 _24258_ (.a(net641),
    .b(_15177_),
    .c(_15474_),
    .o(_15475_));
 b15aoi122an1n04x5 _24259_ (.a(net641),
    .b(_12570_),
    .c(_12720_),
    .d(_12611_),
    .e(_13616_),
    .o1(_15476_));
 b15aoi022al1n12x5 _24260_ (.a(_12570_),
    .b(_14811_),
    .c(_12752_),
    .d(_12545_),
    .o1(_15477_));
 b15oai122an1n12x5 _24261_ (.a(_13629_),
    .b(_15475_),
    .c(_15476_),
    .d(_15477_),
    .e(_12581_),
    .o1(_15478_));
 b15nor004as1n12x5 _24262_ (.a(_15453_),
    .b(_15459_),
    .c(_15473_),
    .d(_15478_),
    .o1(_15479_));
 b15aoi022ar1n04x5 _24263_ (.a(_12511_),
    .b(_13683_),
    .c(_12718_),
    .d(_13565_),
    .o1(_15480_));
 b15oai022al1n06x5 _24264_ (.a(_12683_),
    .b(_12684_),
    .c(_15480_),
    .d(net635),
    .o1(_15481_));
 b15aob012aq1n02x5 _24265_ (.a(net642),
    .b(_12677_),
    .c(_13710_),
    .out0(_15482_));
 b15aoi012an1n02x5 _24266_ (.a(_13628_),
    .b(_13607_),
    .c(_12511_),
    .o1(_15483_));
 b15oai112aq1n08x5 _24267_ (.a(net639),
    .b(_15482_),
    .c(_15483_),
    .d(net635),
    .o1(_15484_));
 b15nano22ar1n02x5 _24268_ (.a(net642),
    .b(net624),
    .c(\us03.a[5] ),
    .out0(_15485_));
 b15oai112ar1n02x5 _24269_ (.a(\us03.a[2] ),
    .b(_12662_),
    .c(_13717_),
    .d(_15485_),
    .o1(_15486_));
 b15aoi022ar1n02x5 _24270_ (.a(\us03.a[2] ),
    .b(_13717_),
    .c(_12687_),
    .d(_12541_),
    .o1(_15487_));
 b15oaoi13ar1n02x5 _24271_ (.a(\us03.a[7] ),
    .b(_15486_),
    .c(_15487_),
    .d(net642),
    .o1(_15488_));
 b15orn003ah1n03x5 _24272_ (.a(net639),
    .b(_12697_),
    .c(_15488_),
    .o(_15489_));
 b15aoai13al1n08x5 _24273_ (.a(net631),
    .b(_15481_),
    .c(_15484_),
    .d(_15489_),
    .o1(_15490_));
 b15nand04as1n16x5 _24274_ (.a(_15432_),
    .b(_15448_),
    .c(_15479_),
    .d(_15490_),
    .o1(_15491_));
 b15xnr002as1n12x5 _24275_ (.a(_15428_),
    .b(_15491_),
    .out0(_15492_));
 b15oai013aq1n02x5 _24276_ (.a(_13910_),
    .b(_13306_),
    .c(_14377_),
    .d(net666),
    .o1(_15493_));
 b15obai22aq1n12x5 _24277_ (.a(_15493_),
    .b(_15081_),
    .c(_13500_),
    .d(_13345_),
    .out0(_15494_));
 b15oai022ar1n08x5 _24278_ (.a(net667),
    .b(_13336_),
    .c(_13510_),
    .d(_14388_),
    .o1(_15495_));
 b15oai022an1n04x5 _24279_ (.a(net655),
    .b(_13324_),
    .c(_13306_),
    .d(_13499_),
    .o1(_15496_));
 b15aoi122ar1n06x5 _24280_ (.a(_15494_),
    .b(_15495_),
    .c(net655),
    .d(_14573_),
    .e(_15496_),
    .o1(_15497_));
 b15oai012as1n02x5 _24281_ (.a(_13416_),
    .b(_15060_),
    .c(net655),
    .o1(_15498_));
 b15aoi022ar1n08x5 _24282_ (.a(_13415_),
    .b(_13403_),
    .c(_13371_),
    .d(_15498_),
    .o1(_15499_));
 b15oai022ah1n08x5 _24283_ (.a(_13340_),
    .b(_15497_),
    .c(_15499_),
    .d(net667),
    .o1(_15500_));
 b15oai012ar1n02x5 _24284_ (.a(net665),
    .b(_15298_),
    .c(_14366_),
    .o1(_15501_));
 b15aoi012aq1n02x5 _24285_ (.a(_13330_),
    .b(_13499_),
    .c(_15501_),
    .o1(_15502_));
 b15inv040al1n03x5 _24286_ (.a(_13403_),
    .o1(_15503_));
 b15oai122ar1n12x5 _24287_ (.a(net659),
    .b(_13531_),
    .c(_15503_),
    .d(_13454_),
    .e(_15060_),
    .o1(_15504_));
 b15oai022aq1n06x5 _24288_ (.a(_15503_),
    .b(_13390_),
    .c(_13454_),
    .d(_13500_),
    .o1(_15505_));
 b15oaoi13al1n08x5 _24289_ (.a(_15502_),
    .b(_15504_),
    .c(_15505_),
    .d(net659),
    .o1(_15506_));
 b15norp03ar1n03x5 _24290_ (.a(\us32.a[1] ),
    .b(net658),
    .c(net647),
    .o1(_15507_));
 b15aoi022as1n06x5 _24291_ (.a(net658),
    .b(_15320_),
    .c(_15507_),
    .d(_14511_),
    .o1(_15508_));
 b15aoi022ar1n12x5 _24292_ (.a(net647),
    .b(_13515_),
    .c(_13478_),
    .d(_14499_),
    .o1(_15509_));
 b15nandp2ah1n03x5 _24293_ (.a(net644),
    .b(_13417_),
    .o1(_15510_));
 b15oai122as1n16x5 _24294_ (.a(net661),
    .b(_15065_),
    .c(_15508_),
    .d(_15509_),
    .e(_15510_),
    .o1(_15511_));
 b15nand03ar1n03x5 _24295_ (.a(net657),
    .b(_13388_),
    .c(_13375_),
    .o1(_15512_));
 b15oaoi13al1n02x5 _24296_ (.a(net665),
    .b(_15512_),
    .c(_13510_),
    .d(net657),
    .o1(_15513_));
 b15norp02ar1n02x5 _24297_ (.a(_13355_),
    .b(_15512_),
    .o1(_15514_));
 b15oai013ah1n03x5 _24298_ (.a(_15511_),
    .b(_15513_),
    .c(_15514_),
    .d(net661),
    .o1(_15515_));
 b15oai022ah1n02x5 _24299_ (.a(net661),
    .b(_13509_),
    .c(_13510_),
    .d(_13514_),
    .o1(_15516_));
 b15nand02as1n02x5 _24300_ (.a(_13488_),
    .b(_14511_),
    .o1(_15517_));
 b15oai012ar1n12x5 _24301_ (.a(_15517_),
    .b(_14400_),
    .c(_13488_),
    .o1(_15518_));
 b15aoi013as1n06x5 _24302_ (.a(_15516_),
    .b(_15518_),
    .c(_13534_),
    .d(net661),
    .o1(_15519_));
 b15oai112al1n12x5 _24303_ (.a(_15506_),
    .b(_15515_),
    .c(_15519_),
    .d(net657),
    .o1(_15520_));
 b15aoi022an1n06x5 _24304_ (.a(net663),
    .b(_13442_),
    .c(_13980_),
    .d(net666),
    .o1(_15521_));
 b15oaoi13an1n04x5 _24305_ (.a(_13362_),
    .b(_13355_),
    .c(_13421_),
    .d(_13916_),
    .o1(_15522_));
 b15oai022al1n12x5 _24306_ (.a(_13347_),
    .b(_15521_),
    .c(_15522_),
    .d(_14560_),
    .o1(_15523_));
 b15norp02ar1n02x5 _24307_ (.a(net659),
    .b(_15060_),
    .o1(_15524_));
 b15oaoi13ar1n02x5 _24308_ (.a(net663),
    .b(_15060_),
    .c(_13531_),
    .d(net659),
    .o1(_15525_));
 b15oab012al1n06x5 _24309_ (.a(_13310_),
    .b(_15524_),
    .c(_15525_),
    .out0(_15526_));
 b15oai013al1n03x5 _24310_ (.a(net659),
    .b(_13315_),
    .c(_13417_),
    .d(_13350_),
    .o1(_15527_));
 b15oai112aq1n06x5 _24311_ (.a(_13925_),
    .b(_15527_),
    .c(net659),
    .d(_13442_),
    .o1(_15528_));
 b15aoi013ar1n03x5 _24312_ (.a(_14517_),
    .b(_13488_),
    .c(_13442_),
    .d(net659),
    .o1(_15529_));
 b15oai013aq1n06x5 _24313_ (.a(_15528_),
    .b(_15529_),
    .c(_13939_),
    .d(_13313_),
    .o1(_15530_));
 b15oab012an1n02x5 _24314_ (.a(net655),
    .b(_14387_),
    .c(_14389_),
    .out0(_15531_));
 b15xor002ar1n04x5 _24315_ (.a(net664),
    .b(net649),
    .out0(_15532_));
 b15oai112aq1n08x5 _24316_ (.a(_13362_),
    .b(_13955_),
    .c(_15532_),
    .d(net666),
    .o1(_15533_));
 b15nand04as1n02x5 _24317_ (.a(_13505_),
    .b(_13423_),
    .c(_13506_),
    .d(_13958_),
    .o1(_15534_));
 b15oai112ah1n08x5 _24318_ (.a(_15533_),
    .b(_15534_),
    .c(_13960_),
    .d(_13390_),
    .o1(_15535_));
 b15norp02al1n02x5 _24319_ (.a(_13355_),
    .b(_13447_),
    .o1(_15536_));
 b15oai112aq1n02x5 _24320_ (.a(net663),
    .b(_13500_),
    .c(_13350_),
    .d(_13315_),
    .o1(_15537_));
 b15oai112aq1n06x5 _24321_ (.a(_15536_),
    .b(_15537_),
    .c(net663),
    .d(_13442_),
    .o1(_15538_));
 b15nand04al1n02x5 _24322_ (.a(_13313_),
    .b(_13505_),
    .c(_13506_),
    .d(_13367_),
    .o1(_15539_));
 b15aob012ar1n04x5 _24323_ (.a(_13423_),
    .b(_13491_),
    .c(_15539_),
    .out0(_15540_));
 b15nona23ar1n12x5 _24324_ (.a(_15531_),
    .b(_15535_),
    .c(_15538_),
    .d(_15540_),
    .out0(_15541_));
 b15nor004as1n12x5 _24325_ (.a(_15523_),
    .b(_15526_),
    .c(_15530_),
    .d(_15541_),
    .o1(_15542_));
 b15nand02al1n12x5 _24326_ (.a(_13402_),
    .b(_13385_),
    .o1(_15543_));
 b15oai012ar1n02x5 _24327_ (.a(_13336_),
    .b(_13306_),
    .c(_13302_),
    .o1(_15544_));
 b15aoi022aq1n04x5 _24328_ (.a(net667),
    .b(_13928_),
    .c(_15544_),
    .d(net659),
    .o1(_15545_));
 b15oai122ar1n12x5 _24329_ (.a(_13313_),
    .b(_15543_),
    .c(_13367_),
    .d(_15545_),
    .e(net665),
    .o1(_15546_));
 b15oaoi13al1n03x5 _24330_ (.a(net665),
    .b(_13367_),
    .c(_13361_),
    .d(_14388_),
    .o1(_15547_));
 b15aoi012al1n02x5 _24331_ (.a(_13924_),
    .b(_13361_),
    .c(net667),
    .o1(_15548_));
 b15oai012ar1n08x5 _24332_ (.a(_15543_),
    .b(_15547_),
    .c(_15548_),
    .o1(_15549_));
 b15oai112as1n12x5 _24333_ (.a(_13494_),
    .b(_13523_),
    .c(_13398_),
    .d(_13479_),
    .o1(_15550_));
 b15aoai13as1n08x5 _24334_ (.a(_15546_),
    .b(_13313_),
    .c(_15549_),
    .d(_15550_),
    .o1(_15551_));
 b15nona23as1n32x5 _24335_ (.a(_15500_),
    .b(_15520_),
    .c(_15542_),
    .d(_15551_),
    .out0(_15552_));
 b15xor002an1n06x5 _24336_ (.a(_15231_),
    .b(_15552_),
    .out0(_15553_));
 b15aoi012an1n06x5 _24337_ (.a(_14058_),
    .b(_13092_),
    .c(_13066_),
    .o1(_15554_));
 b15nand02ar1n02x5 _24338_ (.a(net776),
    .b(net796),
    .o1(_15555_));
 b15oai022ar1n04x5 _24339_ (.a(net786),
    .b(_14034_),
    .c(_15554_),
    .d(_15555_),
    .o1(_15556_));
 b15oai122aq1n02x5 _24340_ (.a(_13130_),
    .b(_14296_),
    .c(_13277_),
    .d(_13086_),
    .e(_13067_),
    .o1(_15557_));
 b15aoi022ar1n02x5 _24341_ (.a(net791),
    .b(_15556_),
    .c(_15557_),
    .d(_13114_),
    .o1(_15558_));
 b15oai122ah1n02x5 _24342_ (.a(net791),
    .b(_13114_),
    .c(_14296_),
    .d(_14114_),
    .e(_13033_),
    .o1(_15559_));
 b15nanb02aq1n02x5 _24343_ (.a(net768),
    .b(\us21.a[0] ),
    .out0(_15560_));
 b15aoi012al1n06x5 _24344_ (.a(_13066_),
    .b(_13206_),
    .c(_15560_),
    .o1(_15561_));
 b15oai012al1n06x5 _24345_ (.a(_13259_),
    .b(_13176_),
    .c(_13092_),
    .o1(_15562_));
 b15oai022ah1n12x5 _24346_ (.a(_13033_),
    .b(_14288_),
    .c(_15561_),
    .d(_15562_),
    .o1(_15563_));
 b15oai012ar1n02x5 _24347_ (.a(_13130_),
    .b(_13086_),
    .c(net796),
    .o1(_15564_));
 b15oai013al1n02x5 _24348_ (.a(_15559_),
    .b(_15563_),
    .c(_15564_),
    .d(net791),
    .o1(_15565_));
 b15aob012aq1n04x5 _24349_ (.a(net782),
    .b(_15558_),
    .c(_15565_),
    .out0(_15566_));
 b15nonb03an1n02x5 _24350_ (.a(net796),
    .b(net786),
    .c(net781),
    .out0(_15567_));
 b15aoai13al1n06x5 _24351_ (.a(_15567_),
    .b(_13147_),
    .c(net791),
    .d(_13213_),
    .o1(_15568_));
 b15nano23as1n03x5 _24352_ (.a(net768),
    .b(net795),
    .c(net787),
    .d(net775),
    .out0(_15569_));
 b15oai112as1n16x5 _24353_ (.a(_14757_),
    .b(_14254_),
    .c(_14695_),
    .d(_15569_),
    .o1(_15570_));
 b15nand04ah1n06x5 _24354_ (.a(_13184_),
    .b(_13128_),
    .c(_13124_),
    .d(_13228_),
    .o1(_15571_));
 b15nand04ah1n06x5 _24355_ (.a(_13129_),
    .b(_13244_),
    .c(_13222_),
    .d(_14103_),
    .o1(_15572_));
 b15nand04as1n12x5 _24356_ (.a(_15568_),
    .b(_15570_),
    .c(_15571_),
    .d(_15572_),
    .o1(_15573_));
 b15aoai13ar1n04x5 _24357_ (.a(_13262_),
    .b(_13171_),
    .c(_13222_),
    .d(_13129_),
    .o1(_15574_));
 b15nand02ar1n02x5 _24358_ (.a(net796),
    .b(_15574_),
    .o1(_15575_));
 b15oai122as1n02x5 _24359_ (.a(_13067_),
    .b(net791),
    .c(_14702_),
    .d(_14114_),
    .e(net786),
    .o1(_15576_));
 b15and003al1n02x5 _24360_ (.a(_13022_),
    .b(_15575_),
    .c(_15576_),
    .o(_15577_));
 b15aoi022al1n02x5 _24361_ (.a(_14030_),
    .b(_13244_),
    .c(_13090_),
    .d(_13124_),
    .o1(_15578_));
 b15oai112al1n08x5 _24362_ (.a(_14316_),
    .b(_15578_),
    .c(_14288_),
    .d(_13211_),
    .o1(_15579_));
 b15aoi112aq1n06x5 _24363_ (.a(_15573_),
    .b(_15577_),
    .c(_15579_),
    .d(net796),
    .o1(_15580_));
 b15oai112an1n02x5 _24364_ (.a(net781),
    .b(_13100_),
    .c(_14089_),
    .d(_14090_),
    .o1(_15581_));
 b15oai112al1n04x5 _24365_ (.a(_13067_),
    .b(_13215_),
    .c(_14249_),
    .d(_14099_),
    .o1(_15582_));
 b15nor004as1n08x5 _24366_ (.a(_13140_),
    .b(_13072_),
    .c(_14687_),
    .d(_14075_),
    .o1(_15583_));
 b15aoai13ah1n03x5 _24367_ (.a(_15583_),
    .b(net774),
    .c(net773),
    .d(_13277_),
    .o1(_15584_));
 b15nand04al1n06x5 _24368_ (.a(_13124_),
    .b(_13176_),
    .c(_13208_),
    .d(_13217_),
    .o1(_15585_));
 b15nand04an1n06x5 _24369_ (.a(_15581_),
    .b(_15582_),
    .c(_15584_),
    .d(_15585_),
    .o1(_15586_));
 b15norp02ar1n03x5 _24370_ (.a(net769),
    .b(_13078_),
    .o1(_15587_));
 b15nor003ah1n02x5 _24371_ (.a(net772),
    .b(net782),
    .c(_14313_),
    .o1(_15588_));
 b15aoai13an1n08x5 _24372_ (.a(_15587_),
    .b(_15588_),
    .c(_14029_),
    .d(_13203_),
    .o1(_15589_));
 b15oab012aq1n03x5 _24373_ (.a(_15276_),
    .b(_13283_),
    .c(_13141_),
    .out0(_15590_));
 b15oai112al1n16x5 _24374_ (.a(_14832_),
    .b(_15589_),
    .c(_15590_),
    .d(net781),
    .o1(_15591_));
 b15norp03ar1n02x5 _24375_ (.a(net786),
    .b(_13161_),
    .c(_14103_),
    .o1(_15592_));
 b15aoi012ar1n02x5 _24376_ (.a(_15592_),
    .b(_14712_),
    .c(_13100_),
    .o1(_15593_));
 b15norp02an1n03x5 _24377_ (.a(net781),
    .b(_15593_),
    .o1(_15594_));
 b15rm6013el1n02x5 _24378_ (.a(_13114_),
    .b(_13072_),
    .c(_14702_),
    .carryb(_15595_));
 b15norp02ar1n02x5 _24379_ (.a(_13050_),
    .b(_14702_),
    .o1(_15596_));
 b15oai112aq1n02x5 _24380_ (.a(net781),
    .b(_15595_),
    .c(_15596_),
    .d(_13046_),
    .o1(_15597_));
 b15nona22ar1n02x5 _24381_ (.a(net796),
    .b(net786),
    .c(net781),
    .out0(_15598_));
 b15oai122as1n02x5 _24382_ (.a(net791),
    .b(_14288_),
    .c(_13211_),
    .d(_15598_),
    .e(_13161_),
    .o1(_15599_));
 b15norp02ar1n02x5 _24383_ (.a(net781),
    .b(_13086_),
    .o1(_15600_));
 b15oai013ar1n02x5 _24384_ (.a(_15599_),
    .b(_14725_),
    .c(_15600_),
    .d(net791),
    .o1(_15601_));
 b15aoi022ar1n02x5 _24385_ (.a(_14099_),
    .b(_13251_),
    .c(_13215_),
    .d(_13046_),
    .o1(_15602_));
 b15oai112aq1n04x5 _24386_ (.a(_15597_),
    .b(_15601_),
    .c(_15602_),
    .d(net795),
    .o1(_15603_));
 b15ornc04as1n12x5 _24387_ (.a(_15586_),
    .b(_15591_),
    .c(_15594_),
    .d(_15603_),
    .o(_15604_));
 b15aoi012al1n02x5 _24388_ (.a(net781),
    .b(_13130_),
    .c(_13227_),
    .o1(_15605_));
 b15aoi022ah1n06x5 _24389_ (.a(_13063_),
    .b(_13162_),
    .c(_15605_),
    .d(_13072_),
    .o1(_15606_));
 b15aoi112ar1n03x5 _24390_ (.a(net791),
    .b(net781),
    .c(_13130_),
    .d(_13227_),
    .o1(_15607_));
 b15oai012al1n06x5 _24391_ (.a(net796),
    .b(_13162_),
    .c(_15607_),
    .o1(_15608_));
 b15oai012ar1n02x5 _24392_ (.a(net781),
    .b(_13277_),
    .c(_13227_),
    .o1(_15609_));
 b15nand02ar1n02x5 _24393_ (.a(net796),
    .b(_13213_),
    .o1(_15610_));
 b15oai112as1n02x5 _24394_ (.a(_13161_),
    .b(_15610_),
    .c(net796),
    .d(_13185_),
    .o1(_15611_));
 b15oai012ah1n04x5 _24395_ (.a(_15609_),
    .b(_15611_),
    .c(net781),
    .o1(_15612_));
 b15aoi013aq1n08x5 _24396_ (.a(_13114_),
    .b(_15606_),
    .c(_15608_),
    .d(_15612_),
    .o1(_15613_));
 b15nano23as1n24x5 _24397_ (.a(_15566_),
    .b(_15580_),
    .c(_15604_),
    .d(_15613_),
    .out0(_15614_));
 b15xor002as1n08x5 _24398_ (.a(_15553_),
    .b(_15614_),
    .out0(_15615_));
 b15xor002ah1n16x5 _24399_ (.a(_15492_),
    .b(_15615_),
    .out0(_15616_));
 b15mdn022as1n12x5 _24400_ (.a(_15356_),
    .b(_15616_),
    .o1(_15617_),
    .sa(net533));
 b15xor002ar1n02x5 _24401_ (.a(net496),
    .b(_15617_),
    .out0(_00127_));
 b15inv040aq1n05x5 _24402_ (.a(net533),
    .o1(_15618_));
 b15norp02al1n04x5 _24403_ (.a(_15618_),
    .b(\text_in_r[7] ),
    .o1(_15619_));
 b15nandp2al1n02x5 _24404_ (.a(_13171_),
    .b(_14051_),
    .o1(_15620_));
 b15oai112ah1n06x5 _24405_ (.a(_13063_),
    .b(_15620_),
    .c(_14293_),
    .d(_13114_),
    .o1(_15621_));
 b15nona23ar1n02x5 _24406_ (.a(_13078_),
    .b(_14874_),
    .c(_13251_),
    .d(_13291_),
    .out0(_15622_));
 b15oai012ah1n02x5 _24407_ (.a(_15622_),
    .b(_13127_),
    .c(_13142_),
    .o1(_15623_));
 b15oaoi13aq1n03x5 _24408_ (.a(_15573_),
    .b(_15621_),
    .c(_15623_),
    .d(_13063_),
    .o1(_15624_));
 b15nano22aq1n03x5 _24409_ (.a(net778),
    .b(net773),
    .c(net784),
    .out0(_15625_));
 b15nonb03al1n04x5 _24410_ (.a(net784),
    .b(net773),
    .c(net778),
    .out0(_15626_));
 b15oai112aq1n16x5 _24411_ (.a(_13063_),
    .b(_14107_),
    .c(_15625_),
    .d(_15626_),
    .o1(_15627_));
 b15nandp3al1n03x5 _24412_ (.a(net791),
    .b(_13181_),
    .c(_14051_),
    .o1(_15628_));
 b15nandp3as1n08x5 _24413_ (.a(_14316_),
    .b(_15627_),
    .c(_15628_),
    .o1(_15629_));
 b15norp02ar1n02x5 _24414_ (.a(net768),
    .b(net785),
    .o1(_15630_));
 b15nona23ah1n02x5 _24415_ (.a(_14063_),
    .b(_15630_),
    .c(_14124_),
    .d(_13210_),
    .out0(_15631_));
 b15aoi022aq1n02x5 _24416_ (.a(net794),
    .b(_13244_),
    .c(_14874_),
    .d(_13124_),
    .o1(_15632_));
 b15oai013aq1n08x5 _24417_ (.a(_15631_),
    .b(_15632_),
    .c(_13156_),
    .d(_13078_),
    .o1(_15633_));
 b15aoi012al1n02x5 _24418_ (.a(_13208_),
    .b(_13217_),
    .c(_13174_),
    .o1(_15634_));
 b15norp03ar1n08x5 _24419_ (.a(_13140_),
    .b(_14025_),
    .c(_15634_),
    .o1(_15635_));
 b15nor004al1n12x5 _24420_ (.a(_14841_),
    .b(_15629_),
    .c(_15633_),
    .d(_15635_),
    .o1(_15636_));
 b15oaoi13al1n04x5 _24421_ (.a(_15246_),
    .b(_13209_),
    .c(_14296_),
    .d(net781),
    .o1(_15637_));
 b15nandp3ar1n02x5 _24422_ (.a(net782),
    .b(_13091_),
    .c(_14281_),
    .o1(_15638_));
 b15nandp3as1n02x5 _24423_ (.a(net772),
    .b(_13208_),
    .c(_14051_),
    .o1(_15639_));
 b15aoi012aq1n02x5 _24424_ (.a(_14123_),
    .b(_15638_),
    .c(_15639_),
    .o1(_15640_));
 b15nor004ar1n06x5 _24425_ (.a(_14121_),
    .b(_14310_),
    .c(_15637_),
    .d(_15640_),
    .o1(_15641_));
 b15nand03ar1n12x5 _24426_ (.a(_15624_),
    .b(_15636_),
    .c(_15641_),
    .o1(_15642_));
 b15oai012ar1n02x5 _24427_ (.a(_13217_),
    .b(_13090_),
    .c(_14030_),
    .o1(_15643_));
 b15oaoi13ar1n02x5 _24428_ (.a(net786),
    .b(_15643_),
    .c(_13040_),
    .d(_13141_),
    .o1(_15644_));
 b15aoai13an1n03x5 _24429_ (.a(net781),
    .b(_15644_),
    .c(_13262_),
    .d(_13090_),
    .o1(_15645_));
 b15oaoi13al1n08x5 _24430_ (.a(_13091_),
    .b(net776),
    .c(net792),
    .d(_14055_),
    .o1(_15646_));
 b15oai022ar1n02x5 _24431_ (.a(_13078_),
    .b(_13040_),
    .c(_15646_),
    .d(net772),
    .o1(_15647_));
 b15nandp2ah1n02x5 _24432_ (.a(_13215_),
    .b(_15647_),
    .o1(_15648_));
 b15aoai13as1n06x5 _24433_ (.a(_15645_),
    .b(net769),
    .c(_14896_),
    .d(_15648_),
    .o1(_15649_));
 b15aoai13ar1n02x5 _24434_ (.a(_13146_),
    .b(_13100_),
    .c(_13208_),
    .d(_13176_),
    .o1(_15650_));
 b15oaoi13an1n02x5 _24435_ (.a(_13114_),
    .b(_15650_),
    .c(_14114_),
    .d(_14095_),
    .o1(_15651_));
 b15aoi013an1n04x5 _24436_ (.a(_15651_),
    .b(_13124_),
    .c(_14030_),
    .d(net791),
    .o1(_15652_));
 b15aoai13as1n02x5 _24437_ (.a(net781),
    .b(_14098_),
    .c(_13171_),
    .d(net791),
    .o1(_15653_));
 b15aoi112an1n04x5 _24438_ (.a(net795),
    .b(_14096_),
    .c(_13181_),
    .d(_13244_),
    .o1(_15654_));
 b15aoi022as1n08x5 _24439_ (.a(net795),
    .b(_15652_),
    .c(_15653_),
    .d(_15654_),
    .o1(_15655_));
 b15nand02ar1n02x5 _24440_ (.a(net787),
    .b(_14249_),
    .o1(_15656_));
 b15oaoi13as1n02x5 _24441_ (.a(_15245_),
    .b(_15656_),
    .c(net787),
    .d(_14066_),
    .o1(_15657_));
 b15oai012ar1n02x5 _24442_ (.a(_13063_),
    .b(_13215_),
    .c(_13267_),
    .o1(_15658_));
 b15nandp3ar1n02x5 _24443_ (.a(net792),
    .b(_13022_),
    .c(_14129_),
    .o1(_15659_));
 b15aob012aq1n02x5 _24444_ (.a(_13234_),
    .b(_15658_),
    .c(_15659_),
    .out0(_15660_));
 b15oa0022ar1n02x5 _24445_ (.a(_14288_),
    .b(_13230_),
    .c(_14114_),
    .d(_13211_),
    .o(_15661_));
 b15norp02ar1n02x5 _24446_ (.a(_13067_),
    .b(_13127_),
    .o1(_15662_));
 b15aoi022ar1n02x5 _24447_ (.a(_13124_),
    .b(_13054_),
    .c(_14249_),
    .d(_15662_),
    .o1(_15663_));
 b15aoai13an1n02x5 _24448_ (.a(_15660_),
    .b(net792),
    .c(_15661_),
    .d(_15663_),
    .o1(_15664_));
 b15nandp3ar1n02x5 _24449_ (.a(_13067_),
    .b(_13213_),
    .c(_13262_),
    .o1(_15665_));
 b15oai112an1n04x5 _24450_ (.a(_13022_),
    .b(_15665_),
    .c(_13254_),
    .d(_13130_),
    .o1(_15666_));
 b15oai022ar1n02x5 _24451_ (.a(_14029_),
    .b(_13227_),
    .c(_15246_),
    .d(_13159_),
    .o1(_15667_));
 b15oai012as1n03x5 _24452_ (.a(_15666_),
    .b(_15667_),
    .c(_13022_),
    .o1(_15668_));
 b15nona23an1n12x5 _24453_ (.a(_15657_),
    .b(_15664_),
    .c(_15668_),
    .d(_13274_),
    .out0(_15669_));
 b15nor004as1n12x5 _24454_ (.a(_15642_),
    .b(_15649_),
    .c(_15655_),
    .d(_15669_),
    .o1(_15670_));
 b15nand03aq1n02x5 _24455_ (.a(net665),
    .b(_13385_),
    .c(_13375_),
    .o1(_15671_));
 b15nandp2aq1n05x5 _24456_ (.a(net661),
    .b(_13928_),
    .o1(_15672_));
 b15oaoi13ar1n08x5 _24457_ (.a(_13355_),
    .b(_15671_),
    .c(_15672_),
    .d(net665),
    .o1(_15673_));
 b15oai022ar1n02x5 _24458_ (.a(_13421_),
    .b(_13510_),
    .c(_13949_),
    .d(_13336_),
    .o1(_15674_));
 b15aoi112ah1n03x5 _24459_ (.a(_13313_),
    .b(_15673_),
    .c(_15674_),
    .d(_13340_),
    .o1(_15675_));
 b15nor004ar1n08x5 _24460_ (.a(net663),
    .b(_13459_),
    .c(_13306_),
    .d(_14522_),
    .o1(_15676_));
 b15aoi112as1n08x5 _24461_ (.a(net656),
    .b(_15676_),
    .c(_13528_),
    .d(_13361_),
    .o1(_15677_));
 b15oaoi13aq1n03x5 _24462_ (.a(_13949_),
    .b(_14406_),
    .c(_14012_),
    .d(net665),
    .o1(_15678_));
 b15mdn022ah1n03x5 _24463_ (.a(_14406_),
    .b(_14012_),
    .o1(_15679_),
    .sa(net661));
 b15aoai13ah1n06x5 _24464_ (.a(_13534_),
    .b(_15678_),
    .c(_15679_),
    .d(_13950_),
    .o1(_15680_));
 b15nanb02ar1n02x5 _24465_ (.a(net654),
    .b(\us32.a[1] ),
    .out0(_15681_));
 b15xor002ar1n02x5 _24466_ (.a(_13355_),
    .b(_15681_),
    .out0(_15682_));
 b15aoai13as1n02x5 _24467_ (.a(net647),
    .b(_13432_),
    .c(_15682_),
    .d(_14377_),
    .o1(_15683_));
 b15nand02an1n02x5 _24468_ (.a(_13355_),
    .b(_13897_),
    .o1(_15684_));
 b15aob012ah1n12x5 _24469_ (.a(_13920_),
    .b(_15683_),
    .c(_15684_),
    .out0(_15685_));
 b15aoi013ah1n06x5 _24470_ (.a(_15675_),
    .b(_15677_),
    .c(_15680_),
    .d(_15685_),
    .o1(_15686_));
 b15oai022ar1n04x5 _24471_ (.a(_13315_),
    .b(_13318_),
    .c(_14560_),
    .d(_13355_),
    .o1(_15687_));
 b15aoai13ar1n03x5 _24472_ (.a(_13421_),
    .b(_14354_),
    .c(_15687_),
    .d(_13340_),
    .o1(_15688_));
 b15aoi013ah1n02x5 _24473_ (.a(net657),
    .b(net661),
    .c(_13950_),
    .d(_13938_),
    .o1(_15689_));
 b15and002al1n02x5 _24474_ (.a(_15688_),
    .b(_15689_),
    .o(_15690_));
 b15norp02al1n02x5 _24475_ (.a(_13330_),
    .b(_13488_),
    .o1(_15691_));
 b15aoi013ah1n03x5 _24476_ (.a(_15691_),
    .b(_13996_),
    .c(_13421_),
    .d(_13355_),
    .o1(_15692_));
 b15aoai13an1n06x5 _24477_ (.a(_13965_),
    .b(_13412_),
    .c(_13996_),
    .d(net667),
    .o1(_15693_));
 b15aoi013ar1n08x5 _24478_ (.a(_15690_),
    .b(_15692_),
    .c(_15693_),
    .d(net657),
    .o1(_15694_));
 b15oai012al1n02x5 _24479_ (.a(net663),
    .b(_13390_),
    .c(_13450_),
    .o1(_15695_));
 b15aoi012aq1n04x5 _24480_ (.a(_15695_),
    .b(_13958_),
    .c(_14000_),
    .o1(_15696_));
 b15oai012an1n03x5 _24481_ (.a(_13500_),
    .b(_13390_),
    .c(net660),
    .o1(_15697_));
 b15nor003ar1n03x5 _24482_ (.a(net652),
    .b(_13302_),
    .c(_13399_),
    .o1(_15698_));
 b15nor003ah1n04x5 _24483_ (.a(_13392_),
    .b(_15697_),
    .c(_15698_),
    .o1(_15699_));
 b15oai022ar1n04x5 _24484_ (.a(_13421_),
    .b(_13494_),
    .c(_13390_),
    .d(net666),
    .o1(_15700_));
 b15aoi012ar1n06x5 _24485_ (.a(_15700_),
    .b(_13999_),
    .c(net666),
    .o1(_15701_));
 b15aoi112as1n08x5 _24486_ (.a(_15696_),
    .b(_15699_),
    .c(_13403_),
    .d(_15701_),
    .o1(_15702_));
 b15oai112al1n06x5 _24487_ (.a(net658),
    .b(_15346_),
    .c(_13382_),
    .d(_13505_),
    .o1(_15703_));
 b15oaoi13aq1n08x5 _24488_ (.a(net649),
    .b(_15703_),
    .c(_15081_),
    .d(_14378_),
    .o1(_15704_));
 b15aoai13ah1n08x5 _24489_ (.a(_13355_),
    .b(_15704_),
    .c(_13999_),
    .d(_13916_),
    .o1(_15705_));
 b15oaoi13aq1n04x5 _24490_ (.a(_13421_),
    .b(_13497_),
    .c(_13511_),
    .d(_15543_),
    .o1(_15706_));
 b15oaoi13aq1n03x5 _24491_ (.a(net657),
    .b(_13896_),
    .c(_14388_),
    .d(_13330_),
    .o1(_15707_));
 b15nand02ar1n02x5 _24492_ (.a(_13421_),
    .b(_13486_),
    .o1(_15708_));
 b15aoi112ah1n02x5 _24493_ (.a(net657),
    .b(_13939_),
    .c(_15672_),
    .d(_15708_),
    .o1(_15709_));
 b15nandp2al1n02x5 _24494_ (.a(_13415_),
    .b(_14366_),
    .o1(_15710_));
 b15oaoi13ar1n08x5 _24495_ (.a(net665),
    .b(_15710_),
    .c(_13507_),
    .d(_13313_),
    .o1(_15711_));
 b15nor004ah1n06x5 _24496_ (.a(_15706_),
    .b(_15707_),
    .c(_15709_),
    .d(_15711_),
    .o1(_15712_));
 b15oai012ah1n04x5 _24497_ (.a(\us32.a[4] ),
    .b(_15068_),
    .c(\us32.a[1] ),
    .o1(_15713_));
 b15oai012an1n04x5 _24498_ (.a(_15068_),
    .b(_13523_),
    .c(_13340_),
    .o1(_15714_));
 b15aoi022as1n08x5 _24499_ (.a(_13421_),
    .b(_15713_),
    .c(_15714_),
    .d(_13489_),
    .o1(_15715_));
 b15nandp3aq1n02x5 _24500_ (.a(net657),
    .b(_13949_),
    .c(_13540_),
    .o1(_15716_));
 b15oaoi13al1n04x5 _24501_ (.a(_15716_),
    .b(_13390_),
    .c(_13371_),
    .d(_15100_),
    .o1(_15717_));
 b15aoi022ar1n16x5 _24502_ (.a(_13362_),
    .b(_13430_),
    .c(_13518_),
    .d(_13410_),
    .o1(_15718_));
 b15oai013as1n08x5 _24503_ (.a(_14578_),
    .b(_15718_),
    .c(_13423_),
    .d(_14363_),
    .o1(_15719_));
 b15nor004as1n08x5 _24504_ (.a(_13964_),
    .b(_15715_),
    .c(_15717_),
    .d(_15719_),
    .o1(_15720_));
 b15oaoi13ar1n02x5 _24505_ (.a(_13340_),
    .b(_13421_),
    .c(_13938_),
    .d(net667),
    .o1(_15721_));
 b15oai012ar1n02x5 _24506_ (.a(net657),
    .b(_13361_),
    .c(_13938_),
    .o1(_15722_));
 b15oaoi13ar1n02x5 _24507_ (.a(_13355_),
    .b(_13421_),
    .c(_13361_),
    .d(_13340_),
    .o1(_15723_));
 b15nor003aq1n03x5 _24508_ (.a(_15721_),
    .b(_15722_),
    .c(_15723_),
    .o1(_15724_));
 b15nano23al1n03x5 _24509_ (.a(_14527_),
    .b(_14528_),
    .c(_15724_),
    .d(_13527_),
    .out0(_15725_));
 b15nand04aq1n08x5 _24510_ (.a(_15705_),
    .b(_15712_),
    .c(_15720_),
    .d(_15725_),
    .o1(_15726_));
 b15nor004as1n12x5 _24511_ (.a(_15686_),
    .b(_15694_),
    .c(_15702_),
    .d(_15726_),
    .o1(_15727_));
 b15xor002ah1n04x5 _24512_ (.a(_15670_),
    .b(_15727_),
    .out0(_15728_));
 b15aoi012ar1n02x5 _24513_ (.a(net898),
    .b(_12789_),
    .c(net903),
    .o1(_15729_));
 b15oai012ar1n02x5 _24514_ (.a(_14177_),
    .b(_12789_),
    .c(_13809_),
    .o1(_15730_));
 b15aoai13ar1n02x5 _24515_ (.a(net907),
    .b(_15729_),
    .c(_15730_),
    .d(_12875_),
    .o1(_15731_));
 b15norp02ar1n02x5 _24516_ (.a(net912),
    .b(_14658_),
    .o1(_15732_));
 b15and002an1n02x5 _24517_ (.a(_15731_),
    .b(_15732_),
    .o(_15733_));
 b15oai112an1n04x5 _24518_ (.a(_13798_),
    .b(_14143_),
    .c(_13835_),
    .d(net912),
    .o1(_15734_));
 b15aoi122ar1n06x5 _24519_ (.a(_12950_),
    .b(net905),
    .c(_14153_),
    .d(_12825_),
    .e(_13794_),
    .o1(_15735_));
 b15nor003al1n02x5 _24520_ (.a(net903),
    .b(_14152_),
    .c(_13011_),
    .o1(_15736_));
 b15aoi112ar1n03x5 _24521_ (.a(net912),
    .b(_15736_),
    .c(_12825_),
    .d(net903),
    .o1(_15737_));
 b15oai112aq1n08x5 _24522_ (.a(net898),
    .b(_15734_),
    .c(_15735_),
    .d(_15737_),
    .o1(_15738_));
 b15aob012aq1n02x5 _24523_ (.a(net907),
    .b(_12924_),
    .c(_13793_),
    .out0(_15739_));
 b15oai012an1n08x5 _24524_ (.a(_15739_),
    .b(_13769_),
    .c(_12827_),
    .o1(_15740_));
 b15oaoi13as1n08x5 _24525_ (.a(_15733_),
    .b(_15738_),
    .c(_15740_),
    .d(net898),
    .o1(_15741_));
 b15nand04as1n02x5 _24526_ (.a(_12904_),
    .b(_12879_),
    .c(_12940_),
    .d(_14233_),
    .o1(_15742_));
 b15oai013ah1n06x5 _24527_ (.a(_15742_),
    .b(_13015_),
    .c(_12973_),
    .d(_14628_),
    .o1(_15743_));
 b15oai013ah1n04x5 _24528_ (.a(_14639_),
    .b(_12922_),
    .c(_12870_),
    .d(net887),
    .o1(_15744_));
 b15nano23al1n06x5 _24529_ (.a(_12998_),
    .b(_15744_),
    .c(net900),
    .d(_12877_),
    .out0(_15745_));
 b15aoi012as1n02x5 _24530_ (.a(_14956_),
    .b(_12987_),
    .c(_13882_),
    .o1(_15746_));
 b15nona23aq1n04x5 _24531_ (.a(_13009_),
    .b(_15746_),
    .c(_12986_),
    .d(_12864_),
    .out0(_15747_));
 b15nand04ah1n12x5 _24532_ (.a(_13882_),
    .b(_12964_),
    .c(_12798_),
    .d(_13871_),
    .o1(_15748_));
 b15norp02ar1n04x5 _24533_ (.a(net894),
    .b(_13015_),
    .o1(_15749_));
 b15aoi022an1n06x5 _24534_ (.a(_12968_),
    .b(_13013_),
    .c(_13809_),
    .d(_12863_),
    .o1(_15750_));
 b15oai122as1n12x5 _24535_ (.a(_15747_),
    .b(_15748_),
    .c(_15749_),
    .d(_15750_),
    .e(_12782_),
    .o1(_15751_));
 b15nor004al1n03x5 _24536_ (.a(_12870_),
    .b(_12877_),
    .c(_12922_),
    .d(_14198_),
    .o1(_15752_));
 b15aoai13aq1n04x5 _24537_ (.a(_13827_),
    .b(_15752_),
    .c(_14210_),
    .d(_12796_),
    .o1(_15753_));
 b15nandp3ar1n02x5 _24538_ (.a(_12863_),
    .b(_12922_),
    .c(_12789_),
    .o1(_15754_));
 b15oai112ar1n02x5 _24539_ (.a(_12968_),
    .b(_12922_),
    .c(_12789_),
    .d(_13809_),
    .o1(_15755_));
 b15and002aq1n02x5 _24540_ (.a(_15754_),
    .b(_15755_),
    .o(_15756_));
 b15nor004ah1n03x5 _24541_ (.a(net892),
    .b(_13797_),
    .c(_13860_),
    .d(_14184_),
    .o1(_15757_));
 b15oai012al1n06x5 _24542_ (.a(_12913_),
    .b(_12827_),
    .c(_12950_),
    .o1(_15758_));
 b15aoi013aq1n08x5 _24543_ (.a(_15757_),
    .b(_15758_),
    .c(net892),
    .d(net899),
    .o1(_15759_));
 b15oai112as1n12x5 _24544_ (.a(_15753_),
    .b(_15756_),
    .c(_14899_),
    .d(_15759_),
    .o1(_15760_));
 b15nor004as1n12x5 _24545_ (.a(_15743_),
    .b(_15745_),
    .c(_15751_),
    .d(_15760_),
    .o1(_15761_));
 b15aoai13ar1n02x5 _24546_ (.a(_12820_),
    .b(_12851_),
    .c(_12883_),
    .d(_12798_),
    .o1(_15762_));
 b15aoi112ar1n02x5 _24547_ (.a(net898),
    .b(_12959_),
    .c(_13809_),
    .d(net912),
    .o1(_15763_));
 b15oaoi13al1n02x5 _24548_ (.a(_15762_),
    .b(_15763_),
    .c(_13801_),
    .d(_13007_),
    .o1(_15764_));
 b15nand03aq1n02x5 _24549_ (.a(_12874_),
    .b(_12904_),
    .c(_12879_),
    .o1(_15765_));
 b15oaoi13al1n02x5 _24550_ (.a(_13783_),
    .b(_15765_),
    .c(_13015_),
    .d(_14173_),
    .o1(_15766_));
 b15norp03ar1n02x5 _24551_ (.a(net898),
    .b(_12857_),
    .c(_12879_),
    .o1(_15767_));
 b15oaoi13ah1n02x5 _24552_ (.a(_15764_),
    .b(net903),
    .c(_15766_),
    .d(_15767_),
    .o1(_15768_));
 b15nonb03al1n02x5 _24553_ (.a(net908),
    .b(net894),
    .c(net892),
    .out0(_15769_));
 b15aoai13as1n04x5 _24554_ (.a(_13844_),
    .b(_15769_),
    .c(_12796_),
    .d(_13015_),
    .o1(_15770_));
 b15oai112an1n04x5 _24555_ (.a(net899),
    .b(_15770_),
    .c(_14910_),
    .d(_12917_),
    .o1(_15771_));
 b15norp02ar1n02x5 _24556_ (.a(_12865_),
    .b(_12977_),
    .o1(_15772_));
 b15aob012as1n02x5 _24557_ (.a(_14963_),
    .b(_15362_),
    .c(_15772_),
    .out0(_15773_));
 b15aoi022ar1n02x5 _24558_ (.a(net894),
    .b(_13859_),
    .c(_12940_),
    .d(_12971_),
    .o1(_15774_));
 b15nand02ar1n02x5 _24559_ (.a(_12782_),
    .b(_12983_),
    .o1(_15775_));
 b15oai022aq1n02x5 _24560_ (.a(_12877_),
    .b(_13805_),
    .c(_15774_),
    .d(_15775_),
    .o1(_15776_));
 b15oai013as1n06x5 _24561_ (.a(_15771_),
    .b(_15773_),
    .c(_15776_),
    .d(net899),
    .o1(_15777_));
 b15norp02aq1n02x5 _24562_ (.a(_12857_),
    .b(_12913_),
    .o1(_15778_));
 b15aoi112as1n04x5 _24563_ (.a(net898),
    .b(_15778_),
    .c(_13786_),
    .d(_14942_),
    .o1(_15779_));
 b15aoi022ar1n08x5 _24564_ (.a(_12877_),
    .b(_13013_),
    .c(_12789_),
    .d(_14591_),
    .o1(_15780_));
 b15aoi122ah1n02x5 _24565_ (.a(_12851_),
    .b(_12922_),
    .c(_13013_),
    .d(_13817_),
    .e(_12950_),
    .o1(_15781_));
 b15nona22al1n02x5 _24566_ (.a(net893),
    .b(net909),
    .c(net886),
    .out0(_15782_));
 b15nanb02ar1n04x5 _24567_ (.a(net886),
    .b(net893),
    .out0(_15783_));
 b15oaoi13al1n04x5 _24568_ (.a(_15368_),
    .b(_15782_),
    .c(_15783_),
    .d(_12910_),
    .o1(_15784_));
 b15nanb03ar1n03x5 _24569_ (.a(net896),
    .b(net886),
    .c(net893),
    .out0(_15785_));
 b15oai013ar1n06x5 _24570_ (.a(_15785_),
    .b(_13770_),
    .c(_12820_),
    .d(net886),
    .o1(_15786_));
 b15aoi022an1n12x5 _24571_ (.a(\us10.a[6] ),
    .b(_15784_),
    .c(_15786_),
    .d(_13850_),
    .o1(_15787_));
 b15aoi022ah1n06x5 _24572_ (.a(_15779_),
    .b(_15780_),
    .c(_15781_),
    .d(_15787_),
    .o1(_15788_));
 b15nand03aq1n03x5 _24573_ (.a(net898),
    .b(_13794_),
    .c(_12957_),
    .o1(_15789_));
 b15aoi012ar1n02x5 _24574_ (.a(net886),
    .b(net889),
    .c(net901),
    .o1(_15790_));
 b15aoi022al1n02x5 _24575_ (.a(_12881_),
    .b(_13786_),
    .c(_15790_),
    .d(net911),
    .o1(_15791_));
 b15nand02ar1n02x5 _24576_ (.a(net901),
    .b(_13843_),
    .o1(_15792_));
 b15oa0022al1n04x5 _24577_ (.a(_12865_),
    .b(_15791_),
    .c(_15792_),
    .d(_13007_),
    .o(_15793_));
 b15aoai13aq1n03x5 _24578_ (.a(_13794_),
    .b(_12825_),
    .c(_13817_),
    .d(_12950_),
    .o1(_15794_));
 b15aoai13ah1n06x5 _24579_ (.a(_15789_),
    .b(net898),
    .c(_15793_),
    .d(_15794_),
    .o1(_15795_));
 b15nano23ar1n12x5 _24580_ (.a(_15768_),
    .b(_15777_),
    .c(_15788_),
    .d(_15795_),
    .out0(_15796_));
 b15nandp3as1n24x5 _24581_ (.a(_15741_),
    .b(_15761_),
    .c(_15796_),
    .o1(_15797_));
 b15xor002as1n16x5 _24582_ (.a(_13663_),
    .b(_15797_),
    .out0(_15798_));
 b15xor002ar1n12x5 _24583_ (.a(_15728_),
    .b(_15798_),
    .out0(_15799_));
 b15orn002as1n02x5 _24584_ (.a(_15491_),
    .b(_15799_),
    .o(_15800_));
 b15nandp2al1n04x5 _24585_ (.a(_15491_),
    .b(_15799_),
    .o1(_15801_));
 b15aoi013as1n08x5 _24586_ (.a(_15619_),
    .b(_15800_),
    .c(_15801_),
    .d(_15618_),
    .o1(_15802_));
 b15xor002ar1n02x5 _24587_ (.a(net492),
    .b(_15802_),
    .out0(_00128_));
 b15bfn001as1n64x5 load_slew406 (.a(\u0.tmp_w[31] ),
    .o(net406));
 b15xor002as1n12x5 _24589_ (.a(_13546_),
    .b(_15670_),
    .out0(_15804_));
 b15xor003aq1n16x5 _24590_ (.a(_13020_),
    .b(net402),
    .c(_15804_),
    .out0(_15805_));
 b15norp02ah1n04x5 _24591_ (.a(ld_r),
    .b(_15805_),
    .o1(_15806_));
 b15inv000al1n06x5 _24592_ (.a(\text_in_r[8] ),
    .o1(_15807_));
 b15bfn001ah1n64x5 load_slew405 (.a(\u0.tmp_w[31] ),
    .o(net405));
 b15aoi012ah1n12x5 _24594_ (.a(_15806_),
    .b(_15807_),
    .c(ld_r),
    .o1(_15809_));
 b15xor002aq1n16x5 _24595_ (.a(net490),
    .b(_15809_),
    .out0(_00089_));
 b15inv000ah1n03x5 _24596_ (.a(\text_in_r[9] ),
    .o1(_15810_));
 b15xnr002as1n12x5 _24597_ (.a(_13297_),
    .b(net402),
    .out0(_15811_));
 b15xor002an1n04x5 _24598_ (.a(_15804_),
    .b(_15811_),
    .out0(_15812_));
 b15qgbxo2an1n05x5 _24599_ (.a(_13892_),
    .b(_14424_),
    .out0(_15813_));
 b15xor002al1n06x5 _24600_ (.a(_15812_),
    .b(_15813_),
    .out0(_15814_));
 b15mdn022aq1n08x5 _24601_ (.a(_15810_),
    .b(_15814_),
    .o1(_15815_),
    .sa(net533));
 b15xor002as1n12x5 _24602_ (.a(\u0.tmp_w[9] ),
    .b(_15815_),
    .out0(_00090_));
 b15inv040ah1n02x5 _24603_ (.a(\text_in_r[10] ),
    .o1(_15816_));
 b15xnr002ah1n12x5 _24604_ (.a(_14136_),
    .b(_14424_),
    .out0(_15817_));
 b15xor002ah1n03x5 _24605_ (.a(_14247_),
    .b(_15817_),
    .out0(_15818_));
 b15xor002ar1n08x5 _24606_ (.a(_14586_),
    .b(_15818_),
    .out0(_15819_));
 b15mdn022al1n02x5 _24607_ (.a(_15816_),
    .b(_15819_),
    .o1(_15820_),
    .sa(net534));
 b15xor002ar1n02x5 _24608_ (.a(\u0.tmp_w[10] ),
    .b(_15820_),
    .out0(_00091_));
 b15nanb02aq1n06x5 _24609_ (.a(\text_in_r[11] ),
    .b(net534),
    .out0(_15821_));
 b15xor002al1n12x5 _24610_ (.a(_14826_),
    .b(_15670_),
    .out0(_15822_));
 b15xor002as1n12x5 _24611_ (.a(_14337_),
    .b(_15822_),
    .out0(_15823_));
 b15xor002ar1n02x5 _24612_ (.a(_14585_),
    .b(_14673_),
    .out0(_15824_));
 b15xor002aq1n02x5 _24613_ (.a(_15107_),
    .b(_15824_),
    .out0(_15825_));
 b15xor002aq1n03x5 _24614_ (.a(_15823_),
    .b(_15825_),
    .out0(_15826_));
 b15oai012ar1n12x5 _24615_ (.a(_15821_),
    .b(_15826_),
    .c(net534),
    .o1(_15827_));
 b15xor002as1n02x5 _24616_ (.a(_10939_),
    .b(_15827_),
    .out0(_00092_));
 b15inv000aq1n04x5 _24617_ (.a(\text_in_r[12] ),
    .o1(_15828_));
 b15xor002ar1n08x5 _24618_ (.a(_14973_),
    .b(_15107_),
    .out0(_15829_));
 b15xor002as1n06x5 _24619_ (.a(_14763_),
    .b(_15670_),
    .out0(_15830_));
 b15xor002ar1n16x5 _24620_ (.a(_15352_),
    .b(_15830_),
    .out0(_15831_));
 b15xor002as1n06x5 _24621_ (.a(_15829_),
    .b(_15831_),
    .out0(_15832_));
 b15bfn001as1n48x5 wire404 (.a(net406),
    .o(net404));
 b15bfn001ah1n24x5 wire403 (.a(_08706_),
    .o(net403));
 b15mdn022al1n12x5 _24624_ (.a(_15828_),
    .b(_15832_),
    .o1(_15835_),
    .sa(net534));
 b15xor002as1n12x5 _24625_ (.a(net475),
    .b(_15835_),
    .out0(_00093_));
 b15xor003ar1n03x5 _24626_ (.a(_14898_),
    .b(_15351_),
    .c(_15552_),
    .out0(_15836_));
 b15xor002ar1n02x5 _24627_ (.a(_15232_),
    .b(_15836_),
    .out0(_15837_));
 b15nor002ar1n03x5 _24628_ (.a(net534),
    .b(_15837_),
    .o1(_15838_));
 b15inv040ah1n02x5 _24629_ (.a(\text_in_r[13] ),
    .o1(_15839_));
 b15aoi012as1n06x5 _24630_ (.a(_15838_),
    .b(_15839_),
    .c(net534),
    .o1(_15840_));
 b15xor002as1n12x5 _24631_ (.a(\u0.tmp_w[13] ),
    .b(_15840_),
    .out0(_00094_));
 b15xnr002ah1n08x5 _24632_ (.a(_15288_),
    .b(_15552_),
    .out0(_15841_));
 b15xor003an1n02x5 _24633_ (.a(_15492_),
    .b(_15727_),
    .c(_15841_),
    .out0(_15842_));
 b15nor002aq1n03x5 _24634_ (.a(net534),
    .b(_15842_),
    .o1(_15843_));
 b15inv040ah1n03x5 _24635_ (.a(\text_in_r[14] ),
    .o1(_15844_));
 b15aoi012al1n12x5 _24636_ (.a(_15843_),
    .b(_15844_),
    .c(net534),
    .o1(_15845_));
 b15xor002ah1n16x5 _24637_ (.a(\u0.tmp_w[14] ),
    .b(_15845_),
    .out0(_00095_));
 b15xor002as1n12x5 _24638_ (.a(_15614_),
    .b(_15727_),
    .out0(_15846_));
 b15xor003al1n03x5 _24639_ (.a(_13546_),
    .b(_15798_),
    .c(_15846_),
    .out0(_15847_));
 b15nor002as1n03x5 _24640_ (.a(net533),
    .b(_15847_),
    .o1(_15848_));
 b15inv020as1n04x5 _24641_ (.a(\text_in_r[15] ),
    .o1(_15849_));
 b15aoi012al1n12x5 _24642_ (.a(_15848_),
    .b(_15849_),
    .c(net533),
    .o1(_15850_));
 b15xor002ah1n16x5 _24643_ (.a(\u0.tmp_w[15] ),
    .b(_15850_),
    .out0(_00096_));
 b15bfn001ah1n32x5 wire402 (.a(_14019_),
    .o(net402));
 b15inv040ah1n02x5 _24645_ (.a(\text_in_r[16] ),
    .o1(_15852_));
 b15nand02ar1n02x5 _24646_ (.a(net541),
    .b(_15852_),
    .o1(_15853_));
 b15xor002as1n16x5 _24647_ (.a(_15670_),
    .b(_15797_),
    .out0(_15854_));
 b15xor002aq1n12x5 _24648_ (.a(_12776_),
    .b(_15854_),
    .out0(_15855_));
 b15xor002as1n16x5 _24649_ (.a(_15811_),
    .b(_15855_),
    .out0(_15856_));
 b15oai012as1n03x5 _24650_ (.a(_15853_),
    .b(_15856_),
    .c(net541),
    .o1(_15857_));
 b15qgbxo2an1n05x5 _24651_ (.a(_11579_),
    .b(_15857_),
    .out0(_00057_));
 b15nanb02an1n12x5 _24652_ (.a(\text_in_r[17] ),
    .b(net542),
    .out0(_15858_));
 b15xor002an1n12x5 _24653_ (.a(_15817_),
    .b(_15854_),
    .out0(_15859_));
 b15xor002ah1n04x5 _24654_ (.a(_13019_),
    .b(_13768_),
    .out0(_15860_));
 b15xor002as1n08x5 _24655_ (.a(_13297_),
    .b(_15860_),
    .out0(_15861_));
 b15xor002as1n16x5 _24656_ (.a(_15859_),
    .b(_15861_),
    .out0(_15862_));
 b15oai012ar1n02x5 _24657_ (.a(_15858_),
    .b(_15862_),
    .c(net541),
    .o1(_15863_));
 b15xor002ar1n02x5 _24658_ (.a(_11696_),
    .b(_15863_),
    .out0(_00058_));
 b15inv040as1n02x5 _24659_ (.a(\text_in_r[18] ),
    .o1(_15864_));
 b15nandp2ar1n12x5 _24660_ (.a(net542),
    .b(_15864_),
    .o1(_15865_));
 b15xor002as1n06x5 _24661_ (.a(_14136_),
    .b(_14337_),
    .out0(_15866_));
 b15xor002as1n08x5 _24662_ (.a(_14586_),
    .b(_15866_),
    .out0(_15867_));
 b15xor002as1n12x5 _24663_ (.a(_13891_),
    .b(_15867_),
    .out0(_15868_));
 b15oai012ar1n02x5 _24664_ (.a(_15865_),
    .b(_15868_),
    .c(net541),
    .o1(_15869_));
 b15xor002al1n02x5 _24665_ (.a(_11603_),
    .b(_15869_),
    .out0(_00059_));
 b15nanb02aq1n12x5 _24666_ (.a(\text_in_r[19] ),
    .b(net542),
    .out0(_15870_));
 b15xnr002as1n06x5 _24667_ (.a(_14247_),
    .b(_15106_),
    .out0(_15871_));
 b15xor002ah1n04x5 _24668_ (.a(_14763_),
    .b(_15797_),
    .out0(_15872_));
 b15xor002as1n08x5 _24669_ (.a(_15871_),
    .b(_15872_),
    .out0(_15873_));
 b15xor002as1n16x5 _24670_ (.a(_15823_),
    .b(_15873_),
    .out0(_15874_));
 b15oai012ar1n02x5 _24671_ (.a(_15870_),
    .b(_15874_),
    .c(net541),
    .o1(_15875_));
 b15xor002ar1n02x5 _24672_ (.a(_11666_),
    .b(_15875_),
    .out0(_00060_));
 b15inv040ah1n02x5 _24673_ (.a(\text_in_r[20] ),
    .o1(_15876_));
 b15xnr002aq1n12x5 _24674_ (.a(_15352_),
    .b(_15854_),
    .out0(_15877_));
 b15xor002aq1n12x5 _24675_ (.a(_14764_),
    .b(_14898_),
    .out0(_15878_));
 b15xor002as1n16x5 _24676_ (.a(_15877_),
    .b(_15878_),
    .out0(_15879_));
 b15mdn022ah1n03x5 _24677_ (.a(_15876_),
    .b(_15879_),
    .o1(_15880_),
    .sa(net542));
 b15xor002ar1n06x5 _24678_ (.a(\u0.tmp_w[20] ),
    .b(_15880_),
    .out0(_00061_));
 b15xor003ah1n06x5 _24679_ (.a(_14974_),
    .b(_15231_),
    .c(_15841_),
    .out0(_15881_));
 b15norp02aq1n24x5 _24680_ (.a(net534),
    .b(_15881_),
    .o1(_15882_));
 b15inv040as1n10x5 _24681_ (.a(\text_in_r[21] ),
    .o1(_15883_));
 b15aoi012ar1n02x5 _24682_ (.a(_15882_),
    .b(_15883_),
    .c(net541),
    .o1(_15884_));
 b15xor002ar1n02x5 _24683_ (.a(\u0.tmp_w[21] ),
    .b(_15884_),
    .out0(_00062_));
 b15inv040ah1n06x5 _24684_ (.a(\text_in_r[22] ),
    .o1(_15885_));
 b15xor002ah1n04x5 _24685_ (.a(_15288_),
    .b(_15491_),
    .out0(_15886_));
 b15xor002as1n08x5 _24686_ (.a(_15173_),
    .b(_15886_),
    .out0(_15887_));
 b15xor002as1n16x5 _24687_ (.a(_15846_),
    .b(_15887_),
    .out0(_15888_));
 b15mdn022al1n02x5 _24688_ (.a(_15885_),
    .b(_15888_),
    .o1(_15889_),
    .sa(net542));
 b15xor002ar1n02x5 _24689_ (.a(\u0.tmp_w[22] ),
    .b(_15889_),
    .out0(_00063_));
 b15xor003ah1n06x5 _24690_ (.a(_15614_),
    .b(_15428_),
    .c(_15670_),
    .out0(_15890_));
 b15xor002as1n06x5 _24691_ (.a(_13664_),
    .b(_15890_),
    .out0(_15891_));
 b15nor002aq1n16x5 _24692_ (.a(net534),
    .b(_15891_),
    .o1(_15892_));
 b15inv040ah1n02x5 _24693_ (.a(\text_in_r[23] ),
    .o1(_15893_));
 b15aoi012ar1n02x5 _24694_ (.a(_15892_),
    .b(_15893_),
    .c(net542),
    .o1(_15894_));
 b15xor002ar1n02x5 _24695_ (.a(\u0.tmp_w[23] ),
    .b(_15894_),
    .out0(_00064_));
 b15inv040ah1n05x5 _24696_ (.a(\text_in_r[24] ),
    .o1(_15895_));
 b15xor002ah1n02x5 _24697_ (.a(_13019_),
    .b(_15811_),
    .out0(_15896_));
 b15xor002ar1n06x5 _24698_ (.a(_15798_),
    .b(_15896_),
    .out0(_15897_));
 b15mdn022ah1n06x5 _24699_ (.a(_15895_),
    .b(_15897_),
    .o1(_15898_),
    .sa(net534));
 b15xor002an1n12x5 _24700_ (.a(net429),
    .b(_15898_),
    .out0(_00025_));
 b15nanb02ar1n02x5 _24701_ (.a(\text_in_r[25] ),
    .b(net533),
    .out0(_15899_));
 b15xor002aq1n02x5 _24702_ (.a(_13020_),
    .b(_15798_),
    .out0(_15900_));
 b15xor002al1n03x5 _24703_ (.a(_13891_),
    .b(_15817_),
    .out0(_15901_));
 b15xor002as1n03x5 _24704_ (.a(_15900_),
    .b(_15901_),
    .out0(_15902_));
 b15oai012as1n04x5 _24705_ (.a(_15899_),
    .b(_15902_),
    .c(net533),
    .o1(_15903_));
 b15xor002an1n08x5 _24706_ (.a(_03026_),
    .b(_15903_),
    .out0(_00026_));
 b15norp02as1n02x5 _24707_ (.a(_15618_),
    .b(\text_in_r[26] ),
    .o1(_15904_));
 b15xor002ah1n03x5 _24708_ (.a(_13892_),
    .b(_14338_),
    .out0(_15905_));
 b15and002ah1n02x5 _24709_ (.a(_14585_),
    .b(_15905_),
    .o(_15906_));
 b15norp02al1n04x5 _24710_ (.a(_14585_),
    .b(_15905_),
    .o1(_15907_));
 b15oaoi13an1n08x5 _24711_ (.a(_15904_),
    .b(_15618_),
    .c(_15906_),
    .d(_15907_),
    .o1(_15908_));
 b15xor002an1n12x5 _24712_ (.a(net422),
    .b(_15908_),
    .out0(_00027_));
 b15inv000an1n05x5 _24713_ (.a(\text_in_r[27] ),
    .o1(_15909_));
 b15xor002as1n02x5 _24714_ (.a(_14493_),
    .b(_15871_),
    .out0(_15910_));
 b15xor002ah1n02x5 _24715_ (.a(_14764_),
    .b(_15798_),
    .out0(_15911_));
 b15xor002ah1n04x5 _24716_ (.a(_15910_),
    .b(_15911_),
    .out0(_15912_));
 b15mdn022al1n12x5 _24717_ (.a(_15909_),
    .b(_15912_),
    .o1(_15913_),
    .sa(net534));
 b15xor002aq1n16x5 _24718_ (.a(net417),
    .b(_15913_),
    .out0(_00028_));
 b15nanb02ar1n02x5 _24719_ (.a(\text_in_r[28] ),
    .b(net534),
    .out0(_15914_));
 b15xor002al1n02x5 _24720_ (.a(_15351_),
    .b(_15797_),
    .out0(_15915_));
 b15xor002al1n02x5 _24721_ (.a(_14673_),
    .b(_15915_),
    .out0(_15916_));
 b15xor002ar1n03x5 _24722_ (.a(_14976_),
    .b(_15916_),
    .out0(_15917_));
 b15oai012aq1n04x5 _24723_ (.a(_15914_),
    .b(_15917_),
    .c(net534),
    .o1(_15918_));
 b15xor002aq1n06x5 _24724_ (.a(_07818_),
    .b(_15918_),
    .out0(_00029_));
 b15xor002ar1n02x5 _24725_ (.a(_14973_),
    .b(_15173_),
    .out0(_15919_));
 b15xor002al1n02x5 _24726_ (.a(_15034_),
    .b(_15919_),
    .out0(_15920_));
 b15xor002ar1n02x5 _24727_ (.a(_15841_),
    .b(_15920_),
    .out0(_15921_));
 b15bfn001ah1n32x5 wire401 (.a(_02505_),
    .o(net401));
 b15cmbn22ar1n02x5 _24729_ (.clk1(\text_in_r[29] ),
    .clk2(_15921_),
    .clkout(_15923_),
    .s(net534));
 b15xor002an1n04x5 _24730_ (.a(net413),
    .b(_15923_),
    .out0(_00030_));
 b15xor003an1n03x5 _24731_ (.a(_15232_),
    .b(_15428_),
    .c(_15846_),
    .out0(_15924_));
 b15nor002al1n02x5 _24732_ (.a(net534),
    .b(_15924_),
    .o1(_15925_));
 b15inv040ah1n02x5 _24733_ (.a(\text_in_r[30] ),
    .o1(_15926_));
 b15aoi012al1n04x5 _24734_ (.a(_15925_),
    .b(_15926_),
    .c(net534),
    .o1(_15927_));
 b15xor002an1n08x5 _24735_ (.a(net408),
    .b(_15927_),
    .out0(_00031_));
 b15xor003ar1n03x5 _24736_ (.a(_15492_),
    .b(_15797_),
    .c(_15804_),
    .out0(_15928_));
 b15norp02al1n02x5 _24737_ (.a(net534),
    .b(_15928_),
    .o1(_15929_));
 b15inv000ah1n03x5 _24738_ (.a(\text_in_r[31] ),
    .o1(_15930_));
 b15aoi012aq1n04x5 _24739_ (.a(_15929_),
    .b(_15930_),
    .c(net534),
    .o1(_15931_));
 b15qgbxo2an1n10x5 _24740_ (.a(net406),
    .b(_15931_),
    .out0(_00032_));
 b15bfn001as1n32x5 wire400 (.a(_03294_),
    .o(net400));
 b15bfn001ah1n32x5 wire399 (.a(_04133_),
    .o(net399));
 b15bfn001ah1n32x5 wire398 (.a(_04404_),
    .o(net398));
 b15bfn001as1n32x5 wire397 (.a(_04643_),
    .o(net397));
 b15bfn001as1n32x5 wire396 (.a(_05607_),
    .o(net396));
 b15bfn001ah1n48x5 wire395 (.a(_05679_),
    .o(net395));
 b15bfn001ah1n32x5 wire394 (.a(_08321_),
    .o(net394));
 b15nor002aq1n06x5 _24748_ (.a(net864),
    .b(\us20.a[6] ),
    .o1(_15939_));
 b15bfn001as1n24x5 wire393 (.a(_03931_),
    .o(net393));
 b15bfn001as1n32x5 wire392 (.a(_04015_),
    .o(net392));
 b15bfn001ah1n24x5 wire391 (.a(_11548_),
    .o(net391));
 b15nonb02as1n16x5 _24752_ (.a(net869),
    .b(\us20.a[4] ),
    .out0(_15943_));
 b15bfn001as1n16x5 wire390 (.a(_00119_),
    .o(net390));
 b15bfn001as1n16x5 wire389 (.a(_00046_),
    .o(net389));
 b15bfn001as1n16x5 wire388 (.a(_00047_),
    .o(net388));
 b15nandp2ar1n24x5 _24756_ (.a(net884),
    .b(net881),
    .o1(_15947_));
 b15aoi013aq1n08x5 _24757_ (.a(net874),
    .b(_15939_),
    .c(_15943_),
    .d(_15947_),
    .o1(_15948_));
 b15bfn000ar1n02x5 output387 (.a(net387),
    .o(text_out[9]));
 b15bfn000ar1n02x5 output386 (.a(net386),
    .o(text_out[99]));
 b15bfn000ar1n02x5 output385 (.a(net385),
    .o(text_out[98]));
 b15norp02ah1n48x5 _24761_ (.a(net868),
    .b(net870),
    .o1(_15952_));
 b15bfn000ar1n02x5 output384 (.a(net384),
    .o(text_out[97]));
 b15bfn000ar1n02x5 output383 (.a(net383),
    .o(text_out[96]));
 b15nonb02as1n16x5 _24764_ (.a(net864),
    .b(\us20.a[6] ),
    .out0(_15955_));
 b15nand03as1n06x5 _24765_ (.a(\us20.a[2] ),
    .b(_15952_),
    .c(_15955_),
    .o1(_15956_));
 b15bfn000ar1n02x5 output382 (.a(net382),
    .o(text_out[95]));
 b15bfn000ar1n02x5 output381 (.a(net381),
    .o(text_out[94]));
 b15inv040ah1n24x5 _24768_ (.a(net882),
    .o1(_15959_));
 b15bfn000ar1n02x5 output380 (.a(net380),
    .o(text_out[93]));
 b15bfn000ar1n02x5 output379 (.a(net379),
    .o(text_out[92]));
 b15bfn000ar1n02x5 output378 (.a(net378),
    .o(text_out[91]));
 b15nonb02ah1n08x5 _24772_ (.a(\us20.a[2] ),
    .b(net880),
    .out0(_15963_));
 b15aoi122al1n02x5 _24773_ (.a(_15948_),
    .b(_15956_),
    .c(net872),
    .d(_15959_),
    .e(_15963_),
    .o1(_15964_));
 b15bfn000ar1n02x5 output377 (.a(net377),
    .o(text_out[90]));
 b15bfn000ar1n02x5 output376 (.a(net376),
    .o(text_out[8]));
 b15bfn000ar1n02x5 output375 (.a(net375),
    .o(text_out[89]));
 b15bfn000ar1n02x5 output374 (.a(net374),
    .o(text_out[88]));
 b15and002as1n08x5 _24778_ (.a(net869),
    .b(\us20.a[7] ),
    .o(_15969_));
 b15norp02aq1n24x5 _24779_ (.a(net877),
    .b(net873),
    .o1(_15970_));
 b15nand03ar1n03x5 _24780_ (.a(net866),
    .b(_15969_),
    .c(_15970_),
    .o1(_15971_));
 b15bfn000ar1n02x5 output373 (.a(net373),
    .o(text_out[87]));
 b15bfn000ar1n02x5 output372 (.a(net372),
    .o(text_out[86]));
 b15nonb02as1n16x5 _24783_ (.a(net874),
    .b(net875),
    .out0(_15974_));
 b15nonb02an1n16x5 _24784_ (.a(net877),
    .b(net873),
    .out0(_15975_));
 b15nor002ah1n02x5 _24785_ (.a(net866),
    .b(\us20.a[1] ),
    .o1(_15976_));
 b15aoi022an1n02x5 _24786_ (.a(net866),
    .b(_15974_),
    .c(_15975_),
    .d(_15976_),
    .o1(_15977_));
 b15bfn000ar1n02x5 output371 (.a(net371),
    .o(text_out[85]));
 b15bfn000ar1n02x5 output370 (.a(net370),
    .o(text_out[84]));
 b15oai013ah1n04x5 _24789_ (.a(_15971_),
    .b(_15977_),
    .c(net863),
    .d(net869),
    .o1(_15980_));
 b15bfn000ar1n02x5 output369 (.a(net369),
    .o(text_out[83]));
 b15bfn000ar1n02x5 output368 (.a(net368),
    .o(text_out[82]));
 b15bfn000ar1n02x5 output367 (.a(net367),
    .o(text_out[81]));
 b15bfn000ar1n02x5 output366 (.a(net366),
    .o(text_out[80]));
 b15aoi013al1n02x5 _24794_ (.a(_15964_),
    .b(_15980_),
    .c(net883),
    .d(\us20.a[4] ),
    .o1(_15985_));
 b15bfn000ar1n02x5 output365 (.a(net365),
    .o(text_out[7]));
 b15nandp2as1n48x5 _24796_ (.a(net867),
    .b(net871),
    .o1(_15987_));
 b15nanb02as1n24x5 _24797_ (.a(net863),
    .b(net865),
    .out0(_15988_));
 b15norp02as1n12x5 _24798_ (.a(_15987_),
    .b(_15988_),
    .o1(_15989_));
 b15bfn000ar1n02x5 output364 (.a(net364),
    .o(text_out[79]));
 b15bfn000ar1n02x5 output363 (.a(net363),
    .o(text_out[78]));
 b15bfn000ar1n02x5 output362 (.a(net362),
    .o(text_out[77]));
 b15orn002ah1n32x5 _24802_ (.a(net878),
    .b(\us20.a[3] ),
    .o(_15993_));
 b15bfn000ar1n02x5 output361 (.a(net361),
    .o(text_out[76]));
 b15nand02ah1n48x5 _24804_ (.a(net878),
    .b(\us20.a[3] ),
    .o1(_15995_));
 b15bfn000ar1n02x5 output360 (.a(net360),
    .o(text_out[75]));
 b15nanb02as1n24x5 _24806_ (.a(net885),
    .b(net881),
    .out0(_15997_));
 b15bfn000ar1n02x5 output359 (.a(net359),
    .o(text_out[74]));
 b15oai022ah1n02x5 _24808_ (.a(net880),
    .b(_15993_),
    .c(_15995_),
    .d(_15997_),
    .o1(_15999_));
 b15nanb02as1n24x5 _24809_ (.a(net876),
    .b(net879),
    .out0(_16000_));
 b15oai012aq1n04x5 _24810_ (.a(_16000_),
    .b(_15995_),
    .c(net880),
    .o1(_16001_));
 b15aoai13as1n06x5 _24811_ (.a(_15989_),
    .b(_15999_),
    .c(_16001_),
    .d(net885),
    .o1(_16002_));
 b15bfn000ar1n02x5 output358 (.a(net358),
    .o(text_out[73]));
 b15ornc04as1n24x5 _24813_ (.a(net868),
    .b(net870),
    .c(net864),
    .d(\us20.a[6] ),
    .o(_16004_));
 b15bfn000ar1n02x5 output357 (.a(net357),
    .o(text_out[72]));
 b15nor002ah1n32x5 _24815_ (.a(net884),
    .b(net881),
    .o1(_16006_));
 b15nand02al1n06x5 _24816_ (.a(_15970_),
    .b(_16006_),
    .o1(_16007_));
 b15nonb02as1n16x5 _24817_ (.a(net865),
    .b(net864),
    .out0(_16008_));
 b15nandp3ah1n12x5 _24818_ (.o1(_16009_),
    .a(net872),
    .b(_15952_),
    .c(_16008_));
 b15nonb02aq1n16x5 _24819_ (.a(net877),
    .b(net884),
    .out0(_16010_));
 b15nand02an1n32x5 _24820_ (.a(net881),
    .b(net878),
    .o1(_16011_));
 b15bfn000ar1n02x5 output356 (.a(net356),
    .o(text_out[71]));
 b15aoi012as1n02x5 _24822_ (.a(_16010_),
    .b(_16011_),
    .c(net883),
    .o1(_16013_));
 b15oai022aq1n12x5 _24823_ (.a(_16004_),
    .b(_16007_),
    .c(_16009_),
    .d(_16013_),
    .o1(_16014_));
 b15bfn000ar1n02x5 output355 (.a(net355),
    .o(text_out[70]));
 b15bfn000ar1n02x5 output354 (.a(net354),
    .o(text_out[6]));
 b15bfn000ar1n02x5 output353 (.a(net353),
    .o(text_out[69]));
 b15inv020ar1n64x5 _24827_ (.a(net875),
    .o1(_16018_));
 b15bfn000ar1n02x5 output352 (.a(net352),
    .o(text_out[68]));
 b15bfn000ar1n02x5 output351 (.a(net351),
    .o(text_out[67]));
 b15nanb02as1n24x5 _24830_ (.a(net866),
    .b(net863),
    .out0(_16021_));
 b15bfn000ar1n02x5 output350 (.a(net350),
    .o(text_out[66]));
 b15nor004an1n04x5 _24832_ (.a(net885),
    .b(_16018_),
    .c(_15987_),
    .d(_16021_),
    .o1(_16023_));
 b15bfn000ar1n02x5 output349 (.a(net349),
    .o(text_out[65]));
 b15nanb02al1n12x5 _24834_ (.a(net875),
    .b(net885),
    .out0(_16025_));
 b15norp02an1n03x5 _24835_ (.a(_16004_),
    .b(_16025_),
    .o1(_16026_));
 b15oaoi13an1n04x5 _24836_ (.a(net879),
    .b(net874),
    .c(_16023_),
    .d(_16026_),
    .o1(_16027_));
 b15inv020ah1n64x5 _24837_ (.a(net874),
    .o1(_16028_));
 b15bfn000ar1n02x5 output348 (.a(net348),
    .o(text_out[64]));
 b15bfn000ar1n02x5 output347 (.a(net347),
    .o(text_out[63]));
 b15nand04as1n16x5 _24840_ (.a(net868),
    .b(net870),
    .c(net864),
    .d(\us20.a[6] ),
    .o1(_16031_));
 b15aoai13al1n02x5 _24841_ (.a(_16028_),
    .b(net875),
    .c(_16031_),
    .d(_16004_),
    .o1(_16032_));
 b15nor002ar1n08x5 _24842_ (.a(net885),
    .b(_16031_),
    .o1(_16033_));
 b15nano23ah1n24x5 _24843_ (.a(net870),
    .b(\us20.a[6] ),
    .c(net864),
    .d(net868),
    .out0(_16034_));
 b15and002ar1n02x5 _24844_ (.a(net885),
    .b(_16034_),
    .o(_16035_));
 b15bfn000ar1n02x5 output346 (.a(net346),
    .o(text_out[62]));
 b15oai013ah1n04x5 _24846_ (.a(_16032_),
    .b(_16033_),
    .c(_16035_),
    .d(_16028_),
    .o1(_16037_));
 b15bfn000ar1n02x5 output345 (.a(net345),
    .o(text_out[61]));
 b15bfn000ar1n02x5 output344 (.a(net344),
    .o(text_out[60]));
 b15nona23as1n32x5 _24849_ (.a(net868),
    .b(\us20.a[6] ),
    .c(net864),
    .d(net870),
    .out0(_16040_));
 b15bfn000ar1n02x5 output343 (.a(net343),
    .o(text_out[5]));
 b15nor002ar1n08x5 _24851_ (.a(_16040_),
    .b(_15995_),
    .o1(_16042_));
 b15bfn000ar1n02x5 output342 (.a(net342),
    .o(text_out[59]));
 b15nor003as1n08x5 _24853_ (.a(net885),
    .b(net876),
    .c(net873),
    .o1(_16044_));
 b15nano23as1n24x5 _24854_ (.a(net870),
    .b(net864),
    .c(\us20.a[6] ),
    .d(net868),
    .out0(_16045_));
 b15bfn000ar1n02x5 output341 (.a(net341),
    .o(text_out[58]));
 b15nano23as1n24x5 _24856_ (.a(net864),
    .b(\us20.a[6] ),
    .c(net868),
    .d(net870),
    .out0(_16047_));
 b15bfn000ar1n02x5 output340 (.a(net340),
    .o(text_out[57]));
 b15oaoi13as1n08x5 _24858_ (.a(_16042_),
    .b(_16044_),
    .c(_16045_),
    .d(_16047_),
    .o1(_16049_));
 b15bfn000ar1n02x5 output339 (.a(net339),
    .o(text_out[56]));
 b15bfn000ar1n02x5 output338 (.a(net338),
    .o(text_out[55]));
 b15aoi013ar1n08x5 _24861_ (.a(_16027_),
    .b(_16037_),
    .c(_16049_),
    .d(net879),
    .o1(_16052_));
 b15nano23ah1n06x5 _24862_ (.a(_15985_),
    .b(_16002_),
    .c(_16014_),
    .d(_16052_),
    .out0(_16053_));
 b15bfn000ar1n02x5 output337 (.a(net337),
    .o(text_out[54]));
 b15bfn000ar1n02x5 output336 (.a(net336),
    .o(text_out[53]));
 b15bfn000ar1n02x5 output335 (.a(net335),
    .o(text_out[52]));
 b15bfn000ar1n02x5 output334 (.a(net334),
    .o(text_out[51]));
 b15nano23as1n24x5 _24867_ (.a(net868),
    .b(\us20.a[6] ),
    .c(net864),
    .d(net870),
    .out0(_16058_));
 b15bfn000ar1n02x5 output333 (.a(net333),
    .o(text_out[50]));
 b15nona23aq1n16x5 _24869_ (.a(\us20.a[4] ),
    .b(net864),
    .c(net866),
    .d(net869),
    .out0(_16060_));
 b15nanb02as1n24x5 _24870_ (.a(net879),
    .b(net875),
    .out0(_16061_));
 b15oai012an1n02x5 _24871_ (.a(_16060_),
    .b(_16061_),
    .c(_16004_),
    .o1(_16062_));
 b15bfn000ar1n02x5 output332 (.a(net332),
    .o(text_out[4]));
 b15aoi022al1n06x5 _24873_ (.a(\us20.a[2] ),
    .b(_16058_),
    .c(_16062_),
    .d(net883),
    .o1(_16064_));
 b15and002as1n16x5 _24874_ (.a(net868),
    .b(net870),
    .o(_16065_));
 b15nor002an1n24x5 _24875_ (.a(net882),
    .b(net875),
    .o1(_16066_));
 b15nand03ar1n24x5 _24876_ (.a(_16065_),
    .b(_15955_),
    .c(_16066_),
    .o1(_16067_));
 b15nor003ar1n12x5 _24877_ (.a(\us20.a[2] ),
    .b(_15987_),
    .c(_16021_),
    .o1(_16068_));
 b15nor004as1n12x5 _24878_ (.a(net869),
    .b(\us20.a[4] ),
    .c(\us20.a[7] ),
    .d(net866),
    .o1(_16069_));
 b15bfn000ar1n02x5 output331 (.a(net331),
    .o(text_out[49]));
 b15aoai13as1n02x5 _24880_ (.a(net880),
    .b(_16068_),
    .c(_16069_),
    .d(\us20.a[2] ),
    .o1(_16071_));
 b15aoi013an1n04x5 _24881_ (.a(net872),
    .b(_16064_),
    .c(_16067_),
    .d(_16071_),
    .o1(_16072_));
 b15bfn000ar1n02x5 output330 (.a(net330),
    .o(text_out[48]));
 b15and002aq1n04x5 _24883_ (.a(_16028_),
    .b(_16034_),
    .o(_16074_));
 b15norp02an1n16x5 _24884_ (.a(_16028_),
    .b(_16060_),
    .o1(_16075_));
 b15oai112aq1n16x5 _24885_ (.a(_16018_),
    .b(_15997_),
    .c(_16074_),
    .d(_16075_),
    .o1(_16076_));
 b15nand02ah1n32x5 _24886_ (.a(net884),
    .b(net877),
    .o1(_16077_));
 b15inv040aq1n60x5 _24887_ (.a(net879),
    .o1(_16078_));
 b15bfn000ar1n02x5 output329 (.a(net329),
    .o(text_out[47]));
 b15orn002as1n32x5 _24889_ (.a(net863),
    .b(net865),
    .o(_16080_));
 b15bfn000ar1n02x5 output328 (.a(net328),
    .o(text_out[46]));
 b15nanb02as1n24x5 _24891_ (.a(net868),
    .b(net870),
    .out0(_16082_));
 b15bfn000ar1n02x5 output327 (.a(net327),
    .o(text_out[45]));
 b15nor003ah1n06x5 _24893_ (.a(_16078_),
    .b(_16080_),
    .c(_16082_),
    .o1(_16084_));
 b15orn002aq1n24x5 _24894_ (.a(net867),
    .b(net871),
    .o(_16085_));
 b15norp03ah1n08x5 _24895_ (.a(net880),
    .b(_16085_),
    .c(_15988_),
    .o1(_16086_));
 b15oai112as1n08x5 _24896_ (.a(_16028_),
    .b(_16077_),
    .c(_16084_),
    .d(_16086_),
    .o1(_16087_));
 b15inv000an1n24x5 _24897_ (.a(net871),
    .o1(_16088_));
 b15orn002al1n08x5 _24898_ (.a(net884),
    .b(net881),
    .o(_16089_));
 b15nanb02al1n24x5 _24899_ (.a(net866),
    .b(net884),
    .out0(_16090_));
 b15aoi012al1n02x5 _24900_ (.a(_16088_),
    .b(_16089_),
    .c(_16090_),
    .o1(_16091_));
 b15inv040al1n12x5 _24901_ (.a(net866),
    .o1(_16092_));
 b15aoi012ah1n04x5 _24902_ (.a(_16091_),
    .b(_16006_),
    .c(_16092_),
    .o1(_16093_));
 b15nandp2al1n02x5 _24903_ (.a(_15969_),
    .b(_15975_),
    .o1(_16094_));
 b15oai112an1n08x5 _24904_ (.a(_16076_),
    .b(_16087_),
    .c(_16093_),
    .d(_16094_),
    .o1(_16095_));
 b15and002aq1n16x5 _24905_ (.a(\us20.a[7] ),
    .b(net866),
    .o(_16096_));
 b15bfn000ar1n02x5 output326 (.a(net326),
    .o(text_out[44]));
 b15bfn000ar1n02x5 output325 (.a(net325),
    .o(text_out[43]));
 b15bfn000ar1n02x5 output324 (.a(net324),
    .o(text_out[42]));
 b15nand02ar1n16x5 _24909_ (.a(net871),
    .b(\us20.a[3] ),
    .o1(_16100_));
 b15norp02ar1n02x5 _24910_ (.a(net867),
    .b(_16100_),
    .o1(_16101_));
 b15nor002ar1n02x5 _24911_ (.a(net871),
    .b(\us20.a[3] ),
    .o1(_16102_));
 b15aoai13ah1n03x5 _24912_ (.a(_16096_),
    .b(_16101_),
    .c(_16102_),
    .d(net867),
    .o1(_16103_));
 b15nanb02an1n16x5 _24913_ (.a(\us20.a[3] ),
    .b(\us20.a[1] ),
    .out0(_16104_));
 b15bfn000ar1n02x5 output323 (.a(net323),
    .o(text_out[41]));
 b15oai112ah1n06x5 _24915_ (.a(_15959_),
    .b(_16104_),
    .c(_15995_),
    .d(\us20.a[1] ),
    .o1(_16106_));
 b15bfn000ar1n02x5 output322 (.a(net322),
    .o(text_out[40]));
 b15oai112al1n08x5 _24917_ (.a(net884),
    .b(_16011_),
    .c(_15993_),
    .d(\us20.a[1] ),
    .o1(_16108_));
 b15aoi012ar1n08x5 _24918_ (.a(_16103_),
    .b(_16106_),
    .c(_16108_),
    .o1(_16109_));
 b15and002ar1n24x5 _24919_ (.a(net879),
    .b(net875),
    .o(_16110_));
 b15nand02al1n06x5 _24920_ (.a(_16008_),
    .b(_16110_),
    .o1(_16111_));
 b15nanb02al1n24x5 _24921_ (.a(net884),
    .b(net873),
    .out0(_16112_));
 b15nanb02as1n24x5 _24922_ (.a(net870),
    .b(net869),
    .out0(_16113_));
 b15oa0022an1n03x5 _24923_ (.a(net873),
    .b(_16082_),
    .c(_16112_),
    .d(_16113_),
    .o(_16114_));
 b15bfn000ar1n02x5 output321 (.a(net321),
    .o(text_out[3]));
 b15qgbna2an1n05x5 _24925_ (.o1(_16116_),
    .a(net863),
    .b(net873));
 b15orn002aq1n04x5 _24926_ (.a(_16113_),
    .b(_16116_),
    .o(_16117_));
 b15rm6013eq1n08x5 _24927_ (.a(net885),
    .b(net878),
    .c(_15976_),
    .carryb(_16118_));
 b15oai022aq1n16x5 _24928_ (.a(_16111_),
    .b(_16114_),
    .c(_16117_),
    .d(_16118_),
    .o1(_16119_));
 b15nor004as1n08x5 _24929_ (.a(_16072_),
    .b(_16095_),
    .c(_16109_),
    .d(_16119_),
    .o1(_16120_));
 b15bfn000ar1n02x5 output320 (.a(net320),
    .o(text_out[39]));
 b15xor002as1n03x5 _24931_ (.a(\us20.a[0] ),
    .b(net881),
    .out0(_16122_));
 b15nandp3ar1n02x5 _24932_ (.a(net878),
    .b(_16069_),
    .c(_16122_),
    .o1(_16123_));
 b15oai013ar1n02x5 _24933_ (.a(_16031_),
    .b(_16082_),
    .c(_16080_),
    .d(_16122_),
    .o1(_16124_));
 b15nona23aq1n24x5 _24934_ (.a(net864),
    .b(\us20.a[6] ),
    .c(net868),
    .d(\us20.a[4] ),
    .out0(_16125_));
 b15nandp2ah1n48x5 _24935_ (.a(net863),
    .b(net865),
    .o1(_16126_));
 b15bfn000ar1n02x5 output319 (.a(net319),
    .o(text_out[38]));
 b15oai022ar1n02x5 _24937_ (.a(\us20.a[1] ),
    .b(_16125_),
    .c(_16126_),
    .d(_16113_),
    .o1(_16128_));
 b15nanb02as1n24x5 _24938_ (.a(net881),
    .b(\us20.a[0] ),
    .out0(_16129_));
 b15aoai13ar1n02x5 _24939_ (.a(_16018_),
    .b(_16124_),
    .c(_16128_),
    .d(_16129_),
    .o1(_16130_));
 b15aob012ar1n02x5 _24940_ (.a(\us20.a[3] ),
    .b(_16123_),
    .c(_16130_),
    .out0(_16131_));
 b15nona23as1n32x5 _24941_ (.a(net868),
    .b(net870),
    .c(net864),
    .d(\us20.a[6] ),
    .out0(_16132_));
 b15norp03as1n08x5 _24942_ (.a(_16028_),
    .b(_16132_),
    .c(_16110_),
    .o1(_16133_));
 b15nanb02as1n24x5 _24943_ (.a(net878),
    .b(\us20.a[3] ),
    .out0(_16134_));
 b15nand02as1n24x5 _24944_ (.a(_15952_),
    .b(_15955_),
    .o1(_16135_));
 b15nand02al1n12x5 _24945_ (.a(_16065_),
    .b(_16008_),
    .o1(_16136_));
 b15nanb02as1n24x5 _24946_ (.a(net872),
    .b(net876),
    .out0(_16137_));
 b15oai022an1n08x5 _24947_ (.a(_16134_),
    .b(_16135_),
    .c(_16136_),
    .d(_16137_),
    .o1(_16138_));
 b15nor003aq1n03x5 _24948_ (.a(net880),
    .b(_15993_),
    .c(_16040_),
    .o1(_16139_));
 b15oai013al1n08x5 _24949_ (.a(net883),
    .b(_16133_),
    .c(_16138_),
    .d(_16139_),
    .o1(_16140_));
 b15nor002as1n06x5 _24950_ (.a(\us20.a[3] ),
    .b(_16125_),
    .o1(_16141_));
 b15aoai13an1n02x5 _24951_ (.a(\us20.a[1] ),
    .b(_16141_),
    .c(_16069_),
    .d(\us20.a[3] ),
    .o1(_16142_));
 b15aoi012al1n02x5 _24952_ (.a(\us20.a[2] ),
    .b(_16141_),
    .c(net885),
    .o1(_16143_));
 b15norp03ar1n02x5 _24953_ (.a(net885),
    .b(_16028_),
    .c(_16132_),
    .o1(_16144_));
 b15nor002ar1n16x5 _24954_ (.a(net885),
    .b(_16078_),
    .o1(_16145_));
 b15aoi012an1n02x5 _24955_ (.a(_16144_),
    .b(_16141_),
    .c(_16145_),
    .o1(_16146_));
 b15nano23as1n24x5 _24956_ (.a(net868),
    .b(net870),
    .c(net864),
    .d(\us20.a[6] ),
    .out0(_16147_));
 b15aoi013aq1n02x5 _24957_ (.a(_16018_),
    .b(\us20.a[3] ),
    .c(_15997_),
    .d(_16147_),
    .o1(_16148_));
 b15aoi022an1n06x5 _24958_ (.a(_16142_),
    .b(_16143_),
    .c(_16146_),
    .d(_16148_),
    .o1(_16149_));
 b15orn002aq1n04x5 _24959_ (.a(net871),
    .b(net866),
    .o(_16150_));
 b15bfn000ar1n02x5 output318 (.a(net318),
    .o(text_out[37]));
 b15nanb03an1n02x5 _24961_ (.a(\us20.a[7] ),
    .b(\us20.a[3] ),
    .c(net867),
    .out0(_16152_));
 b15nanb02aq1n12x5 _24962_ (.a(\us20.a[3] ),
    .b(\us20.a[7] ),
    .out0(_16153_));
 b15bfn000ar1n02x5 output317 (.a(net317),
    .o(text_out[36]));
 b15oaoi13an1n04x5 _24964_ (.a(_16150_),
    .b(_16152_),
    .c(_16153_),
    .d(net867),
    .o1(_16155_));
 b15aoi012as1n02x5 _24965_ (.a(_16089_),
    .b(_16155_),
    .c(_16134_),
    .o1(_16156_));
 b15bfn000ar1n02x5 output316 (.a(net316),
    .o(text_out[35]));
 b15norp02aq1n04x5 _24967_ (.a(net884),
    .b(_15975_),
    .o1(_16158_));
 b15aoi112an1n04x5 _24968_ (.a(_16078_),
    .b(_16158_),
    .c(_16155_),
    .d(net884),
    .o1(_16159_));
 b15and002ah1n12x5 _24969_ (.a(net877),
    .b(net873),
    .o(_16160_));
 b15aoai13al1n02x5 _24970_ (.a(net884),
    .b(_15970_),
    .c(_16160_),
    .d(_16078_),
    .o1(_16161_));
 b15nand02as1n08x5 _24971_ (.a(net871),
    .b(net866),
    .o1(_16162_));
 b15aoi112al1n03x5 _24972_ (.a(net867),
    .b(_16153_),
    .c(_16162_),
    .d(_16150_),
    .o1(_16163_));
 b15nor002as1n24x5 _24973_ (.a(_16080_),
    .b(_16113_),
    .o1(_16164_));
 b15aoai13ah1n03x5 _24974_ (.a(_16161_),
    .b(_16163_),
    .c(\us20.a[3] ),
    .d(_16164_),
    .o1(_16165_));
 b15norp03ar1n12x5 _24975_ (.a(_16156_),
    .b(_16159_),
    .c(_16165_),
    .o1(_16166_));
 b15nano23aq1n08x5 _24976_ (.a(_16131_),
    .b(_16140_),
    .c(_16149_),
    .d(_16166_),
    .out0(_16167_));
 b15nandp3as1n24x5 _24977_ (.a(_16053_),
    .b(_16120_),
    .c(_16167_),
    .o1(_16168_));
 b15bfn000ar1n02x5 output315 (.a(net315),
    .o(text_out[34]));
 b15bfn000ar1n02x5 output314 (.a(net314),
    .o(text_out[33]));
 b15bfn000ar1n02x5 output313 (.a(net313),
    .o(text_out[32]));
 b15bfn000ar1n02x5 output312 (.a(net312),
    .o(text_out[31]));
 b15bfn000ar1n02x5 output311 (.a(net311),
    .o(text_out[30]));
 b15bfn000ar1n02x5 output310 (.a(net310),
    .o(text_out[2]));
 b15bfn000ar1n02x5 output309 (.a(net309),
    .o(text_out[29]));
 b15bfn000ar1n02x5 output308 (.a(net308),
    .o(text_out[28]));
 b15bfn000ar1n02x5 output307 (.a(net307),
    .o(text_out[27]));
 b15bfn000ar1n02x5 output306 (.a(net306),
    .o(text_out[26]));
 b15bfn000ar1n02x5 output305 (.a(net305),
    .o(text_out[25]));
 b15bfn000ar1n02x5 output304 (.a(net304),
    .o(text_out[24]));
 b15and003aq1n16x5 _24990_ (.a(net725),
    .b(net716),
    .c(net720),
    .o(_16181_));
 b15bfn000ar1n02x5 output303 (.a(net303),
    .o(text_out[23]));
 b15bfn000ar1n02x5 output302 (.a(net302),
    .o(text_out[22]));
 b15bfn000ar1n02x5 output301 (.a(net301),
    .o(text_out[21]));
 b15nonb02aq1n06x5 _24994_ (.a(net722),
    .b(net742),
    .out0(_16185_));
 b15nandp2aq1n05x5 _24995_ (.a(_16181_),
    .b(_16185_),
    .o1(_16186_));
 b15bfn000ar1n02x5 output300 (.a(net300),
    .o(text_out[20]));
 b15bfn000ar1n02x5 output299 (.a(net299),
    .o(text_out[1]));
 b15nonb02aq1n06x5 _24998_ (.a(net722),
    .b(net733),
    .out0(_16189_));
 b15bfn000ar1n02x5 output298 (.a(net298),
    .o(text_out[19]));
 b15nor002al1n16x5 _25000_ (.a(net727),
    .b(net720),
    .o1(_16191_));
 b15bfn000ar1n02x5 output297 (.a(net297),
    .o(text_out[18]));
 b15nonb02as1n16x5 _25002_ (.a(net742),
    .b(net722),
    .out0(_16193_));
 b15and002an1n12x5 _25003_ (.a(net726),
    .b(net720),
    .o(_16194_));
 b15aoi022ar1n12x5 _25004_ (.a(_16189_),
    .b(_16191_),
    .c(_16193_),
    .d(_16194_),
    .o1(_16195_));
 b15bfn000ar1n02x5 output296 (.a(net296),
    .o(text_out[17]));
 b15bfn000ar1n02x5 output295 (.a(net295),
    .o(text_out[16]));
 b15bfn000ar1n02x5 output294 (.a(net294),
    .o(text_out[15]));
 b15oai112ah1n16x5 _25008_ (.a(net729),
    .b(_16186_),
    .c(_16195_),
    .d(net718),
    .o1(_16199_));
 b15bfn000ar1n02x5 output293 (.a(net293),
    .o(text_out[14]));
 b15bfn000ar1n02x5 output292 (.a(net292),
    .o(text_out[13]));
 b15nor003ar1n12x5 _25011_ (.a(net734),
    .b(net723),
    .c(net719),
    .o1(_16202_));
 b15orn002al1n16x5 _25012_ (.a(net728),
    .b(net716),
    .o(_16203_));
 b15bfn000ar1n02x5 output291 (.a(net291),
    .o(text_out[12]));
 b15bfn000ar1n02x5 output290 (.a(net290),
    .o(text_out[127]));
 b15nand02ah1n16x5 _25015_ (.a(net728),
    .b(net716),
    .o1(_16206_));
 b15bfn000ar1n02x5 output289 (.a(net289),
    .o(text_out[126]));
 b15bfn000ar1n02x5 output288 (.a(net288),
    .o(text_out[125]));
 b15oai012ar1n02x5 _25018_ (.a(_16203_),
    .b(_16206_),
    .c(net740),
    .o1(_16209_));
 b15bfn000ar1n02x5 output287 (.a(net287),
    .o(text_out[124]));
 b15bfn000ar1n02x5 output286 (.a(net286),
    .o(text_out[123]));
 b15bfn000ar1n02x5 output285 (.a(net285),
    .o(text_out[122]));
 b15nano23as1n24x5 _25022_ (.a(net724),
    .b(net727),
    .c(net718),
    .d(net721),
    .out0(_16213_));
 b15nonb02as1n16x5 _25023_ (.a(net735),
    .b(net741),
    .out0(_16214_));
 b15ao0022ar1n04x5 _25024_ (.a(_16202_),
    .b(_16209_),
    .c(_16213_),
    .d(_16214_),
    .o(_16215_));
 b15bfn000ar1n02x5 output284 (.a(net284),
    .o(text_out[121]));
 b15bfn000ar1n02x5 output283 (.a(net283),
    .o(text_out[120]));
 b15bfn000ar1n02x5 output282 (.a(net282),
    .o(text_out[11]));
 b15oai112aq1n16x5 _25028_ (.a(net738),
    .b(_16199_),
    .c(_16215_),
    .d(net730),
    .o1(_16219_));
 b15bfn000ar1n02x5 output281 (.a(net281),
    .o(text_out[119]));
 b15nanb02as1n24x5 _25030_ (.a(\us02.a[0] ),
    .b(net736),
    .out0(_16221_));
 b15norp02as1n08x5 _25031_ (.a(net739),
    .b(_16221_),
    .o1(_16222_));
 b15norp02as1n48x5 _25032_ (.a(net716),
    .b(net719),
    .o1(_16223_));
 b15nonb02as1n16x5 _25033_ (.a(net723),
    .b(net728),
    .out0(_16224_));
 b15nand02ar1n32x5 _25034_ (.a(_16223_),
    .b(_16224_),
    .o1(_16225_));
 b15inv000an1n64x5 _25035_ (.a(net732),
    .o1(_16226_));
 b15bfn000ar1n02x5 output280 (.a(net280),
    .o(text_out[118]));
 b15oai012an1n02x5 _25037_ (.a(_16222_),
    .b(_16225_),
    .c(_16226_),
    .o1(_16228_));
 b15and002ah1n24x5 _25038_ (.a(net716),
    .b(net719),
    .o(_16229_));
 b15nonb02as1n16x5 _25039_ (.a(net728),
    .b(net723),
    .out0(_16230_));
 b15nand02an1n32x5 _25040_ (.a(_16229_),
    .b(_16230_),
    .o1(_16231_));
 b15bfn000ar1n02x5 output279 (.a(net279),
    .o(text_out[117]));
 b15nonb02ah1n16x5 _25042_ (.a(\us02.a[3] ),
    .b(net736),
    .out0(_16233_));
 b15oai012ar1n03x5 _25043_ (.a(_16231_),
    .b(_16233_),
    .c(_16225_),
    .o1(_16234_));
 b15orn002aq1n32x5 _25044_ (.a(net717),
    .b(net720),
    .o(_16235_));
 b15bfn000ar1n02x5 output278 (.a(net278),
    .o(text_out[116]));
 b15nanb02as1n24x5 _25046_ (.a(net726),
    .b(net722),
    .out0(_16237_));
 b15bfn000ar1n02x5 output277 (.a(net277),
    .o(text_out[115]));
 b15nor002ah1n12x5 _25048_ (.a(_16235_),
    .b(_16237_),
    .o1(_16239_));
 b15oai112an1n08x5 _25049_ (.a(_16228_),
    .b(_16234_),
    .c(net730),
    .d(_16239_),
    .o1(_16240_));
 b15bfn000ar1n02x5 output276 (.a(net276),
    .o(text_out[114]));
 b15bfn000ar1n02x5 output275 (.a(net275),
    .o(text_out[113]));
 b15bfn000ar1n02x5 output274 (.a(net274),
    .o(text_out[112]));
 b15aoi012ar1n02x5 _25053_ (.a(net739),
    .b(net730),
    .c(_16231_),
    .o1(_16244_));
 b15bfn000ar1n02x5 output273 (.a(net273),
    .o(text_out[111]));
 b15bfn000ar1n02x5 output272 (.a(net272),
    .o(text_out[110]));
 b15and002aq1n12x5 _25056_ (.a(net738),
    .b(net730),
    .o(_16247_));
 b15inv000an1n64x5 _25057_ (.a(\us02.a[2] ),
    .o1(_16248_));
 b15bfn000ar1n02x5 output271 (.a(net271),
    .o(text_out[10]));
 b15oaoi13aq1n03x5 _25059_ (.a(_16244_),
    .b(_16247_),
    .c(_16248_),
    .d(_16239_),
    .o1(_16250_));
 b15aoai13as1n06x5 _25060_ (.a(_16219_),
    .b(_16240_),
    .c(\us02.a[0] ),
    .d(_16250_),
    .o1(_16251_));
 b15bfn000ar1n02x5 output270 (.a(net270),
    .o(text_out[109]));
 b15bfn000ar1n02x5 output269 (.a(net269),
    .o(text_out[108]));
 b15bfn000ar1n02x5 output268 (.a(net268),
    .o(text_out[107]));
 b15bfn000ar1n02x5 output267 (.a(net267),
    .o(text_out[106]));
 b15bfn000ar1n02x5 output266 (.a(net266),
    .o(text_out[105]));
 b15nand04ar1n02x5 _25066_ (.a(\us02.a[0] ),
    .b(net734),
    .c(_16223_),
    .d(_16230_),
    .o1(_16257_));
 b15nor002as1n24x5 _25067_ (.a(net724),
    .b(net727),
    .o1(_16258_));
 b15nonb02as1n16x5 _25068_ (.a(net720),
    .b(net717),
    .out0(_16259_));
 b15nandp2ar1n32x5 _25069_ (.a(_16258_),
    .b(_16259_),
    .o1(_16260_));
 b15bfn000ar1n02x5 output265 (.a(net265),
    .o(text_out[104]));
 b15bfn000ar1n02x5 output264 (.a(net264),
    .o(text_out[103]));
 b15oaoi13al1n02x5 _25072_ (.a(net738),
    .b(_16257_),
    .c(_16260_),
    .d(net734),
    .o1(_16263_));
 b15bfn000ar1n02x5 output263 (.a(net263),
    .o(text_out[102]));
 b15bfn000ar1n02x5 output262 (.a(net262),
    .o(text_out[101]));
 b15nand04ar1n02x5 _25075_ (.a(net738),
    .b(net734),
    .c(_16223_),
    .d(_16230_),
    .o1(_16266_));
 b15bfn000ar1n02x5 output261 (.a(net261),
    .o(text_out[100]));
 b15bfn000ar1n02x5 output260 (.a(net260),
    .o(text_out[0]));
 b15oaoi13al1n02x5 _25078_ (.a(\us02.a[0] ),
    .b(_16266_),
    .c(_16260_),
    .d(net738),
    .o1(_16269_));
 b15oai012ah1n03x5 _25079_ (.a(_16226_),
    .b(_16263_),
    .c(_16269_),
    .o1(_16270_));
 b15bfn000ar1n02x5 output259 (.a(net259),
    .o(done));
 b15bfn001ah1n08x5 input258 (.a(text_in[9]),
    .o(net258));
 b15nonb03ah1n08x5 _25082_ (.a(net726),
    .b(net717),
    .c(net720),
    .out0(_16273_));
 b15nor002ar1n08x5 _25083_ (.a(net737),
    .b(net722),
    .o1(_16274_));
 b15aoi022aq1n02x5 _25084_ (.a(net722),
    .b(_16229_),
    .c(_16273_),
    .d(_16274_),
    .o1(_16275_));
 b15inv020as1n08x5 _25085_ (.a(net726),
    .o1(_16276_));
 b15aoi013an1n03x5 _25086_ (.a(_16181_),
    .b(_16223_),
    .c(_16276_),
    .d(net740),
    .o1(_16277_));
 b15inv020aq1n28x5 _25087_ (.a(net723),
    .o1(_16278_));
 b15oai022as1n08x5 _25088_ (.a(net740),
    .b(_16275_),
    .c(_16277_),
    .d(_16278_),
    .o1(_16279_));
 b15nandp2an1n48x5 _25089_ (.a(net718),
    .b(net721),
    .o1(_16280_));
 b15bfn000ar1n02x5 input257 (.a(text_in[99]),
    .o(net257));
 b15nand02as1n16x5 _25091_ (.a(_16223_),
    .b(_16230_),
    .o1(_16282_));
 b15inv020an1n64x5 _25092_ (.a(net740),
    .o1(_16283_));
 b15bfn000ar1n02x5 input256 (.a(text_in[98]),
    .o(net256));
 b15oai022aq1n04x5 _25094_ (.a(_16278_),
    .b(_16280_),
    .c(_16282_),
    .d(_16283_),
    .o1(_16285_));
 b15bfm201ah1n02x5 input255 (.a(text_in[97]),
    .o(net255));
 b15aoai13an1n08x5 _25096_ (.a(_16233_),
    .b(_16279_),
    .c(_16285_),
    .d(net738),
    .o1(_16287_));
 b15bfn000al1n02x5 input254 (.a(text_in[96]),
    .o(net254));
 b15norp02an1n24x5 _25098_ (.a(net730),
    .b(net725),
    .o1(_16289_));
 b15nandp3ar1n02x5 _25099_ (.a(net723),
    .b(_16229_),
    .c(_16289_),
    .o1(_16290_));
 b15nonb02al1n16x5 _25100_ (.a(net716),
    .b(net728),
    .out0(_16291_));
 b15nor002ah1n12x5 _25101_ (.a(net730),
    .b(net723),
    .o1(_16292_));
 b15nonb02aq1n12x5 _25102_ (.a(net728),
    .b(net716),
    .out0(_16293_));
 b15bfn001ah1n16x5 input253 (.a(text_in[95]),
    .o(net253));
 b15and002al1n08x5 _25104_ (.a(net730),
    .b(net723),
    .o(_16295_));
 b15aoi022ar1n02x5 _25105_ (.a(_16291_),
    .b(_16292_),
    .c(_16293_),
    .d(_16295_),
    .o1(_16296_));
 b15bfn001ah1n16x5 input252 (.a(text_in[94]),
    .o(net252));
 b15bfn001ah1n16x5 input251 (.a(text_in[93]),
    .o(net251));
 b15oaoi13ah1n02x5 _25108_ (.a(net738),
    .b(_16290_),
    .c(_16296_),
    .d(net719),
    .o1(_16299_));
 b15bfn001ah1n16x5 input250 (.a(text_in[92]),
    .o(net250));
 b15and002ar1n24x5 _25110_ (.a(net723),
    .b(net728),
    .o(_16301_));
 b15aoai13ar1n02x5 _25111_ (.a(net716),
    .b(_16258_),
    .c(_16301_),
    .d(_16226_),
    .o1(_16302_));
 b15aob012ar1n03x5 _25112_ (.a(_16302_),
    .b(_16295_),
    .c(_16293_),
    .out0(_16303_));
 b15bfn000al1n02x5 input249 (.a(text_in[91]),
    .o(net249));
 b15inv000an1n32x5 _25114_ (.a(net719),
    .o1(_16305_));
 b15bfn000as1n06x5 input248 (.a(text_in[90]),
    .o(net248));
 b15aoi013an1n04x5 _25116_ (.a(_16299_),
    .b(_16303_),
    .c(\us02.a[0] ),
    .d(_16305_),
    .o1(_16307_));
 b15oai112as1n12x5 _25117_ (.a(_16270_),
    .b(_16287_),
    .c(_16248_),
    .d(_16307_),
    .o1(_16308_));
 b15bfn001as1n06x5 input247 (.a(text_in[8]),
    .o(net247));
 b15nanb02as1n24x5 _25119_ (.a(net722),
    .b(net726),
    .out0(_16310_));
 b15nandp2ar1n48x5 _25120_ (.a(\us02.a[0] ),
    .b(\us02.a[2] ),
    .o1(_16311_));
 b15nor004as1n02x5 _25121_ (.a(net737),
    .b(_16280_),
    .c(_16310_),
    .d(_16311_),
    .o1(_16312_));
 b15orn002aq1n24x5 _25122_ (.a(net724),
    .b(net727),
    .o(_16313_));
 b15nanb02as1n24x5 _25123_ (.a(net720),
    .b(net717),
    .out0(_16314_));
 b15nor002ah1n16x5 _25124_ (.a(_16313_),
    .b(_16314_),
    .o1(_16315_));
 b15norp02an1n24x5 _25125_ (.a(net743),
    .b(net735),
    .o1(_16316_));
 b15aoai13an1n02x5 _25126_ (.a(_16226_),
    .b(_16312_),
    .c(_16315_),
    .d(_16316_),
    .o1(_16317_));
 b15nand02as1n32x5 _25127_ (.a(net732),
    .b(net736),
    .o1(_16318_));
 b15norp03al1n02x5 _25128_ (.a(_16313_),
    .b(_16314_),
    .c(_16318_),
    .o1(_16319_));
 b15norp03as1n24x5 _25129_ (.a(net741),
    .b(net731),
    .c(net735),
    .o1(_16320_));
 b15nor002an1n32x5 _25130_ (.a(_16280_),
    .b(_16310_),
    .o1(_16321_));
 b15aoai13aq1n03x5 _25131_ (.a(net737),
    .b(_16319_),
    .c(_16320_),
    .d(_16321_),
    .o1(_16322_));
 b15nand02as1n16x5 _25132_ (.a(net741),
    .b(net731),
    .o1(_16323_));
 b15bfn001aq1n06x5 input246 (.a(text_in[89]),
    .o(net246));
 b15nano23as1n24x5 _25134_ (.a(net724),
    .b(net721),
    .c(net718),
    .d(net727),
    .out0(_16325_));
 b15nandp2ar1n08x5 _25135_ (.a(_16248_),
    .b(_16325_),
    .o1(_16326_));
 b15nandp3ar1n12x5 _25136_ (.o1(_16327_),
    .a(net734),
    .b(_16224_),
    .c(_16229_));
 b15nonb02as1n16x5 _25137_ (.a(net717),
    .b(net720),
    .out0(_16328_));
 b15nandp2al1n08x5 _25138_ (.a(_16258_),
    .b(_16328_),
    .o1(_16329_));
 b15aoi013al1n03x5 _25139_ (.a(_16323_),
    .b(_16326_),
    .c(_16327_),
    .d(_16329_),
    .o1(_16330_));
 b15bfn001as1n06x5 input245 (.a(text_in[88]),
    .o(net245));
 b15nano23aq1n24x5 _25141_ (.a(net724),
    .b(\us02.a[7] ),
    .c(\us02.a[6] ),
    .d(net727),
    .out0(_16332_));
 b15and002aq1n24x5 _25142_ (.a(net743),
    .b(net736),
    .o(_16333_));
 b15oab012ar1n06x5 _25143_ (.a(\us02.a[1] ),
    .b(net741),
    .c(net735),
    .out0(_16334_));
 b15oai112as1n02x5 _25144_ (.a(net731),
    .b(_16332_),
    .c(_16333_),
    .d(_16334_),
    .o1(_16335_));
 b15nona23as1n32x5 _25145_ (.a(net724),
    .b(net718),
    .c(net721),
    .d(net727),
    .out0(_16336_));
 b15nanb02ah1n08x5 _25146_ (.a(net731),
    .b(net739),
    .out0(_16337_));
 b15oai013an1n08x5 _25147_ (.a(_16335_),
    .b(_16336_),
    .c(_16337_),
    .d(_16248_),
    .o1(_16338_));
 b15nano23aq1n08x5 _25148_ (.a(_16317_),
    .b(_16322_),
    .c(_16330_),
    .d(_16338_),
    .out0(_16339_));
 b15andc04ah1n16x5 _25149_ (.a(\us02.a[5] ),
    .b(net728),
    .c(\us02.a[7] ),
    .d(\us02.a[6] ),
    .o(_16340_));
 b15nandp3ar1n02x5 _25150_ (.a(_16226_),
    .b(_16248_),
    .c(_16340_),
    .o1(_16341_));
 b15inv020as1n64x5 _25151_ (.a(net739),
    .o1(_16342_));
 b15nor004as1n12x5 _25152_ (.a(net722),
    .b(net725),
    .c(net716),
    .d(net720),
    .o1(_16343_));
 b15aoi013ar1n02x5 _25153_ (.a(_16342_),
    .b(\us02.a[3] ),
    .c(_16311_),
    .d(_16343_),
    .o1(_16344_));
 b15nor002al1n02x5 _25154_ (.a(net742),
    .b(net732),
    .o1(_16345_));
 b15nand03ar1n02x5 _25155_ (.a(net736),
    .b(_16340_),
    .c(_16345_),
    .o1(_16346_));
 b15and002aq1n12x5 _25156_ (.a(net740),
    .b(net730),
    .o(_16347_));
 b15aoi012ar1n02x5 _25157_ (.a(net739),
    .b(_16347_),
    .c(_16343_),
    .o1(_16348_));
 b15ao0022an1n02x5 _25158_ (.a(_16341_),
    .b(_16344_),
    .c(_16346_),
    .d(_16348_),
    .o(_16349_));
 b15norp02al1n32x5 _25159_ (.a(net738),
    .b(net734),
    .o1(_16350_));
 b15nano22ah1n08x5 _25160_ (.a(net723),
    .b(net720),
    .c(net716),
    .out0(_16351_));
 b15bfn001ah1n06x5 input244 (.a(text_in[87]),
    .o(net244));
 b15nonb02al1n04x5 _25162_ (.a(net730),
    .b(net725),
    .out0(_16353_));
 b15nonb02as1n08x5 _25163_ (.a(net725),
    .b(net730),
    .out0(_16354_));
 b15oai112as1n12x5 _25164_ (.a(_16350_),
    .b(_16351_),
    .c(_16353_),
    .d(_16354_),
    .o1(_16355_));
 b15nonb02aq1n16x5 _25165_ (.a(net734),
    .b(net738),
    .out0(_16356_));
 b15nanb02ah1n24x5 _25166_ (.a(\us02.a[0] ),
    .b(\us02.a[3] ),
    .out0(_16357_));
 b15nandp3al1n12x5 _25167_ (.o1(_16358_),
    .a(net723),
    .b(net728),
    .c(net716));
 b15norp02as1n03x5 _25168_ (.a(_16357_),
    .b(_16358_),
    .o1(_16359_));
 b15bfn001ah1n16x5 input243 (.a(text_in[86]),
    .o(net243));
 b15nanb02as1n24x5 _25170_ (.a(net730),
    .b(net740),
    .out0(_16361_));
 b15norp03an1n04x5 _25171_ (.a(net723),
    .b(_16203_),
    .c(_16361_),
    .o1(_16362_));
 b15oai112ah1n12x5 _25172_ (.a(_16305_),
    .b(_16356_),
    .c(_16359_),
    .d(_16362_),
    .o1(_16363_));
 b15and003al1n03x5 _25173_ (.a(_16349_),
    .b(_16355_),
    .c(_16363_),
    .o(_16364_));
 b15nonb02al1n12x5 _25174_ (.a(net732),
    .b(net743),
    .out0(_16365_));
 b15nandp3al1n03x5 _25175_ (.a(net733),
    .b(_16293_),
    .c(_16365_),
    .o1(_16366_));
 b15nandp2as1n16x5 _25176_ (.a(\us02.a[0] ),
    .b(_16248_),
    .o1(_16367_));
 b15aoi022al1n02x5 _25177_ (.a(net716),
    .b(_16289_),
    .c(_16293_),
    .d(net729),
    .o1(_16368_));
 b15oai112as1n06x5 _25178_ (.a(net738),
    .b(_16366_),
    .c(_16367_),
    .d(_16368_),
    .o1(_16369_));
 b15and002ar1n08x5 _25179_ (.a(net722),
    .b(net719),
    .o(_16370_));
 b15nandp2ar1n02x5 _25180_ (.a(_16291_),
    .b(_16320_),
    .o1(_16371_));
 b15nanb02as1n12x5 _25181_ (.a(net718),
    .b(net725),
    .out0(_16372_));
 b15oai013aq1n06x5 _25182_ (.a(_16371_),
    .b(_16323_),
    .c(_16372_),
    .d(_16248_),
    .o1(_16373_));
 b15oai112as1n16x5 _25183_ (.a(_16369_),
    .b(_16370_),
    .c(net738),
    .d(_16373_),
    .o1(_16374_));
 b15bfn001ah1n16x5 input242 (.a(text_in[85]),
    .o(net242));
 b15oai112as1n04x5 _25185_ (.a(net721),
    .b(_16258_),
    .c(net731),
    .d(net718),
    .o1(_16376_));
 b15nandp2ah1n12x5 _25186_ (.a(net737),
    .b(net735),
    .o1(_16377_));
 b15aoai13as1n02x5 _25187_ (.a(net731),
    .b(_16214_),
    .c(_16377_),
    .d(net741),
    .o1(_16378_));
 b15nanb02as1n24x5 _25188_ (.a(net743),
    .b(\us02.a[1] ),
    .out0(_16379_));
 b15bfn001aq1n06x5 input241 (.a(text_in[84]),
    .o(net241));
 b15orn002as1n24x5 _25190_ (.a(net732),
    .b(net735),
    .o(_16381_));
 b15oaoi13as1n08x5 _25191_ (.a(_16376_),
    .b(_16378_),
    .c(_16379_),
    .d(_16381_),
    .o1(_16382_));
 b15nona23an1n32x5 _25192_ (.a(net718),
    .b(net721),
    .c(net724),
    .d(net727),
    .out0(_16383_));
 b15aoi012aq1n02x5 _25193_ (.a(_16381_),
    .b(_16336_),
    .c(_16383_),
    .o1(_16384_));
 b15bfn000an1n02x5 input240 (.a(text_in[83]),
    .o(net240));
 b15nand02ar1n02x5 _25195_ (.a(net739),
    .b(_16213_),
    .o1(_16386_));
 b15oai112ah1n04x5 _25196_ (.a(_16283_),
    .b(_16386_),
    .c(_16336_),
    .d(net739),
    .o1(_16387_));
 b15nanb02as1n12x5 _25197_ (.a(net739),
    .b(net734),
    .out0(_16388_));
 b15nand02as1n16x5 _25198_ (.a(_16301_),
    .b(_16328_),
    .o1(_16389_));
 b15norp02al1n48x5 _25199_ (.a(\us02.a[1] ),
    .b(net743),
    .o1(_16390_));
 b15nandp2al1n08x5 _25200_ (.a(_16390_),
    .b(_16343_),
    .o1(_16391_));
 b15bfn000ar1n02x5 input239 (.a(text_in[82]),
    .o(net239));
 b15oai022al1n02x5 _25202_ (.a(_16388_),
    .b(_16389_),
    .c(_16391_),
    .d(net734),
    .o1(_16393_));
 b15aoi122an1n04x5 _25203_ (.a(_16382_),
    .b(_16384_),
    .c(_16387_),
    .d(_16226_),
    .e(_16393_),
    .o1(_16394_));
 b15nand04ar1n16x5 _25204_ (.a(_16339_),
    .b(_16364_),
    .c(_16374_),
    .d(_16394_),
    .o1(_16395_));
 b15nona23al1n32x5 _25205_ (.a(net727),
    .b(net717),
    .c(net720),
    .d(net724),
    .out0(_16396_));
 b15norp03as1n04x5 _25206_ (.a(_16318_),
    .b(_16396_),
    .c(_16379_),
    .o1(_16397_));
 b15nand02aq1n24x5 _25207_ (.a(net724),
    .b(net727),
    .o1(_16398_));
 b15nonb02ah1n04x5 _25208_ (.a(net741),
    .b(net737),
    .out0(_16399_));
 b15nor004ar1n08x5 _25209_ (.a(_16398_),
    .b(_16314_),
    .c(_16399_),
    .d(_16381_),
    .o1(_16400_));
 b15norp02an1n24x5 _25210_ (.a(_16342_),
    .b(\us02.a[3] ),
    .o1(_16401_));
 b15ornc04aq1n24x5 _25211_ (.a(net724),
    .b(net727),
    .c(\us02.a[7] ),
    .d(\us02.a[6] ),
    .o(_16402_));
 b15norp02ar1n24x5 _25212_ (.a(_16248_),
    .b(_16402_),
    .o1(_16403_));
 b15aoi112as1n08x5 _25213_ (.a(_16397_),
    .b(_16400_),
    .c(_16401_),
    .d(_16403_),
    .o1(_16404_));
 b15nonb02as1n16x5 _25214_ (.a(net738),
    .b(net734),
    .out0(_16405_));
 b15aoi013al1n06x5 _25215_ (.a(net731),
    .b(_16223_),
    .c(_16230_),
    .d(_16405_),
    .o1(_16406_));
 b15bfn000as1n04x5 input238 (.a(text_in[81]),
    .o(net238));
 b15bfn000ar1n02x5 input237 (.a(text_in[80]),
    .o(net237));
 b15nand02ar1n02x5 _25218_ (.a(net734),
    .b(net718),
    .o1(_16409_));
 b15nand04ah1n04x5 _25219_ (.a(net742),
    .b(net724),
    .c(_16194_),
    .d(_16409_),
    .o1(_16410_));
 b15aoi012an1n02x5 _25220_ (.a(_16325_),
    .b(_16332_),
    .c(_16390_),
    .o1(_16411_));
 b15oai112ah1n08x5 _25221_ (.a(_16406_),
    .b(_16410_),
    .c(_16248_),
    .d(_16411_),
    .o1(_16412_));
 b15nandp3al1n04x5 _25222_ (.a(_16248_),
    .b(_16390_),
    .c(_16213_),
    .o1(_16413_));
 b15nona23as1n32x5 _25223_ (.a(net724),
    .b(net721),
    .c(net718),
    .d(net727),
    .out0(_16414_));
 b15oai112ar1n16x5 _25224_ (.a(net731),
    .b(_16413_),
    .c(_16414_),
    .d(_16377_),
    .o1(_16415_));
 b15nano23aq1n24x5 _25225_ (.a(net728),
    .b(\us02.a[7] ),
    .c(\us02.a[6] ),
    .d(\us02.a[5] ),
    .out0(_16416_));
 b15aoi112al1n02x5 _25226_ (.a(net731),
    .b(_16325_),
    .c(_16350_),
    .d(_16416_),
    .o1(_16417_));
 b15norp02ah1n24x5 _25227_ (.a(net734),
    .b(net722),
    .o1(_16418_));
 b15nano22an1n24x5 _25228_ (.a(net726),
    .b(net720),
    .c(net718),
    .out0(_16419_));
 b15nandp2ah1n12x5 _25229_ (.a(_16418_),
    .b(_16419_),
    .o1(_16420_));
 b15aoi012al1n02x5 _25230_ (.a(_16417_),
    .b(_16420_),
    .c(net731),
    .o1(_16421_));
 b15aoi022ah1n06x5 _25231_ (.a(_16412_),
    .b(_16415_),
    .c(_16421_),
    .d(net741),
    .o1(_16422_));
 b15nand02an1n08x5 _25232_ (.a(_16404_),
    .b(_16422_),
    .o1(_16423_));
 b15nor004as1n12x5 _25233_ (.a(_16251_),
    .b(_16308_),
    .c(_16395_),
    .d(_16423_),
    .o1(_16424_));
 b15bfn001al1n08x5 input236 (.a(text_in[7]),
    .o(net236));
 b15bfn001as1n12x5 input235 (.a(text_in[79]),
    .o(net235));
 b15bfn001ah1n08x5 input234 (.a(text_in[78]),
    .o(net234));
 b15bfn001ah1n08x5 input233 (.a(text_in[77]),
    .o(net233));
 b15nano23as1n12x5 _25238_ (.a(net602),
    .b(net609),
    .c(net613),
    .d(net605),
    .out0(_16429_));
 b15bfn001ah1n12x5 input232 (.a(text_in[76]),
    .o(net232));
 b15bfn000ah1n03x5 input231 (.a(text_in[75]),
    .o(net231));
 b15nand02an1n24x5 _25241_ (.a(net598),
    .b(net600),
    .o1(_16432_));
 b15bfn000as1n02x5 input230 (.a(text_in[74]),
    .o(net230));
 b15bfn001aq1n06x5 input229 (.a(text_in[73]),
    .o(net229));
 b15nonb02as1n16x5 _25244_ (.a(net620),
    .b(net616),
    .out0(_16435_));
 b15bfn001as1n06x5 input228 (.a(text_in[72]),
    .o(net228));
 b15bfn001as1n08x5 input227 (.a(text_in[71]),
    .o(net227));
 b15orn002an1n12x5 _25247_ (.a(net597),
    .b(net601),
    .o(_16438_));
 b15norp02aq1n48x5 _25248_ (.a(net619),
    .b(net615),
    .o1(_16439_));
 b15bfn001as1n06x5 input226 (.a(text_in[70]),
    .o(net226));
 b15oai022ar1n02x5 _25250_ (.a(_16432_),
    .b(_16435_),
    .c(_16438_),
    .d(_16439_),
    .o1(_16441_));
 b15and002al1n02x5 _25251_ (.a(_16429_),
    .b(_16441_),
    .o(_16442_));
 b15bfn001aq1n06x5 input225 (.a(text_in[6]),
    .o(net225));
 b15bfn001as1n06x5 input224 (.a(text_in[69]),
    .o(net224));
 b15bfn001ah1n06x5 input223 (.a(text_in[68]),
    .o(net223));
 b15nonb02aq1n16x5 _25255_ (.a(net603),
    .b(net600),
    .out0(_16446_));
 b15bfn001as1n06x5 input222 (.a(text_in[67]),
    .o(net222));
 b15bfn001as1n06x5 input221 (.a(text_in[66]),
    .o(net221));
 b15bfn000as1n02x5 input220 (.a(text_in[65]),
    .o(net220));
 b15bfn001as1n06x5 input219 (.a(text_in[64]),
    .o(net219));
 b15bfn000as1n02x5 input218 (.a(text_in[63]),
    .o(net218));
 b15bfn000as1n02x5 input217 (.a(text_in[62]),
    .o(net217));
 b15nanb02as1n24x5 _25262_ (.a(net618),
    .b(net615),
    .out0(_16453_));
 b15nand04ar1n04x5 _25263_ (.a(net605),
    .b(net597),
    .c(\us13.a[2] ),
    .d(_16453_),
    .o1(_16454_));
 b15bfn000ah1n02x5 input216 (.a(text_in[61]),
    .o(net216));
 b15and002aq1n32x5 _25265_ (.a(net620),
    .b(net617),
    .o(_16456_));
 b15bfn000ah1n04x5 input215 (.a(text_in[60]),
    .o(net215));
 b15inv020ah1n24x5 _25267_ (.a(\us13.a[7] ),
    .o1(_16458_));
 b15bfn001ah1n16x5 input214 (.a(text_in[5]),
    .o(net214));
 b15inv040al1n40x5 _25269_ (.a(net612),
    .o1(_16460_));
 b15qbfna2bn1n16x5 _25270_ (.a(_16458_),
    .b(_16460_),
    .o1(_16461_));
 b15bfn001as1n08x5 input213 (.a(text_in[59]),
    .o(net213));
 b15bfn000ar1n02x5 input212 (.a(text_in[58]),
    .o(net212));
 b15oai013al1n06x5 _25273_ (.a(_16454_),
    .b(_16456_),
    .c(_16461_),
    .d(net605),
    .o1(_16464_));
 b15bfn000al1n02x5 input211 (.a(text_in[57]),
    .o(net211));
 b15inv020an1n64x5 _25275_ (.a(net608),
    .o1(_16466_));
 b15bfn000ar1n02x5 input210 (.a(text_in[56]),
    .o(net210));
 b15aoi013aq1n08x5 _25277_ (.a(_16442_),
    .b(_16446_),
    .c(_16464_),
    .d(_16466_),
    .o1(_16468_));
 b15bfn000ar1n02x5 input209 (.a(text_in[55]),
    .o(net209));
 b15bfn000ar1n02x5 input208 (.a(text_in[54]),
    .o(net208));
 b15bfn000aq1n02x5 input207 (.a(text_in[53]),
    .o(net207));
 b15bfn000ar1n02x5 input206 (.a(text_in[52]),
    .o(net206));
 b15nonb02as1n16x5 _25282_ (.a(net600),
    .b(net596),
    .out0(_16473_));
 b15bfn001as1n06x5 input205 (.a(text_in[51]),
    .o(net205));
 b15norp02as1n48x5 _25284_ (.a(net602),
    .b(net607),
    .o1(_16475_));
 b15bfn000as1n02x5 input204 (.a(text_in[50]),
    .o(net204));
 b15nandp3ar1n12x5 _25286_ (.o1(_16477_),
    .a(net609),
    .b(_16473_),
    .c(_16475_));
 b15and002ar1n24x5 _25287_ (.a(net615),
    .b(net611),
    .o(_16478_));
 b15orn002aq1n32x5 _25288_ (.a(net611),
    .b(net608),
    .o(_16479_));
 b15bfn001aq1n06x5 input203 (.a(text_in[4]),
    .o(net203));
 b15nonb02as1n16x5 _25290_ (.a(net602),
    .b(net605),
    .out0(_16481_));
 b15nandp2ah1n24x5 _25291_ (.a(_16481_),
    .b(_16473_),
    .o1(_16482_));
 b15oai022as1n06x5 _25292_ (.a(_16477_),
    .b(_16478_),
    .c(_16479_),
    .d(_16482_),
    .o1(_16483_));
 b15nandp2an1n02x5 _25293_ (.a(net619),
    .b(_16483_),
    .o1(_16484_));
 b15bfn000ar1n02x5 input202 (.a(text_in[49]),
    .o(net202));
 b15bfn001aq1n06x5 input201 (.a(text_in[48]),
    .o(net201));
 b15bfn000as1n02x5 input200 (.a(text_in[47]),
    .o(net200));
 b15bfn000ah1n02x5 input199 (.a(text_in[46]),
    .o(net199));
 b15bfn000ar1n02x5 input198 (.a(text_in[45]),
    .o(net198));
 b15nonb02ah1n16x5 _25299_ (.a(net615),
    .b(net619),
    .out0(_16490_));
 b15nandp2ah1n08x5 _25300_ (.a(net612),
    .b(_16490_),
    .o1(_16491_));
 b15nanb02aq1n24x5 _25301_ (.a(net611),
    .b(net619),
    .out0(_16492_));
 b15bfn000ar1n02x5 input197 (.a(text_in[44]),
    .o(net197));
 b15nor002as1n08x5 _25303_ (.a(net599),
    .b(\us13.a[3] ),
    .o1(_16494_));
 b15and003ar1n02x5 _25304_ (.a(_16492_),
    .b(_16475_),
    .c(_16494_),
    .o(_16495_));
 b15bfn000ar1n02x5 input196 (.a(text_in[43]),
    .o(net196));
 b15nanb02as1n24x5 _25306_ (.a(net605),
    .b(net603),
    .out0(_16497_));
 b15nanb02as1n24x5 _25307_ (.a(net609),
    .b(\us13.a[0] ),
    .out0(_16498_));
 b15bfn000ar1n02x5 input195 (.a(text_in[42]),
    .o(net195));
 b15nand02ar1n16x5 _25309_ (.a(net606),
    .b(net610),
    .o1(_16500_));
 b15bfn000ar1n02x5 input194 (.a(text_in[41]),
    .o(net194));
 b15bfn000ar1n02x5 input193 (.a(text_in[40]),
    .o(net193));
 b15oai022ar1n02x5 _25312_ (.a(_16497_),
    .b(_16498_),
    .c(_16500_),
    .d(net603),
    .o1(_16503_));
 b15nonb02as1n16x5 _25313_ (.a(net615),
    .b(net611),
    .out0(_16504_));
 b15bfn001ah1n08x5 input192 (.a(text_in[3]),
    .o(net192));
 b15and003ar1n02x5 _25315_ (.a(net599),
    .b(_16503_),
    .c(_16504_),
    .o(_16506_));
 b15oai112as1n04x5 _25316_ (.a(net598),
    .b(_16491_),
    .c(_16495_),
    .d(_16506_),
    .o1(_16507_));
 b15inv040ah1n36x5 _25317_ (.a(net615),
    .o1(_16508_));
 b15bfn000aq1n02x5 input191 (.a(text_in[39]),
    .o(net191));
 b15nor002al1n24x5 _25319_ (.a(net602),
    .b(net596),
    .o1(_16510_));
 b15nor002as1n04x5 _25320_ (.a(net599),
    .b(net613),
    .o1(_16511_));
 b15bfn000ah1n02x5 input190 (.a(text_in[38]),
    .o(net190));
 b15orn002ar1n12x5 _25322_ (.a(net605),
    .b(net610),
    .o(_16513_));
 b15aoi012ar1n02x5 _25323_ (.a(net618),
    .b(_16500_),
    .c(_16513_),
    .o1(_16514_));
 b15nano22aq1n02x5 _25324_ (.a(_16510_),
    .b(_16511_),
    .c(_16514_),
    .out0(_16515_));
 b15orn002aq1n16x5 _25325_ (.a(net620),
    .b(net612),
    .o(_16516_));
 b15nonb02as1n16x5 _25326_ (.a(net605),
    .b(\us13.a[5] ),
    .out0(_16517_));
 b15nonb03as1n12x5 _25327_ (.a(\us13.a[3] ),
    .b(net599),
    .c(net598),
    .out0(_16518_));
 b15nandp2ar1n24x5 _25328_ (.a(_16517_),
    .b(_16518_),
    .o1(_16519_));
 b15and002ah1n32x5 _25329_ (.a(net596),
    .b(net599),
    .o(_16520_));
 b15nandp2ah1n48x5 _25330_ (.a(_16520_),
    .b(_16517_),
    .o1(_16521_));
 b15nanb02as1n24x5 _25331_ (.a(net613),
    .b(net609),
    .out0(_16522_));
 b15oai122aq1n16x5 _25332_ (.a(_16508_),
    .b(_16516_),
    .c(_16519_),
    .d(_16521_),
    .e(_16522_),
    .o1(_16523_));
 b15nanb02as1n24x5 _25333_ (.a(net608),
    .b(net611),
    .out0(_16524_));
 b15bfn000as1n02x5 input189 (.a(text_in[37]),
    .o(net189));
 b15nor004as1n12x5 _25335_ (.a(net604),
    .b(net607),
    .c(net597),
    .d(net601),
    .o1(_16526_));
 b15nand02al1n02x5 _25336_ (.a(net618),
    .b(_16526_),
    .o1(_16527_));
 b15nand04as1n16x5 _25337_ (.a(net604),
    .b(net607),
    .c(net597),
    .d(net601),
    .o1(_16528_));
 b15oaoi13aq1n02x5 _25338_ (.a(_16524_),
    .b(_16527_),
    .c(_16528_),
    .d(net618),
    .o1(_16529_));
 b15oai022an1n06x5 _25339_ (.a(_16508_),
    .b(_16515_),
    .c(_16523_),
    .d(_16529_),
    .o1(_16530_));
 b15nand04as1n08x5 _25340_ (.a(_16468_),
    .b(_16484_),
    .c(_16507_),
    .d(_16530_),
    .o1(_16531_));
 b15bfn000aq1n02x5 input188 (.a(text_in[36]),
    .o(net188));
 b15bfn000ah1n02x5 input187 (.a(text_in[35]),
    .o(net187));
 b15bfn000ar1n02x5 input186 (.a(text_in[34]),
    .o(net186));
 b15nanb02al1n08x5 _25344_ (.a(net616),
    .b(net601),
    .out0(_16535_));
 b15nandp2as1n08x5 _25345_ (.a(net620),
    .b(\us13.a[3] ),
    .o1(_16536_));
 b15bfn000al1n02x5 input185 (.a(text_in[33]),
    .o(net185));
 b15nanb02as1n24x5 _25347_ (.a(\us13.a[5] ),
    .b(net605),
    .out0(_16538_));
 b15norp02as1n03x5 _25348_ (.a(\us13.a[7] ),
    .b(_16538_),
    .o1(_16539_));
 b15nanb02ar1n02x5 _25349_ (.a(_16536_),
    .b(_16539_),
    .out0(_16540_));
 b15bfn000ah1n03x5 input184 (.a(text_in[32]),
    .o(net184));
 b15nonb02an1n08x5 _25351_ (.a(\us13.a[3] ),
    .b(\us13.a[7] ),
    .out0(_16542_));
 b15aoi112ar1n02x5 _25352_ (.a(net604),
    .b(_16542_),
    .c(_16536_),
    .d(\us13.a[7] ),
    .o1(_16543_));
 b15norp02ah1n16x5 _25353_ (.a(\us13.a[0] ),
    .b(\us13.a[3] ),
    .o1(_16544_));
 b15bfn001aq1n06x5 input183 (.a(text_in[31]),
    .o(net183));
 b15aoi013al1n02x5 _25355_ (.a(_16543_),
    .b(_16544_),
    .c(net597),
    .d(net604),
    .o1(_16546_));
 b15oaoi13al1n02x5 _25356_ (.a(_16535_),
    .b(_16540_),
    .c(net606),
    .d(_16546_),
    .o1(_16547_));
 b15norp02ar1n02x5 _25357_ (.a(net606),
    .b(_16536_),
    .o1(_16548_));
 b15nanb02as1n24x5 _25358_ (.a(net601),
    .b(net597),
    .out0(_16549_));
 b15nor002an1n08x5 _25359_ (.a(net604),
    .b(_16549_),
    .o1(_16550_));
 b15aoai13ar1n02x5 _25360_ (.a(_16548_),
    .b(_16550_),
    .c(_16473_),
    .d(net604),
    .o1(_16551_));
 b15bfn000ah1n06x5 input182 (.a(text_in[30]),
    .o(net182));
 b15bfn001aq1n06x5 input181 (.a(text_in[2]),
    .o(net181));
 b15bfn001ah1n16x5 input180 (.a(text_in[29]),
    .o(net180));
 b15bfn001aq1n06x5 input179 (.a(text_in[28]),
    .o(net179));
 b15oai013ar1n02x5 _25365_ (.a(_16551_),
    .b(_16521_),
    .c(_16453_),
    .d(net610),
    .o1(_16556_));
 b15oab012an1n04x5 _25366_ (.a(net612),
    .b(_16547_),
    .c(_16556_),
    .out0(_16557_));
 b15inv000as1n48x5 _25367_ (.a(net620),
    .o1(_16558_));
 b15bfn001as1n12x5 input178 (.a(text_in[27]),
    .o(net178));
 b15bfn001aq1n06x5 input177 (.a(text_in[26]),
    .o(net177));
 b15nor002al1n04x5 _25370_ (.a(net599),
    .b(net614),
    .o1(_16561_));
 b15bfn000ah1n06x5 input176 (.a(text_in[25]),
    .o(net176));
 b15nandp2al1n08x5 _25372_ (.a(net605),
    .b(net599),
    .o1(_16563_));
 b15orn002an1n08x5 _25373_ (.a(net599),
    .b(net614),
    .o(_16564_));
 b15bfn001as1n12x5 input175 (.a(text_in[24]),
    .o(net175));
 b15oai012an1n02x5 _25375_ (.a(_16563_),
    .b(_16564_),
    .c(net605),
    .o1(_16566_));
 b15aoi022al1n06x5 _25376_ (.a(_16517_),
    .b(_16561_),
    .c(_16566_),
    .d(net603),
    .o1(_16567_));
 b15nor004aq1n03x5 _25377_ (.a(net598),
    .b(_16558_),
    .c(_16524_),
    .d(_16567_),
    .o1(_16568_));
 b15bfn001as1n06x5 input174 (.a(text_in[23]),
    .o(net174));
 b15bfn000ar1n02x5 input173 (.a(text_in[22]),
    .o(net173));
 b15norp02as1n08x5 _25380_ (.a(_16497_),
    .b(_16432_),
    .o1(_16571_));
 b15nandp3ar1n02x5 _25381_ (.a(net613),
    .b(_16466_),
    .c(_16571_),
    .o1(_16572_));
 b15oaoi13aq1n02x5 _25382_ (.a(net617),
    .b(_16572_),
    .c(_16527_),
    .d(_16466_),
    .o1(_16573_));
 b15bfn000ar1n02x5 input172 (.a(text_in[21]),
    .o(net172));
 b15nanb02aq1n24x5 _25384_ (.a(net618),
    .b(net611),
    .out0(_16575_));
 b15nand02aq1n32x5 _25385_ (.a(_16473_),
    .b(_16475_),
    .o1(_16576_));
 b15norp02ah1n48x5 _25386_ (.a(net596),
    .b(net600),
    .o1(_16577_));
 b15bfn000ah1n06x5 input171 (.a(text_in[20]),
    .o(net171));
 b15and002aq1n32x5 _25388_ (.a(net603),
    .b(net606),
    .o(_16579_));
 b15bfn001aq1n06x5 input170 (.a(text_in[1]),
    .o(net170));
 b15nand02aq1n12x5 _25390_ (.a(_16577_),
    .b(_16579_),
    .o1(_16581_));
 b15nandp2an1n12x5 _25391_ (.a(_16460_),
    .b(_16439_),
    .o1(_16582_));
 b15oai022aq1n02x5 _25392_ (.a(_16575_),
    .b(_16576_),
    .c(_16581_),
    .d(_16582_),
    .o1(_16583_));
 b15bfn001aq1n06x5 input169 (.a(text_in[19]),
    .o(net169));
 b15nand02an1n24x5 _25394_ (.a(net620),
    .b(net616),
    .o1(_16585_));
 b15nanb02al1n12x5 _25395_ (.a(net598),
    .b(net606),
    .out0(_16586_));
 b15nandp2al1n04x5 _25396_ (.a(net602),
    .b(net613),
    .o1(_16587_));
 b15xor002ah1n03x5 _25397_ (.a(net600),
    .b(_16587_),
    .out0(_16588_));
 b15norp03aq1n03x5 _25398_ (.a(_16585_),
    .b(_16586_),
    .c(_16588_),
    .o1(_16589_));
 b15oai012as1n06x5 _25399_ (.a(net610),
    .b(_16583_),
    .c(_16589_),
    .o1(_16590_));
 b15and002as1n16x5 _25400_ (.a(net611),
    .b(net609),
    .o(_16591_));
 b15nanb02as1n24x5 _25401_ (.a(net615),
    .b(net618),
    .out0(_16592_));
 b15nor002ar1n02x5 _25402_ (.a(_16592_),
    .b(_16521_),
    .o1(_16593_));
 b15nanb02ah1n12x5 _25403_ (.a(net596),
    .b(net602),
    .out0(_16594_));
 b15nanb02al1n04x5 _25404_ (.a(net614),
    .b(net598),
    .out0(_16595_));
 b15oai022ar1n06x5 _25405_ (.a(_16453_),
    .b(_16594_),
    .c(_16595_),
    .d(net603),
    .o1(_16596_));
 b15inv000al1n48x5 _25406_ (.a(net599),
    .o1(_16597_));
 b15nor002al1n02x5 _25407_ (.a(net605),
    .b(_16597_),
    .o1(_16598_));
 b15aoai13as1n04x5 _25408_ (.a(_16591_),
    .b(_16593_),
    .c(_16596_),
    .d(_16598_),
    .o1(_16599_));
 b15nona23ah1n08x5 _25409_ (.a(_16568_),
    .b(_16573_),
    .c(_16590_),
    .d(_16599_),
    .out0(_16600_));
 b15norp03as1n24x5 _25410_ (.a(net596),
    .b(net600),
    .c(net608),
    .o1(_16601_));
 b15nandp3ar1n02x5 _25411_ (.a(_16475_),
    .b(_16478_),
    .c(_16601_),
    .o1(_16602_));
 b15nandp3ar1n02x5 _25412_ (.a(_16429_),
    .b(_16439_),
    .c(_16473_),
    .o1(_16603_));
 b15norp02ar1n32x5 _25413_ (.a(net613),
    .b(net609),
    .o1(_16604_));
 b15nonb02as1n16x5 _25414_ (.a(net596),
    .b(net600),
    .out0(_16605_));
 b15nand04ah1n03x5 _25415_ (.a(_16592_),
    .b(_16604_),
    .c(_16579_),
    .d(_16605_),
    .o1(_16606_));
 b15and003an1n04x5 _25416_ (.a(_16602_),
    .b(_16603_),
    .c(_16606_),
    .o(_16607_));
 b15nandp3ah1n16x5 _25417_ (.a(net608),
    .b(_16579_),
    .c(_16605_),
    .o1(_16608_));
 b15orn002al1n16x5 _25418_ (.a(net618),
    .b(net614),
    .o(_16609_));
 b15oai022ar1n02x5 _25419_ (.a(net609),
    .b(_16482_),
    .c(_16608_),
    .d(_16609_),
    .o1(_16610_));
 b15bfn001al1n08x5 input168 (.a(text_in[18]),
    .o(net168));
 b15aob012ar1n02x5 _25421_ (.a(_16607_),
    .b(_16610_),
    .c(net613),
    .out0(_16612_));
 b15nonb02as1n16x5 _25422_ (.a(net611),
    .b(net615),
    .out0(_16613_));
 b15and003al1n08x5 _25423_ (.a(_16518_),
    .b(_16579_),
    .c(_16613_),
    .o(_16614_));
 b15nanb02al1n02x5 _25424_ (.a(net599),
    .b(net614),
    .out0(_16615_));
 b15nand02an1n08x5 _25425_ (.a(net599),
    .b(\us13.a[0] ),
    .o1(_16616_));
 b15oai022ar1n02x5 _25426_ (.a(_16538_),
    .b(_16615_),
    .c(_16616_),
    .d(_16497_),
    .o1(_16617_));
 b15aoi013an1n02x5 _25427_ (.a(_16614_),
    .b(_16591_),
    .c(_16617_),
    .d(net598),
    .o1(_16618_));
 b15nonb02as1n16x5 _25428_ (.a(\us13.a[2] ),
    .b(\us13.a[0] ),
    .out0(_16619_));
 b15norp02ah1n08x5 _25429_ (.a(net605),
    .b(net598),
    .o1(_16620_));
 b15nonb02aq1n16x5 _25430_ (.a(\us13.a[3] ),
    .b(net599),
    .out0(_16621_));
 b15xor002ar1n02x5 _25431_ (.a(net603),
    .b(net614),
    .out0(_16622_));
 b15nand04aq1n04x5 _25432_ (.a(_16619_),
    .b(_16620_),
    .c(_16621_),
    .d(_16622_),
    .o1(_16623_));
 b15bfn001al1n08x5 input167 (.a(text_in[17]),
    .o(net167));
 b15and003ar1n02x5 _25434_ (.a(_16508_),
    .b(_16481_),
    .c(_16494_),
    .o(_16625_));
 b15nandp2an1n24x5 _25435_ (.a(net614),
    .b(\us13.a[3] ),
    .o1(_16626_));
 b15norp03ar1n02x5 _25436_ (.a(_16597_),
    .b(_16538_),
    .c(_16626_),
    .o1(_16627_));
 b15oai112as1n02x5 _25437_ (.a(net598),
    .b(_16619_),
    .c(_16625_),
    .d(_16627_),
    .o1(_16628_));
 b15nano23an1n12x5 _25438_ (.a(net606),
    .b(net596),
    .c(net600),
    .d(net602),
    .out0(_16629_));
 b15nand03aq1n12x5 _25439_ (.a(_16490_),
    .b(_16604_),
    .c(_16629_),
    .o1(_16630_));
 b15nand04ar1n06x5 _25440_ (.a(_16481_),
    .b(_16577_),
    .c(_16478_),
    .d(_16544_),
    .o1(_16631_));
 b15nandp2al1n24x5 _25441_ (.a(net613),
    .b(\us13.a[3] ),
    .o1(_16632_));
 b15nor004al1n02x5 _25442_ (.a(net605),
    .b(_16615_),
    .c(_16632_),
    .d(_16594_),
    .o1(_16633_));
 b15nano22ah1n02x5 _25443_ (.a(_16630_),
    .b(_16631_),
    .c(_16633_),
    .out0(_16634_));
 b15nand04ah1n06x5 _25444_ (.a(_16618_),
    .b(_16623_),
    .c(_16628_),
    .d(_16634_),
    .o1(_16635_));
 b15bfn001ah1n12x5 input166 (.a(text_in[16]),
    .o(net166));
 b15aoai13ar1n02x5 _25446_ (.a(net614),
    .b(_16460_),
    .c(net609),
    .d(_16558_),
    .o1(_16637_));
 b15oaoi13aq1n02x5 _25447_ (.a(_16528_),
    .b(_16637_),
    .c(_16544_),
    .d(net613),
    .o1(_16638_));
 b15bfn000ah1n06x5 input165 (.a(text_in[15]),
    .o(net165));
 b15nonb02as1n08x5 _25449_ (.a(net612),
    .b(net610),
    .out0(_16640_));
 b15nand04an1n08x5 _25450_ (.a(_16520_),
    .b(_16435_),
    .c(_16517_),
    .d(_16640_),
    .o1(_16641_));
 b15nanb02al1n16x5 _25451_ (.a(_16522_),
    .b(_16456_),
    .out0(_16642_));
 b15nona23as1n32x5 _25452_ (.a(net604),
    .b(net607),
    .c(net597),
    .d(net601),
    .out0(_16643_));
 b15nand02an1n08x5 _25453_ (.a(_16609_),
    .b(_16604_),
    .o1(_16644_));
 b15oai122as1n16x5 _25454_ (.a(_16641_),
    .b(_16642_),
    .c(_16643_),
    .d(_16581_),
    .e(_16644_),
    .o1(_16645_));
 b15nano23aq1n24x5 _25455_ (.a(net607),
    .b(net600),
    .c(net597),
    .d(net602),
    .out0(_16646_));
 b15bfn001as1n06x5 input164 (.a(text_in[14]),
    .o(net164));
 b15norp03as1n04x5 _25457_ (.a(net615),
    .b(net611),
    .c(net608),
    .o1(_16648_));
 b15nandp2ah1n03x5 _25458_ (.a(_16646_),
    .b(_16648_),
    .o1(_16649_));
 b15nano23as1n24x5 _25459_ (.a(net602),
    .b(net597),
    .c(net600),
    .d(net607),
    .out0(_16650_));
 b15nand02aq1n06x5 _25460_ (.a(net608),
    .b(_16650_),
    .o1(_16651_));
 b15nanb02as1n24x5 _25461_ (.a(\us13.a[2] ),
    .b(net617),
    .out0(_16652_));
 b15aoi012al1n04x5 _25462_ (.a(_16613_),
    .b(_16652_),
    .c(net619),
    .o1(_16653_));
 b15oai012as1n12x5 _25463_ (.a(_16649_),
    .b(_16651_),
    .c(_16653_),
    .o1(_16654_));
 b15bfn001ah1n08x5 input163 (.a(text_in[13]),
    .o(net163));
 b15nonb02ah1n08x5 _25465_ (.a(net606),
    .b(net596),
    .out0(_16656_));
 b15nonb03aq1n12x5 _25466_ (.a(net613),
    .b(net609),
    .c(net599),
    .out0(_16657_));
 b15nandp2as1n02x5 _25467_ (.a(_16656_),
    .b(_16657_),
    .o1(_16658_));
 b15inv020ah1n28x5 _25468_ (.a(net605),
    .o1(_16659_));
 b15oai112al1n08x5 _25469_ (.a(_16659_),
    .b(_16520_),
    .c(_16604_),
    .d(_16591_),
    .o1(_16660_));
 b15aoi112ar1n06x5 _25470_ (.a(net602),
    .b(_16453_),
    .c(_16658_),
    .d(_16660_),
    .o1(_16661_));
 b15nor004aq1n04x5 _25471_ (.a(_16638_),
    .b(_16645_),
    .c(_16654_),
    .d(_16661_),
    .o1(_16662_));
 b15orn002al1n02x5 _25472_ (.a(net602),
    .b(net614),
    .o(_16663_));
 b15norp02ar1n03x5 _25473_ (.a(net609),
    .b(_16663_),
    .o1(_16664_));
 b15nandp2ar1n08x5 _25474_ (.a(net605),
    .b(net596),
    .o1(_16665_));
 b15norp03ar1n02x5 _25475_ (.a(net600),
    .b(_16492_),
    .c(_16665_),
    .o1(_16666_));
 b15nanb02as1n24x5 _25476_ (.a(\us13.a[7] ),
    .b(net601),
    .out0(_16667_));
 b15norp03ar1n02x5 _25477_ (.a(net606),
    .b(_16575_),
    .c(_16667_),
    .o1(_16668_));
 b15oai012aq1n02x5 _25478_ (.a(_16664_),
    .b(_16666_),
    .c(_16668_),
    .o1(_16669_));
 b15norp02as1n08x5 _25479_ (.a(_16439_),
    .b(_16632_),
    .o1(_16670_));
 b15orn002ar1n24x5 _25480_ (.a(\us13.a[5] ),
    .b(net605),
    .o(_16671_));
 b15norp02ar1n12x5 _25481_ (.a(_16671_),
    .b(_16549_),
    .o1(_16672_));
 b15nandp2aq1n32x5 _25482_ (.a(\us13.a[5] ),
    .b(net605),
    .o1(_16673_));
 b15norp02aq1n24x5 _25483_ (.a(_16667_),
    .b(_16673_),
    .o1(_16674_));
 b15aoai13al1n04x5 _25484_ (.a(_16670_),
    .b(_16672_),
    .c(_16674_),
    .d(_16585_),
    .o1(_16675_));
 b15bfn001as1n06x5 input162 (.a(text_in[12]),
    .o(net162));
 b15nonb02ah1n04x5 _25486_ (.a(net617),
    .b(net601),
    .out0(_16677_));
 b15nonb02ar1n08x5 _25487_ (.a(net603),
    .b(net598),
    .out0(_16678_));
 b15nand04ah1n02x5 _25488_ (.a(net606),
    .b(_16619_),
    .c(_16677_),
    .d(_16678_),
    .o1(_16679_));
 b15nandp2aq1n24x5 _25489_ (.a(_16473_),
    .b(_16579_),
    .o1(_16680_));
 b15oaoi13al1n03x5 _25490_ (.a(net610),
    .b(_16679_),
    .c(_16680_),
    .d(_16582_),
    .o1(_16681_));
 b15nor002ah1n24x5 _25491_ (.a(net619),
    .b(net611),
    .o1(_16682_));
 b15nand03al1n03x5 _25492_ (.a(_16475_),
    .b(_16682_),
    .c(_16601_),
    .o1(_16683_));
 b15nonb02ar1n12x5 _25493_ (.a(net600),
    .b(net609),
    .out0(_16684_));
 b15nand04an1n06x5 _25494_ (.a(_16656_),
    .b(_16587_),
    .c(_16663_),
    .d(_16684_),
    .o1(_16685_));
 b15oai012al1n06x5 _25495_ (.a(_16683_),
    .b(_16685_),
    .c(_16682_),
    .o1(_16686_));
 b15nano23al1n06x5 _25496_ (.a(_16669_),
    .b(_16675_),
    .c(_16681_),
    .d(_16686_),
    .out0(_16687_));
 b15nona23as1n08x5 _25497_ (.a(_16612_),
    .b(_16635_),
    .c(_16662_),
    .d(_16687_),
    .out0(_16688_));
 b15nor004as1n12x5 _25498_ (.a(_16531_),
    .b(_16557_),
    .c(_16600_),
    .d(_16688_),
    .o1(_16689_));
 b15xor002as1n12x5 _25499_ (.a(_16424_),
    .b(_16689_),
    .out0(_16690_));
 b15bfn000as1n02x5 input161 (.a(text_in[127]),
    .o(net161));
 b15bfn000ar1n02x5 input160 (.a(text_in[126]),
    .o(net160));
 b15inv000as1n48x5 _25502_ (.a(net764),
    .o1(_16693_));
 b15bfn000ar1n02x5 input159 (.a(text_in[125]),
    .o(net159));
 b15bfn000ar1n02x5 input158 (.a(text_in[124]),
    .o(net158));
 b15bfn000ar1n02x5 input157 (.a(text_in[123]),
    .o(net157));
 b15bfn000ar1n02x5 input156 (.a(text_in[122]),
    .o(net156));
 b15bfn000as1n02x5 input155 (.a(text_in[121]),
    .o(net155));
 b15bfn000ar1n02x5 input154 (.a(text_in[120]),
    .o(net154));
 b15bfn001as1n06x5 input153 (.a(text_in[11]),
    .o(net153));
 b15bfn000ah1n02x5 input152 (.a(text_in[119]),
    .o(net152));
 b15and002aq1n32x5 _25511_ (.a(net749),
    .b(net752),
    .o(_16702_));
 b15bfn000ar1n02x5 input151 (.a(text_in[118]),
    .o(net151));
 b15bfn001aq1n06x5 input150 (.a(text_in[117]),
    .o(net150));
 b15bfn001aq1n06x5 input149 (.a(text_in[116]),
    .o(net149));
 b15bfn000al1n02x5 input148 (.a(text_in[115]),
    .o(net148));
 b15bfn000ah1n02x5 input147 (.a(text_in[114]),
    .o(net147));
 b15nonb02as1n16x5 _25517_ (.a(net746),
    .b(net745),
    .out0(_16708_));
 b15nand04an1n02x5 _25518_ (.a(net754),
    .b(net757),
    .c(_16702_),
    .d(_16708_),
    .o1(_16709_));
 b15norp02as1n48x5 _25519_ (.a(net744),
    .b(net747),
    .o1(_16710_));
 b15nand02ah1n24x5 _25520_ (.a(_16702_),
    .b(_16710_),
    .o1(_16711_));
 b15bfn000as1n03x5 input146 (.a(text_in[113]),
    .o(net146));
 b15orn002aq1n32x5 _25522_ (.a(net756),
    .b(net757),
    .o(_16713_));
 b15bfn000ar1n02x5 input145 (.a(text_in[112]),
    .o(net145));
 b15oaoi13ar1n04x5 _25524_ (.a(_16693_),
    .b(_16709_),
    .c(_16711_),
    .d(_16713_),
    .o1(_16715_));
 b15bfn001as1n06x5 input144 (.a(text_in[111]),
    .o(net144));
 b15bfn001ah1n12x5 input143 (.a(text_in[110]),
    .o(net143));
 b15bfn001ah1n12x5 input142 (.a(text_in[10]),
    .o(net142));
 b15nano22as1n05x5 _25528_ (.a(net760),
    .b(net756),
    .c(net767),
    .out0(_16719_));
 b15bfn001as1n08x5 input141 (.a(text_in[109]),
    .o(net141));
 b15aoi013as1n06x5 _25530_ (.a(_16715_),
    .b(_16719_),
    .c(_16702_),
    .d(_16708_),
    .o1(_16721_));
 b15bfn001as1n08x5 input140 (.a(text_in[108]),
    .o(net140));
 b15bfn001as1n06x5 input139 (.a(text_in[107]),
    .o(net139));
 b15bfn001as1n06x5 input138 (.a(text_in[106]),
    .o(net138));
 b15nonb02as1n16x5 _25534_ (.a(net749),
    .b(net752),
    .out0(_16725_));
 b15and002as1n32x5 _25535_ (.a(net745),
    .b(net746),
    .o(_16726_));
 b15bfn000ar1n02x5 input137 (.a(text_in[105]),
    .o(net137));
 b15nandp2ar1n32x5 _25537_ (.a(net767),
    .b(net756),
    .o1(_16728_));
 b15aoi013ar1n02x5 _25538_ (.a(net761),
    .b(_16725_),
    .c(_16726_),
    .d(_16728_),
    .o1(_16729_));
 b15bfn000ar1n02x5 input136 (.a(text_in[104]),
    .o(net136));
 b15inv000an1n24x5 _25540_ (.a(net749),
    .o1(_16731_));
 b15bfn000ah1n03x5 input135 (.a(text_in[103]),
    .o(net135));
 b15bfn000as1n02x5 input134 (.a(text_in[102]),
    .o(net134));
 b15bfn000an1n02x5 input133 (.a(text_in[101]),
    .o(net133));
 b15norp02as1n02x5 _25544_ (.a(net754),
    .b(net745),
    .o1(_16735_));
 b15bfm201ah1n02x5 input132 (.a(text_in[100]),
    .o(net132));
 b15bfn001al1n08x5 input131 (.a(text_in[0]),
    .o(net131));
 b15bfn000as1n03x5 input130 (.a(rst),
    .o(net130));
 b15nanb02al1n08x5 _25548_ (.a(net752),
    .b(net747),
    .out0(_16739_));
 b15orn003ar1n02x5 _25549_ (.a(_16731_),
    .b(_16735_),
    .c(_16739_),
    .o(_16740_));
 b15inv020as1n64x5 _25550_ (.a(net755),
    .o1(_16741_));
 b15nano23as1n24x5 _25551_ (.a(net753),
    .b(net744),
    .c(net747),
    .d(net751),
    .out0(_16742_));
 b15nand02as1n02x5 _25552_ (.a(_16741_),
    .b(_16742_),
    .o1(_16743_));
 b15aoi012as1n02x5 _25553_ (.a(_16729_),
    .b(_16740_),
    .c(_16743_),
    .o1(_16744_));
 b15bfn001as1n80x5 input129 (.a(ld),
    .o(net129));
 b15nor002aq1n08x5 _25555_ (.a(net761),
    .b(net754),
    .o1(_16746_));
 b15bfn000al1n02x5 input128 (.a(key[9]),
    .o(net128));
 b15nona23as1n32x5 _25557_ (.a(net752),
    .b(net745),
    .c(net746),
    .d(net749),
    .out0(_16748_));
 b15bfn000ah1n02x5 input127 (.a(key[99]),
    .o(net127));
 b15and002aq1n12x5 _25559_ (.a(net760),
    .b(net756),
    .o(_16750_));
 b15aoi012an1n02x5 _25560_ (.a(_16746_),
    .b(_16748_),
    .c(_16750_),
    .o1(_16751_));
 b15bfn000as1n02x5 input126 (.a(key[98]),
    .o(net126));
 b15bfn001ah1n06x5 input125 (.a(key[97]),
    .o(net125));
 b15bfn000ar1n02x5 input124 (.a(key[96]),
    .o(net124));
 b15oai112ah1n06x5 _25564_ (.a(net757),
    .b(_16744_),
    .c(_16751_),
    .d(net765),
    .o1(_16755_));
 b15bfn001as1n06x5 input123 (.a(key[95]),
    .o(net123));
 b15bfn001as1n06x5 input122 (.a(key[94]),
    .o(net122));
 b15nano23as1n24x5 _25567_ (.a(net745),
    .b(net746),
    .c(net749),
    .d(net752),
    .out0(_16758_));
 b15bfn001as1n08x5 input121 (.a(key[93]),
    .o(net121));
 b15nanb02as1n24x5 _25569_ (.a(net766),
    .b(net758),
    .out0(_16760_));
 b15nanb02aq1n24x5 _25570_ (.a(net754),
    .b(net766),
    .out0(_16761_));
 b15nand03al1n02x5 _25571_ (.a(_16758_),
    .b(_16760_),
    .c(_16761_),
    .o1(_16762_));
 b15xnr002as1n16x5 _25572_ (.a(net754),
    .b(net758),
    .out0(_16763_));
 b15nand02ar1n32x5 _25573_ (.a(_16702_),
    .b(_16708_),
    .o1(_16764_));
 b15oaoi13aq1n04x5 _25574_ (.a(net761),
    .b(_16762_),
    .c(_16763_),
    .d(_16764_),
    .o1(_16765_));
 b15bfn000ah1n03x5 input120 (.a(key[92]),
    .o(net120));
 b15bfn000as1n02x5 input119 (.a(key[91]),
    .o(net119));
 b15nonb02ah1n08x5 _25577_ (.a(net755),
    .b(net751),
    .out0(_16768_));
 b15nandp3ar1n08x5 _25578_ (.a(\us31.a[4] ),
    .b(_16708_),
    .c(_16768_),
    .o1(_16769_));
 b15inv000as1n48x5 _25579_ (.a(net761),
    .o1(_16770_));
 b15bfn000ar1n02x5 input118 (.a(key[90]),
    .o(net118));
 b15xor002as1n16x5 _25581_ (.a(net764),
    .b(net759),
    .out0(_16772_));
 b15orn002ar1n02x5 _25582_ (.a(_16770_),
    .b(_16772_),
    .o(_16773_));
 b15inv000al1n80x5 _25583_ (.a(\us31.a[2] ),
    .o1(_16774_));
 b15nand02aq1n24x5 _25584_ (.a(net764),
    .b(_16774_),
    .o1(_16775_));
 b15bfn000ar1n02x5 input117 (.a(key[8]),
    .o(net117));
 b15bfn000al1n02x5 input116 (.a(key[89]),
    .o(net116));
 b15oaoi13an1n04x5 _25587_ (.a(_16769_),
    .b(_16773_),
    .c(_16775_),
    .d(net762),
    .o1(_16778_));
 b15bfm201ah1n02x5 input115 (.a(key[88]),
    .o(net115));
 b15nanb02as1n24x5 _25589_ (.a(net767),
    .b(net760),
    .out0(_16780_));
 b15oai012ar1n02x5 _25590_ (.a(net754),
    .b(_16774_),
    .c(_16780_),
    .o1(_16781_));
 b15nonb03as1n12x5 _25591_ (.a(net747),
    .b(net745),
    .c(net752),
    .out0(_16782_));
 b15and002aq1n16x5 _25592_ (.a(net764),
    .b(net759),
    .o(_16783_));
 b15oai112ar1n04x5 _25593_ (.a(_16731_),
    .b(_16782_),
    .c(_16783_),
    .d(net761),
    .o1(_16784_));
 b15nonb02as1n16x5 _25594_ (.a(net752),
    .b(net749),
    .out0(_16785_));
 b15nandp2aq1n32x5 _25595_ (.a(_16710_),
    .b(_16785_),
    .o1(_16786_));
 b15aoi012al1n02x5 _25596_ (.a(_16781_),
    .b(_16784_),
    .c(_16786_),
    .o1(_16787_));
 b15and002an1n24x5 _25597_ (.a(net763),
    .b(\us31.a[0] ),
    .o(_16788_));
 b15nano23as1n24x5 _25598_ (.a(net749),
    .b(net745),
    .c(net746),
    .d(net752),
    .out0(_16789_));
 b15nandp2aq1n16x5 _25599_ (.a(net754),
    .b(_16789_),
    .o1(_16790_));
 b15bfn000an1n02x5 input114 (.a(key[87]),
    .o(net114));
 b15bfn001ah1n16x5 input113 (.a(key[86]),
    .o(net113));
 b15nand04as1n16x5 _25602_ (.a(net749),
    .b(net752),
    .c(net745),
    .d(net746),
    .o1(_16793_));
 b15oaoi13ar1n03x5 _25603_ (.a(_16788_),
    .b(_16790_),
    .c(_16793_),
    .d(_16713_),
    .o1(_16794_));
 b15nor004ar1n06x5 _25604_ (.a(_16765_),
    .b(_16778_),
    .c(_16787_),
    .d(_16794_),
    .o1(_16795_));
 b15nandp3an1n08x5 _25605_ (.a(_16721_),
    .b(_16755_),
    .c(_16795_),
    .o1(_16796_));
 b15bfn000ah1n03x5 input112 (.a(key[85]),
    .o(net112));
 b15norp02as1n48x5 _25607_ (.a(\us31.a[3] ),
    .b(\us31.a[2] ),
    .o1(_16798_));
 b15bfn000ah1n04x5 input111 (.a(key[84]),
    .o(net111));
 b15nandp3ar1n02x5 _25609_ (.a(_16710_),
    .b(_16798_),
    .c(_16725_),
    .o1(_16800_));
 b15bfn000as1n04x5 input110 (.a(key[83]),
    .o(net110));
 b15nandp3ah1n08x5 _25611_ (.a(net755),
    .b(_16785_),
    .c(_16726_),
    .o1(_16802_));
 b15oaoi13an1n03x5 _25612_ (.a(net762),
    .b(_16800_),
    .c(_16802_),
    .d(_16774_),
    .o1(_16803_));
 b15and002ah1n16x5 _25613_ (.a(net759),
    .b(\us31.a[5] ),
    .o(_16804_));
 b15bfn000ah1n02x5 input109 (.a(key[82]),
    .o(net109));
 b15norp03as1n12x5 _25615_ (.a(net752),
    .b(net745),
    .c(net746),
    .o1(_16806_));
 b15nand02aq1n06x5 _25616_ (.a(_16804_),
    .b(_16806_),
    .o1(_16807_));
 b15bfn000ah1n03x5 input108 (.a(key[81]),
    .o(net108));
 b15bfn000ar1n02x5 input107 (.a(key[80]),
    .o(net107));
 b15nand02ar1n32x5 _25619_ (.a(_16710_),
    .b(_16725_),
    .o1(_16810_));
 b15qbfna2bn1n16x5 _25620_ (.a(_16785_),
    .b(_16726_),
    .o1(_16811_));
 b15aoai13al1n04x5 _25621_ (.a(_16807_),
    .b(net766),
    .c(_16810_),
    .d(_16811_),
    .o1(_16812_));
 b15nonb02ah1n16x5 _25622_ (.a(net761),
    .b(net754),
    .out0(_16813_));
 b15aoi012al1n06x5 _25623_ (.a(_16803_),
    .b(_16812_),
    .c(_16813_),
    .o1(_16814_));
 b15nonb02aq1n16x5 _25624_ (.a(net765),
    .b(net754),
    .out0(_16815_));
 b15bfn000ah1n03x5 input106 (.a(key[7]),
    .o(net106));
 b15bfn000ah1n02x5 input105 (.a(key[79]),
    .o(net105));
 b15bfn000al1n02x5 input104 (.a(key[78]),
    .o(net104));
 b15bfn000an1n02x5 input103 (.a(key[77]),
    .o(net103));
 b15nonb02ah1n12x5 _25629_ (.a(net750),
    .b(net748),
    .out0(_16820_));
 b15bfn000ah1n03x5 input102 (.a(key[76]),
    .o(net102));
 b15bfn000ah1n02x5 input101 (.a(key[75]),
    .o(net101));
 b15nonb02al1n02x5 _25632_ (.a(net760),
    .b(net750),
    .out0(_16823_));
 b15nonb02as1n12x5 _25633_ (.a(net748),
    .b(net753),
    .out0(_16824_));
 b15aoi022ar1n08x5 _25634_ (.a(net753),
    .b(_16820_),
    .c(_16823_),
    .d(_16824_),
    .o1(_16825_));
 b15nor003al1n08x5 _25635_ (.a(_16774_),
    .b(net744),
    .c(_16825_),
    .o1(_16826_));
 b15and002ar1n08x5 _25636_ (.a(\us31.a[4] ),
    .b(_16708_),
    .o(_16827_));
 b15bfn000an1n02x5 input100 (.a(key[74]),
    .o(net100));
 b15aoai13ar1n08x5 _25638_ (.a(_16815_),
    .b(_16826_),
    .c(_16827_),
    .d(_16774_),
    .o1(_16829_));
 b15nonb02as1n16x5 _25639_ (.a(net745),
    .b(net746),
    .out0(_16830_));
 b15norp02ah1n32x5 _25640_ (.a(net749),
    .b(net752),
    .o1(_16831_));
 b15nandp2al1n48x5 _25641_ (.a(_16830_),
    .b(_16831_),
    .o1(_16832_));
 b15bfn000aq1n02x5 input99 (.a(key[73]),
    .o(net99));
 b15nonb02aq1n16x5 _25643_ (.a(net755),
    .b(net763),
    .out0(_16834_));
 b15nand02ah1n24x5 _25644_ (.a(_16774_),
    .b(_16834_),
    .o1(_16835_));
 b15nonb02as1n16x5 _25645_ (.a(net767),
    .b(net760),
    .out0(_16836_));
 b15bfn000al1n02x5 input98 (.a(key[72]),
    .o(net98));
 b15xor002al1n02x5 _25647_ (.a(net753),
    .b(_16836_),
    .out0(_16838_));
 b15nanb02as1n24x5 _25648_ (.a(\us31.a[2] ),
    .b(\us31.a[3] ),
    .out0(_16839_));
 b15bfn000as1n02x5 input97 (.a(key[71]),
    .o(net97));
 b15nand03an1n06x5 _25650_ (.a(net750),
    .b(net744),
    .c(net748),
    .o1(_16841_));
 b15orn002al1n02x5 _25651_ (.a(_16839_),
    .b(_16841_),
    .o(_16842_));
 b15oai022an1n06x5 _25652_ (.a(_16832_),
    .b(_16835_),
    .c(_16838_),
    .d(_16842_),
    .o1(_16843_));
 b15and002al1n32x5 _25653_ (.a(net756),
    .b(net757),
    .o(_16844_));
 b15nonb02ah1n03x5 _25654_ (.a(net766),
    .b(net749),
    .out0(_16845_));
 b15nonb02an1n06x5 _25655_ (.a(net749),
    .b(net766),
    .out0(_16846_));
 b15aoi022an1n04x5 _25656_ (.a(_16726_),
    .b(_16845_),
    .c(_16846_),
    .d(_16710_),
    .o1(_16847_));
 b15nano22ah1n06x5 _25657_ (.a(\us31.a[4] ),
    .b(_16844_),
    .c(_16847_),
    .out0(_16848_));
 b15nanb02as1n24x5 _25658_ (.a(net753),
    .b(net750),
    .out0(_16849_));
 b15nandp2as1n12x5 _25659_ (.a(net744),
    .b(net748),
    .o1(_16850_));
 b15nor003ar1n12x5 _25660_ (.a(_16713_),
    .b(_16849_),
    .c(_16850_),
    .o1(_16851_));
 b15nand02ar1n24x5 _25661_ (.a(net762),
    .b(net766),
    .o1(_16852_));
 b15aoi112aq1n08x5 _25662_ (.a(_16843_),
    .b(_16848_),
    .c(_16851_),
    .d(_16852_),
    .o1(_16853_));
 b15norp03an1n03x5 _25663_ (.a(net751),
    .b(\us31.a[7] ),
    .c(net748),
    .o1(_16854_));
 b15nanb02as1n24x5 _25664_ (.a(net763),
    .b(net764),
    .out0(_16855_));
 b15nanb02as1n24x5 _25665_ (.a(\us31.a[3] ),
    .b(\us31.a[2] ),
    .out0(_16856_));
 b15oai012aq1n02x5 _25666_ (.a(_16854_),
    .b(_16855_),
    .c(_16856_),
    .o1(_16857_));
 b15bfn000ar1n02x5 input96 (.a(key[70]),
    .o(net96));
 b15oaoi13ar1n04x5 _25668_ (.a(_16857_),
    .b(net755),
    .c(\us31.a[4] ),
    .d(_16788_),
    .o1(_16859_));
 b15nonb02as1n16x5 _25669_ (.a(\us31.a[0] ),
    .b(\us31.a[2] ),
    .out0(_16860_));
 b15nonb02as1n16x5 _25670_ (.a(net757),
    .b(net756),
    .out0(_16861_));
 b15bfn000as1n02x5 input95 (.a(key[6]),
    .o(net95));
 b15bfn000ar1n02x5 input94 (.a(key[69]),
    .o(net94));
 b15aoai13al1n06x5 _25673_ (.a(net763),
    .b(_16860_),
    .c(_16861_),
    .d(_16693_),
    .o1(_16864_));
 b15oai112an1n16x5 _25674_ (.a(_16859_),
    .b(_16864_),
    .c(net759),
    .d(\us31.a[4] ),
    .o1(_16865_));
 b15nand04aq1n16x5 _25675_ (.a(_16814_),
    .b(_16829_),
    .c(_16853_),
    .d(_16865_),
    .o1(_16866_));
 b15nona23an1n32x5 _25676_ (.a(net749),
    .b(net747),
    .c(net745),
    .d(net752),
    .out0(_16867_));
 b15oai012ar1n02x5 _25677_ (.a(_16774_),
    .b(_16867_),
    .c(_16761_),
    .o1(_16868_));
 b15bfn000ah1n02x5 input93 (.a(key[68]),
    .o(net93));
 b15nor003al1n03x5 _25679_ (.a(net765),
    .b(net756),
    .c(net749),
    .o1(_16870_));
 b15nand02an1n04x5 _25680_ (.a(_16830_),
    .b(_16870_),
    .o1(_16871_));
 b15norp02as1n12x5 _25681_ (.a(net756),
    .b(net751),
    .o1(_16872_));
 b15and002aq1n16x5 _25682_ (.a(net754),
    .b(net749),
    .o(_16873_));
 b15oai112an1n08x5 _25683_ (.a(net765),
    .b(_16708_),
    .c(_16872_),
    .d(_16873_),
    .o1(_16874_));
 b15aoi112aq1n08x5 _25684_ (.a(net761),
    .b(net752),
    .c(_16871_),
    .d(_16874_),
    .o1(_16875_));
 b15bfn000ar1n02x5 input92 (.a(key[67]),
    .o(net92));
 b15oai022ar1n02x5 _25686_ (.a(_16741_),
    .b(_16711_),
    .c(_16761_),
    .d(_16832_),
    .o1(_16877_));
 b15bfn000an1n02x5 input91 (.a(key[66]),
    .o(net91));
 b15bfn000al1n02x5 input90 (.a(key[65]),
    .o(net90));
 b15aoi112al1n02x5 _25689_ (.a(_16868_),
    .b(_16875_),
    .c(_16877_),
    .d(net761),
    .o1(_16880_));
 b15inv040aq1n05x5 _25690_ (.a(net747),
    .o1(_16881_));
 b15aoi022ar1n04x5 _25691_ (.a(_16702_),
    .b(_16735_),
    .c(_16831_),
    .d(net745),
    .o1(_16882_));
 b15nor003as1n04x5 _25692_ (.a(_16693_),
    .b(_16881_),
    .c(_16882_),
    .o1(_16883_));
 b15bfn000ar1n02x5 input89 (.a(key[64]),
    .o(net89));
 b15bfn000ah1n04x5 input88 (.a(key[63]),
    .o(net88));
 b15bfn000ar1n02x5 input87 (.a(key[62]),
    .o(net87));
 b15nona22al1n16x5 _25696_ (.a(net763),
    .b(net755),
    .c(net764),
    .out0(_16887_));
 b15nona23ah1n32x5 _25697_ (.a(\us31.a[5] ),
    .b(\us31.a[4] ),
    .c(\us31.a[7] ),
    .d(\us31.a[6] ),
    .out0(_16888_));
 b15bfn001as1n06x5 input86 (.a(key[61]),
    .o(net86));
 b15oai122an1n08x5 _25699_ (.a(net758),
    .b(_16832_),
    .c(_16887_),
    .d(_16888_),
    .e(_16770_),
    .o1(_16890_));
 b15oab012ah1n03x5 _25700_ (.a(_16880_),
    .b(_16883_),
    .c(_16890_),
    .out0(_16891_));
 b15nonb02ah1n16x5 _25701_ (.a(net756),
    .b(net757),
    .out0(_16892_));
 b15nand04aq1n02x5 _25702_ (.a(_16785_),
    .b(_16726_),
    .c(_16892_),
    .d(_16788_),
    .o1(_16893_));
 b15norp02al1n48x5 _25703_ (.a(net760),
    .b(net767),
    .o1(_16894_));
 b15nand03an1n02x5 _25704_ (.a(_16798_),
    .b(_16789_),
    .c(_16894_),
    .o1(_16895_));
 b15nano22as1n24x5 _25705_ (.a(\us31.a[4] ),
    .b(\us31.a[7] ),
    .c(\us31.a[6] ),
    .out0(_16896_));
 b15nand02as1n32x5 _25706_ (.a(net749),
    .b(_16896_),
    .o1(_16897_));
 b15nandp2an1n48x5 _25707_ (.a(net764),
    .b(net759),
    .o1(_16898_));
 b15nandp2al1n08x5 _25708_ (.a(_16750_),
    .b(_16898_),
    .o1(_16899_));
 b15oai112al1n06x5 _25709_ (.a(_16893_),
    .b(_16895_),
    .c(_16897_),
    .d(_16899_),
    .o1(_16900_));
 b15bfn001ah1n08x5 input85 (.a(key[60]),
    .o(net85));
 b15andc04ah1n12x5 _25711_ (.a(net750),
    .b(net753),
    .c(net744),
    .d(net748),
    .o(_16902_));
 b15nand02an1n16x5 _25712_ (.a(net757),
    .b(_16902_),
    .o1(_16903_));
 b15nonb03al1n03x5 _25713_ (.a(_16728_),
    .b(_16813_),
    .c(_16903_),
    .out0(_16904_));
 b15nano23as1n24x5 _25714_ (.a(net752),
    .b(net746),
    .c(net745),
    .d(net749),
    .out0(_16905_));
 b15aoi022ar1n02x5 _25715_ (.a(_16742_),
    .b(_16892_),
    .c(_16861_),
    .d(_16905_),
    .o1(_16906_));
 b15nonb02as1n16x5 _25716_ (.a(net760),
    .b(net767),
    .out0(_16907_));
 b15nor002ah1n06x5 _25717_ (.a(_16907_),
    .b(_16836_),
    .o1(_16908_));
 b15nor002ar1n02x5 _25718_ (.a(_16906_),
    .b(_16908_),
    .o1(_16909_));
 b15orn003ah1n08x5 _25719_ (.a(_16900_),
    .b(_16904_),
    .c(_16909_),
    .o(_16910_));
 b15bfn000ar1n02x5 input84 (.a(key[5]),
    .o(net84));
 b15norp02ar1n03x5 _25721_ (.a(net758),
    .b(_16748_),
    .o1(_16912_));
 b15bfn000aq1n02x5 input83 (.a(key[59]),
    .o(net83));
 b15oab012ar1n02x5 _25723_ (.a(_16912_),
    .b(_16897_),
    .c(net761),
    .out0(_16914_));
 b15nano23an1n24x5 _25724_ (.a(net749),
    .b(net746),
    .c(net745),
    .d(net752),
    .out0(_16915_));
 b15bfn000an1n02x5 input82 (.a(key[58]),
    .o(net82));
 b15aoi022ar1n02x5 _25726_ (.a(net761),
    .b(_16915_),
    .c(_16896_),
    .d(_16804_),
    .o1(_16917_));
 b15oaoi13al1n02x5 _25727_ (.a(net754),
    .b(_16914_),
    .c(_16917_),
    .d(_16693_),
    .o1(_16918_));
 b15nandp3ar1n12x5 _25728_ (.o1(_16919_),
    .a(_16774_),
    .b(_16710_),
    .c(_16725_));
 b15bfn000ar1n02x5 input81 (.a(key[57]),
    .o(net81));
 b15oai112ar1n04x5 _25730_ (.a(net761),
    .b(_16919_),
    .c(_16898_),
    .d(_16867_),
    .o1(_16921_));
 b15oai022ar1n02x5 _25731_ (.a(_16867_),
    .b(_16760_),
    .c(_16810_),
    .d(_16693_),
    .o1(_16922_));
 b15bfn000an1n02x5 input80 (.a(key[56]),
    .o(net80));
 b15oai112ah1n04x5 _25733_ (.a(net754),
    .b(_16921_),
    .c(_16922_),
    .d(net761),
    .o1(_16924_));
 b15nona22ah1n04x5 _25734_ (.a(_16910_),
    .b(_16918_),
    .c(_16924_),
    .out0(_16925_));
 b15nor004as1n12x5 _25735_ (.a(_16796_),
    .b(_16866_),
    .c(_16891_),
    .d(_16925_),
    .o1(_16926_));
 b15and002as1n04x5 _25736_ (.a(net722),
    .b(net717),
    .o(_16927_));
 b15nanb02as1n24x5 _25737_ (.a(net726),
    .b(net720),
    .out0(_16928_));
 b15nanb02ah1n16x5 _25738_ (.a(net720),
    .b(net726),
    .out0(_16929_));
 b15oai022ar1n02x5 _25739_ (.a(_16283_),
    .b(_16928_),
    .c(_16929_),
    .d(_16221_),
    .o1(_16930_));
 b15and003ar1n02x5 _25740_ (.a(net737),
    .b(_16927_),
    .c(_16930_),
    .o(_16931_));
 b15nano22ah1n16x5 _25741_ (.a(net717),
    .b(net720),
    .c(net726),
    .out0(_16932_));
 b15and003ar1n02x5 _25742_ (.a(_16283_),
    .b(_16189_),
    .c(_16932_),
    .o(_16933_));
 b15orn003an1n04x5 _25743_ (.a(_16226_),
    .b(_16931_),
    .c(_16933_),
    .o(_16934_));
 b15nonb02ar1n12x5 _25744_ (.a(net733),
    .b(net722),
    .out0(_16935_));
 b15nandp2ah1n32x5 _25745_ (.a(\us02.a[1] ),
    .b(net741),
    .o1(_16936_));
 b15bfn001ah1n06x5 input79 (.a(key[55]),
    .o(net79));
 b15norp03ar1n02x5 _25747_ (.a(_16276_),
    .b(_16314_),
    .c(_16936_),
    .o1(_16938_));
 b15nonb02ah1n06x5 _25748_ (.a(net719),
    .b(net738),
    .out0(_16939_));
 b15oai012ar1n08x5 _25749_ (.a(_16206_),
    .b(_16203_),
    .c(_16283_),
    .o1(_16940_));
 b15aoai13ar1n03x5 _25750_ (.a(_16935_),
    .b(_16938_),
    .c(_16939_),
    .d(_16940_),
    .o1(_16941_));
 b15xor002an1n04x5 _25751_ (.a(net738),
    .b(_16193_),
    .out0(_16942_));
 b15bfn000as1n03x5 input78 (.a(key[54]),
    .o(net78));
 b15aoi022ah1n08x5 _25753_ (.a(_16351_),
    .b(_16936_),
    .c(_16942_),
    .d(_16328_),
    .o1(_16944_));
 b15bfn001aq1n06x5 input77 (.a(key[53]),
    .o(net77));
 b15oai013as1n06x5 _25755_ (.a(_16941_),
    .b(_16944_),
    .c(net733),
    .d(_16276_),
    .o1(_16946_));
 b15nandp2ah1n04x5 _25756_ (.a(_16342_),
    .b(_16214_),
    .o1(_16947_));
 b15oai022aq1n16x5 _25757_ (.a(_16947_),
    .b(_16282_),
    .c(_16420_),
    .d(_16283_),
    .o1(_16948_));
 b15bfn001ah1n06x5 input76 (.a(key[52]),
    .o(net76));
 b15oai022ah1n12x5 _25759_ (.a(_16934_),
    .b(_16946_),
    .c(_16948_),
    .d(net729),
    .o1(_16950_));
 b15nona22ar1n32x5 _25760_ (.a(net726),
    .b(net717),
    .c(net719),
    .out0(_16951_));
 b15nanb02ah1n24x5 _25761_ (.a(net730),
    .b(net723),
    .out0(_16952_));
 b15orn002al1n02x5 _25762_ (.a(_16951_),
    .b(_16952_),
    .o(_16953_));
 b15aoi022aq1n06x5 _25763_ (.a(_16223_),
    .b(_16354_),
    .c(_16932_),
    .d(net729),
    .o1(_16954_));
 b15inv040aq1n04x5 _25764_ (.a(_16274_),
    .o1(_16955_));
 b15oaoi13al1n08x5 _25765_ (.a(net733),
    .b(_16953_),
    .c(_16954_),
    .d(_16955_),
    .o1(_16956_));
 b15norp02an1n16x5 _25766_ (.a(net730),
    .b(_16248_),
    .o1(_16957_));
 b15nand02ah1n32x5 _25767_ (.a(_16301_),
    .b(_16259_),
    .o1(_16958_));
 b15oai012aq1n06x5 _25768_ (.a(_16391_),
    .b(_16958_),
    .c(net739),
    .o1(_16959_));
 b15and002an1n24x5 _25769_ (.a(net738),
    .b(net740),
    .o(_16960_));
 b15nandp2an1n04x5 _25770_ (.a(_16351_),
    .b(_16960_),
    .o1(_16961_));
 b15bfn000ah1n02x5 input75 (.a(key[51]),
    .o(net75));
 b15oai012as1n03x5 _25772_ (.a(_16961_),
    .b(_16225_),
    .c(_16342_),
    .o1(_16963_));
 b15oaoi13al1n04x5 _25773_ (.a(_16956_),
    .b(_16957_),
    .c(_16959_),
    .d(_16963_),
    .o1(_16964_));
 b15orn002al1n12x5 _25774_ (.a(net739),
    .b(net741),
    .o(_16965_));
 b15nanb02as1n08x5 _25775_ (.a(net723),
    .b(net738),
    .out0(_16966_));
 b15nanb02al1n16x5 _25776_ (.a(net725),
    .b(net718),
    .out0(_16967_));
 b15oai022an1n02x5 _25777_ (.a(_16278_),
    .b(_16372_),
    .c(_16966_),
    .d(_16967_),
    .o1(_16968_));
 b15nand04al1n02x5 _25778_ (.a(net732),
    .b(net719),
    .c(_16965_),
    .d(_16968_),
    .o1(_16969_));
 b15nonb02as1n16x5 _25779_ (.a(net737),
    .b(net740),
    .out0(_16970_));
 b15nor004al1n02x5 _25780_ (.a(_16276_),
    .b(_16314_),
    .c(_16970_),
    .d(_16952_),
    .o1(_16971_));
 b15nanb02an1n16x5 _25781_ (.a(net738),
    .b(net730),
    .out0(_16972_));
 b15oai022ar1n02x5 _25782_ (.a(_16280_),
    .b(_16337_),
    .c(_16972_),
    .d(_16235_),
    .o1(_16973_));
 b15aoi012ar1n02x5 _25783_ (.a(_16971_),
    .b(_16973_),
    .c(_16258_),
    .o1(_16974_));
 b15aob012as1n02x5 _25784_ (.a(net733),
    .b(_16969_),
    .c(_16974_),
    .out0(_16975_));
 b15oai013ar1n02x5 _25785_ (.a(_16283_),
    .b(_16318_),
    .c(_16414_),
    .d(net737),
    .o1(_16976_));
 b15norp02ah1n24x5 _25786_ (.a(_16237_),
    .b(_16280_),
    .o1(_16977_));
 b15aoi013an1n02x5 _25787_ (.a(_16976_),
    .b(_16977_),
    .c(_16401_),
    .d(_16248_),
    .o1(_16978_));
 b15nanb02as1n24x5 _25788_ (.a(net718),
    .b(net719),
    .out0(_16979_));
 b15nor002al1n24x5 _25789_ (.a(_16313_),
    .b(_16979_),
    .o1(_16980_));
 b15inv040aq1n04x5 _25790_ (.a(_16377_),
    .o1(_16981_));
 b15qgbxo2an1n05x5 _25791_ (.a(net733),
    .b(net719),
    .out0(_16982_));
 b15norp02aq1n03x5 _25792_ (.a(_16372_),
    .b(_16952_),
    .o1(_16983_));
 b15aoi022ah1n06x5 _25793_ (.a(_16980_),
    .b(_16981_),
    .c(_16982_),
    .d(_16983_),
    .o1(_16984_));
 b15bfn000ar1n02x5 input74 (.a(key[50]),
    .o(net74));
 b15nandp2ar1n24x5 _25795_ (.a(\us02.a[1] ),
    .b(net731),
    .o1(_16986_));
 b15oai022ar1n02x5 _25796_ (.a(_16280_),
    .b(_16986_),
    .c(_16979_),
    .d(_16972_),
    .o1(_16987_));
 b15norp02al1n12x5 _25797_ (.a(net739),
    .b(net730),
    .o1(_16988_));
 b15and002as1n04x5 _25798_ (.a(_16328_),
    .b(_16988_),
    .o(_16989_));
 b15oai112ah1n04x5 _25799_ (.a(net726),
    .b(_16418_),
    .c(_16987_),
    .d(_16989_),
    .o1(_16990_));
 b15aoi013ar1n04x5 _25800_ (.a(_16978_),
    .b(_16984_),
    .c(_16990_),
    .d(net742),
    .o1(_16991_));
 b15bfn000ah1n06x5 input73 (.a(key[4]),
    .o(net73));
 b15nanb02as1n24x5 _25802_ (.a(net732),
    .b(net736),
    .out0(_16993_));
 b15bfn000ar1n02x5 input72 (.a(key[49]),
    .o(net72));
 b15nanb02as1n24x5 _25804_ (.a(net736),
    .b(net732),
    .out0(_16995_));
 b15aoi112ar1n02x5 _25805_ (.a(net742),
    .b(_16336_),
    .c(_16993_),
    .d(_16995_),
    .o1(_16996_));
 b15nonb02ah1n16x5 _25806_ (.a(\us02.a[0] ),
    .b(net732),
    .out0(_16997_));
 b15aoi013as1n03x5 _25807_ (.a(_16996_),
    .b(_16935_),
    .c(_16997_),
    .d(_16223_),
    .o1(_16998_));
 b15nor002as1n06x5 _25808_ (.a(_16235_),
    .b(_16310_),
    .o1(_16999_));
 b15nor002an1n03x5 _25809_ (.a(_16248_),
    .b(_16323_),
    .o1(_17000_));
 b15oai012aq1n03x5 _25810_ (.a(_16999_),
    .b(_16320_),
    .c(_17000_),
    .o1(_17001_));
 b15nanb02ah1n02x5 _25811_ (.a(_16327_),
    .b(_16226_),
    .out0(_17002_));
 b15aoi013ar1n04x5 _25812_ (.a(_16342_),
    .b(_16998_),
    .c(_17001_),
    .d(_17002_),
    .o1(_17003_));
 b15nano23al1n08x5 _25813_ (.a(_16964_),
    .b(_16975_),
    .c(_16991_),
    .d(_17003_),
    .out0(_17004_));
 b15nand04as1n16x5 _25814_ (.a(net724),
    .b(net727),
    .c(net718),
    .d(net721),
    .o1(_17005_));
 b15nor003al1n04x5 _25815_ (.a(net735),
    .b(_17005_),
    .c(_16379_),
    .o1(_17006_));
 b15bfn000ar1n02x5 input71 (.a(key[48]),
    .o(net71));
 b15nano23as1n24x5 _25817_ (.a(\us02.a[7] ),
    .b(\us02.a[6] ),
    .c(\us02.a[5] ),
    .d(net728),
    .out0(_17008_));
 b15xnr002as1n12x5 _25818_ (.a(net743),
    .b(net736),
    .out0(_17009_));
 b15aoi013ah1n06x5 _25819_ (.a(_17006_),
    .b(_17008_),
    .c(_17009_),
    .d(_16342_),
    .o1(_17010_));
 b15nor004ar1n02x5 _25820_ (.a(net717),
    .b(_16986_),
    .c(_16398_),
    .d(_16333_),
    .o1(_17011_));
 b15nor004ar1n03x5 _25821_ (.a(net724),
    .b(_16203_),
    .c(_16318_),
    .d(_16379_),
    .o1(_17012_));
 b15nor002an1n02x5 _25822_ (.a(_17011_),
    .b(_17012_),
    .o1(_17013_));
 b15oai022as1n06x5 _25823_ (.a(net731),
    .b(_17010_),
    .c(_17013_),
    .d(net721),
    .o1(_17014_));
 b15nanb02an1n24x5 _25824_ (.a(net737),
    .b(net742),
    .out0(_17015_));
 b15nor004ah1n03x5 _25825_ (.a(_16237_),
    .b(_16280_),
    .c(_17015_),
    .d(_16993_),
    .o1(_17016_));
 b15nanb02al1n06x5 _25826_ (.a(net735),
    .b(net719),
    .out0(_17017_));
 b15nor004an1n03x5 _25827_ (.a(net724),
    .b(_16986_),
    .c(_16203_),
    .d(_17017_),
    .o1(_17018_));
 b15nor003an1n06x5 _25828_ (.a(_16381_),
    .b(_16414_),
    .c(_16936_),
    .o1(_17019_));
 b15norp03al1n04x5 _25829_ (.a(_16995_),
    .b(_17015_),
    .c(_16396_),
    .o1(_17020_));
 b15nor004al1n06x5 _25830_ (.a(_17016_),
    .b(_17018_),
    .c(_17019_),
    .d(_17020_),
    .o1(_17021_));
 b15nanb03al1n12x5 _25831_ (.a(net724),
    .b(net727),
    .c(net717),
    .out0(_17022_));
 b15nand03al1n02x5 _25832_ (.a(net742),
    .b(net729),
    .c(net720),
    .o1(_17023_));
 b15orn002ar1n03x5 _25833_ (.a(net729),
    .b(net720),
    .o(_17024_));
 b15aoi112ah1n03x5 _25834_ (.a(_16377_),
    .b(_17022_),
    .c(_17023_),
    .d(_17024_),
    .o1(_17025_));
 b15norp02aq1n03x5 _25835_ (.a(net726),
    .b(net718),
    .o1(_17026_));
 b15aob012an1n03x5 _25836_ (.a(_16358_),
    .b(_17026_),
    .c(_16193_),
    .out0(_17027_));
 b15norp02ah1n12x5 _25837_ (.a(net729),
    .b(net733),
    .o1(_17028_));
 b15aoi013an1n03x5 _25838_ (.a(_17025_),
    .b(_17027_),
    .c(_17028_),
    .d(_16939_),
    .o1(_17029_));
 b15and002an1n02x5 _25839_ (.a(_16291_),
    .b(_16350_),
    .o(_17030_));
 b15nor002aq1n12x5 _25840_ (.a(net723),
    .b(net719),
    .o1(_17031_));
 b15cmbn22as1n02x5 _25841_ (.clk1(_17031_),
    .clk2(_16370_),
    .clkout(_17032_),
    .s(net729));
 b15norp02ar1n08x5 _25842_ (.a(_17015_),
    .b(_16993_),
    .o1(_17033_));
 b15oai012ar1n02x5 _25843_ (.a(_16336_),
    .b(_16314_),
    .c(_16313_),
    .o1(_17034_));
 b15aoi022aq1n02x5 _25844_ (.a(_17030_),
    .b(_17032_),
    .c(_17033_),
    .d(_17034_),
    .o1(_17035_));
 b15nor004ar1n04x5 _25845_ (.a(net737),
    .b(net729),
    .c(_16358_),
    .d(_16982_),
    .o1(_17036_));
 b15oab012al1n03x5 _25846_ (.a(_17036_),
    .b(_16318_),
    .c(_16186_),
    .out0(_17037_));
 b15nand04ah1n08x5 _25847_ (.a(_17021_),
    .b(_17029_),
    .c(_17035_),
    .d(_17037_),
    .o1(_17038_));
 b15nandp3ar1n04x5 _25848_ (.a(_16233_),
    .b(_16340_),
    .c(_16399_),
    .o1(_17039_));
 b15nandp3aq1n03x5 _25849_ (.a(net734),
    .b(_16247_),
    .c(_16325_),
    .o1(_17040_));
 b15and002ah1n16x5 _25850_ (.a(net729),
    .b(net733),
    .o(_17041_));
 b15nand04ah1n06x5 _25851_ (.a(_16223_),
    .b(_16224_),
    .c(_16399_),
    .d(_17041_),
    .o1(_17042_));
 b15nandp3ar1n12x5 _25852_ (.o1(_17043_),
    .a(_17039_),
    .b(_17040_),
    .c(_17042_));
 b15and002ah1n04x5 _25853_ (.a(_16202_),
    .b(_16293_),
    .o(_17044_));
 b15nona23an1n16x5 _25854_ (.a(net727),
    .b(net721),
    .c(net718),
    .d(net724),
    .out0(_17045_));
 b15norp02as1n03x5 _25855_ (.a(net737),
    .b(_17045_),
    .o1(_17046_));
 b15oab012ar1n02x5 _25856_ (.a(_16226_),
    .b(_17044_),
    .c(_17046_),
    .out0(_17047_));
 b15nor002ah1n04x5 _25857_ (.a(_16383_),
    .b(_16361_),
    .o1(_17048_));
 b15aoi012as1n02x5 _25858_ (.a(net731),
    .b(_16965_),
    .c(_16936_),
    .o1(_17049_));
 b15aoai13aq1n08x5 _25859_ (.a(_16248_),
    .b(_17048_),
    .c(_17049_),
    .d(_16315_),
    .o1(_17050_));
 b15oai013as1n03x5 _25860_ (.a(net737),
    .b(_16235_),
    .c(_16237_),
    .d(_16997_),
    .o1(_17051_));
 b15nanb02al1n12x5 _25861_ (.a(net733),
    .b(net722),
    .out0(_17052_));
 b15orn002aq1n04x5 _25862_ (.a(net726),
    .b(net720),
    .o(_17053_));
 b15aoi112an1n04x5 _25863_ (.a(_17052_),
    .b(_17053_),
    .c(net729),
    .d(_16390_),
    .o1(_17054_));
 b15inv020as1n16x5 _25864_ (.a(net717),
    .o1(_17055_));
 b15oai112as1n12x5 _25865_ (.a(_17051_),
    .b(_17054_),
    .c(_16283_),
    .d(_17055_),
    .o1(_17056_));
 b15nona23ah1n05x5 _25866_ (.a(_17043_),
    .b(_17047_),
    .c(_17050_),
    .d(_17056_),
    .out0(_17057_));
 b15nano22ar1n02x5 _25867_ (.a(net737),
    .b(net740),
    .c(net722),
    .out0(_17058_));
 b15aoi022ar1n02x5 _25868_ (.a(_16390_),
    .b(_16273_),
    .c(_16419_),
    .d(_17058_),
    .o1(_17059_));
 b15aoai13ar1n02x5 _25869_ (.a(_16274_),
    .b(_16273_),
    .c(net740),
    .d(_16932_),
    .o1(_17060_));
 b15aob012an1n06x5 _25870_ (.a(_17041_),
    .b(_17059_),
    .c(_17060_),
    .out0(_17061_));
 b15nor002ah1n06x5 _25871_ (.a(\us02.a[1] ),
    .b(_16318_),
    .o1(_17062_));
 b15ao0022ar1n02x5 _25872_ (.a(_16194_),
    .b(_16292_),
    .c(_16295_),
    .d(_16191_),
    .o(_17063_));
 b15norp02ar1n02x5 _25873_ (.a(_16342_),
    .b(_17055_),
    .o1(_17064_));
 b15aoi022al1n02x5 _25874_ (.a(_16977_),
    .b(_17062_),
    .c(_17063_),
    .d(_17064_),
    .o1(_17065_));
 b15oai012an1n06x5 _25875_ (.a(_17061_),
    .b(_17065_),
    .c(net742),
    .o1(_17066_));
 b15nor004an1n12x5 _25876_ (.a(_17014_),
    .b(_17038_),
    .c(_17057_),
    .d(_17066_),
    .o1(_17067_));
 b15nandp3as1n24x5 _25877_ (.a(_16950_),
    .b(_17004_),
    .c(_17067_),
    .o1(_17068_));
 b15xnr002aq1n16x5 _25878_ (.a(_16926_),
    .b(_17068_),
    .out0(_17069_));
 b15xor003aq1n04x5 _25879_ (.a(_16168_),
    .b(_16690_),
    .c(_17069_),
    .out0(_17070_));
 b15norp02an1n12x5 _25880_ (.a(net540),
    .b(_17070_),
    .o1(_17071_));
 b15inv020ah1n12x5 _25881_ (.a(\text_in_r[32] ),
    .o1(_17072_));
 b15aoi012aq1n08x5 _25882_ (.a(_17071_),
    .b(_17072_),
    .c(ld_r),
    .o1(_17073_));
 b15xor002as1n16x5 _25883_ (.a(\u0.w[2][0] ),
    .b(_17073_),
    .out0(_00113_));
 b15bfn001as1n06x5 input70 (.a(key[47]),
    .o(net70));
 b15bfn000as1n03x5 input69 (.a(key[46]),
    .o(net69));
 b15norp02ar1n04x5 _25886_ (.a(_16460_),
    .b(_16643_),
    .o1(_17076_));
 b15norp02ar1n16x5 _25887_ (.a(_16438_),
    .b(_16538_),
    .o1(_17077_));
 b15bfn001as1n06x5 input68 (.a(key[45]),
    .o(net68));
 b15aoai13ar1n02x5 _25889_ (.a(net616),
    .b(_17076_),
    .c(_17077_),
    .d(_16460_),
    .o1(_17079_));
 b15nand02ah1n12x5 _25890_ (.a(net605),
    .b(\us13.a[2] ),
    .o1(_17080_));
 b15oai022aq1n04x5 _25891_ (.a(net606),
    .b(_16667_),
    .c(_16549_),
    .d(_17080_),
    .o1(_17081_));
 b15bfn001as1n08x5 input67 (.a(key[44]),
    .o(net67));
 b15aoi013al1n02x5 _25893_ (.a(_17076_),
    .b(_17081_),
    .c(net604),
    .d(net616),
    .o1(_17083_));
 b15oai012as1n04x5 _25894_ (.a(_17079_),
    .b(_17083_),
    .c(net620),
    .o1(_17084_));
 b15nandp2aq1n16x5 _25895_ (.a(_16577_),
    .b(_16475_),
    .o1(_17085_));
 b15nonb03ah1n08x5 _25896_ (.a(net614),
    .b(net613),
    .c(net618),
    .out0(_17086_));
 b15norp02ah1n12x5 _25897_ (.a(_16432_),
    .b(_16673_),
    .o1(_17087_));
 b15nandp2aq1n48x5 _25898_ (.a(net619),
    .b(net611),
    .o1(_17088_));
 b15nor004an1n03x5 _25899_ (.a(net604),
    .b(net598),
    .c(_16563_),
    .d(_17088_),
    .o1(_17089_));
 b15oai013al1n06x5 _25900_ (.a(net617),
    .b(_16526_),
    .c(_17087_),
    .d(_17089_),
    .o1(_17090_));
 b15nona23aq1n32x5 _25901_ (.a(net606),
    .b(net600),
    .c(net596),
    .d(net602),
    .out0(_17091_));
 b15norp02ar1n02x5 _25902_ (.a(net611),
    .b(_17091_),
    .o1(_17092_));
 b15orn002al1n16x5 _25903_ (.a(net606),
    .b(net599),
    .o(_17093_));
 b15oai012ar1n04x5 _25904_ (.a(_17093_),
    .b(_16563_),
    .c(_16609_),
    .o1(_17094_));
 b15aoi013an1n03x5 _25905_ (.a(_17092_),
    .b(_17094_),
    .c(_16510_),
    .d(net611),
    .o1(_17095_));
 b15aoi022aq1n12x5 _25906_ (.a(_17085_),
    .b(_17086_),
    .c(_17090_),
    .d(_17095_),
    .o1(_17096_));
 b15nand02aq1n04x5 _25907_ (.a(net607),
    .b(_16460_),
    .o1(_17097_));
 b15aoi112ar1n02x5 _25908_ (.a(net620),
    .b(_16667_),
    .c(_16508_),
    .d(net604),
    .o1(_17098_));
 b15inv000as1n28x5 _25909_ (.a(\us13.a[5] ),
    .o1(_17099_));
 b15bfn000as1n02x5 input66 (.a(key[43]),
    .o(net66));
 b15bfn000as1n02x5 input65 (.a(key[42]),
    .o(net65));
 b15nand02ar1n02x5 _25912_ (.a(_16435_),
    .b(_16473_),
    .o1(_17102_));
 b15oabi12ar1n02x5 _25913_ (.a(net620),
    .b(net616),
    .c(\us13.a[7] ),
    .out0(_17103_));
 b15aoi022ar1n02x5 _25914_ (.a(\us13.a[7] ),
    .b(net620),
    .c(_17103_),
    .d(net607),
    .o1(_17104_));
 b15oaoi13ar1n02x5 _25915_ (.a(_17099_),
    .b(_17102_),
    .c(_17104_),
    .d(net601),
    .o1(_17105_));
 b15oab012aq1n03x5 _25916_ (.a(_17097_),
    .b(_17098_),
    .c(_17105_),
    .out0(_17106_));
 b15oai013ar1n12x5 _25917_ (.a(net610),
    .b(_17084_),
    .c(_17096_),
    .d(_17106_),
    .o1(_17107_));
 b15bfn001ah1n06x5 input64 (.a(key[41]),
    .o(net64));
 b15bfn000ar1n02x5 input63 (.a(key[40]),
    .o(net63));
 b15norp02aq1n04x5 _25920_ (.a(net600),
    .b(net618),
    .o1(_17110_));
 b15nandp3an1n03x5 _25921_ (.a(net611),
    .b(_16510_),
    .c(_17110_),
    .o1(_17111_));
 b15nor002as1n06x5 _25922_ (.a(net603),
    .b(net600),
    .o1(_17112_));
 b15nanb02as1n16x5 _25923_ (.a(net606),
    .b(net596),
    .out0(_17113_));
 b15nand04an1n06x5 _25924_ (.a(_17112_),
    .b(_16586_),
    .c(_16613_),
    .d(_17113_),
    .o1(_17114_));
 b15oai112an1n12x5 _25925_ (.a(_17111_),
    .b(_17114_),
    .c(_16609_),
    .d(_17085_),
    .o1(_17115_));
 b15nona23as1n32x5 _25926_ (.a(net604),
    .b(net601),
    .c(net597),
    .d(net607),
    .out0(_17116_));
 b15norp02an1n02x5 _25927_ (.a(net612),
    .b(_17116_),
    .o1(_17117_));
 b15nand02ar1n02x5 _25928_ (.a(net616),
    .b(_17117_),
    .o1(_17118_));
 b15nand03as1n12x5 _25929_ (.a(net612),
    .b(_16473_),
    .c(_16579_),
    .o1(_17119_));
 b15oaoi13an1n03x5 _25930_ (.a(net620),
    .b(_17118_),
    .c(_17119_),
    .d(net616),
    .o1(_17120_));
 b15nor002aq1n02x5 _25931_ (.a(_16492_),
    .b(_16680_),
    .o1(_17121_));
 b15oai013aq1n06x5 _25932_ (.a(_16466_),
    .b(_17115_),
    .c(_17120_),
    .d(_17121_),
    .o1(_17122_));
 b15bfm201ah1n02x5 input62 (.a(key[3]),
    .o(net62));
 b15nand02ar1n02x5 _25934_ (.a(net620),
    .b(_16646_),
    .o1(_17124_));
 b15nand02ah1n32x5 _25935_ (.a(_16481_),
    .b(_16520_),
    .o1(_17125_));
 b15bfn000as1n02x5 input61 (.a(key[39]),
    .o(net61));
 b15oaoi13as1n03x5 _25937_ (.a(_16524_),
    .b(_17124_),
    .c(_17125_),
    .d(net620),
    .o1(_17127_));
 b15nano23as1n24x5 _25938_ (.a(net602),
    .b(net600),
    .c(net597),
    .d(net607),
    .out0(_17128_));
 b15aoai13as1n08x5 _25939_ (.a(net616),
    .b(_17127_),
    .c(_17128_),
    .d(_16460_),
    .o1(_17129_));
 b15bfn000ah1n02x5 input60 (.a(key[38]),
    .o(net60));
 b15nand03as1n12x5 _25941_ (.a(net608),
    .b(_16473_),
    .c(_16579_),
    .o1(_17131_));
 b15oai022ah1n02x5 _25942_ (.a(_16498_),
    .b(_16643_),
    .c(_17131_),
    .d(_16439_),
    .o1(_17132_));
 b15aoai13ar1n04x5 _25943_ (.a(net620),
    .b(net616),
    .c(_16466_),
    .d(_16528_),
    .o1(_17133_));
 b15nandp3ar1n08x5 _25944_ (.a(_16586_),
    .b(_17113_),
    .c(_16684_),
    .o1(_17134_));
 b15oaoi13an1n04x5 _25945_ (.a(_17099_),
    .b(_17134_),
    .c(_16500_),
    .d(_16438_),
    .o1(_17135_));
 b15aoai13an1n06x5 _25946_ (.a(net612),
    .b(_17132_),
    .c(_17133_),
    .d(_17135_),
    .o1(_17136_));
 b15bfn000as1n02x5 input59 (.a(key[37]),
    .o(net59));
 b15oaoi13aq1n03x5 _25948_ (.a(_17088_),
    .b(_16608_),
    .c(net610),
    .d(_17091_),
    .o1(_17138_));
 b15nand02aq1n24x5 _25949_ (.a(net597),
    .b(net608),
    .o1(_17139_));
 b15oai012ah1n04x5 _25950_ (.a(_17139_),
    .b(_16461_),
    .c(net610),
    .o1(_17140_));
 b15bfn001ah1n08x5 input58 (.a(key[36]),
    .o(net58));
 b15bfn000aq1n02x5 input57 (.a(key[35]),
    .o(net57));
 b15aoi013ah1n06x5 _25953_ (.a(_17138_),
    .b(_17140_),
    .c(_16517_),
    .d(_16597_),
    .o1(_17143_));
 b15bfn001as1n12x5 input56 (.a(key[34]),
    .o(net56));
 b15oai112as1n16x5 _25955_ (.a(_17129_),
    .b(_17136_),
    .c(_17143_),
    .d(net616),
    .o1(_17145_));
 b15nano23as1n16x5 _25956_ (.a(net596),
    .b(net600),
    .c(net602),
    .d(net607),
    .out0(_17146_));
 b15nand04ar1n08x5 _25957_ (.a(_16592_),
    .b(_16453_),
    .c(_16604_),
    .d(_17146_),
    .o1(_17147_));
 b15nor004an1n04x5 _25958_ (.a(net606),
    .b(net596),
    .c(net600),
    .d(net609),
    .o1(_17148_));
 b15aoi022al1n08x5 _25959_ (.a(_16591_),
    .b(_16629_),
    .c(_17148_),
    .d(_16504_),
    .o1(_17149_));
 b15nand02aq1n04x5 _25960_ (.a(_16558_),
    .b(_16577_),
    .o1(_17150_));
 b15norp02an1n03x5 _25961_ (.a(net606),
    .b(net609),
    .o1(_17151_));
 b15and002an1n08x5 _25962_ (.a(net615),
    .b(net609),
    .o(_17152_));
 b15aoi022ah1n04x5 _25963_ (.a(net602),
    .b(_17151_),
    .c(_16517_),
    .d(_17152_),
    .o1(_17153_));
 b15oai112an1n16x5 _25964_ (.a(_17147_),
    .b(_17149_),
    .c(_17150_),
    .d(_17153_),
    .o1(_17154_));
 b15oai112as1n04x5 _25965_ (.a(_16475_),
    .b(_16605_),
    .c(_16613_),
    .d(_17086_),
    .o1(_17155_));
 b15nanb02ar1n06x5 _25966_ (.a(_17088_),
    .b(_16597_),
    .out0(_17156_));
 b15nonb02as1n03x5 _25967_ (.a(net596),
    .b(net606),
    .out0(_17157_));
 b15mdn022ar1n08x5 _25968_ (.a(_16656_),
    .b(_17157_),
    .o1(_17158_),
    .sa(net603));
 b15oaoi13as1n08x5 _25969_ (.a(net609),
    .b(_17155_),
    .c(_17156_),
    .d(_17158_),
    .o1(_17159_));
 b15bfn001al1n08x5 input55 (.a(key[33]),
    .o(net55));
 b15nano22al1n12x5 _25971_ (.a(net599),
    .b(net609),
    .c(net613),
    .out0(_17161_));
 b15aoi022ar1n12x5 _25972_ (.a(_16481_),
    .b(_16657_),
    .c(_17161_),
    .d(_16517_),
    .o1(_17162_));
 b15nor003aq1n06x5 _25973_ (.a(net596),
    .b(net614),
    .c(_17162_),
    .o1(_17163_));
 b15nandp3ar1n08x5 _25974_ (.a(net609),
    .b(_16520_),
    .c(_16517_),
    .o1(_17164_));
 b15nandp3ar1n16x5 _25975_ (.a(net618),
    .b(net614),
    .c(net613),
    .o1(_17165_));
 b15nor002aq1n03x5 _25976_ (.a(_16504_),
    .b(_16613_),
    .o1(_17166_));
 b15oaoi13aq1n04x5 _25977_ (.a(_17164_),
    .b(_17165_),
    .c(_17166_),
    .d(net618),
    .o1(_17167_));
 b15nor004as1n12x5 _25978_ (.a(_17154_),
    .b(_17159_),
    .c(_17163_),
    .d(_17167_),
    .o1(_17168_));
 b15oai012ah1n02x5 _25979_ (.a(net619),
    .b(_17128_),
    .c(_16650_),
    .o1(_17169_));
 b15bfn000ar1n02x5 input54 (.a(key[32]),
    .o(net54));
 b15mdn022an1n06x5 _25981_ (.a(_16646_),
    .b(_16650_),
    .o1(_17171_),
    .sa(_16508_));
 b15oaoi13ah1n08x5 _25982_ (.a(_16479_),
    .b(_17169_),
    .c(_17171_),
    .d(net619),
    .o1(_17172_));
 b15nandp3al1n08x5 _25983_ (.a(net608),
    .b(_16475_),
    .c(_16605_),
    .o1(_17173_));
 b15bfn000ah1n06x5 input53 (.a(key[31]),
    .o(net53));
 b15nanb02as1n24x5 _25985_ (.a(net615),
    .b(net611),
    .out0(_17175_));
 b15nandp3ar1n12x5 _25986_ (.o1(_17176_),
    .a(net619),
    .b(_16652_),
    .c(_17175_));
 b15nand02ah1n03x5 _25987_ (.a(_16558_),
    .b(_16504_),
    .o1(_17177_));
 b15aoi012al1n06x5 _25988_ (.a(_17173_),
    .b(_17176_),
    .c(_17177_),
    .o1(_17178_));
 b15nonb02an1n04x5 _25989_ (.a(net600),
    .b(net603),
    .out0(_17179_));
 b15aoi012as1n02x5 _25990_ (.a(_17179_),
    .b(_17110_),
    .c(net603),
    .o1(_17180_));
 b15and002as1n08x5 _25991_ (.a(net606),
    .b(net596),
    .o(_17181_));
 b15nandp3ah1n02x5 _25992_ (.a(_16466_),
    .b(_17181_),
    .c(_17175_),
    .o1(_17182_));
 b15nandp2as1n16x5 _25993_ (.a(_16579_),
    .b(_16605_),
    .o1(_17183_));
 b15aoi112ah1n04x5 _25994_ (.a(_17180_),
    .b(_17182_),
    .c(_16682_),
    .d(_17183_),
    .o1(_17184_));
 b15nor004aq1n12x5 _25995_ (.a(_16645_),
    .b(_17172_),
    .c(_17178_),
    .d(_17184_),
    .o1(_17185_));
 b15bfn000an1n02x5 input52 (.a(key[30]),
    .o(net52));
 b15bfn001ah1n06x5 input51 (.a(key[2]),
    .o(net51));
 b15aoi022aq1n08x5 _25998_ (.a(_16473_),
    .b(_16475_),
    .c(_16571_),
    .d(net610),
    .o1(_17188_));
 b15aoi112an1n02x5 _25999_ (.a(net611),
    .b(_16544_),
    .c(_16576_),
    .d(_16456_),
    .o1(_17189_));
 b15nonb02ar1n12x5 _26000_ (.a(net608),
    .b(net616),
    .out0(_17190_));
 b15aoi122ah1n08x5 _26001_ (.a(net620),
    .b(net616),
    .c(_16576_),
    .d(_17125_),
    .e(_17190_),
    .o1(_17191_));
 b15nand04ar1n02x5 _26002_ (.a(net615),
    .b(net610),
    .c(_16481_),
    .d(_16520_),
    .o1(_17192_));
 b15oaoi13aq1n03x5 _26003_ (.a(_16558_),
    .b(_17192_),
    .c(_16576_),
    .d(net615),
    .o1(_17193_));
 b15oaoi13an1n04x5 _26004_ (.a(_17189_),
    .b(net611),
    .c(_17191_),
    .d(_17193_),
    .o1(_17194_));
 b15oai112as1n16x5 _26005_ (.a(_17168_),
    .b(_17185_),
    .c(_17188_),
    .d(_17194_),
    .o1(_17195_));
 b15nano23as1n24x5 _26006_ (.a(_17107_),
    .b(_17122_),
    .c(_17145_),
    .d(_17195_),
    .out0(_17196_));
 b15nand03an1n03x5 _26007_ (.a(net719),
    .b(_16230_),
    .c(_17033_),
    .o1(_17197_));
 b15oai022ar1n02x5 _26008_ (.a(_16986_),
    .b(_16316_),
    .c(_16993_),
    .d(net737),
    .o1(_17198_));
 b15aoi022ah1n04x5 _26009_ (.a(_16191_),
    .b(_17033_),
    .c(_17198_),
    .d(_16194_),
    .o1(_17199_));
 b15oaoi13ar1n08x5 _26010_ (.a(_17055_),
    .b(_17197_),
    .c(_17199_),
    .d(_16278_),
    .o1(_17200_));
 b15oai022ar1n02x5 _26011_ (.a(_16995_),
    .b(_16383_),
    .c(_16414_),
    .d(_16993_),
    .o1(_17201_));
 b15aoi112as1n02x5 _26012_ (.a(\us02.a[1] ),
    .b(_17201_),
    .c(_16980_),
    .d(net743),
    .o1(_17202_));
 b15nanb02ar1n12x5 _26013_ (.a(net717),
    .b(net722),
    .out0(_17203_));
 b15aoi012as1n06x5 _26014_ (.a(_17203_),
    .b(_16928_),
    .c(_16929_),
    .o1(_17204_));
 b15aoi022ah1n06x5 _26015_ (.a(_16977_),
    .b(_17000_),
    .c(_17204_),
    .d(_17028_),
    .o1(_17205_));
 b15nor003ar1n12x5 _26016_ (.a(_16235_),
    .b(_16237_),
    .c(_16381_),
    .o1(_17206_));
 b15aoi013al1n02x5 _26017_ (.a(_17206_),
    .b(_16311_),
    .c(_16999_),
    .d(net731),
    .o1(_17207_));
 b15aoi013as1n02x5 _26018_ (.a(_17202_),
    .b(_17205_),
    .c(_17207_),
    .d(net737),
    .o1(_17208_));
 b15nandp3ar1n02x5 _26019_ (.a(net735),
    .b(_16213_),
    .c(_16936_),
    .o1(_17209_));
 b15nandp2ar1n03x5 _26020_ (.a(\us02.a[1] ),
    .b(_17009_),
    .o1(_17210_));
 b15aob012ar1n02x5 _26021_ (.a(_16321_),
    .b(_17210_),
    .c(_16947_),
    .out0(_17211_));
 b15aoi012aq1n02x5 _26022_ (.a(_16226_),
    .b(_17209_),
    .c(_17211_),
    .o1(_17212_));
 b15nor003ah1n04x5 _26023_ (.a(_17200_),
    .b(_17208_),
    .c(_17212_),
    .o1(_17213_));
 b15aoi022ar1n02x5 _26024_ (.a(net740),
    .b(_16273_),
    .c(_16970_),
    .d(_16932_),
    .o1(_17214_));
 b15oai012aq1n03x5 _26025_ (.a(net722),
    .b(_16993_),
    .c(_17214_),
    .o1(_17215_));
 b15nand03ar1n02x5 _26026_ (.a(net726),
    .b(_16328_),
    .c(_17028_),
    .o1(_17216_));
 b15oai012as1n04x5 _26027_ (.a(_17216_),
    .b(_16951_),
    .c(_16226_),
    .o1(_17217_));
 b15aoai13as1n08x5 _26028_ (.a(_17215_),
    .b(net722),
    .c(_16970_),
    .d(_17217_),
    .o1(_17218_));
 b15oai012ar1n02x5 _26029_ (.a(_16361_),
    .b(_16365_),
    .c(_16342_),
    .o1(_17219_));
 b15oa0022al1n03x5 _26030_ (.a(_16995_),
    .b(_16260_),
    .c(_16420_),
    .d(_17219_),
    .o(_17220_));
 b15norp02al1n04x5 _26031_ (.a(net735),
    .b(_16402_),
    .o1(_17221_));
 b15aoai13al1n04x5 _26032_ (.a(_16401_),
    .b(_17221_),
    .c(net735),
    .d(_16321_),
    .o1(_17222_));
 b15norp02ar1n12x5 _26033_ (.a(_16310_),
    .b(_16979_),
    .o1(_17223_));
 b15nonb02as1n16x5 _26034_ (.a(\us02.a[0] ),
    .b(net736),
    .out0(_17224_));
 b15norp02ah1n12x5 _26035_ (.a(_16398_),
    .b(_16314_),
    .o1(_17225_));
 b15aoi022al1n08x5 _26036_ (.a(_16222_),
    .b(_17223_),
    .c(_17224_),
    .d(_17225_),
    .o1(_17226_));
 b15oai112ar1n16x5 _26037_ (.a(_17220_),
    .b(_17222_),
    .c(_16226_),
    .d(_17226_),
    .o1(_17227_));
 b15nandp3ah1n02x5 _26038_ (.a(net729),
    .b(net717),
    .c(net719),
    .o1(_17228_));
 b15oaoi13ah1n08x5 _26039_ (.a(_16313_),
    .b(_17228_),
    .c(net729),
    .d(_16235_),
    .o1(_17229_));
 b15aob012al1n12x5 _26040_ (.a(net740),
    .b(net729),
    .c(net737),
    .out0(_17230_));
 b15nand03as1n08x5 _26041_ (.a(net733),
    .b(_17229_),
    .c(_17230_),
    .o1(_17231_));
 b15oai112an1n02x5 _26042_ (.a(_16283_),
    .b(_17005_),
    .c(_16951_),
    .d(net724),
    .o1(_17232_));
 b15oai112ah1n04x5 _26043_ (.a(_16957_),
    .b(_17232_),
    .c(_16283_),
    .d(_16315_),
    .o1(_17233_));
 b15norp03ar1n02x5 _26044_ (.a(net731),
    .b(_16390_),
    .c(_17045_),
    .o1(_17234_));
 b15aoi013aq1n02x5 _26045_ (.a(_17234_),
    .b(_16936_),
    .c(_16977_),
    .d(net731),
    .o1(_17235_));
 b15oai112an1n06x5 _26046_ (.a(_17231_),
    .b(_17233_),
    .c(_17235_),
    .d(net735),
    .o1(_17236_));
 b15oai022ar1n04x5 _26047_ (.a(_16995_),
    .b(_16383_),
    .c(_16336_),
    .d(_16377_),
    .o1(_17237_));
 b15bfn000as1n06x5 input50 (.a(key[29]),
    .o(net50));
 b15xor002as1n03x5 _26049_ (.a(net733),
    .b(net717),
    .out0(_17239_));
 b15nor004as1n12x5 _26050_ (.a(net729),
    .b(net722),
    .c(_16928_),
    .d(_17239_),
    .o1(_17240_));
 b15oai012al1n06x5 _26051_ (.a(net741),
    .b(_17237_),
    .c(_17240_),
    .o1(_17241_));
 b15oai012ar1n02x5 _26052_ (.a(net731),
    .b(net735),
    .c(_16936_),
    .o1(_17242_));
 b15oaoi13an1n02x5 _26053_ (.a(_17242_),
    .b(_16958_),
    .c(_16329_),
    .d(_16214_),
    .o1(_17243_));
 b15nandp2aq1n02x5 _26054_ (.a(net735),
    .b(_16958_),
    .o1(_17244_));
 b15aoai13an1n06x5 _26055_ (.a(_17243_),
    .b(\us02.a[1] ),
    .c(net741),
    .d(_17244_),
    .o1(_17245_));
 b15nona23as1n12x5 _26056_ (.a(_17227_),
    .b(_17236_),
    .c(_17241_),
    .d(_17245_),
    .out0(_17246_));
 b15nandp2al1n08x5 _26057_ (.a(net730),
    .b(net716),
    .o1(_17247_));
 b15nanb03ar1n02x5 _26058_ (.a(net720),
    .b(net725),
    .c(net740),
    .out0(_17248_));
 b15oaoi13an1n03x5 _26059_ (.a(_17247_),
    .b(_17248_),
    .c(net740),
    .d(_16928_),
    .o1(_17249_));
 b15aoai13aq1n03x5 _26060_ (.a(net722),
    .b(_17249_),
    .c(_16289_),
    .d(_16223_),
    .o1(_17250_));
 b15nonb03as1n06x5 _26061_ (.a(net716),
    .b(net719),
    .c(net725),
    .out0(_17251_));
 b15nand02al1n02x5 _26062_ (.a(_16292_),
    .b(_17251_),
    .o1(_17252_));
 b15aob012ar1n12x5 _26063_ (.a(_16356_),
    .b(_17250_),
    .c(_17252_),
    .out0(_17253_));
 b15aoai13ar1n02x5 _26064_ (.a(_17026_),
    .b(_17031_),
    .c(_16311_),
    .d(_16370_),
    .o1(_17254_));
 b15oab012an1n02x5 _26065_ (.a(_17254_),
    .b(_16403_),
    .c(net738),
    .out0(_17255_));
 b15nandp3an1n02x5 _26066_ (.a(_16193_),
    .b(_16405_),
    .c(_16932_),
    .o1(_17256_));
 b15oai112an1n06x5 _26067_ (.a(net729),
    .b(_17256_),
    .c(_16414_),
    .d(_16405_),
    .o1(_17257_));
 b15nona23ah1n32x5 _26068_ (.a(\us02.a[5] ),
    .b(net728),
    .c(\us02.a[7] ),
    .d(\us02.a[6] ),
    .out0(_17258_));
 b15oaoi13aq1n04x5 _26069_ (.a(_16367_),
    .b(_16958_),
    .c(_17258_),
    .d(_16342_),
    .o1(_17259_));
 b15nand02al1n06x5 _26070_ (.a(net738),
    .b(net725),
    .o1(_17260_));
 b15aoi013ah1n02x5 _26071_ (.a(net730),
    .b(_16214_),
    .c(_16351_),
    .d(_17260_),
    .o1(_17261_));
 b15nano22ar1n03x5 _26072_ (.a(net716),
    .b(net719),
    .c(net723),
    .out0(_17262_));
 b15aoi022ar1n08x5 _26073_ (.a(net723),
    .b(_16223_),
    .c(_16350_),
    .d(_17262_),
    .o1(_17263_));
 b15oai013aq1n08x5 _26074_ (.a(_17261_),
    .b(_17263_),
    .c(net725),
    .d(net740),
    .o1(_17264_));
 b15oai022as1n08x5 _26075_ (.a(_17255_),
    .b(_17257_),
    .c(_17259_),
    .d(_17264_),
    .o1(_17265_));
 b15nandp3ar1n02x5 _26076_ (.a(_16342_),
    .b(net733),
    .c(_17229_),
    .o1(_17266_));
 b15oai012ah1n02x5 _26077_ (.a(_17224_),
    .b(_17204_),
    .c(_16321_),
    .o1(_17267_));
 b15aob012al1n06x5 _26078_ (.a(_16226_),
    .b(_17266_),
    .c(_17267_),
    .out0(_17268_));
 b15norp02ah1n02x5 _26079_ (.a(net735),
    .b(net727),
    .o1(_17269_));
 b15and003aq1n04x5 _26080_ (.a(net731),
    .b(net724),
    .c(net718),
    .o(_17270_));
 b15nor004as1n08x5 _26081_ (.a(net741),
    .b(net731),
    .c(net724),
    .d(net718),
    .o1(_17271_));
 b15oai112an1n12x5 _26082_ (.a(_16379_),
    .b(_17269_),
    .c(_17270_),
    .d(_17271_),
    .o1(_17272_));
 b15aoi022an1n04x5 _26083_ (.a(_16258_),
    .b(_17028_),
    .c(_17041_),
    .d(_16301_),
    .o1(_17273_));
 b15oai013an1n08x5 _26084_ (.a(_17272_),
    .b(_17273_),
    .c(_16379_),
    .d(_17055_),
    .o1(_17274_));
 b15norp02aq1n04x5 _26085_ (.a(net722),
    .b(net717),
    .o1(_17275_));
 b15aoi022ar1n08x5 _26086_ (.a(_16283_),
    .b(_16927_),
    .c(_17275_),
    .d(_16342_),
    .o1(_17276_));
 b15aoi022ar1n08x5 _26087_ (.a(net737),
    .b(_16927_),
    .c(_17275_),
    .d(net733),
    .o1(_17277_));
 b15oai022ar1n12x5 _26088_ (.a(net733),
    .b(_17276_),
    .c(_17277_),
    .d(net740),
    .o1(_17278_));
 b15aoai13as1n06x5 _26089_ (.a(_16305_),
    .b(_17274_),
    .c(_17278_),
    .d(_16354_),
    .o1(_17279_));
 b15nand04as1n16x5 _26090_ (.a(_17253_),
    .b(_17265_),
    .c(_17268_),
    .d(_17279_),
    .o1(_17280_));
 b15nano23as1n24x5 _26091_ (.a(_17213_),
    .b(_17218_),
    .c(_17246_),
    .d(_17280_),
    .out0(_17281_));
 b15xor002as1n08x5 _26092_ (.a(_17196_),
    .b(_17281_),
    .out0(_17282_));
 b15xor002ar1n04x5 _26093_ (.a(_17069_),
    .b(_17282_),
    .out0(_17283_));
 b15bfn001ah1n06x5 input49 (.a(key[28]),
    .o(net49));
 b15nanb02ah1n24x5 _26095_ (.a(net750),
    .b(net753),
    .out0(_17285_));
 b15aoi013ar1n02x5 _26096_ (.a(\us31.a[2] ),
    .b(_16708_),
    .c(_16849_),
    .d(_17285_),
    .o1(_17286_));
 b15norp02as1n12x5 _26097_ (.a(net762),
    .b(\us31.a[2] ),
    .o1(_17287_));
 b15and002as1n02x5 _26098_ (.a(net767),
    .b(net750),
    .o(_17288_));
 b15aoi012ar1n02x5 _26099_ (.a(_17287_),
    .b(_17288_),
    .c(_16827_),
    .o1(_17289_));
 b15bfn000ah1n02x5 input48 (.a(key[27]),
    .o(net48));
 b15bfn000ah1n04x5 input47 (.a(key[26]),
    .o(net47));
 b15and003as1n04x5 _26102_ (.a(net750),
    .b(\us31.a[4] ),
    .c(\us31.a[7] ),
    .o(_17292_));
 b15bfn000ar1n02x5 input46 (.a(key[25]),
    .o(net46));
 b15nor003ah1n02x5 _26104_ (.a(net750),
    .b(\us31.a[4] ),
    .c(\us31.a[7] ),
    .o1(_17294_));
 b15oai112an1n06x5 _26105_ (.a(net748),
    .b(_16894_),
    .c(_17292_),
    .d(_17294_),
    .o1(_17295_));
 b15aoi012ar1n02x5 _26106_ (.a(_17286_),
    .b(_17289_),
    .c(_17295_),
    .o1(_17296_));
 b15nand02al1n24x5 _26107_ (.a(net753),
    .b(net744),
    .o1(_17297_));
 b15and002aq1n08x5 _26108_ (.a(net750),
    .b(net748),
    .o(_17298_));
 b15norp02aq1n04x5 _26109_ (.a(net750),
    .b(net748),
    .o1(_17299_));
 b15aoi012ar1n02x5 _26110_ (.a(_17298_),
    .b(_16852_),
    .c(_17299_),
    .o1(_17300_));
 b15nor004an1n02x5 _26111_ (.a(\us31.a[2] ),
    .b(_17297_),
    .c(_16894_),
    .d(_17300_),
    .o1(_17301_));
 b15oab012ah1n06x5 _26112_ (.a(net755),
    .b(_17296_),
    .c(_17301_),
    .out0(_17302_));
 b15nano23aq1n24x5 _26113_ (.a(net749),
    .b(net752),
    .c(net745),
    .d(net746),
    .out0(_17303_));
 b15nand03ah1n02x5 _26114_ (.a(net761),
    .b(_17303_),
    .c(_16798_),
    .o1(_17304_));
 b15bfn000aq1n02x5 input45 (.a(key[24]),
    .o(net45));
 b15bfn000aq1n02x5 input44 (.a(key[23]),
    .o(net44));
 b15nandp3ar1n03x5 _26117_ (.a(_16798_),
    .b(_16907_),
    .c(_16758_),
    .o1(_17307_));
 b15bfn001al1n08x5 input43 (.a(key[22]),
    .o(net43));
 b15nonb02ar1n12x5 _26119_ (.a(net767),
    .b(net753),
    .out0(_17309_));
 b15bfn000as1n02x5 input42 (.a(key[21]),
    .o(net42));
 b15nand04aq1n03x5 _26121_ (.a(net749),
    .b(_16780_),
    .c(_16830_),
    .d(_16861_),
    .o1(_17311_));
 b15oai112as1n06x5 _26122_ (.a(_17304_),
    .b(_17307_),
    .c(_17309_),
    .d(_17311_),
    .o1(_17312_));
 b15nand02ah1n06x5 _26123_ (.a(net765),
    .b(_16798_),
    .o1(_17313_));
 b15nand02as1n32x5 _26124_ (.a(_16725_),
    .b(_16726_),
    .o1(_17314_));
 b15oai022aq1n04x5 _26125_ (.a(_16748_),
    .b(_16760_),
    .c(_17313_),
    .d(_17314_),
    .o1(_17315_));
 b15aoi012aq1n08x5 _26126_ (.a(_17312_),
    .b(_17315_),
    .c(net761),
    .o1(_17316_));
 b15nanb02aq1n12x5 _26127_ (.a(net763),
    .b(net759),
    .out0(_17317_));
 b15bfn001ah1n06x5 input41 (.a(key[20]),
    .o(net41));
 b15nandp3al1n16x5 _26129_ (.a(_16785_),
    .b(_16726_),
    .c(_16815_),
    .o1(_17319_));
 b15nand02an1n08x5 _26130_ (.a(net755),
    .b(_16758_),
    .o1(_17320_));
 b15aoi012ar1n02x5 _26131_ (.a(_17317_),
    .b(_17319_),
    .c(_17320_),
    .o1(_17321_));
 b15bfn000ah1n06x5 input40 (.a(key[1]),
    .o(net40));
 b15oai012an1n02x5 _26133_ (.a(_17320_),
    .b(_16711_),
    .c(net755),
    .o1(_17323_));
 b15aoi012al1n04x5 _26134_ (.a(_17321_),
    .b(_17323_),
    .c(_16860_),
    .o1(_17324_));
 b15nand04al1n02x5 _26135_ (.a(net749),
    .b(_16798_),
    .c(_16896_),
    .d(_16855_),
    .o1(_17325_));
 b15nandp2ar1n05x5 _26136_ (.a(net766),
    .b(_16713_),
    .o1(_17326_));
 b15oai012aq1n04x5 _26137_ (.a(_17325_),
    .b(_17326_),
    .c(_16832_),
    .o1(_17327_));
 b15nonb02as1n08x5 _26138_ (.a(\us31.a[7] ),
    .b(net753),
    .out0(_17328_));
 b15aoi013as1n02x5 _26139_ (.a(_17327_),
    .b(_17328_),
    .c(_16873_),
    .d(_16783_),
    .o1(_17329_));
 b15nandp3ar1n02x5 _26140_ (.a(_16896_),
    .b(_16804_),
    .c(_16834_),
    .o1(_17330_));
 b15nand04ar1n03x5 _26141_ (.a(net763),
    .b(_16798_),
    .c(_16785_),
    .d(_16726_),
    .o1(_17331_));
 b15aoi012al1n02x5 _26142_ (.a(net766),
    .b(_17330_),
    .c(_17331_),
    .o1(_17332_));
 b15norp02ar1n02x5 _26143_ (.a(net764),
    .b(net755),
    .o1(_17333_));
 b15oai112an1n04x5 _26144_ (.a(_16725_),
    .b(_16726_),
    .c(_16783_),
    .d(_17333_),
    .o1(_17334_));
 b15norp02ar1n24x5 _26145_ (.a(net766),
    .b(net759),
    .o1(_17335_));
 b15oaoi13al1n04x5 _26146_ (.a(net763),
    .b(_17334_),
    .c(_16790_),
    .d(_17335_),
    .o1(_17336_));
 b15nor004as1n12x5 _26147_ (.a(net751),
    .b(net753),
    .c(net744),
    .d(net748),
    .o1(_17337_));
 b15nand03ah1n06x5 _26148_ (.a(_16798_),
    .b(_16894_),
    .c(_17337_),
    .o1(_17338_));
 b15orn002aq1n12x5 _26149_ (.a(net765),
    .b(net757),
    .o(_17339_));
 b15bfn000ar1n02x5 input39 (.a(key[19]),
    .o(net39));
 b15nandp3ar1n03x5 _26151_ (.a(net762),
    .b(net765),
    .c(net758),
    .o1(_17341_));
 b15nand04aq1n08x5 _26152_ (.a(_17339_),
    .b(_16768_),
    .c(_16782_),
    .d(_17341_),
    .o1(_17342_));
 b15aoi022as1n06x5 _26153_ (.a(net762),
    .b(_16772_),
    .c(_16836_),
    .d(net758),
    .o1(_17343_));
 b15nand03ar1n08x5 _26154_ (.a(\us31.a[4] ),
    .b(_16708_),
    .c(_16873_),
    .o1(_17344_));
 b15oai112as1n16x5 _26155_ (.a(_17338_),
    .b(_17342_),
    .c(_17343_),
    .d(_17344_),
    .o1(_17345_));
 b15nand03ar1n03x5 _26156_ (.a(net759),
    .b(_17303_),
    .c(_16834_),
    .o1(_17346_));
 b15aoai13ar1n04x5 _26157_ (.a(_17346_),
    .b(_16748_),
    .c(_16775_),
    .d(_16835_),
    .o1(_17347_));
 b15nor004ar1n06x5 _26158_ (.a(_17332_),
    .b(_17336_),
    .c(_17345_),
    .d(_17347_),
    .o1(_17348_));
 b15nand04as1n08x5 _26159_ (.a(_17316_),
    .b(_17324_),
    .c(_17329_),
    .d(_17348_),
    .o1(_17349_));
 b15bfn000ar1n02x5 input38 (.a(key[18]),
    .o(net38));
 b15nand04ah1n06x5 _26161_ (.a(_16741_),
    .b(_16774_),
    .c(_16830_),
    .d(_16831_),
    .o1(_17351_));
 b15nand03ah1n03x5 _26162_ (.a(net761),
    .b(_16830_),
    .c(_16831_),
    .o1(_17352_));
 b15aob012as1n03x5 _26163_ (.a(_16844_),
    .b(_17352_),
    .c(_16888_),
    .out0(_17353_));
 b15nor002ah1n06x5 _26164_ (.a(net758),
    .b(_16711_),
    .o1(_17354_));
 b15nand02ar1n16x5 _26165_ (.a(net758),
    .b(_17303_),
    .o1(_17355_));
 b15oai012aq1n02x5 _26166_ (.a(_16802_),
    .b(_17355_),
    .c(net754),
    .o1(_17356_));
 b15aoi022ah1n06x5 _26167_ (.a(_17354_),
    .b(_16834_),
    .c(_17356_),
    .d(net761),
    .o1(_17357_));
 b15aoi013aq1n08x5 _26168_ (.a(net766),
    .b(_17351_),
    .c(_17353_),
    .d(_17357_),
    .o1(_17358_));
 b15nonb02an1n08x5 _26169_ (.a(net750),
    .b(net759),
    .out0(_17359_));
 b15nand04as1n04x5 _26170_ (.a(net748),
    .b(_17328_),
    .c(_16855_),
    .d(_17359_),
    .o1(_17360_));
 b15nand03an1n06x5 _26171_ (.a(\us31.a[4] ),
    .b(net748),
    .c(_17317_),
    .o1(_17361_));
 b15and002ar1n02x5 _26172_ (.a(net751),
    .b(\us31.a[7] ),
    .o(_17362_));
 b15nor002an1n03x5 _26173_ (.a(net750),
    .b(\us31.a[7] ),
    .o1(_17363_));
 b15aoi022ah1n04x5 _26174_ (.a(_16898_),
    .b(_17362_),
    .c(_17363_),
    .d(\us31.a[0] ),
    .o1(_17364_));
 b15oai122as1n12x5 _26175_ (.a(_17360_),
    .b(_17361_),
    .c(_17364_),
    .d(_16711_),
    .e(_16898_),
    .o1(_17365_));
 b15aoai13ah1n02x5 _26176_ (.a(net763),
    .b(_16725_),
    .c(_16785_),
    .d(net766),
    .o1(_17366_));
 b15orn002aq1n24x5 _26177_ (.a(net760),
    .b(net767),
    .o(_17367_));
 b15oai122ah1n08x5 _26178_ (.a(_17366_),
    .b(_17367_),
    .c(_17285_),
    .d(_16693_),
    .e(_16849_),
    .o1(_17368_));
 b15norp03ah1n12x5 _26179_ (.a(\us31.a[2] ),
    .b(net744),
    .c(net748),
    .o1(_17369_));
 b15aoai13ah1n06x5 _26180_ (.a(net755),
    .b(_17365_),
    .c(_17368_),
    .d(_17369_),
    .o1(_17370_));
 b15ornc04as1n24x5 _26181_ (.a(net749),
    .b(net752),
    .c(net745),
    .d(net746),
    .o(_17371_));
 b15bfn000ah1n03x5 input37 (.a(key[17]),
    .o(net37));
 b15nand02ah1n32x5 _26183_ (.a(_16708_),
    .b(_16785_),
    .o1(_17373_));
 b15oai012an1n02x5 _26184_ (.a(_17371_),
    .b(_17373_),
    .c(net755),
    .o1(_17374_));
 b15and003an1n08x5 _26185_ (.a(net766),
    .b(net754),
    .c(net758),
    .o(_17375_));
 b15aoai13as1n02x5 _26186_ (.a(net763),
    .b(_17375_),
    .c(_17371_),
    .d(_17335_),
    .o1(_17376_));
 b15nand02ar1n02x5 _26187_ (.a(_16798_),
    .b(_16905_),
    .o1(_17377_));
 b15aoi022an1n02x5 _26188_ (.a(net759),
    .b(_17371_),
    .c(_17377_),
    .d(_17326_),
    .o1(_17378_));
 b15oai112ah1n06x5 _26189_ (.a(_17374_),
    .b(_17376_),
    .c(_17378_),
    .d(net763),
    .o1(_17379_));
 b15nandp3ar1n08x5 _26190_ (.a(_16830_),
    .b(_16831_),
    .c(_16894_),
    .o1(_17380_));
 b15oai112an1n04x5 _26191_ (.a(_16741_),
    .b(_17380_),
    .c(_16748_),
    .d(_16774_),
    .o1(_17381_));
 b15nandp2ar1n12x5 _26192_ (.a(net761),
    .b(net757),
    .o1(_17382_));
 b15nor002ah1n06x5 _26193_ (.a(_16867_),
    .b(_17382_),
    .o1(_17383_));
 b15bfn000ar1n02x5 input36 (.a(key[16]),
    .o(net36));
 b15aoi012al1n02x5 _26195_ (.a(_16811_),
    .b(_16855_),
    .c(net758),
    .o1(_17385_));
 b15oai013aq1n06x5 _26196_ (.a(_17381_),
    .b(_17383_),
    .c(_17385_),
    .d(_16741_),
    .o1(_17386_));
 b15oai012ar1n02x5 _26197_ (.a(_16741_),
    .b(_16725_),
    .c(_16785_),
    .o1(_17387_));
 b15oai012ar1n03x5 _26198_ (.a(_17387_),
    .b(_16849_),
    .c(_16774_),
    .o1(_17388_));
 b15orn002al1n16x5 _26199_ (.a(net744),
    .b(net748),
    .o(_17389_));
 b15orn002as1n08x5 _26200_ (.a(net765),
    .b(net754),
    .o(_17390_));
 b15aoi012al1n02x5 _26201_ (.a(net761),
    .b(net758),
    .c(_17390_),
    .o1(_17391_));
 b15aoi012aq1n06x5 _26202_ (.a(_17389_),
    .b(_16919_),
    .c(_17391_),
    .o1(_17392_));
 b15oaoi13an1n02x5 _26203_ (.a(_16834_),
    .b(_16813_),
    .c(_16786_),
    .d(net759),
    .o1(_17393_));
 b15oai112an1n06x5 _26204_ (.a(_17388_),
    .b(_17392_),
    .c(_17393_),
    .d(_16693_),
    .o1(_17394_));
 b15nand04as1n08x5 _26205_ (.a(_17370_),
    .b(_17379_),
    .c(_17386_),
    .d(_17394_),
    .o1(_17395_));
 b15nor004as1n12x5 _26206_ (.a(_17302_),
    .b(_17349_),
    .c(_17358_),
    .d(_17395_),
    .o1(_17396_));
 b15bfn001aq1n06x5 input35 (.a(key[15]),
    .o(net35));
 b15nor002ah1n03x5 _26208_ (.a(net870),
    .b(net863),
    .o1(_17398_));
 b15nand04ah1n08x5 _26209_ (.a(net865),
    .b(_15959_),
    .c(_17398_),
    .d(_16160_),
    .o1(_17399_));
 b15nandp2as1n05x5 _26210_ (.a(net883),
    .b(_15970_),
    .o1(_17400_));
 b15nand02as1n24x5 _26211_ (.a(_15952_),
    .b(_16008_),
    .o1(_17401_));
 b15oai112ah1n12x5 _26212_ (.a(net879),
    .b(_17399_),
    .c(_17400_),
    .d(_17401_),
    .o1(_17402_));
 b15bfn000al1n02x5 input34 (.a(key[14]),
    .o(net34));
 b15aoi122ar1n02x5 _26214_ (.a(net875),
    .b(net874),
    .c(_16058_),
    .d(_16047_),
    .e(net882),
    .o1(_17404_));
 b15nand02ar1n16x5 _26215_ (.a(net874),
    .b(_16047_),
    .o1(_17405_));
 b15aoi012ar1n02x5 _26216_ (.a(_17404_),
    .b(_17405_),
    .c(net875),
    .o1(_17406_));
 b15nand02ar1n16x5 _26217_ (.a(_16096_),
    .b(_15943_),
    .o1(_17407_));
 b15oai022ar1n02x5 _26218_ (.a(_17407_),
    .b(_16134_),
    .c(_16137_),
    .d(_16135_),
    .o1(_17408_));
 b15oa0022an1n04x5 _26219_ (.a(_17402_),
    .b(_17406_),
    .c(_17408_),
    .d(net879),
    .o(_17409_));
 b15nonb02as1n16x5 _26220_ (.a(net881),
    .b(\us20.a[2] ),
    .out0(_17410_));
 b15bfn001al1n08x5 input33 (.a(key[13]),
    .o(net33));
 b15bfn000ah1n06x5 input32 (.a(key[12]),
    .o(net32));
 b15nor002al1n04x5 _26223_ (.a(\us20.a[4] ),
    .b(\us20.a[6] ),
    .o1(_17413_));
 b15nanb02ah1n24x5 _26224_ (.a(net863),
    .b(net867),
    .out0(_17414_));
 b15nanb02as1n12x5 _26225_ (.a(\us20.a[0] ),
    .b(\us20.a[7] ),
    .out0(_17415_));
 b15oai012aq1n08x5 _26226_ (.a(_17414_),
    .b(_17415_),
    .c(net869),
    .o1(_17416_));
 b15aoi013al1n06x5 _26227_ (.a(\us20.a[3] ),
    .b(_17410_),
    .c(_17413_),
    .d(_17416_),
    .o1(_17417_));
 b15nand02ar1n02x5 _26228_ (.a(_16018_),
    .b(_16058_),
    .o1(_17418_));
 b15aob012an1n03x5 _26229_ (.a(net885),
    .b(_15956_),
    .c(_17418_),
    .out0(_17419_));
 b15norp02al1n48x5 _26230_ (.a(\us20.a[1] ),
    .b(net875),
    .o1(_17420_));
 b15aoi022al1n06x5 _26231_ (.a(_16034_),
    .b(_17420_),
    .c(_16058_),
    .d(net880),
    .o1(_17421_));
 b15bfn000an1n02x5 input31 (.a(key[127]),
    .o(net31));
 b15oai112an1n12x5 _26233_ (.a(_17417_),
    .b(_17419_),
    .c(_17421_),
    .d(net885),
    .o1(_17423_));
 b15nor003ar1n06x5 _26234_ (.a(_15997_),
    .b(_15987_),
    .c(_16021_),
    .o1(_17424_));
 b15oai012an1n04x5 _26235_ (.a(_16040_),
    .b(_16125_),
    .c(net880),
    .o1(_17425_));
 b15oai012ar1n04x5 _26236_ (.a(net875),
    .b(_17424_),
    .c(_17425_),
    .o1(_17426_));
 b15norp02aq1n16x5 _26237_ (.a(_15987_),
    .b(_16021_),
    .o1(_17427_));
 b15aoi022ar1n04x5 _26238_ (.a(net885),
    .b(_17427_),
    .c(_16045_),
    .d(_16078_),
    .o1(_17428_));
 b15oai112ah1n06x5 _26239_ (.a(net874),
    .b(_17426_),
    .c(_17428_),
    .d(_16110_),
    .o1(_17429_));
 b15aoi012ar1n08x5 _26240_ (.a(_17409_),
    .b(_17423_),
    .c(_17429_),
    .o1(_17430_));
 b15oai012ar1n02x5 _26241_ (.a(net883),
    .b(_15970_),
    .c(_16160_),
    .o1(_17431_));
 b15nand02ah1n12x5 _26242_ (.a(net879),
    .b(net872),
    .o1(_17432_));
 b15oaoi13ah1n02x5 _26243_ (.a(_16136_),
    .b(_17431_),
    .c(_17432_),
    .d(net883),
    .o1(_17433_));
 b15norp03ah1n12x5 _26244_ (.a(net873),
    .b(_16031_),
    .c(_16061_),
    .o1(_17434_));
 b15norp02ar1n02x5 _26245_ (.a(_16132_),
    .b(_16007_),
    .o1(_17435_));
 b15nor003an1n03x5 _26246_ (.a(_17433_),
    .b(_17434_),
    .c(_17435_),
    .o1(_17436_));
 b15nor002ah1n12x5 _26247_ (.a(_16085_),
    .b(_15988_),
    .o1(_17437_));
 b15bfn000ah1n02x5 input30 (.a(key[126]),
    .o(net30));
 b15bfn000aq1n02x5 input29 (.a(key[125]),
    .o(net29));
 b15xor002ar1n02x5 _26250_ (.a(net883),
    .b(_15975_),
    .out0(_17440_));
 b15aoai13ar1n02x5 _26251_ (.a(_17437_),
    .b(_15974_),
    .c(_16078_),
    .d(_17440_),
    .o1(_17441_));
 b15nona22an1n08x5 _26252_ (.a(\us20.a[7] ),
    .b(\us20.a[3] ),
    .c(net866),
    .out0(_17442_));
 b15nor002ah1n04x5 _26253_ (.a(_15987_),
    .b(_17442_),
    .o1(_17443_));
 b15and002as1n04x5 _26254_ (.a(net873),
    .b(_16034_),
    .o(_17444_));
 b15aoi022al1n04x5 _26255_ (.a(_15963_),
    .b(_17443_),
    .c(_17444_),
    .d(_17410_),
    .o1(_17445_));
 b15nor002aq1n24x5 _26256_ (.a(_16080_),
    .b(_16082_),
    .o1(_17446_));
 b15and002ah1n12x5 _26257_ (.a(net879),
    .b(net872),
    .o(_17447_));
 b15norp02aq1n04x5 _26258_ (.a(net879),
    .b(net872),
    .o1(_17448_));
 b15nor003aq1n04x5 _26259_ (.a(net882),
    .b(_16080_),
    .c(_16113_),
    .o1(_17449_));
 b15aoi022as1n04x5 _26260_ (.a(_17446_),
    .b(_17447_),
    .c(_17448_),
    .d(_17449_),
    .o1(_17450_));
 b15bfn000ar1n02x5 input28 (.a(key[124]),
    .o(net28));
 b15oai022as1n02x5 _26262_ (.a(net883),
    .b(_17445_),
    .c(_17450_),
    .d(net876),
    .o1(_17452_));
 b15nano22al1n05x5 _26263_ (.a(_17436_),
    .b(_17441_),
    .c(_17452_),
    .out0(_17453_));
 b15xor002an1n04x5 _26264_ (.a(net871),
    .b(net878),
    .out0(_17454_));
 b15nandp2al1n12x5 _26265_ (.a(net866),
    .b(net884),
    .o1(_17455_));
 b15nano23ar1n02x5 _26266_ (.a(net863),
    .b(_17454_),
    .c(_17455_),
    .d(net869),
    .out0(_17456_));
 b15nonb02as1n16x5 _26267_ (.a(\us20.a[4] ),
    .b(net869),
    .out0(_17457_));
 b15nand02an1n32x5 _26268_ (.a(_16096_),
    .b(_17457_),
    .o1(_17458_));
 b15oai012ah1n16x5 _26269_ (.a(net877),
    .b(net881),
    .c(net884),
    .o1(_17459_));
 b15oab012aq1n02x5 _26270_ (.a(_17456_),
    .b(_17458_),
    .c(_17459_),
    .out0(_17460_));
 b15aoi012ah1n02x5 _26271_ (.a(net873),
    .b(_16067_),
    .c(_17460_),
    .o1(_17461_));
 b15nanb02an1n12x5 _26272_ (.a(net871),
    .b(net863),
    .out0(_17462_));
 b15inv000as1n20x5 _26273_ (.a(net867),
    .o1(_17463_));
 b15bfn000al1n02x5 input27 (.a(key[123]),
    .o(net27));
 b15oai012ar1n08x5 _26275_ (.a(_16082_),
    .b(_17462_),
    .c(_17463_),
    .o1(_17465_));
 b15nand04ah1n02x5 _26276_ (.a(net866),
    .b(_15997_),
    .c(_16129_),
    .d(_17465_),
    .o1(_17466_));
 b15aoai13aq1n06x5 _26277_ (.a(_15939_),
    .b(_15952_),
    .c(_16065_),
    .d(_16145_),
    .o1(_17467_));
 b15aoi012al1n02x5 _26278_ (.a(_15995_),
    .b(_17466_),
    .c(_17467_),
    .o1(_17468_));
 b15and002as1n16x5 _26279_ (.a(net885),
    .b(\us20.a[1] ),
    .o(_17469_));
 b15norp03ar1n02x5 _26280_ (.a(net878),
    .b(_16028_),
    .c(_16125_),
    .o1(_17470_));
 b15aoai13al1n02x5 _26281_ (.a(_17469_),
    .b(_17470_),
    .c(_16074_),
    .d(net878),
    .o1(_17471_));
 b15mdn022ar1n02x5 _26282_ (.a(_16134_),
    .b(_16137_),
    .o1(_17472_),
    .sa(_16088_));
 b15aoi022ar1n02x5 _26283_ (.a(_17457_),
    .b(_15974_),
    .c(_17472_),
    .d(net869),
    .o1(_17473_));
 b15oai013al1n04x5 _26284_ (.a(_17471_),
    .b(_17473_),
    .c(_16126_),
    .d(_15997_),
    .o1(_17474_));
 b15norp03an1n08x5 _26285_ (.a(_17461_),
    .b(_17468_),
    .c(_17474_),
    .o1(_17475_));
 b15aoi112aq1n03x5 _26286_ (.a(\us20.a[4] ),
    .b(\us20.a[7] ),
    .c(net885),
    .d(\us20.a[1] ),
    .o1(_17476_));
 b15nano23ar1n02x5 _26287_ (.a(\us20.a[4] ),
    .b(\us20.a[7] ),
    .c(\us20.a[1] ),
    .d(net868),
    .out0(_17477_));
 b15oab012al1n02x5 _26288_ (.a(\us20.a[6] ),
    .b(_17476_),
    .c(_17477_),
    .out0(_17478_));
 b15nandp2ar1n24x5 _26289_ (.a(net869),
    .b(\us20.a[7] ),
    .o1(_17479_));
 b15and002ah1n03x5 _26290_ (.a(\us20.a[4] ),
    .b(\us20.a[6] ),
    .o(_17480_));
 b15oai013as1n02x5 _26291_ (.a(\us20.a[2] ),
    .b(_17479_),
    .c(_17413_),
    .d(_17480_),
    .o1(_17481_));
 b15aoi012al1n04x5 _26292_ (.a(_17478_),
    .b(_17481_),
    .c(_16145_),
    .o1(_17482_));
 b15aoi012ar1n04x5 _26293_ (.a(\us20.a[2] ),
    .b(_16145_),
    .c(_16045_),
    .o1(_17483_));
 b15nor003ar1n12x5 _26294_ (.a(\us20.a[3] ),
    .b(_17482_),
    .c(_17483_),
    .o1(_17484_));
 b15bfn000as1n02x5 input26 (.a(key[122]),
    .o(net26));
 b15nand02ar1n02x5 _26296_ (.a(net882),
    .b(net872),
    .o1(_17486_));
 b15andc04aq1n16x5 _26297_ (.a(net868),
    .b(net870),
    .c(net863),
    .d(net865),
    .o(_17487_));
 b15nandp2an1n03x5 _26298_ (.a(net879),
    .b(_17487_),
    .o1(_17488_));
 b15oaoi13aq1n02x5 _26299_ (.a(_17486_),
    .b(_17488_),
    .c(net879),
    .d(_16136_),
    .o1(_17489_));
 b15nor003ah1n08x5 _26300_ (.a(net872),
    .b(_16080_),
    .c(_16082_),
    .o1(_17490_));
 b15and002al1n04x5 _26301_ (.a(_16078_),
    .b(_17490_),
    .o(_17491_));
 b15oab012ah1n08x5 _26302_ (.c(_17491_),
    .a(net875),
    .b(_17489_),
    .out0(_17492_));
 b15nor002aq1n06x5 _26303_ (.a(net883),
    .b(_16137_),
    .o1(_17493_));
 b15aoai13aq1n08x5 _26304_ (.a(_17493_),
    .b(_17446_),
    .c(_16078_),
    .d(_16058_),
    .o1(_17494_));
 b15aoai13as1n02x5 _26305_ (.a(_17410_),
    .b(_16141_),
    .c(\us20.a[3] ),
    .d(_16069_),
    .o1(_17495_));
 b15xor002ar1n02x5 _26306_ (.a(net867),
    .b(net866),
    .out0(_17496_));
 b15nanb02aq1n16x5 _26307_ (.a(net863),
    .b(net871),
    .out0(_17497_));
 b15nano23al1n02x5 _26308_ (.a(_17420_),
    .b(_17496_),
    .c(_17497_),
    .d(_16028_),
    .out0(_17498_));
 b15aoi012an1n02x5 _26309_ (.a(_17498_),
    .b(_16141_),
    .c(net884),
    .o1(_17499_));
 b15nanb02ar1n02x5 _26310_ (.a(\us20.a[3] ),
    .b(net867),
    .out0(_17500_));
 b15oai012an1n04x5 _26311_ (.a(_17500_),
    .b(_16134_),
    .c(net867),
    .o1(_17501_));
 b15nor003aq1n03x5 _26312_ (.a(net881),
    .b(_17462_),
    .c(_16090_),
    .o1(_17502_));
 b15nanb02as1n24x5 _26313_ (.a(net866),
    .b(net881),
    .out0(_17503_));
 b15nanb02as1n06x5 _26314_ (.a(net881),
    .b(net866),
    .out0(_17504_));
 b15oai022aq1n04x5 _26315_ (.a(_17497_),
    .b(_17503_),
    .c(_17504_),
    .d(_17462_),
    .o1(_17505_));
 b15nor003ah1n02x5 _26316_ (.a(net867),
    .b(net884),
    .c(_15995_),
    .o1(_17506_));
 b15aoi022aq1n08x5 _26317_ (.a(_17501_),
    .b(_17502_),
    .c(_17505_),
    .d(_17506_),
    .o1(_17507_));
 b15nand04ah1n08x5 _26318_ (.a(_17494_),
    .b(_17495_),
    .c(_17499_),
    .d(_17507_),
    .o1(_17508_));
 b15nor002ah1n16x5 _26319_ (.a(_16113_),
    .b(_16021_),
    .o1(_17509_));
 b15nandp3ar1n03x5 _26320_ (.a(_15997_),
    .b(_15974_),
    .c(_17509_),
    .o1(_17510_));
 b15oai022aq1n04x5 _26321_ (.a(_15993_),
    .b(_16150_),
    .c(_16162_),
    .d(_15995_),
    .o1(_17511_));
 b15nand03ah1n02x5 _26322_ (.a(\us20.a[1] ),
    .b(_15969_),
    .c(_17511_),
    .o1(_17512_));
 b15nor002ah1n06x5 _26323_ (.a(net866),
    .b(_16085_),
    .o1(_17513_));
 b15nand02ar1n02x5 _26324_ (.a(\us20.a[3] ),
    .b(_17415_),
    .o1(_17514_));
 b15nand04aq1n04x5 _26325_ (.a(_17410_),
    .b(_16153_),
    .c(_17513_),
    .d(_17514_),
    .o1(_17515_));
 b15orn003an1n02x5 _26326_ (.a(net864),
    .b(net882),
    .c(net874),
    .o(_17516_));
 b15nandp3al1n08x5 _26327_ (.a(\us20.a[6] ),
    .b(net879),
    .c(net875),
    .o1(_17517_));
 b15orn002as1n08x5 _26328_ (.a(net879),
    .b(net875),
    .o(_17518_));
 b15oaoi13as1n08x5 _26329_ (.a(_17516_),
    .b(_17517_),
    .c(_17518_),
    .d(\us20.a[6] ),
    .o1(_17519_));
 b15orn002ah1n03x5 _26330_ (.a(net880),
    .b(net872),
    .o(_17520_));
 b15oai022aq1n08x5 _26331_ (.a(_16021_),
    .b(_17432_),
    .c(_17520_),
    .d(_15988_),
    .o1(_17521_));
 b15norp02ar1n08x5 _26332_ (.a(_15959_),
    .b(_16018_),
    .o1(_17522_));
 b15aoai13as1n08x5 _26333_ (.a(_15952_),
    .b(_17519_),
    .c(_17521_),
    .d(_17522_),
    .o1(_17523_));
 b15nand04al1n08x5 _26334_ (.a(_17510_),
    .b(_17512_),
    .c(_17515_),
    .d(_17523_),
    .o1(_17524_));
 b15nor004an1n12x5 _26335_ (.a(_17484_),
    .b(_17492_),
    .c(_17508_),
    .d(_17524_),
    .o1(_17525_));
 b15andc04as1n16x5 _26336_ (.a(_17430_),
    .b(_17453_),
    .c(_17475_),
    .d(_17525_),
    .o(_17526_));
 b15xor002al1n04x5 _26337_ (.a(_16424_),
    .b(_17526_),
    .out0(_17527_));
 b15xnr002al1n04x5 _26338_ (.a(_17396_),
    .b(_17527_),
    .out0(_17528_));
 b15xor002ar1n03x5 _26339_ (.a(_17283_),
    .b(_17528_),
    .out0(_17529_));
 b15cmbn22aq1n08x5 _26340_ (.clk1(\text_in_r[33] ),
    .clk2(_17529_),
    .clkout(_17530_),
    .s(net540));
 b15xor002as1n16x5 _26341_ (.a(net531),
    .b(_17530_),
    .out0(_00114_));
 b15inv000al1n12x5 _26342_ (.a(\text_in_r[34] ),
    .o1(_17531_));
 b15nand04ar1n03x5 _26343_ (.a(_16466_),
    .b(_16609_),
    .c(_16620_),
    .d(_17112_),
    .o1(_17532_));
 b15aoi012al1n02x5 _26344_ (.a(net613),
    .b(_16608_),
    .c(_17532_),
    .o1(_17533_));
 b15aoai13ah1n03x5 _26345_ (.a(_16585_),
    .b(_17533_),
    .c(_16670_),
    .d(_17128_),
    .o1(_17534_));
 b15bfn000ah1n03x5 input25 (.a(key[121]),
    .o(net25));
 b15nand02ah1n06x5 _26347_ (.a(_17152_),
    .b(_16650_),
    .o1(_17536_));
 b15oai112al1n12x5 _26348_ (.a(_16558_),
    .b(_17536_),
    .c(_17183_),
    .d(_16524_),
    .o1(_17537_));
 b15orn003ar1n02x5 _26349_ (.a(net608),
    .b(_16652_),
    .c(_16528_),
    .o(_17538_));
 b15oai013aq1n06x5 _26350_ (.a(_17538_),
    .b(_17125_),
    .c(_16504_),
    .d(_16466_),
    .o1(_17539_));
 b15oai012ar1n16x5 _26351_ (.a(_17537_),
    .b(_17539_),
    .c(_16558_),
    .o1(_17540_));
 b15nand02as1n06x5 _26352_ (.a(_16526_),
    .b(_16591_),
    .o1(_17541_));
 b15nonb02al1n06x5 _26353_ (.a(net598),
    .b(net603),
    .out0(_17542_));
 b15oai112al1n12x5 _26354_ (.a(_16659_),
    .b(_16597_),
    .c(_17542_),
    .d(_16678_),
    .o1(_17543_));
 b15oaoi13aq1n03x5 _26355_ (.a(net614),
    .b(_17541_),
    .c(_17543_),
    .d(net609),
    .o1(_17544_));
 b15and002ar1n24x5 _26356_ (.a(net599),
    .b(\us13.a[2] ),
    .o(_17545_));
 b15nand02an1n02x5 _26357_ (.a(_16481_),
    .b(_17545_),
    .o1(_17546_));
 b15oai012al1n03x5 _26358_ (.a(_16517_),
    .b(_17545_),
    .c(_16511_),
    .o1(_17547_));
 b15aoi112an1n04x5 _26359_ (.a(_16458_),
    .b(net609),
    .c(_17546_),
    .d(_17547_),
    .o1(_17548_));
 b15aoi012ah1n06x5 _26360_ (.a(_17544_),
    .b(_17548_),
    .c(net614),
    .o1(_17549_));
 b15nand02an1n02x5 _26361_ (.a(_16682_),
    .b(_16542_),
    .o1(_17550_));
 b15qgbna2an1n05x5 _26362_ (.o1(_17551_),
    .a(net599),
    .b(_16517_));
 b15oaoi13as1n04x5 _26363_ (.a(_17550_),
    .b(_17551_),
    .c(net599),
    .d(_16497_),
    .o1(_17552_));
 b15nonb03ah1n04x5 _26364_ (.a(net596),
    .b(net609),
    .c(net606),
    .out0(_17553_));
 b15aoai13ah1n02x5 _26365_ (.a(_17553_),
    .b(_17179_),
    .c(_16446_),
    .d(net613),
    .o1(_17554_));
 b15oai122al1n08x5 _26366_ (.a(_17554_),
    .b(_16680_),
    .c(_16498_),
    .d(_16479_),
    .e(_16521_),
    .o1(_17555_));
 b15oai012aq1n06x5 _26367_ (.a(net614),
    .b(_17552_),
    .c(_17555_),
    .o1(_17556_));
 b15nand04aq1n16x5 _26368_ (.a(_17534_),
    .b(_17540_),
    .c(_17549_),
    .d(_17556_),
    .o1(_17557_));
 b15and003ar1n02x5 _26369_ (.a(_16481_),
    .b(_16456_),
    .c(_16518_),
    .o(_17558_));
 b15norp03al1n08x5 _26370_ (.a(_17099_),
    .b(_16458_),
    .c(_16535_),
    .o1(_17559_));
 b15aoi013ah1n02x5 _26371_ (.a(_17558_),
    .b(_17559_),
    .c(_16513_),
    .d(_16500_),
    .o1(_17560_));
 b15oaoi13an1n04x5 _26372_ (.a(_16460_),
    .b(_17560_),
    .c(_16643_),
    .d(net610),
    .o1(_17561_));
 b15nano23an1n24x5 _26373_ (.a(net602),
    .b(net607),
    .c(net596),
    .d(net600),
    .out0(_17562_));
 b15nand02al1n12x5 _26374_ (.a(_17562_),
    .b(_16648_),
    .o1(_17563_));
 b15oai012an1n04x5 _26375_ (.a(_17563_),
    .b(_16477_),
    .c(_16453_),
    .o1(_17564_));
 b15nonb02ah1n08x5 _26376_ (.a(\us13.a[0] ),
    .b(\us13.a[2] ),
    .out0(_17565_));
 b15nano22as1n02x5 _26377_ (.a(net598),
    .b(net599),
    .c(\us13.a[3] ),
    .out0(_17566_));
 b15oai112aq1n12x5 _26378_ (.a(_17565_),
    .b(_16517_),
    .c(_16518_),
    .d(_17566_),
    .o1(_17567_));
 b15oai013ah1n06x5 _26379_ (.a(_17567_),
    .b(_17543_),
    .c(_16682_),
    .d(net609),
    .o1(_17568_));
 b15oai022ah1n08x5 _26380_ (.a(_16498_),
    .b(_17091_),
    .c(_17164_),
    .d(_16435_),
    .o1(_17569_));
 b15aoi112an1n06x5 _26381_ (.a(_17564_),
    .b(_17568_),
    .c(_17569_),
    .d(net613),
    .o1(_17570_));
 b15aoi012ar1n02x5 _26382_ (.a(net613),
    .b(_16671_),
    .c(_16558_),
    .o1(_17571_));
 b15oai112ar1n04x5 _26383_ (.a(_16621_),
    .b(_17542_),
    .c(_17571_),
    .d(_16508_),
    .o1(_17572_));
 b15aoi022ar1n02x5 _26384_ (.a(_16678_),
    .b(_16657_),
    .c(_17161_),
    .d(_17542_),
    .o1(_17573_));
 b15nand02ah1n08x5 _26385_ (.a(_16592_),
    .b(_16453_),
    .o1(_17574_));
 b15nanb03ar1n02x5 _26386_ (.a(_17573_),
    .b(net605),
    .c(_17574_),
    .out0(_17575_));
 b15aoi022aq1n04x5 _26387_ (.a(net610),
    .b(_16650_),
    .c(_16684_),
    .d(_16510_),
    .o1(_17576_));
 b15norp03ar1n03x5 _26388_ (.a(net617),
    .b(_17088_),
    .c(_17576_),
    .o1(_17577_));
 b15nand02ah1n24x5 _26389_ (.a(_16577_),
    .b(_16517_),
    .o1(_17578_));
 b15oaoi13an1n02x5 _26390_ (.a(_16585_),
    .b(_17541_),
    .c(_17578_),
    .d(_16479_),
    .o1(_17579_));
 b15nano23an1n03x5 _26391_ (.a(_17572_),
    .b(_17575_),
    .c(_17577_),
    .d(_17579_),
    .out0(_17580_));
 b15xor002ar1n02x5 _26392_ (.a(net605),
    .b(\us13.a[0] ),
    .out0(_17581_));
 b15nano23al1n03x5 _26393_ (.a(_16504_),
    .b(_16510_),
    .c(_17581_),
    .d(net609),
    .out0(_17582_));
 b15oab012ar1n02x5 _26394_ (.a(net613),
    .b(net614),
    .c(net605),
    .out0(_17583_));
 b15nor003al1n04x5 _26395_ (.a(_16498_),
    .b(_16594_),
    .c(_17583_),
    .o1(_17584_));
 b15oai012ah1n06x5 _26396_ (.a(net599),
    .b(_17582_),
    .c(_17584_),
    .o1(_17585_));
 b15orn002as1n03x5 _26397_ (.a(net605),
    .b(net598),
    .o(_17586_));
 b15oai022ar1n02x5 _26398_ (.a(_16522_),
    .b(_17586_),
    .c(_16524_),
    .d(_16665_),
    .o1(_17587_));
 b15qgbbf1an1n05x5 input24 (.a(key[120]),
    .o(net24));
 b15aoi022as1n04x5 _26400_ (.a(_16517_),
    .b(_16542_),
    .c(_17587_),
    .d(net603),
    .o1(_17589_));
 b15oai112ah1n12x5 _26401_ (.a(_16607_),
    .b(_17585_),
    .c(_17589_),
    .d(_16564_),
    .o1(_17590_));
 b15bfn000aq1n02x5 input23 (.a(key[11]),
    .o(net23));
 b15aob012ar1n02x5 _26403_ (.a(net617),
    .b(_16429_),
    .c(_16520_),
    .out0(_17592_));
 b15oai022ar1n02x5 _26404_ (.a(net605),
    .b(_16522_),
    .c(_17080_),
    .d(net609),
    .o1(_17593_));
 b15aoi013ah1n02x5 _26405_ (.a(_17592_),
    .b(_17593_),
    .c(_16577_),
    .d(_17099_),
    .o1(_17594_));
 b15aoi012al1n02x5 _26406_ (.a(net617),
    .b(_16466_),
    .c(_17087_),
    .o1(_17595_));
 b15norp03ar1n08x5 _26407_ (.a(net618),
    .b(_17594_),
    .c(_17595_),
    .o1(_17596_));
 b15nano23as1n12x5 _26408_ (.a(_17570_),
    .b(_17580_),
    .c(_17590_),
    .d(_17596_),
    .out0(_17597_));
 b15aoi012ar1n02x5 _26409_ (.a(net612),
    .b(_16643_),
    .c(net616),
    .o1(_17598_));
 b15and002ar1n02x5 _26410_ (.a(_16558_),
    .b(_17562_),
    .o(_17599_));
 b15oai013as1n04x5 _26411_ (.a(_17598_),
    .b(_17599_),
    .c(_16674_),
    .d(net616),
    .o1(_17600_));
 b15nandp3al1n04x5 _26412_ (.a(_16619_),
    .b(_16579_),
    .c(_16605_),
    .o1(_17601_));
 b15nand02al1n24x5 _26413_ (.a(net616),
    .b(net612),
    .o1(_17602_));
 b15norp03aq1n02x5 _26414_ (.a(net597),
    .b(_16671_),
    .c(_17602_),
    .o1(_17603_));
 b15nandp2al1n02x5 _26415_ (.a(_16652_),
    .b(_17088_),
    .o1(_17604_));
 b15aoi013an1n04x5 _26416_ (.a(_17603_),
    .b(_17604_),
    .c(net597),
    .d(_16579_),
    .o1(_17605_));
 b15oai112al1n16x5 _26417_ (.a(_17600_),
    .b(_17601_),
    .c(_17605_),
    .d(_16597_),
    .o1(_17606_));
 b15nor002as1n03x5 _26418_ (.a(_16671_),
    .b(_16595_),
    .o1(_17607_));
 b15nanb02ar1n03x5 _26419_ (.a(net614),
    .b(net605),
    .out0(_17608_));
 b15oai112al1n06x5 _26420_ (.a(\us13.a[5] ),
    .b(_17608_),
    .c(_16652_),
    .d(net605),
    .o1(_17609_));
 b15aoi012ar1n02x5 _26421_ (.a(net598),
    .b(_17080_),
    .c(_17099_),
    .o1(_17610_));
 b15aoai13ah1n03x5 _26422_ (.a(net599),
    .b(_17607_),
    .c(_17609_),
    .d(_17610_),
    .o1(_17611_));
 b15nandp2an1n03x5 _26423_ (.a(_16597_),
    .b(\us13.a[2] ),
    .o1(_17612_));
 b15oai013as1n08x5 _26424_ (.a(_17611_),
    .b(_17612_),
    .c(_16673_),
    .d(\us13.a[7] ),
    .o1(_17613_));
 b15aoai13as1n08x5 _26425_ (.a(net610),
    .b(_17606_),
    .c(_17613_),
    .d(net620),
    .o1(_17614_));
 b15nona23as1n32x5 _26426_ (.a(_17557_),
    .b(_17561_),
    .c(_17597_),
    .d(_17614_),
    .out0(_17615_));
 b15nandp2aq1n03x5 _26427_ (.a(_16028_),
    .b(_16069_),
    .o1(_17616_));
 b15aoi112an1n03x5 _26428_ (.a(net882),
    .b(net875),
    .c(_17616_),
    .d(_17401_),
    .o1(_00529_));
 b15aoai13ah1n02x5 _26429_ (.a(net879),
    .b(_00529_),
    .c(_17437_),
    .d(_16160_),
    .o1(_00530_));
 b15nand02an1n06x5 _26430_ (.a(net883),
    .b(_16133_),
    .o1(_00531_));
 b15nand02ar1n02x5 _26431_ (.a(net870),
    .b(net879),
    .o1(_00532_));
 b15oai022ar1n02x5 _26432_ (.a(net879),
    .b(_16113_),
    .c(_00532_),
    .d(net868),
    .o1(_00533_));
 b15and003al1n02x5 _26433_ (.a(_16008_),
    .b(_16066_),
    .c(_00533_),
    .o(_00534_));
 b15xor002ah1n16x5 _26434_ (.a(net880),
    .b(net877),
    .out0(_00535_));
 b15orn002ah1n02x5 _26435_ (.a(_15959_),
    .b(_00535_),
    .o(_00536_));
 b15oaoi13as1n02x5 _26436_ (.a(_17458_),
    .b(_00536_),
    .c(net882),
    .d(_17420_),
    .o1(_00537_));
 b15oai012ar1n08x5 _26437_ (.a(net872),
    .b(_00534_),
    .c(_00537_),
    .o1(_00538_));
 b15oai112al1n02x5 _26438_ (.a(_17410_),
    .b(_16112_),
    .c(_16075_),
    .d(_16045_),
    .o1(_00539_));
 b15norp02an1n08x5 _26439_ (.a(net868),
    .b(net864),
    .o1(_00540_));
 b15nonb02as1n06x5 _26440_ (.a(net885),
    .b(net875),
    .out0(_00541_));
 b15oai012aq1n06x5 _26441_ (.a(_00540_),
    .b(_00541_),
    .c(_16078_),
    .o1(_00542_));
 b15nanb02ah1n16x5 _26442_ (.a(net882),
    .b(net876),
    .out0(_00543_));
 b15oai012ar1n06x5 _26443_ (.a(_00542_),
    .b(_00543_),
    .c(_17479_),
    .o1(_00544_));
 b15nor002aq1n04x5 _26444_ (.a(net865),
    .b(_16100_),
    .o1(_00545_));
 b15aobi12al1n04x5 _26445_ (.a(_00539_),
    .b(_00544_),
    .c(_00545_),
    .out0(_00546_));
 b15nand04aq1n08x5 _26446_ (.a(_00530_),
    .b(_00531_),
    .c(_00538_),
    .d(_00546_),
    .o1(_00547_));
 b15aoi012al1n04x5 _26447_ (.a(_16110_),
    .b(_17420_),
    .c(_16040_),
    .o1(_00548_));
 b15nor002ar1n04x5 _26448_ (.a(_17407_),
    .b(_00541_),
    .o1(_00549_));
 b15norp02ar1n48x5 _26449_ (.a(_16126_),
    .b(_16113_),
    .o1(_00550_));
 b15oai222an1n16x5 _26450_ (.a(net882),
    .b(_00548_),
    .c(_00549_),
    .d(_16078_),
    .e(_00550_),
    .f(_16045_),
    .o1(_00551_));
 b15nor003as1n02x5 _26451_ (.a(net866),
    .b(_15997_),
    .c(_17497_),
    .o1(_00552_));
 b15nor002ar1n03x5 _26452_ (.a(net871),
    .b(_16126_),
    .o1(_00553_));
 b15oaoi13an1n04x5 _26453_ (.a(_16018_),
    .b(_17463_),
    .c(_00552_),
    .d(_00553_),
    .o1(_00554_));
 b15norp03ar1n02x5 _26454_ (.a(\us20.a[7] ),
    .b(_16085_),
    .c(_16129_),
    .o1(_00555_));
 b15norp02ar1n02x5 _26455_ (.a(_15987_),
    .b(_17415_),
    .o1(_00556_));
 b15oaoi13as1n02x5 _26456_ (.a(net878),
    .b(_16092_),
    .c(_00555_),
    .d(_00556_),
    .o1(_00557_));
 b15oab012ah1n08x5 _26457_ (.c(_00557_),
    .a(\us20.a[3] ),
    .b(_00554_),
    .out0(_00558_));
 b15nonb02ar1n02x5 _26458_ (.a(net875),
    .b(net870),
    .out0(_00559_));
 b15aoai13ar1n02x5 _26459_ (.a(_00540_),
    .b(_00559_),
    .c(net870),
    .d(_00541_),
    .o1(_00560_));
 b15nand02ar1n08x5 _26460_ (.a(net864),
    .b(_16065_),
    .o1(_00561_));
 b15oaoi13as1n02x5 _26461_ (.a(\us20.a[6] ),
    .b(_00560_),
    .c(_00561_),
    .d(net875),
    .o1(_00562_));
 b15oai012as1n04x5 _26462_ (.a(net879),
    .b(_16047_),
    .c(_00562_),
    .o1(_00563_));
 b15aoi022an1n12x5 _26463_ (.a(net872),
    .b(_00551_),
    .c(_00558_),
    .d(_00563_),
    .o1(_00564_));
 b15nor003al1n03x5 _26464_ (.a(net873),
    .b(_17455_),
    .c(_17414_),
    .o1(_00565_));
 b15aoai13ar1n04x5 _26465_ (.a(net880),
    .b(_16133_),
    .c(_00565_),
    .d(net871),
    .o1(_00566_));
 b15aoai13aq1n02x5 _26466_ (.a(net880),
    .b(_16044_),
    .c(net873),
    .d(net883),
    .o1(_00567_));
 b15oai012an1n02x5 _26467_ (.a(_16028_),
    .b(_16085_),
    .c(_16021_),
    .o1(_00568_));
 b15bfn000as1n02x5 input22 (.a(key[119]),
    .o(net22));
 b15oai112aq1n06x5 _26469_ (.a(_00567_),
    .b(_00568_),
    .c(_16028_),
    .d(_16068_),
    .o1(_00570_));
 b15nor002aq1n02x5 _26470_ (.a(_16125_),
    .b(_17469_),
    .o1(_00571_));
 b15oaoi13an1n03x5 _26471_ (.a(_17410_),
    .b(_15963_),
    .c(_16113_),
    .d(_16080_),
    .o1(_00572_));
 b15oai122ah1n08x5 _26472_ (.a(_16028_),
    .b(_16164_),
    .c(_00571_),
    .d(_00572_),
    .e(net883),
    .o1(_00573_));
 b15nanb03ar1n02x5 _26473_ (.a(net871),
    .b(net876),
    .c(net869),
    .out0(_00574_));
 b15oaoi13as1n02x5 _26474_ (.a(net873),
    .b(_00574_),
    .c(_16000_),
    .d(_16082_),
    .o1(_00575_));
 b15and003ar1n02x5 _26475_ (.a(net876),
    .b(_17457_),
    .c(_16104_),
    .o(_00576_));
 b15oai112al1n08x5 _26476_ (.a(net885),
    .b(_16008_),
    .c(_00575_),
    .d(_00576_),
    .o1(_00577_));
 b15nand04aq1n12x5 _26477_ (.a(_00566_),
    .b(_00570_),
    .c(_00573_),
    .d(_00577_),
    .o1(_00578_));
 b15nor003aq1n03x5 _26478_ (.a(_16085_),
    .b(_16021_),
    .c(_16134_),
    .o1(_00579_));
 b15orn002ar1n02x5 _26479_ (.a(net871),
    .b(net881),
    .o(_00580_));
 b15nor004ar1n06x5 _26480_ (.a(net873),
    .b(_17455_),
    .c(_17414_),
    .d(_00580_),
    .o1(_00581_));
 b15nor004ar1n06x5 _26481_ (.a(net873),
    .b(_16126_),
    .c(_16113_),
    .d(_16011_),
    .o1(_00582_));
 b15qgbno3an1n05x5 _26482_ (.o1(_00583_),
    .a(_16004_),
    .b(_16000_),
    .c(_16112_));
 b15nor004ar1n08x5 _26483_ (.a(_00579_),
    .b(_00581_),
    .c(_00582_),
    .d(_00583_),
    .o1(_00584_));
 b15nor003al1n08x5 _26484_ (.a(net871),
    .b(net863),
    .c(net865),
    .o1(_00585_));
 b15and003aq1n08x5 _26485_ (.a(net871),
    .b(net863),
    .c(net866),
    .o(_00586_));
 b15aoi022ar1n02x5 _26486_ (.a(_16160_),
    .b(_00585_),
    .c(_00586_),
    .d(_15970_),
    .o1(_00587_));
 b15orn003ah1n02x5 _26487_ (.a(_17463_),
    .b(_15947_),
    .c(_00587_),
    .o(_00588_));
 b15nona23ar1n24x5 _26488_ (.a(net871),
    .b(net865),
    .c(net863),
    .d(net869),
    .out0(_00589_));
 b15norp02an1n02x5 _26489_ (.a(net873),
    .b(_00589_),
    .o1(_00590_));
 b15aoi013ar1n06x5 _26490_ (.a(_00590_),
    .b(_16058_),
    .c(_15947_),
    .d(net873),
    .o1(_00591_));
 b15oai112aq1n16x5 _26491_ (.a(_00584_),
    .b(_00588_),
    .c(_00591_),
    .d(_17459_),
    .o1(_00592_));
 b15nanb02ar1n02x5 _26492_ (.a(\us20.a[7] ),
    .b(net884),
    .out0(_00593_));
 b15aoi112aq1n02x5 _26493_ (.a(_15995_),
    .b(_16150_),
    .c(_00593_),
    .d(net881),
    .o1(_00594_));
 b15norp03aq1n03x5 _26494_ (.a(\us20.a[3] ),
    .b(_16126_),
    .c(_16011_),
    .o1(_00595_));
 b15aoai13aq1n06x5 _26495_ (.a(_17463_),
    .b(_00594_),
    .c(_00595_),
    .d(net871),
    .o1(_00596_));
 b15aoi022ar1n02x5 _26496_ (.a(_15974_),
    .b(_00585_),
    .c(_00586_),
    .d(_15975_),
    .o1(_00597_));
 b15nanb02aq1n12x5 _26497_ (.a(net872),
    .b(net865),
    .out0(_00598_));
 b15nanb02as1n24x5 _26498_ (.a(net879),
    .b(net872),
    .out0(_00599_));
 b15nona22ah1n05x5 _26499_ (.a(net871),
    .b(net866),
    .c(net863),
    .out0(_00600_));
 b15oa0022ar1n02x5 _26500_ (.a(_17497_),
    .b(_00598_),
    .c(_00599_),
    .d(_00600_),
    .o(_00601_));
 b15oai022ar1n02x5 _26501_ (.a(net881),
    .b(_00597_),
    .c(_00601_),
    .d(_16077_),
    .o1(_00602_));
 b15aob012ar1n08x5 _26502_ (.a(_00596_),
    .b(_00602_),
    .c(net869),
    .out0(_00603_));
 b15nor003as1n04x5 _26503_ (.a(_15987_),
    .b(_16021_),
    .c(_16137_),
    .o1(_00604_));
 b15norp03ar1n12x5 _26504_ (.a(_16028_),
    .b(_15987_),
    .c(_15988_),
    .o1(_00605_));
 b15aoai13ar1n04x5 _26505_ (.a(_16078_),
    .b(_00604_),
    .c(_00605_),
    .d(_00543_),
    .o1(_00606_));
 b15aoi012ar1n04x5 _26506_ (.a(_00604_),
    .b(_17447_),
    .c(_17509_),
    .o1(_00607_));
 b15aoi022ah1n06x5 _26507_ (.a(_15974_),
    .b(_16164_),
    .c(_17448_),
    .d(_17487_),
    .o1(_00608_));
 b15aoai13as1n08x5 _26508_ (.a(_00606_),
    .b(net882),
    .c(_00607_),
    .d(_00608_),
    .o1(_00609_));
 b15nor004as1n12x5 _26509_ (.a(_00578_),
    .b(_00592_),
    .c(_00603_),
    .d(_00609_),
    .o1(_00610_));
 b15oaoi13al1n02x5 _26510_ (.a(_16028_),
    .b(_17522_),
    .c(_17487_),
    .d(_16147_),
    .o1(_00611_));
 b15qbfna2bn1n16x5 _26511_ (.a(_16147_),
    .b(_16006_),
    .o1(_00612_));
 b15aoai13ah1n03x5 _26512_ (.a(_00611_),
    .b(net875),
    .c(_00612_),
    .d(_17488_),
    .o1(_00613_));
 b15nor002al1n32x5 _26513_ (.a(_16126_),
    .b(_16082_),
    .o1(_00614_));
 b15oai022ar1n02x5 _26514_ (.a(_16061_),
    .b(_17401_),
    .c(_17458_),
    .d(net875),
    .o1(_00615_));
 b15aoi022ar1n02x5 _26515_ (.a(_17410_),
    .b(_00614_),
    .c(_00615_),
    .d(net882),
    .o1(_00616_));
 b15aob012aq1n12x5 _26516_ (.a(_00613_),
    .b(_00616_),
    .c(_16028_),
    .out0(_00617_));
 b15nona23as1n32x5 _26517_ (.a(_00547_),
    .b(_00564_),
    .c(_00610_),
    .d(_00617_),
    .out0(_00618_));
 b15xnr002as1n12x5 _26518_ (.a(_17615_),
    .b(_00618_),
    .out0(_00619_));
 b15nandp2al1n02x5 _26519_ (.a(_16213_),
    .b(_16997_),
    .o1(_00620_));
 b15nor002aq1n08x5 _26520_ (.a(_16389_),
    .b(_16993_),
    .o1(_00621_));
 b15nor002as1n06x5 _26521_ (.a(_16398_),
    .b(_16979_),
    .o1(_00622_));
 b15oaoi13as1n02x5 _26522_ (.a(_00621_),
    .b(_16233_),
    .c(_16239_),
    .d(_00622_),
    .o1(_00623_));
 b15aoai13an1n03x5 _26523_ (.a(net732),
    .b(_16403_),
    .c(_00622_),
    .d(net742),
    .o1(_00624_));
 b15aoi013as1n04x5 _26524_ (.a(net738),
    .b(_00620_),
    .c(_00623_),
    .d(_00624_),
    .o1(_00625_));
 b15bfn000as1n02x5 input21 (.a(key[118]),
    .o(net21));
 b15aoi022ar1n02x5 _26526_ (.a(_16259_),
    .b(_16316_),
    .c(_16333_),
    .d(_16328_),
    .o1(_00627_));
 b15oaoi13an1n02x5 _26527_ (.a(net737),
    .b(_16414_),
    .c(_00627_),
    .d(_16237_),
    .o1(_00628_));
 b15nand02ar1n02x5 _26528_ (.a(net727),
    .b(_16193_),
    .o1(_00629_));
 b15nand02ar1n02x5 _26529_ (.a(net735),
    .b(_16259_),
    .o1(_00630_));
 b15oaoi13ar1n03x5 _26530_ (.a(_00629_),
    .b(_00630_),
    .c(_16314_),
    .d(net735),
    .o1(_00631_));
 b15aoi012ar1n02x5 _26531_ (.a(_16379_),
    .b(_16420_),
    .c(_17045_),
    .o1(_00632_));
 b15oai013ah1n03x5 _26532_ (.a(net731),
    .b(_00628_),
    .c(_00631_),
    .d(_00632_),
    .o1(_00633_));
 b15nanb02ar1n03x5 _26533_ (.a(net722),
    .b(net717),
    .out0(_00634_));
 b15oai013aq1n02x5 _26534_ (.a(net729),
    .b(_17053_),
    .c(_16981_),
    .d(_00634_),
    .o1(_00635_));
 b15nor003al1n03x5 _26535_ (.a(net722),
    .b(net726),
    .c(net720),
    .o1(_00636_));
 b15aoai13an1n02x5 _26536_ (.a(net717),
    .b(_00636_),
    .c(_16194_),
    .d(_16185_),
    .o1(_00637_));
 b15aobi12ar1n02x5 _26537_ (.a(_17024_),
    .b(net720),
    .c(net742),
    .out0(_00638_));
 b15oai013ah1n02x5 _26538_ (.a(_00637_),
    .b(_00638_),
    .c(net717),
    .d(_16237_),
    .o1(_00639_));
 b15oa0012ar1n02x5 _26539_ (.a(_00634_),
    .b(_17203_),
    .c(net729),
    .o(_00640_));
 b15oai013ah1n02x5 _26540_ (.a(net737),
    .b(_17053_),
    .c(_16320_),
    .d(_00640_),
    .o1(_00641_));
 b15nandp3aq1n08x5 _26541_ (.a(_00635_),
    .b(_00639_),
    .c(_00641_),
    .o1(_00642_));
 b15nand02aq1n12x5 _26542_ (.a(_00633_),
    .b(_00642_),
    .o1(_00643_));
 b15nand02ah1n16x5 _26543_ (.a(net733),
    .b(net722),
    .o1(_00644_));
 b15orn002aq1n08x5 _26544_ (.a(net733),
    .b(net722),
    .o(_00645_));
 b15oai022an1n08x5 _26545_ (.a(_00644_),
    .b(_16928_),
    .c(_16929_),
    .d(_00645_),
    .o1(_00646_));
 b15aoi122ah1n06x5 _26546_ (.a(net730),
    .b(_16214_),
    .c(_16213_),
    .d(_00646_),
    .e(net716),
    .o1(_00647_));
 b15norp03ar1n03x5 _26547_ (.a(_16203_),
    .b(_17031_),
    .c(_17224_),
    .o1(_00648_));
 b15aoai13al1n06x5 _26548_ (.a(_00648_),
    .b(_16278_),
    .c(_16305_),
    .d(_16221_),
    .o1(_00649_));
 b15nandp2ar1n12x5 _26549_ (.a(_16248_),
    .b(_17008_),
    .o1(_00650_));
 b15aoi013an1n06x5 _26550_ (.a(_00647_),
    .b(_00649_),
    .c(_00650_),
    .d(net729),
    .o1(_00651_));
 b15aoi012al1n02x5 _26551_ (.a(net738),
    .b(_16321_),
    .c(_16997_),
    .o1(_00652_));
 b15nanb02al1n12x5 _26552_ (.a(net729),
    .b(net719),
    .out0(_00653_));
 b15oai022ar1n02x5 _26553_ (.a(net728),
    .b(_16235_),
    .c(_16206_),
    .d(_00653_),
    .o1(_00654_));
 b15aoi022an1n02x5 _26554_ (.a(_16295_),
    .b(_16932_),
    .c(_00654_),
    .d(_16278_),
    .o1(_00655_));
 b15oai022aq1n06x5 _26555_ (.a(_16226_),
    .b(_16389_),
    .c(_00652_),
    .d(_00655_),
    .o1(_00656_));
 b15oaoi13al1n04x5 _26556_ (.a(net734),
    .b(_16960_),
    .c(_16231_),
    .d(net729),
    .o1(_00657_));
 b15aoi022as1n12x5 _26557_ (.a(net738),
    .b(_00651_),
    .c(_00656_),
    .d(_00657_),
    .o1(_00658_));
 b15nanb02ah1n08x5 _26558_ (.a(net722),
    .b(net730),
    .out0(_00659_));
 b15oai022as1n06x5 _26559_ (.a(_16280_),
    .b(_16952_),
    .c(_00659_),
    .d(_16235_),
    .o1(_00660_));
 b15nand02an1n02x5 _26560_ (.a(net728),
    .b(_00660_),
    .o1(_00661_));
 b15nor003ar1n06x5 _26561_ (.a(net732),
    .b(net723),
    .c(_16951_),
    .o1(_00662_));
 b15norp02as1n02x5 _26562_ (.a(_16226_),
    .b(_16396_),
    .o1(_00663_));
 b15oai012as1n02x5 _26563_ (.a(net742),
    .b(_00662_),
    .c(_00663_),
    .o1(_00664_));
 b15aoi012aq1n06x5 _26564_ (.a(_16388_),
    .b(_00661_),
    .c(_00664_),
    .o1(_00665_));
 b15nand04an1n06x5 _26565_ (.a(_16248_),
    .b(net728),
    .c(_16960_),
    .d(_00660_),
    .o1(_00666_));
 b15aoai13an1n03x5 _26566_ (.a(_16957_),
    .b(_17008_),
    .c(_16965_),
    .d(_16332_),
    .o1(_00667_));
 b15aoi012as1n02x5 _26567_ (.a(_17044_),
    .b(_16932_),
    .c(_16193_),
    .o1(_00668_));
 b15oai112aq1n12x5 _26568_ (.a(_00666_),
    .b(_00667_),
    .c(_16972_),
    .d(_00668_),
    .o1(_00669_));
 b15nand04an1n06x5 _26569_ (.a(net722),
    .b(_17055_),
    .c(_16194_),
    .d(_16960_),
    .o1(_00670_));
 b15nand02ar1n04x5 _26570_ (.a(net722),
    .b(_16305_),
    .o1(_00671_));
 b15nand04aq1n16x5 _26571_ (.a(net733),
    .b(net726),
    .c(net717),
    .d(_17230_),
    .o1(_00672_));
 b15oaoi13al1n04x5 _26572_ (.a(net729),
    .b(_00670_),
    .c(_00671_),
    .d(_00672_),
    .o1(_00673_));
 b15aobi12al1n06x5 _26573_ (.a(_00644_),
    .b(_16418_),
    .c(_16342_),
    .out0(_00674_));
 b15nandp2ah1n05x5 _26574_ (.a(_16181_),
    .b(_16347_),
    .o1(_00675_));
 b15nandp2aq1n04x5 _26575_ (.a(_17041_),
    .b(_16927_),
    .o1(_00676_));
 b15oa0022al1n04x5 _26576_ (.a(_16970_),
    .b(_16928_),
    .c(_16929_),
    .d(net740),
    .o(_00677_));
 b15orn002ah1n04x5 _26577_ (.a(_16305_),
    .b(_00659_),
    .o(_00678_));
 b15oai222as1n16x5 _26578_ (.a(_00674_),
    .b(_00675_),
    .c(_00676_),
    .d(_00677_),
    .e(_00672_),
    .f(_00678_),
    .o1(_00679_));
 b15nona22al1n04x5 _26579_ (.a(net729),
    .b(net717),
    .c(net733),
    .out0(_00680_));
 b15nona22an1n04x5 _26580_ (.a(net742),
    .b(net720),
    .c(net737),
    .out0(_00681_));
 b15nanb03ah1n04x5 _26581_ (.a(net737),
    .b(net742),
    .c(net720),
    .out0(_00682_));
 b15aoi112ar1n08x5 _26582_ (.a(_16310_),
    .b(_00680_),
    .c(_00681_),
    .d(_00682_),
    .o1(_00683_));
 b15nor004as1n08x5 _26583_ (.a(_16237_),
    .b(_16280_),
    .c(_16995_),
    .d(_17015_),
    .o1(_00684_));
 b15nand04as1n02x5 _26584_ (.a(net733),
    .b(net722),
    .c(net726),
    .d(net720),
    .o1(_00685_));
 b15xor002as1n02x5 _26585_ (.a(net737),
    .b(net726),
    .out0(_00686_));
 b15oai013al1n08x5 _26586_ (.a(_00685_),
    .b(_00686_),
    .c(net720),
    .d(_00645_),
    .o1(_00687_));
 b15norp02an1n04x5 _26587_ (.a(net717),
    .b(_16361_),
    .o1(_00688_));
 b15aoi112as1n08x5 _26588_ (.a(_00683_),
    .b(_00684_),
    .c(_00687_),
    .d(_00688_),
    .o1(_00689_));
 b15nor004ah1n03x5 _26589_ (.a(net733),
    .b(_17203_),
    .c(_16936_),
    .d(_16928_),
    .o1(_00690_));
 b15aoai13aq1n08x5 _26590_ (.a(net729),
    .b(_00690_),
    .c(_16333_),
    .d(_16213_),
    .o1(_00691_));
 b15nona23ar1n32x5 _26591_ (.a(_00673_),
    .b(_00679_),
    .c(_00689_),
    .d(_00691_),
    .out0(_00692_));
 b15nand02ar1n02x5 _26592_ (.a(net738),
    .b(net719),
    .o1(_00693_));
 b15oaoi13aq1n03x5 _26593_ (.a(_00693_),
    .b(net734),
    .c(net730),
    .d(_17258_),
    .o1(_00694_));
 b15and002al1n02x5 _26594_ (.a(_16291_),
    .b(_16292_),
    .o(_00695_));
 b15orn002ar1n04x5 _26595_ (.a(net723),
    .b(net716),
    .o(_00696_));
 b15oai022an1n12x5 _26596_ (.a(_16193_),
    .b(_17247_),
    .c(_00696_),
    .d(_16361_),
    .o1(_00697_));
 b15aoai13al1n08x5 _26597_ (.a(_00694_),
    .b(_00695_),
    .c(net728),
    .d(_00697_),
    .o1(_00698_));
 b15nona23an1n02x5 _26598_ (.a(net725),
    .b(net716),
    .c(net740),
    .d(net723),
    .out0(_00699_));
 b15oaoi13ar1n04x5 _26599_ (.a(_00653_),
    .b(_00699_),
    .c(_16966_),
    .d(_16206_),
    .o1(_00700_));
 b15aoai13as1n06x5 _26600_ (.a(net734),
    .b(_00700_),
    .c(_16343_),
    .d(_16347_),
    .o1(_00701_));
 b15norp02al1n02x5 _26601_ (.a(net739),
    .b(_16383_),
    .o1(_00702_));
 b15aoai13ah1n04x5 _26602_ (.a(_16316_),
    .b(_00702_),
    .c(_00662_),
    .d(net739),
    .o1(_00703_));
 b15nand04al1n12x5 _26603_ (.a(_16404_),
    .b(_00698_),
    .c(_00701_),
    .d(_00703_),
    .o1(_00704_));
 b15nor004ah1n12x5 _26604_ (.a(_00665_),
    .b(_00669_),
    .c(_00692_),
    .d(_00704_),
    .o1(_00705_));
 b15nona23as1n32x5 _26605_ (.a(_00625_),
    .b(_00643_),
    .c(_00658_),
    .d(_00705_),
    .out0(_00706_));
 b15nor003an1n02x5 _26606_ (.a(_16713_),
    .b(_17367_),
    .c(_17371_),
    .o1(_00707_));
 b15nona23ah1n32x5 _26607_ (.a(\us31.a[4] ),
    .b(\us31.a[6] ),
    .c(\us31.a[7] ),
    .d(\us31.a[5] ),
    .out0(_00708_));
 b15oai012aq1n04x5 _26608_ (.a(_00708_),
    .b(_16835_),
    .c(_16867_),
    .o1(_00709_));
 b15aoi013aq1n06x5 _26609_ (.a(_00707_),
    .b(_00709_),
    .c(_16780_),
    .d(_16892_),
    .o1(_00710_));
 b15bfn000ah1n02x5 input20 (.a(key[117]),
    .o(net20));
 b15nandp3al1n03x5 _26611_ (.a(_16830_),
    .b(_16831_),
    .c(_17375_),
    .o1(_00712_));
 b15oaoi13as1n08x5 _26612_ (.a(_16770_),
    .b(_00712_),
    .c(_17390_),
    .d(_16748_),
    .o1(_00713_));
 b15nonb02an1n12x5 _26613_ (.a(net758),
    .b(net750),
    .out0(_00714_));
 b15nand03ah1n03x5 _26614_ (.a(_16746_),
    .b(_16896_),
    .c(_00714_),
    .o1(_00715_));
 b15bfn000an1n02x5 input19 (.a(key[116]),
    .o(net19));
 b15nand03al1n03x5 _26616_ (.a(_16861_),
    .b(_16852_),
    .c(_17337_),
    .o1(_00717_));
 b15oai112aq1n08x5 _26617_ (.a(_00715_),
    .b(_00717_),
    .c(_16786_),
    .d(_16899_),
    .o1(_00718_));
 b15nanb02aq1n24x5 _26618_ (.a(net760),
    .b(net756),
    .out0(_00719_));
 b15oai022ah1n06x5 _26619_ (.a(net754),
    .b(_16748_),
    .c(_00719_),
    .d(_16832_),
    .o1(_00720_));
 b15aoi112as1n08x5 _26620_ (.a(_00713_),
    .b(_00718_),
    .c(_16860_),
    .d(_00720_),
    .o1(_00721_));
 b15nandp2al1n08x5 _26621_ (.a(_16770_),
    .b(_16741_),
    .o1(_00722_));
 b15norp02al1n04x5 _26622_ (.a(_16896_),
    .b(_16782_),
    .o1(_00723_));
 b15nand03as1n04x5 _26623_ (.a(net751),
    .b(_16907_),
    .c(_16844_),
    .o1(_00724_));
 b15nandp2al1n04x5 _26624_ (.a(_16907_),
    .b(_00714_),
    .o1(_00725_));
 b15nonb02ah1n12x5 _26625_ (.a(net753),
    .b(net756),
    .out0(_00726_));
 b15aoi022an1n06x5 _26626_ (.a(net754),
    .b(_16782_),
    .c(_00726_),
    .d(_16710_),
    .o1(_00727_));
 b15oai222aq1n16x5 _26627_ (.a(_00722_),
    .b(_16903_),
    .c(_00723_),
    .d(_00724_),
    .e(_00725_),
    .f(_00727_),
    .o1(_00728_));
 b15aoi013ah1n06x5 _26628_ (.a(_00728_),
    .b(_16788_),
    .c(_16758_),
    .d(_16798_),
    .o1(_00729_));
 b15nandp2aq1n24x5 _26629_ (.a(_16731_),
    .b(_16782_),
    .o1(_00730_));
 b15oaoi13ar1n04x5 _26630_ (.a(_16839_),
    .b(_00730_),
    .c(net761),
    .d(_17314_),
    .o1(_00731_));
 b15nand02ar1n02x5 _26631_ (.a(_16780_),
    .b(_16861_),
    .o1(_00732_));
 b15oai022as1n02x5 _26632_ (.a(_16832_),
    .b(_00732_),
    .c(_17355_),
    .d(_16761_),
    .o1(_00733_));
 b15oai022ah1n06x5 _26633_ (.a(_16693_),
    .b(_00730_),
    .c(_16832_),
    .d(_17390_),
    .o1(_00734_));
 b15nonb02as1n16x5 _26634_ (.a(net761),
    .b(net758),
    .out0(_00735_));
 b15aoi112aq1n08x5 _26635_ (.a(_00731_),
    .b(_00733_),
    .c(_00734_),
    .d(_00735_),
    .o1(_00736_));
 b15nand04as1n08x5 _26636_ (.a(_00710_),
    .b(_00721_),
    .c(_00729_),
    .d(_00736_),
    .o1(_00737_));
 b15nonb02ar1n06x5 _26637_ (.a(net756),
    .b(net753),
    .out0(_00738_));
 b15nonb02aq1n04x5 _26638_ (.a(net750),
    .b(net760),
    .out0(_00739_));
 b15nona23ah1n02x5 _26639_ (.a(_00726_),
    .b(_00738_),
    .c(_00739_),
    .d(_16710_),
    .out0(_00740_));
 b15oa0022ar1n02x5 _26640_ (.a(net756),
    .b(_17285_),
    .c(_16728_),
    .d(_16849_),
    .o(_00741_));
 b15nand02ar1n02x5 _26641_ (.a(net760),
    .b(_16726_),
    .o1(_00742_));
 b15oai112an1n06x5 _26642_ (.a(_17319_),
    .b(_00740_),
    .c(_00741_),
    .d(_00742_),
    .o1(_00743_));
 b15qgbbf1an1n05x5 input18 (.a(key[115]),
    .o(net18));
 b15norp02ar1n08x5 _26644_ (.a(net767),
    .b(_16849_),
    .o1(_00745_));
 b15oai022as1n02x5 _26645_ (.a(net756),
    .b(_17389_),
    .c(_16850_),
    .d(_00719_),
    .o1(_00746_));
 b15aoai13aq1n06x5 _26646_ (.a(net757),
    .b(_00743_),
    .c(_00745_),
    .d(_00746_),
    .o1(_00747_));
 b15aoi013al1n03x5 _26647_ (.a(net760),
    .b(_17288_),
    .c(_17369_),
    .d(_00726_),
    .o1(_00748_));
 b15nano22ar1n02x5 _26648_ (.a(net757),
    .b(net744),
    .c(net767),
    .out0(_00749_));
 b15oai112ah1n04x5 _26649_ (.a(net750),
    .b(_00726_),
    .c(_00749_),
    .d(_17369_),
    .o1(_00750_));
 b15nanb02an1n08x5 _26650_ (.a(net753),
    .b(net744),
    .out0(_00751_));
 b15nonb02al1n12x5 _26651_ (.a(net748),
    .b(net751),
    .out0(_00752_));
 b15aoi022ah1n08x5 _26652_ (.a(_16798_),
    .b(_16820_),
    .c(_16844_),
    .d(_00752_),
    .o1(_00753_));
 b15oaoi13an1n08x5 _26653_ (.a(_00748_),
    .b(_00750_),
    .c(_00751_),
    .d(_00753_),
    .o1(_00754_));
 b15xor002as1n02x5 _26654_ (.a(_16774_),
    .b(net753),
    .out0(_00755_));
 b15bfn000ar1n02x5 input17 (.a(key[114]),
    .o(net17));
 b15nano23aq1n03x5 _26656_ (.a(net767),
    .b(_00755_),
    .c(net750),
    .d(_16850_),
    .out0(_00757_));
 b15oaoi13al1n04x5 _26657_ (.a(net767),
    .b(_17355_),
    .c(_16832_),
    .d(net757),
    .o1(_00758_));
 b15oaoi13ah1n04x5 _26658_ (.a(_00754_),
    .b(_16750_),
    .c(_00757_),
    .d(_00758_),
    .o1(_00759_));
 b15nonb03ar1n12x5 _26659_ (.a(net753),
    .b(\us31.a[2] ),
    .c(net762),
    .out0(_00760_));
 b15oai012ar1n02x5 _26660_ (.a(_00760_),
    .b(_00752_),
    .c(_16820_),
    .o1(_00761_));
 b15nandp2an1n05x5 _26661_ (.a(_16881_),
    .b(_16831_),
    .o1(_00762_));
 b15oaoi13an1n03x5 _26662_ (.a(net744),
    .b(_00761_),
    .c(_00762_),
    .d(_17287_),
    .o1(_00763_));
 b15oai112al1n02x5 _26663_ (.a(_16702_),
    .b(_16708_),
    .c(_16907_),
    .d(_16783_),
    .o1(_00764_));
 b15oai013as1n02x5 _26664_ (.a(_00764_),
    .b(_17373_),
    .c(_17367_),
    .d(_16774_),
    .o1(_00765_));
 b15and003ah1n02x5 _26665_ (.a(net759),
    .b(net753),
    .c(\us31.a[7] ),
    .o(_00766_));
 b15nor003as1n03x5 _26666_ (.a(net759),
    .b(net753),
    .c(\us31.a[7] ),
    .o1(_00767_));
 b15oai012al1n12x5 _26667_ (.a(_17298_),
    .b(_00766_),
    .c(_00767_),
    .o1(_00768_));
 b15oai122ar1n16x5 _26668_ (.a(_00768_),
    .b(_17373_),
    .c(_16898_),
    .d(_17339_),
    .e(_16811_),
    .o1(_00769_));
 b15aoi112ah1n04x5 _26669_ (.a(_00763_),
    .b(_00765_),
    .c(_00769_),
    .d(net760),
    .o1(_00770_));
 b15oai112aq1n16x5 _26670_ (.a(_00747_),
    .b(_00759_),
    .c(_16741_),
    .d(_00770_),
    .o1(_00771_));
 b15nanb02aq1n16x5 _26671_ (.a(net748),
    .b(\us31.a[7] ),
    .out0(_00772_));
 b15nor002an1n06x5 _26672_ (.a(\us31.a[4] ),
    .b(_00772_),
    .o1(_00773_));
 b15aoi022ar1n04x5 _26673_ (.a(net762),
    .b(_16905_),
    .c(_00739_),
    .d(_00773_),
    .o1(_00774_));
 b15oa0022an1n02x5 _26674_ (.a(_16764_),
    .b(_16835_),
    .c(_00774_),
    .d(_16856_),
    .o(_00775_));
 b15oai012as1n03x5 _26675_ (.a(_00730_),
    .b(_16748_),
    .c(net761),
    .o1(_00776_));
 b15oai012ar1n06x5 _26676_ (.a(_16743_),
    .b(_17314_),
    .c(_16741_),
    .o1(_00777_));
 b15aoi022an1n12x5 _26677_ (.a(_16861_),
    .b(_00776_),
    .c(_00777_),
    .d(_00735_),
    .o1(_00778_));
 b15aoi022aq1n12x5 _26678_ (.a(_16710_),
    .b(_00726_),
    .c(_00738_),
    .d(_16726_),
    .o1(_00779_));
 b15oai013ah1n03x5 _26679_ (.a(_16693_),
    .b(net751),
    .c(_17317_),
    .d(_00779_),
    .o1(_00780_));
 b15nanb02al1n16x5 _26680_ (.a(net759),
    .b(net763),
    .out0(_00781_));
 b15bfn000as1n02x5 input16 (.a(key[113]),
    .o(net16));
 b15nand02an1n04x5 _26682_ (.a(net759),
    .b(\us31.a[7] ),
    .o1(_00783_));
 b15oai022ah1n04x5 _26683_ (.a(net745),
    .b(_00781_),
    .c(_00783_),
    .d(net763),
    .o1(_00784_));
 b15and003ar1n03x5 _26684_ (.a(\us31.a[4] ),
    .b(net748),
    .c(_16768_),
    .o(_00785_));
 b15aoi012ar1n08x5 _26685_ (.a(_00780_),
    .b(_00784_),
    .c(_00785_),
    .o1(_00786_));
 b15aoi022as1n06x5 _26686_ (.a(net765),
    .b(_00775_),
    .c(_00778_),
    .d(_00786_),
    .o1(_00787_));
 b15bfn000ar1n02x5 input15 (.a(key[112]),
    .o(net15));
 b15nona22ah1n12x5 _26688_ (.a(net753),
    .b(net744),
    .c(net747),
    .out0(_00789_));
 b15oai022ar1n02x5 _26689_ (.a(net748),
    .b(_17297_),
    .c(_00789_),
    .d(_16855_),
    .o1(_00790_));
 b15aoi012aq1n02x5 _26690_ (.a(_16741_),
    .b(_00714_),
    .c(_00790_),
    .o1(_00791_));
 b15nandp2aq1n05x5 _26691_ (.a(_16770_),
    .b(_16783_),
    .o1(_00792_));
 b15oa0022an1n02x5 _26692_ (.a(_00730_),
    .b(_00792_),
    .c(_00781_),
    .d(_17371_),
    .o(_00793_));
 b15nanb02aq1n12x5 _26693_ (.a(\us31.a[7] ),
    .b(net748),
    .out0(_00794_));
 b15oai022an1n08x5 _26694_ (.a(net759),
    .b(_00772_),
    .c(_17317_),
    .d(_00794_),
    .o1(_00795_));
 b15aoi013al1n03x5 _26695_ (.a(net755),
    .b(_16702_),
    .c(_00795_),
    .d(_16693_),
    .o1(_00796_));
 b15nor003ar1n02x5 _26696_ (.a(net762),
    .b(\us31.a[4] ),
    .c(_00772_),
    .o1(_00797_));
 b15oai112as1n04x5 _26697_ (.a(net751),
    .b(_16860_),
    .c(_00797_),
    .d(_16827_),
    .o1(_00798_));
 b15aoi013ah1n04x5 _26698_ (.a(_00791_),
    .b(_00793_),
    .c(_00796_),
    .d(_00798_),
    .o1(_00799_));
 b15inv020ar1n05x5 _26699_ (.a(net744),
    .o1(_00800_));
 b15and003ar1n08x5 _26700_ (.a(net753),
    .b(_00800_),
    .c(_16881_),
    .o(_00801_));
 b15norp02ah1n04x5 _26701_ (.a(net757),
    .b(net751),
    .o1(_00802_));
 b15nand03aq1n02x5 _26702_ (.a(_16746_),
    .b(_00801_),
    .c(_00802_),
    .o1(_00803_));
 b15norp03al1n02x5 _26703_ (.a(_16839_),
    .b(_16852_),
    .c(_16793_),
    .o1(_00804_));
 b15aoi013ar1n02x5 _26704_ (.a(_00804_),
    .b(_16894_),
    .c(_16758_),
    .d(_16798_),
    .o1(_00805_));
 b15nanb02ar1n02x5 _26705_ (.a(_16728_),
    .b(_17382_),
    .out0(_00806_));
 b15oai112as1n02x5 _26706_ (.a(_00803_),
    .b(_00805_),
    .c(_16897_),
    .d(_00806_),
    .o1(_00807_));
 b15and003ar1n02x5 _26707_ (.a(_16746_),
    .b(_16782_),
    .c(_00802_),
    .o(_00808_));
 b15aoai13ah1n03x5 _26708_ (.a(net765),
    .b(_00808_),
    .c(_16750_),
    .d(_17354_),
    .o1(_00809_));
 b15nano23aq1n02x5 _26709_ (.a(net753),
    .b(net748),
    .c(net760),
    .d(net750),
    .out0(_00810_));
 b15nanb02an1n03x5 _26710_ (.a(net748),
    .b(net750),
    .out0(_00811_));
 b15oab012al1n04x5 _26711_ (.a(_00810_),
    .b(_00811_),
    .c(net753),
    .out0(_00812_));
 b15nor004ar1n06x5 _26712_ (.a(net744),
    .b(_16713_),
    .c(_16836_),
    .d(_00812_),
    .o1(_00813_));
 b15nor004ah1n03x5 _26713_ (.a(net750),
    .b(_16850_),
    .c(_16761_),
    .d(_00755_),
    .o1(_00814_));
 b15norp03an1n12x5 _26714_ (.a(_16849_),
    .b(_16850_),
    .c(_16856_),
    .o1(_00815_));
 b15aoi112aq1n06x5 _26715_ (.a(_00813_),
    .b(_00814_),
    .c(_00815_),
    .d(_16907_),
    .o1(_00816_));
 b15nona23an1n12x5 _26716_ (.a(_00799_),
    .b(_00807_),
    .c(_00809_),
    .d(_00816_),
    .out0(_00817_));
 b15nor004as1n12x5 _26717_ (.a(_00737_),
    .b(_00771_),
    .c(_00787_),
    .d(_00817_),
    .o1(_00818_));
 b15xor002ar1n08x5 _26718_ (.a(_17281_),
    .b(_00818_),
    .out0(_00819_));
 b15qgbxo2an1n05x5 _26719_ (.a(_00706_),
    .b(_00819_),
    .out0(_00820_));
 b15xor002aq1n08x5 _26720_ (.a(_00619_),
    .b(_00820_),
    .out0(_00821_));
 b15mdn022an1n16x5 _26721_ (.a(_17531_),
    .b(_00821_),
    .o1(_00822_),
    .sa(net540));
 b15xor002as1n16x5 _26722_ (.a(\u0.w[2][2] ),
    .b(_00822_),
    .out0(_00115_));
 b15orn002aq1n12x5 _26723_ (.a(net615),
    .b(net611),
    .o(_00823_));
 b15nand04an1n06x5 _26724_ (.a(_16475_),
    .b(_16605_),
    .c(_00823_),
    .d(_17165_),
    .o1(_00824_));
 b15aoai13ar1n04x5 _26725_ (.a(net614),
    .b(net613),
    .c(_16475_),
    .d(_16605_),
    .o1(_00825_));
 b15aoi022al1n08x5 _26726_ (.a(_16482_),
    .b(_00824_),
    .c(_00825_),
    .d(_16558_),
    .o1(_00826_));
 b15nor003an1n12x5 _26727_ (.a(_16616_),
    .b(_17175_),
    .c(_16594_),
    .o1(_00827_));
 b15ao0022al1n03x5 _26728_ (.a(net600),
    .b(_16510_),
    .c(_00827_),
    .d(net606),
    .o(_00828_));
 b15nand02aq1n04x5 _26729_ (.a(_16659_),
    .b(_16575_),
    .o1(_00829_));
 b15aoai13as1n08x5 _26730_ (.a(net609),
    .b(_00826_),
    .c(_00828_),
    .d(_00829_),
    .o1(_00830_));
 b15aoi122ar1n06x5 _26731_ (.a(net619),
    .b(_16504_),
    .c(_16571_),
    .d(_16672_),
    .e(_16508_),
    .o1(_00831_));
 b15aob012as1n02x5 _26732_ (.a(net620),
    .b(_16539_),
    .c(_17545_),
    .out0(_00832_));
 b15nona22ar1n04x5 _26733_ (.a(net607),
    .b(net616),
    .c(net601),
    .out0(_00833_));
 b15nanb02ah1n03x5 _26734_ (.a(net601),
    .b(net607),
    .out0(_00834_));
 b15and003ar1n02x5 _26735_ (.a(net604),
    .b(_00833_),
    .c(_00834_),
    .o(_00835_));
 b15aoi012al1n04x5 _26736_ (.a(_00835_),
    .b(_17093_),
    .c(_17099_),
    .o1(_00836_));
 b15aoi013al1n08x5 _26737_ (.a(_00832_),
    .b(_00836_),
    .c(_16460_),
    .d(\us13.a[7] ),
    .o1(_00837_));
 b15oai013ah1n06x5 _26738_ (.a(_00830_),
    .b(_00831_),
    .c(_00837_),
    .d(net610),
    .o1(_00838_));
 b15nor004ah1n08x5 _26739_ (.a(net610),
    .b(_16453_),
    .c(_16667_),
    .d(_16673_),
    .o1(_00839_));
 b15aoai13ah1n02x5 _26740_ (.a(net612),
    .b(_00839_),
    .c(_17146_),
    .d(net608),
    .o1(_00840_));
 b15norp03ar1n02x5 _26741_ (.a(net608),
    .b(_17116_),
    .c(_17088_),
    .o1(_00841_));
 b15oai012aq1n02x5 _26742_ (.a(_16575_),
    .b(_16652_),
    .c(_16558_),
    .o1(_00842_));
 b15aoi013aq1n02x5 _26743_ (.a(_00841_),
    .b(_00842_),
    .c(_16526_),
    .d(net608),
    .o1(_00843_));
 b15and002ar1n02x5 _26744_ (.a(net597),
    .b(net608),
    .o(_00844_));
 b15aoi112ar1n02x5 _26745_ (.a(net597),
    .b(net608),
    .c(net611),
    .d(net616),
    .o1(_00845_));
 b15oai112as1n02x5 _26746_ (.a(_16597_),
    .b(_16517_),
    .c(_00844_),
    .d(_00845_),
    .o1(_00846_));
 b15nonb02ah1n06x5 _26747_ (.a(net616),
    .b(net608),
    .out0(_00847_));
 b15norp03aq1n02x5 _26748_ (.a(_16492_),
    .b(_17190_),
    .c(_00847_),
    .o1(_00848_));
 b15aoi112aq1n04x5 _26749_ (.a(_00846_),
    .b(_00848_),
    .c(_16682_),
    .d(_17190_),
    .o1(_00849_));
 b15nand04al1n03x5 _26750_ (.a(net608),
    .b(_16435_),
    .c(_16473_),
    .d(_16475_),
    .o1(_00850_));
 b15nanb02ah1n04x5 _26751_ (.a(net608),
    .b(net616),
    .out0(_00851_));
 b15oaoi13aq1n03x5 _26752_ (.a(net612),
    .b(_00850_),
    .c(_00851_),
    .d(_17116_),
    .o1(_00852_));
 b15nano23ar1n08x5 _26753_ (.a(_00840_),
    .b(_00843_),
    .c(_00849_),
    .d(_00852_),
    .out0(_00853_));
 b15nandp3aq1n02x5 _26754_ (.a(_16456_),
    .b(_16591_),
    .c(_16650_),
    .o1(_00854_));
 b15oai013as1n06x5 _26755_ (.a(_00854_),
    .b(_16626_),
    .c(_16521_),
    .d(_16682_),
    .o1(_00855_));
 b15nandp3ar1n03x5 _26756_ (.a(net611),
    .b(_16439_),
    .c(_17562_),
    .o1(_00856_));
 b15oai013as1n06x5 _26757_ (.a(_00856_),
    .b(_16528_),
    .c(_16479_),
    .d(_16435_),
    .o1(_00857_));
 b15nand02an1n16x5 _26758_ (.a(_16597_),
    .b(_16439_),
    .o1(_00858_));
 b15nandp2ah1n05x5 _26759_ (.a(_16458_),
    .b(_16475_),
    .o1(_00859_));
 b15nano23aq1n12x5 _26760_ (.a(_16640_),
    .b(_00858_),
    .c(_00859_),
    .d(_16456_),
    .out0(_00860_));
 b15and002aq1n04x5 _26761_ (.a(_17151_),
    .b(_00827_),
    .o(_00861_));
 b15nor004ah1n12x5 _26762_ (.a(_00855_),
    .b(_00857_),
    .c(_00860_),
    .d(_00861_),
    .o1(_00862_));
 b15norp03ah1n02x5 _26763_ (.a(net619),
    .b(net611),
    .c(_16680_),
    .o1(_00863_));
 b15nand02ar1n02x5 _26764_ (.a(net619),
    .b(_00823_),
    .o1(_00864_));
 b15aoi012ah1n02x5 _26765_ (.a(_17183_),
    .b(_16582_),
    .c(_00864_),
    .o1(_00865_));
 b15oai012aq1n06x5 _26766_ (.a(net608),
    .b(_00863_),
    .c(_00865_),
    .o1(_00866_));
 b15nandp3ar1n02x5 _26767_ (.a(net620),
    .b(_16504_),
    .c(_17146_),
    .o1(_00867_));
 b15oai012aq1n04x5 _26768_ (.a(_00867_),
    .b(_17125_),
    .c(_16491_),
    .o1(_00868_));
 b15oai022an1n08x5 _26769_ (.a(_16576_),
    .b(_16516_),
    .c(_16528_),
    .d(_17165_),
    .o1(_00869_));
 b15oai012ar1n08x5 _26770_ (.a(_16466_),
    .b(_00868_),
    .c(_00869_),
    .o1(_00870_));
 b15nand04as1n16x5 _26771_ (.a(_00853_),
    .b(_00862_),
    .c(_00866_),
    .d(_00870_),
    .o1(_00871_));
 b15norp02ar1n02x5 _26772_ (.a(\us13.a[2] ),
    .b(_17113_),
    .o1(_00872_));
 b15norp02al1n02x5 _26773_ (.a(net604),
    .b(_16535_),
    .o1(_00873_));
 b15aoai13ar1n02x5 _26774_ (.a(_00872_),
    .b(_00873_),
    .c(_16677_),
    .d(net604),
    .o1(_00874_));
 b15nandp3aq1n02x5 _26775_ (.a(net604),
    .b(\us13.a[7] ),
    .c(net612),
    .o1(_00875_));
 b15oaoi13an1n04x5 _26776_ (.a(_00875_),
    .b(_00833_),
    .c(_16435_),
    .d(_00834_),
    .o1(_00876_));
 b15oaoi13ah1n03x5 _26777_ (.a(_16521_),
    .b(_17176_),
    .c(_16460_),
    .d(_16609_),
    .o1(_00877_));
 b15nano23al1n05x5 _26778_ (.a(_16466_),
    .b(_00874_),
    .c(_00876_),
    .d(_00877_),
    .out0(_00878_));
 b15oai012ar1n02x5 _26779_ (.a(net610),
    .b(_16492_),
    .c(_16528_),
    .o1(_00879_));
 b15aoi012aq1n02x5 _26780_ (.a(_00879_),
    .b(_16571_),
    .c(_16478_),
    .o1(_00880_));
 b15aoi022as1n04x5 _26781_ (.a(net617),
    .b(_17087_),
    .c(_16571_),
    .d(\us13.a[2] ),
    .o1(_00881_));
 b15oaoi13al1n08x5 _26782_ (.a(_00878_),
    .b(_00880_),
    .c(net619),
    .d(_00881_),
    .o1(_00882_));
 b15aoi012ar1n02x5 _26783_ (.a(_16609_),
    .b(_16528_),
    .c(_17091_),
    .o1(_00883_));
 b15aoi013aq1n04x5 _26784_ (.a(_00883_),
    .b(_16650_),
    .c(net614),
    .d(net618),
    .o1(_00884_));
 b15oai222as1n12x5 _26785_ (.a(_16482_),
    .b(_16644_),
    .c(_17578_),
    .d(_16642_),
    .e(_00884_),
    .f(_16524_),
    .o1(_00885_));
 b15nor004ar1n02x5 _26786_ (.a(_16497_),
    .b(_16592_),
    .c(_16438_),
    .d(_16632_),
    .o1(_00886_));
 b15nor003ar1n02x5 _26787_ (.a(_16522_),
    .b(_16453_),
    .c(_17091_),
    .o1(_00887_));
 b15norp02ar1n02x5 _26788_ (.a(_16490_),
    .b(_17113_),
    .o1(_00888_));
 b15aoi112aq1n02x5 _26789_ (.a(_00886_),
    .b(_00887_),
    .c(_00888_),
    .d(_17161_),
    .o1(_00889_));
 b15norp03ar1n02x5 _26790_ (.a(net606),
    .b(_16432_),
    .c(_16524_),
    .o1(_00890_));
 b15aoi012ar1n02x5 _26791_ (.a(_00890_),
    .b(_16518_),
    .c(net606),
    .o1(_00891_));
 b15oai013al1n02x5 _26792_ (.a(_00889_),
    .b(_00891_),
    .c(_16609_),
    .d(net604),
    .o1(_00892_));
 b15norp02ar1n03x5 _26793_ (.a(net598),
    .b(_16498_),
    .o1(_00893_));
 b15nano22ar1n05x5 _26794_ (.a(net617),
    .b(net613),
    .c(net599),
    .out0(_00894_));
 b15oaoi13ar1n02x5 _26795_ (.a(_00894_),
    .b(net599),
    .c(_16504_),
    .d(_16613_),
    .o1(_00895_));
 b15norp02aq1n02x5 _26796_ (.a(_16673_),
    .b(_00895_),
    .o1(_00896_));
 b15aoai13ar1n08x5 _26797_ (.a(_00893_),
    .b(_00896_),
    .c(_16475_),
    .d(_16511_),
    .o1(_00897_));
 b15oai022al1n02x5 _26798_ (.a(_16576_),
    .b(_16479_),
    .c(_17183_),
    .d(_16632_),
    .o1(_00898_));
 b15nandp3ar1n02x5 _26799_ (.a(_16481_),
    .b(_16577_),
    .c(_16652_),
    .o1(_00899_));
 b15nandp2al1n08x5 _26800_ (.a(_16473_),
    .b(_16517_),
    .o1(_00900_));
 b15oai012ar1n04x5 _26801_ (.a(_00899_),
    .b(_00900_),
    .c(_16652_),
    .o1(_00901_));
 b15nor002al1n04x5 _26802_ (.a(_16558_),
    .b(net608),
    .o1(_00902_));
 b15aoi022as1n04x5 _26803_ (.a(net615),
    .b(_00898_),
    .c(_00901_),
    .d(_00902_),
    .o1(_00903_));
 b15nona23aq1n05x5 _26804_ (.a(_00885_),
    .b(_00892_),
    .c(_00897_),
    .d(_00903_),
    .out0(_00904_));
 b15nor004as1n12x5 _26805_ (.a(_00838_),
    .b(_00871_),
    .c(_00882_),
    .d(_00904_),
    .o1(_00905_));
 b15aoai13ar1n02x5 _26806_ (.a(net742),
    .b(_16291_),
    .c(_16293_),
    .d(net733),
    .o1(_00906_));
 b15oaoi13an1n02x5 _26807_ (.a(net719),
    .b(_00906_),
    .c(_16967_),
    .d(net733),
    .o1(_00907_));
 b15norp03an1n02x5 _26808_ (.a(_16291_),
    .b(_16293_),
    .c(_17017_),
    .o1(_00908_));
 b15oai112ah1n04x5 _26809_ (.a(net723),
    .b(_16401_),
    .c(_00907_),
    .d(_00908_),
    .o1(_00909_));
 b15aoi022ar1n02x5 _26810_ (.a(_16229_),
    .b(_16189_),
    .c(_16935_),
    .d(_16223_),
    .o1(_00910_));
 b15orn003ar1n02x5 _26811_ (.a(net726),
    .b(_16379_),
    .c(_00910_),
    .o(_00911_));
 b15nonb02ah1n06x5 _26812_ (.a(net725),
    .b(net740),
    .out0(_00912_));
 b15oai112al1n08x5 _26813_ (.a(_16223_),
    .b(_16274_),
    .c(_16333_),
    .d(_00912_),
    .o1(_00913_));
 b15and002ar1n02x5 _26814_ (.a(_16406_),
    .b(_00913_),
    .o(_00914_));
 b15aoi022al1n02x5 _26815_ (.a(_16214_),
    .b(_16321_),
    .c(_16977_),
    .d(_17224_),
    .o1(_00915_));
 b15oai112aq1n08x5 _26816_ (.a(_00911_),
    .b(_00914_),
    .c(net737),
    .d(_00915_),
    .o1(_00916_));
 b15aoi012as1n02x5 _26817_ (.a(_17008_),
    .b(_16977_),
    .c(_17015_),
    .o1(_00917_));
 b15aoi012aq1n02x5 _26818_ (.a(net735),
    .b(_16379_),
    .c(_17008_),
    .o1(_00918_));
 b15oai012ah1n08x5 _26819_ (.a(net731),
    .b(_00917_),
    .c(_00918_),
    .o1(_00919_));
 b15aobi12ah1n08x5 _26820_ (.a(_00909_),
    .b(_00916_),
    .c(_00919_),
    .out0(_00920_));
 b15mdn022as1n02x5 _26821_ (.a(_16206_),
    .b(_16203_),
    .o1(_00921_),
    .sa(_16342_));
 b15aoi022al1n08x5 _26822_ (.a(net716),
    .b(_16289_),
    .c(_00921_),
    .d(net730),
    .o1(_00922_));
 b15oai022al1n12x5 _26823_ (.a(_16206_),
    .b(_16952_),
    .c(_00922_),
    .d(net723),
    .o1(_00923_));
 b15nand03al1n24x5 _26824_ (.a(_16305_),
    .b(_17224_),
    .c(_00923_),
    .o1(_00924_));
 b15oai022ar1n04x5 _26825_ (.a(net741),
    .b(_16233_),
    .c(_16993_),
    .d(net739),
    .o1(_00925_));
 b15aoi022ah1n06x5 _26826_ (.a(_16222_),
    .b(_16213_),
    .c(_16980_),
    .d(_00925_),
    .o1(_00926_));
 b15nonb03ah1n08x5 _26827_ (.a(net720),
    .b(net716),
    .c(net725),
    .out0(_00927_));
 b15nand04as1n02x5 _26828_ (.a(_16248_),
    .b(_00927_),
    .c(_16347_),
    .d(_16966_),
    .o1(_00928_));
 b15aoi022ah1n02x5 _26829_ (.a(net733),
    .b(_17031_),
    .c(_16370_),
    .d(_16405_),
    .o1(_00929_));
 b15nand02as1n06x5 _26830_ (.a(net729),
    .b(net725),
    .o1(_00930_));
 b15oai013ah1n06x5 _26831_ (.a(_00928_),
    .b(_00929_),
    .c(_00930_),
    .d(_17055_),
    .o1(_00931_));
 b15aoai13aq1n08x5 _26832_ (.a(_16340_),
    .b(_16320_),
    .c(_17041_),
    .d(_16970_),
    .o1(_00932_));
 b15mdn022al1n04x5 _26833_ (.a(_16223_),
    .b(_16229_),
    .o1(_00933_),
    .sa(net740));
 b15oai013an1n08x5 _26834_ (.a(_00932_),
    .b(_00933_),
    .c(_16993_),
    .d(_16237_),
    .o1(_00934_));
 b15oai022ah1n02x5 _26835_ (.a(_16206_),
    .b(_16361_),
    .c(_16357_),
    .d(_16203_),
    .o1(_00935_));
 b15nand02an1n03x5 _26836_ (.a(net734),
    .b(_17031_),
    .o1(_00936_));
 b15aoi022an1n04x5 _26837_ (.a(net740),
    .b(_16223_),
    .c(_16229_),
    .d(net734),
    .o1(_00937_));
 b15nandp2as1n04x5 _26838_ (.a(_16224_),
    .b(_16988_),
    .o1(_00938_));
 b15obai22as1n08x5 _26839_ (.a(_00935_),
    .b(_00936_),
    .c(_00937_),
    .d(_00938_),
    .out0(_00939_));
 b15cmbn22al1n02x5 _26840_ (.clk1(_16952_),
    .clk2(_00659_),
    .clkout(_00940_),
    .s(_16283_));
 b15nand03aq1n03x5 _26841_ (.a(_16305_),
    .b(_16291_),
    .c(_16356_),
    .o1(_00941_));
 b15nonb02ah1n02x5 _26842_ (.a(net719),
    .b(net723),
    .out0(_00942_));
 b15nona23an1n04x5 _26843_ (.a(_16353_),
    .b(_00912_),
    .c(_16405_),
    .d(_00942_),
    .out0(_00943_));
 b15oai022an1n08x5 _26844_ (.a(_00940_),
    .b(_00941_),
    .c(_00943_),
    .d(net716),
    .o1(_00944_));
 b15nor004as1n12x5 _26845_ (.a(_00931_),
    .b(_00934_),
    .c(_00939_),
    .d(_00944_),
    .o1(_00945_));
 b15oai022ar1n02x5 _26846_ (.a(net735),
    .b(_16357_),
    .c(_17009_),
    .d(_16337_),
    .o1(_00946_));
 b15aoi012aq1n04x5 _26847_ (.a(_00946_),
    .b(_16333_),
    .c(_16342_),
    .o1(_00947_));
 b15oai112as1n16x5 _26848_ (.a(_00926_),
    .b(_00945_),
    .c(_16958_),
    .d(_00947_),
    .o1(_00948_));
 b15norp03ar1n02x5 _26849_ (.a(net743),
    .b(_16248_),
    .c(_17005_),
    .o1(_00949_));
 b15aoai13ar1n02x5 _26850_ (.a(_16342_),
    .b(_00949_),
    .c(_16325_),
    .d(net743),
    .o1(_00950_));
 b15aoi013ar1n02x5 _26851_ (.a(net732),
    .b(net735),
    .c(_16340_),
    .d(_16960_),
    .o1(_00951_));
 b15and002ar1n02x5 _26852_ (.a(_16332_),
    .b(_17009_),
    .o(_00952_));
 b15aoai13ar1n04x5 _26853_ (.a(\us02.a[1] ),
    .b(_00952_),
    .c(_16315_),
    .d(_16311_),
    .o1(_00953_));
 b15nor002ah1n04x5 _26854_ (.a(net735),
    .b(_16970_),
    .o1(_00954_));
 b15aoi112ar1n03x5 _26855_ (.a(_16226_),
    .b(_17223_),
    .c(_16977_),
    .d(_00954_),
    .o1(_00955_));
 b15ao0022al1n04x5 _26856_ (.a(_00950_),
    .b(_00951_),
    .c(_00953_),
    .d(_00955_),
    .o(_00956_));
 b15oaoi13ar1n02x5 _26857_ (.a(_17225_),
    .b(_16381_),
    .c(_16316_),
    .d(_16321_),
    .o1(_00957_));
 b15oaoi13ar1n02x5 _26858_ (.a(net743),
    .b(net732),
    .c(net736),
    .d(_16416_),
    .o1(_00958_));
 b15orn003ah1n02x5 _26859_ (.a(_16342_),
    .b(_00957_),
    .c(_00958_),
    .o(_00959_));
 b15aoi012al1n04x5 _26860_ (.a(_16283_),
    .b(_17028_),
    .c(_16343_),
    .o1(_00960_));
 b15aoi022an1n06x5 _26861_ (.a(_16342_),
    .b(_00927_),
    .c(_16328_),
    .d(net725),
    .o1(_00961_));
 b15nand02aq1n02x5 _26862_ (.a(net722),
    .b(_17041_),
    .o1(_00962_));
 b15aoi022al1n08x5 _26863_ (.a(_16229_),
    .b(_16289_),
    .c(_16273_),
    .d(_16247_),
    .o1(_00963_));
 b15oai122as1n08x5 _26864_ (.a(_00960_),
    .b(_00961_),
    .c(_00962_),
    .d(_00963_),
    .e(_00645_),
    .o1(_00964_));
 b15orn003al1n02x5 _26865_ (.a(_16226_),
    .b(net718),
    .c(_16929_),
    .o(_00965_));
 b15oaoi13al1n08x5 _26866_ (.a(_16955_),
    .b(_00965_),
    .c(net729),
    .d(_16967_),
    .o1(_00966_));
 b15oai013as1n12x5 _26867_ (.a(_00964_),
    .b(_00966_),
    .c(net740),
    .d(_00621_),
    .o1(_00967_));
 b15nand02al1n03x5 _26868_ (.a(_16405_),
    .b(_16416_),
    .o1(_00968_));
 b15oaoi13ah1n08x5 _26869_ (.a(net730),
    .b(_00968_),
    .c(_16336_),
    .d(_16311_),
    .o1(_00969_));
 b15oai022as1n02x5 _26870_ (.a(_16231_),
    .b(_16361_),
    .c(_16357_),
    .d(_16389_),
    .o1(_00970_));
 b15aoi112ah1n06x5 _26871_ (.a(_17043_),
    .b(_00969_),
    .c(_00970_),
    .d(_16350_),
    .o1(_00971_));
 b15nand04as1n12x5 _26872_ (.a(_00956_),
    .b(_00959_),
    .c(_00967_),
    .d(_00971_),
    .o1(_00972_));
 b15nano23as1n24x5 _26873_ (.a(_00920_),
    .b(_00924_),
    .c(_00948_),
    .d(_00972_),
    .out0(_00973_));
 b15xor002an1n16x5 _26874_ (.a(_00905_),
    .b(_00973_),
    .out0(_00974_));
 b15oaoi13an1n02x5 _26875_ (.a(net879),
    .b(_17616_),
    .c(_16009_),
    .d(net875),
    .o1(_00975_));
 b15oai022al1n02x5 _26876_ (.a(_15993_),
    .b(_16132_),
    .c(_00599_),
    .d(_16040_),
    .o1(_00976_));
 b15aoai13ar1n02x5 _26877_ (.a(net868),
    .b(net874),
    .c(net875),
    .d(net879),
    .o1(_00977_));
 b15nand04ar1n02x5 _26878_ (.a(net870),
    .b(_16008_),
    .c(_17518_),
    .d(_00977_),
    .o1(_00978_));
 b15oai012ar1n02x5 _26879_ (.a(_00978_),
    .b(_17616_),
    .c(net875),
    .o1(_00979_));
 b15oai013aq1n04x5 _26880_ (.a(net882),
    .b(_00975_),
    .c(_00976_),
    .d(_00979_),
    .o1(_00980_));
 b15aoi012an1n02x5 _26881_ (.a(\us20.a[3] ),
    .b(_16045_),
    .c(_17410_),
    .o1(_00981_));
 b15nano22ar1n03x5 _26882_ (.a(net871),
    .b(\us20.a[7] ),
    .c(net878),
    .out0(_00982_));
 b15nor003ah1n02x5 _26883_ (.a(net871),
    .b(\us20.a[7] ),
    .c(net881),
    .o1(_00983_));
 b15oai112ah1n08x5 _26884_ (.a(net867),
    .b(_16092_),
    .c(_00982_),
    .d(_00983_),
    .o1(_00984_));
 b15nand03an1n06x5 _26885_ (.a(_17463_),
    .b(_17420_),
    .c(_00586_),
    .o1(_00985_));
 b15aoai13an1n08x5 _26886_ (.a(_00981_),
    .b(_15959_),
    .c(_00984_),
    .d(_00985_),
    .o1(_00986_));
 b15oai013ar1n04x5 _26887_ (.a(net873),
    .b(_15987_),
    .c(_16021_),
    .d(_17459_),
    .o1(_00987_));
 b15nand03ar1n06x5 _26888_ (.a(net867),
    .b(net866),
    .c(net878),
    .o1(_00988_));
 b15orn003ar1n02x5 _26889_ (.a(net867),
    .b(net866),
    .c(net878),
    .o(_00989_));
 b15aoi112al1n02x5 _26890_ (.a(_16078_),
    .b(_17462_),
    .c(_00988_),
    .d(_00989_),
    .o1(_00990_));
 b15nona22ar1n02x5 _26891_ (.a(net871),
    .b(net884),
    .c(net863),
    .out0(_00991_));
 b15oaoi13as1n02x5 _26892_ (.a(_00991_),
    .b(_00988_),
    .c(_17503_),
    .d(net867),
    .o1(_00992_));
 b15orn003al1n08x5 _26893_ (.a(_00987_),
    .b(_00990_),
    .c(_00992_),
    .o(_00993_));
 b15norp02ar1n03x5 _26894_ (.a(net880),
    .b(_16047_),
    .o1(_00994_));
 b15aoi022aq1n02x5 _26895_ (.a(_15952_),
    .b(_15955_),
    .c(_16008_),
    .d(_16065_),
    .o1(_00995_));
 b15oai112ah1n08x5 _26896_ (.a(_16067_),
    .b(_00994_),
    .c(_00995_),
    .d(_16077_),
    .o1(_00996_));
 b15oai122aq1n08x5 _26897_ (.a(\us20.a[1] ),
    .b(_16018_),
    .c(_16060_),
    .d(_16040_),
    .e(net885),
    .o1(_00997_));
 b15aoai13an1n08x5 _26898_ (.a(_00986_),
    .b(_00993_),
    .c(_00996_),
    .d(_00997_),
    .o1(_00998_));
 b15nor002al1n16x5 _26899_ (.a(net884),
    .b(net872),
    .o1(_00999_));
 b15nano23as1n02x5 _26900_ (.a(net863),
    .b(net865),
    .c(net880),
    .d(net869),
    .out0(_01000_));
 b15oai112ah1n06x5 _26901_ (.a(_00999_),
    .b(_01000_),
    .c(_16088_),
    .d(net877),
    .o1(_01001_));
 b15nonb02an1n16x5 _26902_ (.a(net884),
    .b(net880),
    .out0(_01002_));
 b15oai013ar1n02x5 _26903_ (.a(_01001_),
    .b(_17401_),
    .c(_15993_),
    .d(_01002_),
    .o1(_01003_));
 b15nand04ah1n08x5 _26904_ (.a(_16096_),
    .b(_17457_),
    .c(_15975_),
    .d(_17469_),
    .o1(_01004_));
 b15nona23ar1n12x5 _26905_ (.a(_17479_),
    .b(_16090_),
    .c(_17447_),
    .d(_17454_),
    .out0(_01005_));
 b15oai112aq1n02x5 _26906_ (.a(_01004_),
    .b(_01005_),
    .c(_16066_),
    .d(_17405_),
    .o1(_01006_));
 b15norp02ar1n02x5 _26907_ (.a(_16066_),
    .b(_17432_),
    .o1(_01007_));
 b15aoi012ar1n02x5 _26908_ (.a(_17444_),
    .b(_00614_),
    .c(_01007_),
    .o1(_01008_));
 b15nor002ah1n02x5 _26909_ (.a(_16077_),
    .b(_17414_),
    .o1(_01009_));
 b15norp03aq1n02x5 _26910_ (.a(_16088_),
    .b(net873),
    .c(_17503_),
    .o1(_01010_));
 b15and003ar1n02x5 _26911_ (.a(_16088_),
    .b(net873),
    .c(_17503_),
    .o(_01011_));
 b15oai012aq1n06x5 _26912_ (.a(_01009_),
    .b(_01010_),
    .c(_01011_),
    .o1(_01012_));
 b15nona23aq1n05x5 _26913_ (.a(_01003_),
    .b(_01006_),
    .c(_01008_),
    .d(_01012_),
    .out0(_01013_));
 b15nor002an1n08x5 _26914_ (.a(_16078_),
    .b(_15993_),
    .o1(_01014_));
 b15oaoi13ar1n02x5 _26915_ (.a(net882),
    .b(_16000_),
    .c(_16137_),
    .d(net879),
    .o1(_01015_));
 b15oai012ar1n02x5 _26916_ (.a(_17509_),
    .b(_01014_),
    .c(_01015_),
    .o1(_01016_));
 b15norp02ar1n02x5 _26917_ (.a(_16040_),
    .b(_00999_),
    .o1(_01017_));
 b15aoi012ar1n02x5 _26918_ (.a(_01017_),
    .b(_00999_),
    .c(_16086_),
    .o1(_01018_));
 b15oai012an1n04x5 _26919_ (.a(_01016_),
    .b(_01018_),
    .c(_16018_),
    .o1(_01019_));
 b15nano23ar1n06x5 _26920_ (.a(_00980_),
    .b(_00998_),
    .c(_01013_),
    .d(_01019_),
    .out0(_01020_));
 b15oai012ar1n02x5 _26921_ (.a(_16011_),
    .b(_16058_),
    .c(_17446_),
    .o1(_01021_));
 b15oai112al1n02x5 _26922_ (.a(_15959_),
    .b(_17432_),
    .c(_17446_),
    .d(net879),
    .o1(_01022_));
 b15oai112an1n02x5 _26923_ (.a(net882),
    .b(_15995_),
    .c(_17518_),
    .d(_16058_),
    .o1(_01023_));
 b15aoi012as1n02x5 _26924_ (.a(_01021_),
    .b(_01022_),
    .c(_01023_),
    .o1(_01024_));
 b15nanb03aq1n12x5 _26925_ (.a(net877),
    .b(net873),
    .c(net884),
    .out0(_01025_));
 b15norp02al1n02x5 _26926_ (.a(_16004_),
    .b(_01025_),
    .o1(_01026_));
 b15aoi112an1n03x5 _26927_ (.a(_16078_),
    .b(_01026_),
    .c(_17493_),
    .d(_15989_),
    .o1(_01027_));
 b15aoi022al1n04x5 _26928_ (.a(_00550_),
    .b(_15974_),
    .c(_17493_),
    .d(_17487_),
    .o1(_01028_));
 b15aoi012al1n06x5 _26929_ (.a(_01027_),
    .b(_01028_),
    .c(_16078_),
    .o1(_01029_));
 b15aoi022ar1n02x5 _26930_ (.a(net879),
    .b(_17427_),
    .c(_16164_),
    .d(net883),
    .o1(_01030_));
 b15oaoi13ah1n02x5 _26931_ (.a(_16018_),
    .b(_00612_),
    .c(_01030_),
    .d(net872),
    .o1(_01031_));
 b15aoi022ar1n02x5 _26932_ (.a(_16008_),
    .b(_15974_),
    .c(_15975_),
    .d(_15955_),
    .o1(_01032_));
 b15oai022ar1n02x5 _26933_ (.a(_16004_),
    .b(_15995_),
    .c(_01032_),
    .d(_15987_),
    .o1(_01033_));
 b15oaoi13ar1n03x5 _26934_ (.a(_16018_),
    .b(_16009_),
    .c(_16104_),
    .d(_16004_),
    .o1(_01034_));
 b15oab012al1n02x5 _26935_ (.a(net883),
    .b(_01033_),
    .c(_01034_),
    .out0(_01035_));
 b15nor004aq1n06x5 _26936_ (.a(_01024_),
    .b(_01029_),
    .c(_01031_),
    .d(_01035_),
    .o1(_01036_));
 b15oai012ar1n04x5 _26937_ (.a(_16025_),
    .b(_15997_),
    .c(_16088_),
    .o1(_01037_));
 b15nanb02ar1n24x5 _26938_ (.a(net873),
    .b(net885),
    .out0(_01038_));
 b15xor002al1n04x5 _26939_ (.a(\us20.a[6] ),
    .b(net879),
    .out0(_01039_));
 b15aoi013as1n04x5 _26940_ (.a(_01038_),
    .b(_01039_),
    .c(net864),
    .d(_15943_),
    .o1(_01040_));
 b15oai122as1n12x5 _26941_ (.a(_01040_),
    .b(_00561_),
    .c(_17517_),
    .d(_16061_),
    .e(_17401_),
    .o1(_01041_));
 b15nand04an1n08x5 _26942_ (.a(net865),
    .b(_15969_),
    .c(_01037_),
    .d(_01041_),
    .o1(_01042_));
 b15aoi022ar1n02x5 _26943_ (.a(_00550_),
    .b(_17518_),
    .c(_17437_),
    .d(_16110_),
    .o1(_01043_));
 b15aob012ah1n03x5 _26944_ (.a(_01041_),
    .b(_01043_),
    .c(_00999_),
    .out0(_01044_));
 b15nandp3ah1n02x5 _26945_ (.a(net869),
    .b(_16129_),
    .c(_17480_),
    .o1(_01045_));
 b15oaoi13ar1n04x5 _26946_ (.a(net878),
    .b(_01045_),
    .c(_16090_),
    .d(_16085_),
    .o1(_01046_));
 b15aoai13as1n08x5 _26947_ (.a(\us20.a[7] ),
    .b(_01046_),
    .c(_17513_),
    .d(_16006_),
    .o1(_01047_));
 b15aoi022ah1n12x5 _26948_ (.a(net872),
    .b(_01042_),
    .c(_01044_),
    .d(_01047_),
    .o1(_01048_));
 b15nano22as1n24x5 _26949_ (.a(_01020_),
    .b(_01036_),
    .c(_01048_),
    .out0(_01049_));
 b15xor002ah1n02x5 _26950_ (.a(_00974_),
    .b(_01049_),
    .out0(_01050_));
 b15nonb02ar1n12x5 _26951_ (.a(net754),
    .b(net765),
    .out0(_01051_));
 b15nonb03as1n04x5 _26952_ (.a(net762),
    .b(net758),
    .c(net745),
    .out0(_01052_));
 b15nand04as1n04x5 _26953_ (.a(net747),
    .b(_01051_),
    .c(_16785_),
    .d(_01052_),
    .o1(_01053_));
 b15oai112as1n04x5 _26954_ (.a(_16892_),
    .b(_16894_),
    .c(_17303_),
    .d(_16915_),
    .o1(_01054_));
 b15norp02an1n03x5 _26955_ (.a(_16770_),
    .b(_16815_),
    .o1(_01055_));
 b15oai112aq1n12x5 _26956_ (.a(_01053_),
    .b(_01054_),
    .c(_01055_),
    .d(_16919_),
    .o1(_01056_));
 b15aoi012ar1n02x5 _26957_ (.a(_16713_),
    .b(_16897_),
    .c(_16811_),
    .o1(_01057_));
 b15nandp2al1n04x5 _26958_ (.a(_16896_),
    .b(_16846_),
    .o1(_01058_));
 b15oai012as1n04x5 _26959_ (.a(_01058_),
    .b(_16811_),
    .c(_16693_),
    .o1(_01059_));
 b15oaoi13ah1n04x5 _26960_ (.a(_01056_),
    .b(_01057_),
    .c(_01059_),
    .d(net762),
    .o1(_01060_));
 b15nano22aq1n02x5 _26961_ (.a(net759),
    .b(\us31.a[4] ),
    .c(\us31.a[7] ),
    .out0(_01061_));
 b15aoi012al1n06x5 _26962_ (.a(_01061_),
    .b(_17359_),
    .c(_17328_),
    .o1(_01062_));
 b15nand02ar1n02x5 _26963_ (.a(net747),
    .b(_16834_),
    .o1(_01063_));
 b15oai012ar1n02x5 _26964_ (.a(_16741_),
    .b(_16804_),
    .c(_00735_),
    .o1(_01064_));
 b15nand02ar1n02x5 _26965_ (.a(\us31.a[4] ),
    .b(_16708_),
    .o1(_01065_));
 b15oai022aq1n04x5 _26966_ (.a(_01062_),
    .b(_01063_),
    .c(_01064_),
    .d(_01065_),
    .o1(_01066_));
 b15oai022ar1n04x5 _26967_ (.a(_16774_),
    .b(_16790_),
    .c(_17371_),
    .d(_16713_),
    .o1(_01067_));
 b15aoi022ah1n06x5 _26968_ (.a(net766),
    .b(_01066_),
    .c(_01067_),
    .d(_16836_),
    .o1(_01068_));
 b15nona22al1n08x5 _26969_ (.a(net766),
    .b(net758),
    .c(net763),
    .out0(_01069_));
 b15oai022aq1n02x5 _26970_ (.a(_16888_),
    .b(_16855_),
    .c(_17371_),
    .d(_01069_),
    .o1(_01070_));
 b15nonb02ah1n02x5 _26971_ (.a(_16854_),
    .b(_17317_),
    .out0(_01071_));
 b15nor002ar1n02x5 _26972_ (.a(_16888_),
    .b(_00781_),
    .o1(_01072_));
 b15oai013aq1n06x5 _26973_ (.a(net755),
    .b(_01070_),
    .c(_01071_),
    .d(_01072_),
    .o1(_01073_));
 b15aoi022ar1n08x5 _26974_ (.a(net765),
    .b(_16793_),
    .c(_17371_),
    .d(_16907_),
    .o1(_01074_));
 b15xnr002al1n12x5 _26975_ (.a(net744),
    .b(net747),
    .out0(_01075_));
 b15and003as1n02x5 _26976_ (.a(_16693_),
    .b(_16702_),
    .c(_01075_),
    .o(_01076_));
 b15oai112aq1n16x5 _26977_ (.a(_16798_),
    .b(_01074_),
    .c(_01076_),
    .d(net761),
    .o1(_01077_));
 b15oaoi13an1n03x5 _26978_ (.a(_16887_),
    .b(_00708_),
    .c(_00794_),
    .d(net751),
    .o1(_01078_));
 b15nor002aq1n06x5 _26979_ (.a(_16741_),
    .b(_00708_),
    .o1(_01079_));
 b15aoai13an1n06x5 _26980_ (.a(net759),
    .b(_01078_),
    .c(_01079_),
    .d(_16907_),
    .o1(_01080_));
 b15nano23ar1n02x5 _26981_ (.a(_16741_),
    .b(_01052_),
    .c(net747),
    .d(_17285_),
    .out0(_01081_));
 b15aoai13al1n02x5 _26982_ (.a(net765),
    .b(_01081_),
    .c(_17337_),
    .d(_16844_),
    .o1(_01082_));
 b15andc04ah1n03x5 _26983_ (.a(_01073_),
    .b(_01077_),
    .c(_01080_),
    .d(_01082_),
    .o(_01083_));
 b15aoai13ar1n03x5 _26984_ (.a(_16861_),
    .b(_17337_),
    .c(_16789_),
    .d(net765),
    .o1(_01084_));
 b15nandp3an1n03x5 _26985_ (.a(net758),
    .b(net749),
    .c(_16830_),
    .o1(_01085_));
 b15nandp3an1n03x5 _26986_ (.a(_16774_),
    .b(_16731_),
    .c(_16782_),
    .o1(_01086_));
 b15aoai13aq1n06x5 _26987_ (.a(_01084_),
    .b(_17390_),
    .c(_01085_),
    .d(_01086_),
    .o1(_01087_));
 b15aoi022ar1n04x5 _26988_ (.a(net758),
    .b(_16758_),
    .c(_16836_),
    .d(_17303_),
    .o1(_01088_));
 b15aoi012ah1n02x5 _26989_ (.a(_16758_),
    .b(_17303_),
    .c(net758),
    .o1(_01089_));
 b15oai112as1n08x5 _26990_ (.a(_16741_),
    .b(_01088_),
    .c(_01089_),
    .d(_16780_),
    .o1(_01090_));
 b15nor004ah1n03x5 _26991_ (.a(_16774_),
    .b(_17285_),
    .c(_16850_),
    .d(_17367_),
    .o1(_01091_));
 b15nor004ah1n03x5 _26992_ (.a(_16770_),
    .b(_17389_),
    .c(_16849_),
    .d(_16772_),
    .o1(_01092_));
 b15nano22an1n02x5 _26993_ (.a(net757),
    .b(net753),
    .c(net748),
    .out0(_01093_));
 b15nano22aq1n05x5 _26994_ (.a(net767),
    .b(net750),
    .c(net744),
    .out0(_01094_));
 b15nand02as1n04x5 _26995_ (.a(net767),
    .b(net750),
    .o1(_01095_));
 b15nonb02aq1n02x5 _26996_ (.a(net744),
    .b(net760),
    .out0(_01096_));
 b15aoai13ah1n06x5 _26997_ (.a(_01093_),
    .b(_01094_),
    .c(_01095_),
    .d(_01096_),
    .o1(_01097_));
 b15nona23aq1n16x5 _26998_ (.a(_01091_),
    .b(_01092_),
    .c(_01097_),
    .d(net756),
    .out0(_01098_));
 b15aoi022an1n16x5 _26999_ (.a(net761),
    .b(_01087_),
    .c(_01090_),
    .d(_01098_),
    .o1(_01099_));
 b15nand04as1n16x5 _27000_ (.a(_01060_),
    .b(_01068_),
    .c(_01083_),
    .d(_01099_),
    .o1(_01100_));
 b15nandp3as1n03x5 _27001_ (.a(net758),
    .b(_16725_),
    .c(_16726_),
    .o1(_01101_));
 b15aoi022as1n04x5 _27002_ (.a(_16785_),
    .b(_16726_),
    .c(_16782_),
    .d(_16731_),
    .o1(_01102_));
 b15oai022an1n06x5 _27003_ (.a(net763),
    .b(_01101_),
    .c(_01069_),
    .d(_01102_),
    .o1(_01103_));
 b15nonb02al1n04x5 _27004_ (.a(net762),
    .b(\us31.a[7] ),
    .out0(_01104_));
 b15nonb03ah1n02x5 _27005_ (.a(net753),
    .b(net748),
    .c(\us31.a[2] ),
    .out0(_01105_));
 b15aoai13an1n08x5 _27006_ (.a(_01104_),
    .b(_01105_),
    .c(\us31.a[2] ),
    .d(_16824_),
    .o1(_01106_));
 b15nandp3ar1n08x5 _27007_ (.a(\us31.a[4] ),
    .b(net745),
    .c(net748),
    .o1(_01107_));
 b15nanb02an1n03x5 _27008_ (.a(_01107_),
    .b(_17287_),
    .out0(_01108_));
 b15aoai13an1n06x5 _27009_ (.a(_01101_),
    .b(net751),
    .c(_01106_),
    .d(_01108_),
    .o1(_01109_));
 b15aoai13ah1n08x5 _27010_ (.a(net755),
    .b(_01103_),
    .c(_01109_),
    .d(net766),
    .o1(_01110_));
 b15nand02an1n03x5 _27011_ (.a(net762),
    .b(net755),
    .o1(_01111_));
 b15aoai13ar1n04x5 _27012_ (.a(_16832_),
    .b(_01111_),
    .c(_16793_),
    .d(_01058_),
    .o1(_01112_));
 b15aoi012ah1n02x5 _27013_ (.a(_16844_),
    .b(_16798_),
    .c(_16693_),
    .o1(_01113_));
 b15oai012as1n08x5 _27014_ (.a(_01112_),
    .b(_01113_),
    .c(_16770_),
    .o1(_01114_));
 b15nandp3ar1n02x5 _27015_ (.a(net756),
    .b(net751),
    .c(net753),
    .o1(_01115_));
 b15nand04ar1n02x5 _27016_ (.a(net767),
    .b(net757),
    .c(net744),
    .d(net747),
    .o1(_01116_));
 b15orn002ar1n02x5 _27017_ (.a(net760),
    .b(net757),
    .o(_01117_));
 b15oaoi13as1n02x5 _27018_ (.a(_01115_),
    .b(_01116_),
    .c(_01075_),
    .d(_01117_),
    .o1(_01118_));
 b15nanb02ah1n08x5 _27019_ (.a(net757),
    .b(net751),
    .out0(_01119_));
 b15nor003aq1n04x5 _27020_ (.a(_16728_),
    .b(_00789_),
    .c(_01119_),
    .o1(_01120_));
 b15oaoi13an1n04x5 _27021_ (.a(_01118_),
    .b(net760),
    .c(_00815_),
    .d(_01120_),
    .o1(_01121_));
 b15nano23al1n03x5 _27022_ (.a(_16896_),
    .b(_00802_),
    .c(_16719_),
    .d(_16746_),
    .out0(_01122_));
 b15norp02ar1n02x5 _27023_ (.a(net757),
    .b(_16780_),
    .o1(_01123_));
 b15nor002ah1n04x5 _27024_ (.a(_16849_),
    .b(_16850_),
    .o1(_01124_));
 b15aoi013ah1n02x5 _27025_ (.a(_01122_),
    .b(_01123_),
    .c(_01124_),
    .d(net756),
    .o1(_01125_));
 b15nand03an1n06x5 _27026_ (.a(_16824_),
    .b(_16861_),
    .c(_01094_),
    .o1(_01126_));
 b15nor002ar1n16x5 _27027_ (.a(net753),
    .b(net744),
    .o1(_01127_));
 b15oab012al1n03x5 _27028_ (.a(_01127_),
    .b(_17297_),
    .c(net760),
    .out0(_01128_));
 b15nand02as1n02x5 _27029_ (.a(_16861_),
    .b(_16820_),
    .o1(_01129_));
 b15oai122an1n12x5 _27030_ (.a(_01126_),
    .b(_01128_),
    .c(_01129_),
    .d(_16786_),
    .e(_16835_),
    .o1(_01130_));
 b15aoi013ah1n03x5 _27031_ (.a(net761),
    .b(net766),
    .c(_16915_),
    .d(_16763_),
    .o1(_01131_));
 b15aoi013an1n04x5 _27032_ (.a(_16770_),
    .b(net758),
    .c(_16785_),
    .d(_16726_),
    .o1(_01132_));
 b15nonb03aq1n02x5 _27033_ (.a(net754),
    .b(net758),
    .c(net766),
    .out0(_01133_));
 b15aoi022ah1n06x5 _27034_ (.a(_16905_),
    .b(_17375_),
    .c(_01133_),
    .d(_16789_),
    .o1(_01134_));
 b15aoi012an1n12x5 _27035_ (.a(_01131_),
    .b(_01132_),
    .c(_01134_),
    .o1(_01135_));
 b15nano23an1n12x5 _27036_ (.a(_01121_),
    .b(_01125_),
    .c(_01130_),
    .d(_01135_),
    .out0(_01136_));
 b15nand04as1n16x5 _27037_ (.a(_00729_),
    .b(_01110_),
    .c(_01114_),
    .d(_01136_),
    .o1(_01137_));
 b15nor002ah1n32x5 _27038_ (.a(_01100_),
    .b(_01137_),
    .o1(_01138_));
 b15xor002as1n12x5 _27039_ (.a(_00706_),
    .b(_01138_),
    .out0(_01139_));
 b15xor002al1n03x5 _27040_ (.a(_17069_),
    .b(_01139_),
    .out0(_01140_));
 b15xor002al1n04x5 _27041_ (.a(_01050_),
    .b(_01140_),
    .out0(_01141_));
 b15cmbn22ah1n12x5 _27042_ (.clk1(\text_in_r[35] ),
    .clk2(_01141_),
    .clkout(_01142_),
    .s(net540));
 b15xor002as1n16x5 _27043_ (.a(net530),
    .b(_01142_),
    .out0(_00116_));
 b15aoi012ar1n02x5 _27044_ (.a(net732),
    .b(_16248_),
    .c(_16332_),
    .o1(_01143_));
 b15aoi122ah1n02x5 _27045_ (.a(_16226_),
    .b(_16202_),
    .c(_16293_),
    .d(_16328_),
    .e(_16301_),
    .o1(_01144_));
 b15oai012ah1n02x5 _27046_ (.a(_16342_),
    .b(_01143_),
    .c(_01144_),
    .o1(_01145_));
 b15nand03an1n06x5 _27047_ (.a(_16226_),
    .b(_16223_),
    .c(_16230_),
    .o1(_01146_));
 b15oai122aq1n04x5 _27048_ (.a(_01146_),
    .b(_16993_),
    .c(_17045_),
    .d(_16226_),
    .e(_16225_),
    .o1(_01147_));
 b15oai112ah1n04x5 _27049_ (.a(net742),
    .b(_01145_),
    .c(_01147_),
    .d(_16342_),
    .o1(_01148_));
 b15nand02as1n03x5 _27050_ (.a(_16283_),
    .b(_16226_),
    .o1(_01149_));
 b15oai012ah1n02x5 _27051_ (.a(net739),
    .b(_16231_),
    .c(_01149_),
    .o1(_01150_));
 b15aoi013as1n04x5 _27052_ (.a(_01150_),
    .b(_16416_),
    .c(_16221_),
    .d(net731),
    .o1(_01151_));
 b15oai013ar1n02x5 _27053_ (.a(_16342_),
    .b(net740),
    .c(_16235_),
    .d(_16237_),
    .o1(_01152_));
 b15oai022ar1n02x5 _27054_ (.a(net729),
    .b(_16372_),
    .c(_17247_),
    .d(net725),
    .o1(_01153_));
 b15aoi013an1n02x5 _27055_ (.a(_01152_),
    .b(_01153_),
    .c(_16193_),
    .d(net720),
    .o1(_01154_));
 b15nanb03al1n16x5 _27056_ (.a(net722),
    .b(net725),
    .c(net733),
    .out0(_01155_));
 b15aoi012ar1n02x5 _27057_ (.a(_16235_),
    .b(_16237_),
    .c(_01155_),
    .o1(_01156_));
 b15aoi013al1n02x5 _27058_ (.a(_01156_),
    .b(_16418_),
    .c(net720),
    .d(net725),
    .o1(_01157_));
 b15oa0012aq1n06x5 _27059_ (.a(_01154_),
    .b(_01157_),
    .c(net729),
    .o(_01158_));
 b15norp03ah1n03x5 _27060_ (.a(net722),
    .b(_16381_),
    .c(_16928_),
    .o1(_01159_));
 b15inv000al1n02x5 _27061_ (.a(_16935_),
    .o1(_01160_));
 b15oai022ar1n08x5 _27062_ (.a(_17052_),
    .b(_16928_),
    .c(_16929_),
    .d(_01160_),
    .o1(_01161_));
 b15aoai13as1n08x5 _27063_ (.a(net718),
    .b(_01159_),
    .c(_01161_),
    .d(net729),
    .o1(_01162_));
 b15aoai13as1n06x5 _27064_ (.a(_01148_),
    .b(_01151_),
    .c(_01158_),
    .d(_01162_),
    .o1(_01163_));
 b15oaoi13aq1n03x5 _27065_ (.a(_01149_),
    .b(_16225_),
    .c(_16388_),
    .d(_16402_),
    .o1(_01164_));
 b15oai022an1n02x5 _27066_ (.a(_16986_),
    .b(_16336_),
    .c(_16993_),
    .d(_16260_),
    .o1(_01165_));
 b15aoi112aq1n04x5 _27067_ (.a(_16338_),
    .b(_01164_),
    .c(_01165_),
    .d(_16283_),
    .o1(_01166_));
 b15aoai13ar1n03x5 _27068_ (.a(_01155_),
    .b(net734),
    .c(_16398_),
    .d(_16313_),
    .o1(_01167_));
 b15aoi013aq1n03x5 _27069_ (.a(net731),
    .b(_16328_),
    .c(_16970_),
    .d(_01167_),
    .o1(_01168_));
 b15norp02ar1n02x5 _27070_ (.a(_16278_),
    .b(_16372_),
    .o1(_01169_));
 b15aoi022as1n04x5 _27071_ (.a(_16291_),
    .b(_16935_),
    .c(_01169_),
    .d(_16350_),
    .o1(_01170_));
 b15orn003ar1n03x5 _27072_ (.a(_16283_),
    .b(net719),
    .c(_01170_),
    .o(_01171_));
 b15oai012an1n04x5 _27073_ (.a(_16391_),
    .b(_16388_),
    .c(_16396_),
    .o1(_01172_));
 b15aoi112al1n06x5 _27074_ (.a(_16226_),
    .b(_01172_),
    .c(_17224_),
    .d(_16321_),
    .o1(_01173_));
 b15aoai13as1n06x5 _27075_ (.a(_01166_),
    .b(_01168_),
    .c(_01171_),
    .d(_01173_),
    .o1(_01174_));
 b15aoi022an1n02x5 _27076_ (.a(_16278_),
    .b(_16259_),
    .c(_16328_),
    .d(_16185_),
    .o1(_01175_));
 b15oai013ar1n02x5 _27077_ (.a(_16283_),
    .b(_17052_),
    .c(_16314_),
    .d(_16342_),
    .o1(_01176_));
 b15aob012ar1n02x5 _27078_ (.a(_00930_),
    .b(_01176_),
    .c(_16289_),
    .out0(_01177_));
 b15nanb03as1n03x5 _27079_ (.a(_01175_),
    .b(_16405_),
    .c(_01177_),
    .out0(_01178_));
 b15aoi022an1n06x5 _27080_ (.a(_16343_),
    .b(_16997_),
    .c(_17229_),
    .d(net737),
    .o1(_01179_));
 b15bfn000as1n02x5 input14 (.a(key[111]),
    .o(net14));
 b15oai012an1n12x5 _27082_ (.a(_01178_),
    .b(_01179_),
    .c(net733),
    .o1(_01181_));
 b15oai012ar1n02x5 _27083_ (.a(_16313_),
    .b(_16398_),
    .c(_16283_),
    .o1(_01182_));
 b15aoai13ar1n02x5 _27084_ (.a(net735),
    .b(_17048_),
    .c(_01182_),
    .d(_16989_),
    .o1(_01183_));
 b15xor002ar1n02x5 _27085_ (.a(net729),
    .b(net717),
    .out0(_01184_));
 b15and003ar1n03x5 _27086_ (.a(_16333_),
    .b(_00636_),
    .c(_01184_),
    .o(_01185_));
 b15oai022ar1n02x5 _27087_ (.a(net731),
    .b(_16235_),
    .c(_16280_),
    .d(net742),
    .o1(_01186_));
 b15aoi013an1n02x5 _27088_ (.a(_01185_),
    .b(_01186_),
    .c(_16301_),
    .d(_16356_),
    .o1(_01187_));
 b15nor002an1n03x5 _27089_ (.a(net733),
    .b(_16323_),
    .o1(_01188_));
 b15norp02as1n03x5 _27090_ (.a(_16965_),
    .b(_16952_),
    .o1(_01189_));
 b15aoi222aq1n12x5 _27091_ (.a(_16233_),
    .b(_16980_),
    .c(_16325_),
    .d(_01188_),
    .e(_01189_),
    .f(_16419_),
    .o1(_01190_));
 b15nor003aq1n06x5 _27092_ (.a(_16276_),
    .b(_16979_),
    .c(_00644_),
    .o1(_01191_));
 b15norp03ar1n03x5 _27093_ (.a(_16280_),
    .b(_16310_),
    .c(_16986_),
    .o1(_01192_));
 b15nor004as1n02x5 _27094_ (.a(_16237_),
    .b(_16390_),
    .c(_16280_),
    .d(_16381_),
    .o1(_01193_));
 b15nor004ah1n04x5 _27095_ (.a(_17019_),
    .b(_01191_),
    .c(_01192_),
    .d(_01193_),
    .o1(_01194_));
 b15nand04an1n04x5 _27096_ (.a(_01183_),
    .b(_01187_),
    .c(_01190_),
    .d(_01194_),
    .o1(_01195_));
 b15nona23ah1n08x5 _27097_ (.a(_16185_),
    .b(_16193_),
    .c(_16932_),
    .d(net733),
    .out0(_01196_));
 b15nandp2ah1n02x5 _27098_ (.a(_16325_),
    .b(_17210_),
    .o1(_01197_));
 b15oaoi13an1n04x5 _27099_ (.a(net731),
    .b(_01196_),
    .c(_01197_),
    .d(_16334_),
    .o1(_01198_));
 b15oai022an1n06x5 _27100_ (.a(net723),
    .b(_16967_),
    .c(_16372_),
    .d(_00644_),
    .o1(_01199_));
 b15and003ar1n03x5 _27101_ (.a(net737),
    .b(_16305_),
    .c(_01199_),
    .o(_01200_));
 b15oai022aq1n02x5 _27102_ (.a(_17005_),
    .b(_17015_),
    .c(_16396_),
    .d(_16221_),
    .o1(_01201_));
 b15oai012al1n08x5 _27103_ (.a(net731),
    .b(_01200_),
    .c(_01201_),
    .o1(_01202_));
 b15aoai13ah1n02x5 _27104_ (.a(_16223_),
    .b(_16224_),
    .c(_16230_),
    .d(_16283_),
    .o1(_01203_));
 b15aoi012ar1n02x5 _27105_ (.a(_16318_),
    .b(_01203_),
    .c(_17005_),
    .o1(_01204_));
 b15nand02ar1n02x5 _27106_ (.a(_16248_),
    .b(_16936_),
    .o1(_01205_));
 b15oai022ar1n02x5 _27107_ (.a(_16283_),
    .b(_16327_),
    .c(_16958_),
    .d(_01205_),
    .o1(_01206_));
 b15aoi012ah1n02x5 _27108_ (.a(_01204_),
    .b(_01206_),
    .c(net731),
    .o1(_01207_));
 b15nona23an1n12x5 _27109_ (.a(_01195_),
    .b(_01198_),
    .c(_01202_),
    .d(_01207_),
    .out0(_01208_));
 b15nor004as1n12x5 _27110_ (.a(_01163_),
    .b(_01174_),
    .c(_01181_),
    .d(_01208_),
    .o1(_01209_));
 b15aoi012ar1n02x5 _27111_ (.a(_17553_),
    .b(_16656_),
    .c(net609),
    .o1(_01210_));
 b15nanb03ar1n04x5 _27112_ (.a(_01210_),
    .b(_16446_),
    .c(_16435_),
    .out0(_01211_));
 b15nor003as1n03x5 _27113_ (.a(net618),
    .b(net615),
    .c(net609),
    .o1(_01212_));
 b15aoi022ah1n08x5 _27114_ (.a(_17152_),
    .b(_16646_),
    .c(_01212_),
    .d(_17128_),
    .o1(_01213_));
 b15aoi013an1n04x5 _27115_ (.a(net613),
    .b(_16477_),
    .c(_01211_),
    .d(_01213_),
    .o1(_01214_));
 b15norp02as1n04x5 _27116_ (.a(net596),
    .b(_16439_),
    .o1(_01215_));
 b15nand02as1n12x5 _27117_ (.a(_17099_),
    .b(\us13.a[0] ),
    .o1(_01216_));
 b15aoi022an1n04x5 _27118_ (.a(net606),
    .b(_01215_),
    .c(_17157_),
    .d(_01216_),
    .o1(_01217_));
 b15oai022ah1n06x5 _27119_ (.a(_17586_),
    .b(_00858_),
    .c(_01217_),
    .d(_16597_),
    .o1(_01218_));
 b15nand03aq1n12x5 _27120_ (.a(net618),
    .b(_16481_),
    .c(_16520_),
    .o1(_01219_));
 b15aoi012al1n04x5 _27121_ (.a(_16524_),
    .b(_01219_),
    .c(net603),
    .o1(_01220_));
 b15nand02as1n06x5 _27122_ (.a(_16466_),
    .b(_16620_),
    .o1(_01221_));
 b15aoi012ar1n04x5 _27123_ (.a(_16446_),
    .b(_17545_),
    .c(_17099_),
    .o1(_01222_));
 b15oai122an1n16x5 _27124_ (.a(_16558_),
    .b(_16528_),
    .c(_17175_),
    .d(_01221_),
    .e(_01222_),
    .o1(_01223_));
 b15norp02aq1n16x5 _27125_ (.a(_16673_),
    .b(_16549_),
    .o1(_01224_));
 b15nand03an1n04x5 _27126_ (.a(_16508_),
    .b(_16640_),
    .c(_01224_),
    .o1(_01225_));
 b15oai112an1n12x5 _27127_ (.a(net618),
    .b(_01225_),
    .c(_17116_),
    .d(_16626_),
    .o1(_01226_));
 b15aoi122an1n08x5 _27128_ (.a(_01214_),
    .b(_01218_),
    .c(_01220_),
    .d(_01223_),
    .e(_01226_),
    .o1(_01227_));
 b15orn002ar1n02x5 _27129_ (.a(_16516_),
    .b(_16608_),
    .o(_01228_));
 b15aoi022ar1n02x5 _27130_ (.a(_16659_),
    .b(_16473_),
    .c(_16494_),
    .d(_17181_),
    .o1(_01229_));
 b15oai013ah1n03x5 _27131_ (.a(_01228_),
    .b(_01216_),
    .c(_01229_),
    .d(net613),
    .o1(_01230_));
 b15nandp2ar1n03x5 _27132_ (.a(_16619_),
    .b(_16517_),
    .o1(_01231_));
 b15oai013as1n08x5 _27133_ (.a(_01231_),
    .b(_16619_),
    .c(_17565_),
    .d(_16497_),
    .o1(_01232_));
 b15nor002an1n03x5 _27134_ (.a(net609),
    .b(_16549_),
    .o1(_01233_));
 b15aoai13ar1n08x5 _27135_ (.a(net617),
    .b(_01230_),
    .c(_01232_),
    .d(_01233_),
    .o1(_01234_));
 b15nand02ar1n02x5 _27136_ (.a(net615),
    .b(_17562_),
    .o1(_01235_));
 b15nand02ar1n02x5 _27137_ (.a(_16453_),
    .b(_16526_),
    .o1(_01236_));
 b15aoi013an1n03x5 _27138_ (.a(_16466_),
    .b(_01235_),
    .c(_01219_),
    .d(_01236_),
    .o1(_01237_));
 b15aoai13an1n06x5 _27139_ (.a(net611),
    .b(_01237_),
    .c(_16674_),
    .d(_16466_),
    .o1(_01238_));
 b15nandp2an1n08x5 _27140_ (.a(_16475_),
    .b(_16605_),
    .o1(_01239_));
 b15nano22ar1n02x5 _27141_ (.a(net604),
    .b(net612),
    .c(net597),
    .out0(_01240_));
 b15aoi013al1n04x5 _27142_ (.a(_01240_),
    .b(net615),
    .c(net597),
    .d(_17099_),
    .o1(_01241_));
 b15oai222an1n16x5 _27143_ (.a(_17175_),
    .b(_17116_),
    .c(_01239_),
    .d(_17088_),
    .e(_01241_),
    .f(_17093_),
    .o1(_01242_));
 b15oai012aq1n04x5 _27144_ (.a(_16680_),
    .b(_16682_),
    .c(_16482_),
    .o1(_01243_));
 b15oai112al1n08x5 _27145_ (.a(_16456_),
    .b(_17119_),
    .c(_16482_),
    .d(net611),
    .o1(_01244_));
 b15aoai13aq1n06x5 _27146_ (.a(net608),
    .b(_01242_),
    .c(_01243_),
    .d(_01244_),
    .o1(_01245_));
 b15aoi022ar1n08x5 _27147_ (.a(_16475_),
    .b(_16621_),
    .c(_16579_),
    .d(_16684_),
    .o1(_01246_));
 b15oai012aq1n03x5 _27148_ (.a(_16508_),
    .b(_01246_),
    .c(net598),
    .o1(_01247_));
 b15nandp2aq1n03x5 _27149_ (.a(net608),
    .b(_16646_),
    .o1(_01248_));
 b15oai112al1n06x5 _27150_ (.a(net615),
    .b(_01248_),
    .c(_17183_),
    .d(_16479_),
    .o1(_01249_));
 b15nand03ah1n06x5 _27151_ (.a(_16558_),
    .b(_01247_),
    .c(_01249_),
    .o1(_01250_));
 b15nand02an1n02x5 _27152_ (.a(_17146_),
    .b(_17190_),
    .o1(_01251_));
 b15oai012as1n06x5 _27153_ (.a(_01251_),
    .b(_17125_),
    .c(_16479_),
    .o1(_01252_));
 b15nand03as1n06x5 _27154_ (.a(_16508_),
    .b(_16517_),
    .c(_16621_),
    .o1(_01253_));
 b15nano22an1n03x5 _27155_ (.a(net599),
    .b(net614),
    .c(\us13.a[3] ),
    .out0(_01254_));
 b15nand02aq1n06x5 _27156_ (.a(_16481_),
    .b(_01254_),
    .o1(_01255_));
 b15aoi012al1n12x5 _27157_ (.a(_16461_),
    .b(_01253_),
    .c(_01255_),
    .o1(_01256_));
 b15oai012al1n08x5 _27158_ (.a(net619),
    .b(_01252_),
    .c(_01256_),
    .o1(_01257_));
 b15nand04as1n16x5 _27159_ (.a(_01238_),
    .b(_01245_),
    .c(_01250_),
    .d(_01257_),
    .o1(_01258_));
 b15and002as1n03x5 _27160_ (.a(net599),
    .b(net618),
    .o(_01259_));
 b15nanb02al1n04x5 _27161_ (.a(net609),
    .b(net602),
    .out0(_01260_));
 b15nand04al1n12x5 _27162_ (.a(_16508_),
    .b(_17181_),
    .c(_01259_),
    .d(_01260_),
    .o1(_01261_));
 b15oaoi13ar1n03x5 _27163_ (.a(net613),
    .b(_01261_),
    .c(_17116_),
    .d(_16626_),
    .o1(_01262_));
 b15oai022ah1n06x5 _27164_ (.a(net617),
    .b(_16432_),
    .c(_16438_),
    .d(_16439_),
    .o1(_01263_));
 b15nor002as1n04x5 _27165_ (.a(_16671_),
    .b(_16479_),
    .o1(_01264_));
 b15aoi112ah1n03x5 _27166_ (.a(_16654_),
    .b(_01262_),
    .c(_01263_),
    .d(_01264_),
    .o1(_01265_));
 b15nand03al1n03x5 _27167_ (.a(_16456_),
    .b(_16517_),
    .c(_16601_),
    .o1(_01266_));
 b15oai012ar1n04x5 _27168_ (.a(_16498_),
    .b(_16604_),
    .c(net614),
    .o1(_01267_));
 b15oai012al1n06x5 _27169_ (.a(_01266_),
    .b(_01267_),
    .c(_16521_),
    .o1(_01268_));
 b15aoi022an1n06x5 _27170_ (.a(_16517_),
    .b(_16621_),
    .c(_01254_),
    .d(_16481_),
    .o1(_01269_));
 b15nand03an1n06x5 _27171_ (.a(_16458_),
    .b(_16558_),
    .c(net613),
    .o1(_01270_));
 b15oa0022ar1n03x5 _27172_ (.a(_16671_),
    .b(_16652_),
    .c(_17080_),
    .d(_17099_),
    .o(_01271_));
 b15nand02al1n04x5 _27173_ (.a(\us13.a[3] ),
    .b(_16520_),
    .o1(_01272_));
 b15oai022an1n12x5 _27174_ (.a(_01269_),
    .b(_01270_),
    .c(_01271_),
    .d(_01272_),
    .o1(_01273_));
 b15oai012as1n04x5 _27175_ (.a(_01261_),
    .b(_01221_),
    .c(_16564_),
    .o1(_01274_));
 b15aoi112ar1n08x5 _27176_ (.a(_01268_),
    .b(_01273_),
    .c(_01274_),
    .d(net603),
    .o1(_01275_));
 b15aoi022ar1n02x5 _27177_ (.a(_16429_),
    .b(_16520_),
    .c(_16656_),
    .d(_16657_),
    .o1(_01276_));
 b15nandp2aq1n16x5 _27178_ (.a(_16481_),
    .b(_16518_),
    .o1(_01277_));
 b15oaoi13aq1n03x5 _27179_ (.a(net614),
    .b(_01276_),
    .c(_01277_),
    .d(net618),
    .o1(_01278_));
 b15nano22aq1n03x5 _27180_ (.a(net605),
    .b(net598),
    .c(net614),
    .out0(_01279_));
 b15nonb03al1n04x5 _27181_ (.a(net614),
    .b(net598),
    .c(net605),
    .out0(_01280_));
 b15oai112ah1n12x5 _27182_ (.a(\us13.a[0] ),
    .b(_16621_),
    .c(_01279_),
    .d(_01280_),
    .o1(_01281_));
 b15oai013ah1n08x5 _27183_ (.a(_01281_),
    .b(_16513_),
    .c(_16652_),
    .d(_16432_),
    .o1(_01282_));
 b15aoi112al1n06x5 _27184_ (.a(_17159_),
    .b(_01278_),
    .c(_01282_),
    .d(net603),
    .o1(_01283_));
 b15nand03an1n16x5 _27185_ (.a(_01265_),
    .b(_01275_),
    .c(_01283_),
    .o1(_01284_));
 b15nano23as1n24x5 _27186_ (.a(_01227_),
    .b(_01234_),
    .c(_01258_),
    .d(_01284_),
    .out0(_01285_));
 b15xor002ah1n08x5 _27187_ (.a(_01209_),
    .b(_01285_),
    .out0(_01286_));
 b15xor002an1n02x5 _27188_ (.a(_17069_),
    .b(_01286_),
    .out0(_01287_));
 b15xor002al1n12x5 _27189_ (.a(net758),
    .b(\us31.a[7] ),
    .out0(_01288_));
 b15nand03as1n06x5 _27190_ (.a(_16824_),
    .b(_16873_),
    .c(_01288_),
    .o1(_01289_));
 b15nandp3as1n08x5 _27191_ (.a(net757),
    .b(_16750_),
    .c(_16789_),
    .o1(_01290_));
 b15nand02an1n02x5 _27192_ (.a(_01289_),
    .b(_01290_),
    .o1(_01291_));
 b15nor003aq1n02x5 _27193_ (.a(\us31.a[3] ),
    .b(net759),
    .c(net748),
    .o1(_01292_));
 b15xor002al1n04x5 _27194_ (.a(net759),
    .b(net748),
    .out0(_01293_));
 b15aoai13an1n06x5 _27195_ (.a(_17292_),
    .b(_01292_),
    .c(_01293_),
    .d(\us31.a[3] ),
    .o1(_01294_));
 b15nor002ar1n02x5 _27196_ (.a(\us31.a[4] ),
    .b(_00719_),
    .o1(_01295_));
 b15oai112as1n06x5 _27197_ (.a(_16830_),
    .b(_00714_),
    .c(_00726_),
    .d(_01295_),
    .o1(_01296_));
 b15aoi022aq1n02x5 _27198_ (.a(_16798_),
    .b(_16758_),
    .c(_16789_),
    .d(_16813_),
    .o1(_01297_));
 b15nand03aq1n03x5 _27199_ (.a(_01294_),
    .b(_01296_),
    .c(_01297_),
    .o1(_01298_));
 b15oai012ar1n08x5 _27200_ (.a(net766),
    .b(_01291_),
    .c(_01298_),
    .o1(_01299_));
 b15aoi022ar1n02x5 _27201_ (.a(net766),
    .b(_17299_),
    .c(_17298_),
    .d(_16907_),
    .o1(_01300_));
 b15norp03ar1n04x5 _27202_ (.a(net767),
    .b(net750),
    .c(net748),
    .o1(_01301_));
 b15aoi012ar1n02x5 _27203_ (.a(_01301_),
    .b(_16860_),
    .c(_17298_),
    .o1(_01302_));
 b15oai022ar1n02x5 _27204_ (.a(\us31.a[2] ),
    .b(_01300_),
    .c(_01302_),
    .d(net762),
    .o1(_01303_));
 b15and003aq1n03x5 _27205_ (.a(_16741_),
    .b(_17328_),
    .c(_01303_),
    .o(_01304_));
 b15nand02an1n24x5 _27206_ (.a(_16872_),
    .b(_00801_),
    .o1(_01305_));
 b15nor003ar1n06x5 _27207_ (.a(net762),
    .b(_16860_),
    .c(_01305_),
    .o1(_01306_));
 b15oai022al1n02x5 _27208_ (.a(net767),
    .b(_17285_),
    .c(_01095_),
    .d(net753),
    .o1(_01307_));
 b15nandp2ah1n16x5 _27209_ (.a(net756),
    .b(net757),
    .o1(_01308_));
 b15nano23aq1n08x5 _27210_ (.a(_16710_),
    .b(_01307_),
    .c(_01308_),
    .d(net760),
    .out0(_01309_));
 b15aoi012ah1n02x5 _27211_ (.a(_00738_),
    .b(_00726_),
    .c(_16780_),
    .o1(_01310_));
 b15nor004ah1n06x5 _27212_ (.a(_16774_),
    .b(_16836_),
    .c(_16841_),
    .d(_01310_),
    .o1(_01311_));
 b15nor004as1n08x5 _27213_ (.a(_01304_),
    .b(_01306_),
    .c(_01309_),
    .d(_01311_),
    .o1(_01312_));
 b15aoai13al1n08x5 _27214_ (.a(_16836_),
    .b(_16915_),
    .c(net758),
    .d(_17337_),
    .o1(_01313_));
 b15oai022ar1n02x5 _27215_ (.a(net759),
    .b(_16748_),
    .c(_16760_),
    .d(_17371_),
    .o1(_01314_));
 b15aob012al1n06x5 _27216_ (.a(_01313_),
    .b(_01314_),
    .c(net763),
    .out0(_01315_));
 b15nano23ar1n02x5 _27217_ (.a(net763),
    .b(\us31.a[0] ),
    .c(net759),
    .d(net748),
    .out0(_01316_));
 b15oaoi13as1n02x5 _27218_ (.a(_16741_),
    .b(_01316_),
    .c(_17292_),
    .d(_17363_),
    .o1(_01317_));
 b15xnr002aq1n08x5 _27219_ (.a(net750),
    .b(\us31.a[7] ),
    .out0(_01318_));
 b15aoi022as1n04x5 _27220_ (.a(_01127_),
    .b(_00714_),
    .c(_00760_),
    .d(_01318_),
    .o1(_01319_));
 b15oai013as1n06x5 _27221_ (.a(_01317_),
    .b(_01319_),
    .c(net748),
    .d(\us31.a[0] ),
    .o1(_01320_));
 b15aoai13ah1n03x5 _27222_ (.a(_16770_),
    .b(_16758_),
    .c(_16860_),
    .d(_16742_),
    .o1(_01321_));
 b15oai122an1n12x5 _27223_ (.a(_01321_),
    .b(_17335_),
    .c(_16888_),
    .d(_16867_),
    .e(_01069_),
    .o1(_01322_));
 b15oai022ar1n12x5 _27224_ (.a(net755),
    .b(_01315_),
    .c(_01320_),
    .d(_01322_),
    .o1(_01323_));
 b15nand02ar1n16x5 _27225_ (.a(_16693_),
    .b(_16892_),
    .o1(_01324_));
 b15oai122as1n04x5 _27226_ (.a(net762),
    .b(_00708_),
    .c(_01324_),
    .d(_01289_),
    .e(_16774_),
    .o1(_01325_));
 b15aoi012ah1n02x5 _27227_ (.a(net758),
    .b(_17319_),
    .c(_01289_),
    .o1(_01326_));
 b15nor004ah1n04x5 _27228_ (.a(net755),
    .b(net751),
    .c(_16760_),
    .d(_01107_),
    .o1(_01327_));
 b15oai013ar1n08x5 _27229_ (.a(_01325_),
    .b(_01326_),
    .c(_01327_),
    .d(net762),
    .o1(_01328_));
 b15orn002ar1n02x5 _27230_ (.a(net763),
    .b(\us31.a[4] ),
    .o(_01329_));
 b15oai112aq1n02x5 _27231_ (.a(net750),
    .b(net745),
    .c(net748),
    .d(_16693_),
    .o1(_01330_));
 b15oaoi13ar1n04x5 _27232_ (.a(_01329_),
    .b(_01330_),
    .c(net750),
    .d(_00794_),
    .o1(_01331_));
 b15nor002as1n08x5 _27233_ (.a(net765),
    .b(_16739_),
    .o1(_01332_));
 b15aoi112an1n06x5 _27234_ (.a(net755),
    .b(_01331_),
    .c(_01332_),
    .d(_01318_),
    .o1(_01333_));
 b15oai012al1n06x5 _27235_ (.a(net758),
    .b(_16742_),
    .c(_16741_),
    .o1(_01334_));
 b15oai112as1n16x5 _27236_ (.a(_01323_),
    .b(_01328_),
    .c(_01333_),
    .d(_01334_),
    .o1(_01335_));
 b15aoi012ar1n06x5 _27237_ (.a(_17298_),
    .b(_17299_),
    .c(net762),
    .o1(_01336_));
 b15nor004aq1n06x5 _27238_ (.a(_16713_),
    .b(_17297_),
    .c(_16836_),
    .d(_01336_),
    .o1(_01337_));
 b15nand02ar1n02x5 _27239_ (.a(_16772_),
    .b(_16813_),
    .o1(_01338_));
 b15aoi013as1n02x5 _27240_ (.a(_16764_),
    .b(_00792_),
    .c(_01324_),
    .d(_01338_),
    .o1(_01339_));
 b15oai012ah1n02x5 _27241_ (.a(_16769_),
    .b(_16832_),
    .c(_16899_),
    .o1(_01340_));
 b15aoi022ah1n06x5 _27242_ (.a(_16708_),
    .b(_16845_),
    .c(_16846_),
    .d(_16830_),
    .o1(_01341_));
 b15nand02al1n02x5 _27243_ (.a(\us31.a[4] ),
    .b(_16861_),
    .o1(_01342_));
 b15aoi022ah1n06x5 _27244_ (.a(_16693_),
    .b(_16763_),
    .c(_16836_),
    .d(_16892_),
    .o1(_01343_));
 b15oai022an1n06x5 _27245_ (.a(_01341_),
    .b(_01342_),
    .c(_01343_),
    .d(_00730_),
    .o1(_01344_));
 b15nor004an1n06x5 _27246_ (.a(_01337_),
    .b(_01339_),
    .c(_01340_),
    .d(_01344_),
    .o1(_01345_));
 b15nonb02ar1n04x5 _27247_ (.a(net752),
    .b(net761),
    .out0(_01346_));
 b15nano23an1n03x5 _27248_ (.a(_16815_),
    .b(_16804_),
    .c(_01346_),
    .d(net746),
    .out0(_01347_));
 b15norp03al1n02x5 _27249_ (.a(_16739_),
    .b(_16728_),
    .c(_01119_),
    .o1(_01348_));
 b15oab012ah1n06x5 _27250_ (.a(net745),
    .b(_01347_),
    .c(_01348_),
    .out0(_01349_));
 b15oai022al1n08x5 _27251_ (.a(_16897_),
    .b(_01308_),
    .c(_17373_),
    .d(_16761_),
    .o1(_01350_));
 b15oai022ar1n08x5 _27252_ (.a(_16888_),
    .b(_17367_),
    .c(_17371_),
    .d(_16775_),
    .o1(_01351_));
 b15aoi122an1n08x5 _27253_ (.a(_01349_),
    .b(_01350_),
    .c(net761),
    .d(_01351_),
    .e(_16741_),
    .o1(_01352_));
 b15oai022ah1n02x5 _27254_ (.a(_16761_),
    .b(_16810_),
    .c(_17355_),
    .d(net765),
    .o1(_01353_));
 b15nor002aq1n04x5 _27255_ (.a(net762),
    .b(_01353_),
    .o1(_01354_));
 b15xor002an1n16x5 _27256_ (.a(\us31.a[4] ),
    .b(\us31.a[6] ),
    .out0(_01355_));
 b15norp03ah1n03x5 _27257_ (.a(net759),
    .b(net751),
    .c(\us31.a[7] ),
    .o1(_01356_));
 b15aoi022an1n12x5 _27258_ (.a(_16896_),
    .b(_16804_),
    .c(_01355_),
    .d(_01356_),
    .o1(_01357_));
 b15oai022as1n06x5 _27259_ (.a(_17335_),
    .b(_16802_),
    .c(_01357_),
    .d(net755),
    .o1(_01358_));
 b15nor004aq1n06x5 _27260_ (.a(net755),
    .b(net751),
    .c(_16898_),
    .d(_01107_),
    .o1(_01359_));
 b15nandp2an1n08x5 _27261_ (.a(_16798_),
    .b(_16789_),
    .o1(_01360_));
 b15aob012ar1n08x5 _27262_ (.a(_01360_),
    .b(_16902_),
    .c(_01051_),
    .out0(_01361_));
 b15nor004aq1n06x5 _27263_ (.a(_16770_),
    .b(_01358_),
    .c(_01359_),
    .d(_01361_),
    .o1(_01362_));
 b15oai112as1n16x5 _27264_ (.a(_01345_),
    .b(_01352_),
    .c(_01354_),
    .d(_01362_),
    .o1(_01363_));
 b15nano23as1n24x5 _27265_ (.a(_01299_),
    .b(_01312_),
    .c(_01335_),
    .d(_01363_),
    .out0(_01364_));
 b15nandp3an1n02x5 _27266_ (.a(net880),
    .b(_16034_),
    .c(_16077_),
    .o1(_01365_));
 b15oaoi13an1n04x5 _27267_ (.a(_16028_),
    .b(_01365_),
    .c(_16061_),
    .d(_16040_),
    .o1(_01366_));
 b15aoi022aq1n02x5 _27268_ (.a(\us20.a[1] ),
    .b(_15943_),
    .c(_17420_),
    .d(\us20.a[4] ),
    .o1(_01367_));
 b15nand02an1n02x5 _27269_ (.a(net874),
    .b(_15939_),
    .o1(_01368_));
 b15oai022ah1n06x5 _27270_ (.a(net874),
    .b(_17407_),
    .c(_01367_),
    .d(_01368_),
    .o1(_01369_));
 b15aoi112as1n08x5 _27271_ (.a(_16119_),
    .b(_01366_),
    .c(_01369_),
    .d(net885),
    .o1(_01370_));
 b15oai012ar1n02x5 _27272_ (.a(net876),
    .b(_17448_),
    .c(net882),
    .o1(_01371_));
 b15oai012ar1n02x5 _27273_ (.a(net879),
    .b(net872),
    .c(_16066_),
    .o1(_01372_));
 b15aoi012aq1n02x5 _27274_ (.a(_16135_),
    .b(_01371_),
    .c(_01372_),
    .o1(_01373_));
 b15oaoi13aq1n02x5 _27275_ (.a(_17400_),
    .b(_16004_),
    .c(_16078_),
    .d(_17401_),
    .o1(_01374_));
 b15aob012al1n04x5 _27276_ (.a(_17405_),
    .b(_00999_),
    .c(_17427_),
    .out0(_01375_));
 b15aoi112aq1n04x5 _27277_ (.a(_01373_),
    .b(_01374_),
    .c(_01375_),
    .d(_17410_),
    .o1(_01376_));
 b15nonb02an1n04x5 _27278_ (.a(net866),
    .b(net881),
    .out0(_01377_));
 b15xor002an1n02x5 _27279_ (.a(\us20.a[7] ),
    .b(net878),
    .out0(_01378_));
 b15nand04aq1n08x5 _27280_ (.a(\us20.a[3] ),
    .b(_15943_),
    .c(_01377_),
    .d(_01378_),
    .o1(_01379_));
 b15oai013an1n12x5 _27281_ (.a(_01379_),
    .b(_17458_),
    .c(_16137_),
    .d(_15997_),
    .o1(_01380_));
 b15oai012al1n03x5 _27282_ (.a(_00598_),
    .b(_17432_),
    .c(net865),
    .o1(_01381_));
 b15norp02aq1n03x5 _27283_ (.a(net863),
    .b(_15987_),
    .o1(_01382_));
 b15aoi013ah1n03x5 _27284_ (.a(_01380_),
    .b(_01381_),
    .c(_01382_),
    .d(net876),
    .o1(_01383_));
 b15aoai13ah1n02x5 _27285_ (.a(_01002_),
    .b(_00604_),
    .c(_16047_),
    .d(net872),
    .o1(_01384_));
 b15inv040as1n02x5 _27286_ (.a(net863),
    .o1(_01385_));
 b15nand04ar1n04x5 _27287_ (.a(_01385_),
    .b(_15952_),
    .c(_17493_),
    .d(_17503_),
    .o1(_01386_));
 b15norp03ar1n02x5 _27288_ (.a(_16080_),
    .b(_16113_),
    .c(_15995_),
    .o1(_01387_));
 b15aoi012ar1n02x5 _27289_ (.a(_16134_),
    .b(_15959_),
    .c(net869),
    .o1(_01388_));
 b15aoi013al1n03x5 _27290_ (.a(_01387_),
    .b(_01388_),
    .c(net865),
    .d(_17398_),
    .o1(_01389_));
 b15and003al1n03x5 _27291_ (.a(_01384_),
    .b(_01386_),
    .c(_01389_),
    .o(_01390_));
 b15nand04ah1n12x5 _27292_ (.a(_01370_),
    .b(_01376_),
    .c(_01383_),
    .d(_01390_),
    .o1(_01391_));
 b15nanb02ah1n24x5 _27293_ (.a(net865),
    .b(net877),
    .out0(_01392_));
 b15obai22ar1n02x5 _27294_ (.a(_01382_),
    .b(_01392_),
    .c(net876),
    .d(_16132_),
    .out0(_01393_));
 b15oai012ar1n02x5 _27295_ (.a(_00536_),
    .b(_16000_),
    .c(net882),
    .o1(_01394_));
 b15aoi022an1n02x5 _27296_ (.a(_16078_),
    .b(_01393_),
    .c(_01394_),
    .d(_17509_),
    .o1(_01395_));
 b15orn002al1n08x5 _27297_ (.a(net871),
    .b(net863),
    .o(_01396_));
 b15obai22ah1n04x5 _27298_ (.a(_00586_),
    .b(_17469_),
    .c(_01396_),
    .d(_17503_),
    .out0(_01397_));
 b15aoi022aq1n12x5 _27299_ (.a(net880),
    .b(_00550_),
    .c(_01397_),
    .d(_17463_),
    .o1(_01398_));
 b15oai022an1n08x5 _27300_ (.a(net872),
    .b(_01395_),
    .c(_01398_),
    .d(_15993_),
    .o1(_01399_));
 b15aoi022ar1n02x5 _27301_ (.a(_16078_),
    .b(_17487_),
    .c(_16047_),
    .d(_16028_),
    .o1(_01400_));
 b15oai022ar1n02x5 _27302_ (.a(_16028_),
    .b(_16031_),
    .c(_01400_),
    .d(net882),
    .o1(_01401_));
 b15nandp2ah1n02x5 _27303_ (.a(net876),
    .b(_01401_),
    .o1(_01402_));
 b15oai022al1n02x5 _27304_ (.a(_15995_),
    .b(_17458_),
    .c(_17400_),
    .d(_16040_),
    .o1(_01403_));
 b15nandp2ar1n03x5 _27305_ (.a(net879),
    .b(_01403_),
    .o1(_01404_));
 b15aoi012ah1n02x5 _27306_ (.a(_17449_),
    .b(_17487_),
    .c(net882),
    .o1(_01405_));
 b15oai112aq1n12x5 _27307_ (.a(_01402_),
    .b(_01404_),
    .c(_01405_),
    .d(_00599_),
    .o1(_01406_));
 b15oai012an1n03x5 _27308_ (.a(_16129_),
    .b(_16000_),
    .c(net883),
    .o1(_01407_));
 b15aoi012ah1n04x5 _27309_ (.a(_16028_),
    .b(_17427_),
    .c(_01407_),
    .o1(_01408_));
 b15oai022ar1n02x5 _27310_ (.a(_15987_),
    .b(_15988_),
    .c(_16006_),
    .d(net877),
    .o1(_01409_));
 b15nanb03al1n04x5 _27311_ (.a(net877),
    .b(net880),
    .c(net884),
    .out0(_01410_));
 b15aoai13aq1n02x5 _27312_ (.a(_01409_),
    .b(_00614_),
    .c(_15989_),
    .d(_01410_),
    .o1(_01411_));
 b15mdn022ar1n02x5 _27313_ (.a(_17504_),
    .b(_01392_),
    .o1(_01412_),
    .sa(_17463_));
 b15norp02ar1n02x5 _27314_ (.a(_16010_),
    .b(_17497_),
    .o1(_01413_));
 b15oai012ar1n02x5 _27315_ (.a(_01410_),
    .b(_00535_),
    .c(net884),
    .o1(_01414_));
 b15aoi022an1n04x5 _27316_ (.a(_01412_),
    .b(_01413_),
    .c(_01414_),
    .d(_16058_),
    .o1(_01415_));
 b15nona22an1n05x5 _27317_ (.a(net869),
    .b(net865),
    .c(net863),
    .out0(_01416_));
 b15oai022ar1n02x5 _27318_ (.a(_17504_),
    .b(_17414_),
    .c(_01416_),
    .d(_16011_),
    .o1(_01417_));
 b15aoi013aq1n02x5 _27319_ (.a(net873),
    .b(_01417_),
    .c(net871),
    .d(_15959_),
    .o1(_01418_));
 b15aoi022al1n06x5 _27320_ (.a(_01408_),
    .b(_01411_),
    .c(_01415_),
    .d(_01418_),
    .o1(_01419_));
 b15aoi012ar1n02x5 _27321_ (.a(_16004_),
    .b(_16089_),
    .c(_16077_),
    .o1(_01420_));
 b15aoi012ar1n02x5 _27322_ (.a(_01420_),
    .b(_16010_),
    .c(_17446_),
    .o1(_01421_));
 b15aoi013al1n02x5 _27323_ (.a(_16028_),
    .b(_16045_),
    .c(_00543_),
    .d(net880),
    .o1(_01422_));
 b15oai012al1n02x5 _27324_ (.a(_17446_),
    .b(_15963_),
    .c(_17469_),
    .o1(_01423_));
 b15aoi022al1n04x5 _27325_ (.a(_01421_),
    .b(_01422_),
    .c(_01423_),
    .d(_15948_),
    .o1(_01424_));
 b15orn002as1n04x5 _27326_ (.a(_01419_),
    .b(_01424_),
    .o(_01425_));
 b15nor004as1n12x5 _27327_ (.a(_01391_),
    .b(_01399_),
    .c(_01406_),
    .d(_01425_),
    .o1(_01426_));
 b15xnr002ar1n02x5 _27328_ (.a(_00973_),
    .b(_01426_),
    .out0(_01427_));
 b15xor002an1n02x5 _27329_ (.a(_01364_),
    .b(_01427_),
    .out0(_01428_));
 b15xor002al1n03x5 _27330_ (.a(_01287_),
    .b(_01428_),
    .out0(_01429_));
 b15cmbn22ar1n16x5 _27331_ (.clk1(\text_in_r[36] ),
    .clk2(_01429_),
    .clkout(_01430_),
    .s(net540));
 b15xor002as1n16x5 _27332_ (.a(\u0.w[2][4] ),
    .b(_01430_),
    .out0(_00117_));
 b15inv040as1n03x5 _27333_ (.a(\text_in_r[37] ),
    .o1(_01431_));
 b15oaoi13ar1n02x5 _27334_ (.a(_16100_),
    .b(_15988_),
    .c(_01385_),
    .d(_01392_),
    .o1(_01432_));
 b15oab012ah1n02x5 _27335_ (.a(_01432_),
    .b(_00600_),
    .c(_15993_),
    .out0(_01433_));
 b15aoi013an1n03x5 _27336_ (.a(_16061_),
    .b(_15955_),
    .c(_16065_),
    .d(net872),
    .o1(_01434_));
 b15oai012aq1n04x5 _27337_ (.a(_15959_),
    .b(_17410_),
    .c(_01434_),
    .o1(_01435_));
 b15aob012al1n04x5 _27338_ (.a(net880),
    .b(_16077_),
    .c(_00605_),
    .out0(_01436_));
 b15nona23an1n12x5 _27339_ (.a(_01433_),
    .b(_17463_),
    .c(_01435_),
    .d(_01436_),
    .out0(_01437_));
 b15nand04ar1n02x5 _27340_ (.a(_16028_),
    .b(_15952_),
    .c(_15955_),
    .d(_17410_),
    .o1(_01438_));
 b15oai112ar1n04x5 _27341_ (.a(net882),
    .b(_01438_),
    .c(_17405_),
    .d(_16061_),
    .o1(_01439_));
 b15aoi122ar1n02x5 _27342_ (.a(net882),
    .b(net874),
    .c(_16164_),
    .d(_01014_),
    .e(_16147_),
    .o1(_01440_));
 b15oai013ar1n02x5 _27343_ (.a(_16078_),
    .b(net874),
    .c(_16126_),
    .d(_16113_),
    .o1(_01441_));
 b15norp03ar1n02x5 _27344_ (.a(_16126_),
    .b(_16113_),
    .c(_15995_),
    .o1(_01442_));
 b15norp03ar1n02x5 _27345_ (.a(net874),
    .b(_16126_),
    .c(_16082_),
    .o1(_01443_));
 b15oai013ar1n03x5 _27346_ (.a(_01441_),
    .b(_01442_),
    .c(_01443_),
    .d(_16078_),
    .o1(_01444_));
 b15aob012ar1n02x5 _27347_ (.a(_01439_),
    .b(_01440_),
    .c(_01444_),
    .out0(_01445_));
 b15aoi013ah1n02x5 _27348_ (.a(_16018_),
    .b(_15939_),
    .c(_17457_),
    .d(_15947_),
    .o1(_01446_));
 b15aoi012ar1n02x5 _27349_ (.a(\us20.a[2] ),
    .b(_15952_),
    .c(_15955_),
    .o1(_01447_));
 b15oai013as1n03x5 _27350_ (.a(net874),
    .b(_16006_),
    .c(_01446_),
    .d(_01447_),
    .o1(_01448_));
 b15aoi013an1n03x5 _27351_ (.a(_17476_),
    .b(_17469_),
    .c(_16065_),
    .d(net864),
    .o1(_01449_));
 b15nor004ar1n02x5 _27352_ (.a(net868),
    .b(net870),
    .c(net864),
    .d(net885),
    .o1(_01450_));
 b15aoi012an1n02x5 _27353_ (.a(_01450_),
    .b(_16034_),
    .c(net885),
    .o1(_01451_));
 b15oai022an1n06x5 _27354_ (.a(_01392_),
    .b(_01449_),
    .c(_01451_),
    .d(_16000_),
    .o1(_01452_));
 b15norp03al1n02x5 _27355_ (.a(_16078_),
    .b(_00541_),
    .c(_16010_),
    .o1(_01453_));
 b15nor003al1n08x5 _27356_ (.a(\us20.a[2] ),
    .b(_16080_),
    .c(_16113_),
    .o1(_01454_));
 b15and002ar1n02x5 _27357_ (.a(net875),
    .b(_16034_),
    .o(_01455_));
 b15oab012as1n02x5 _27358_ (.a(_01453_),
    .b(_01454_),
    .c(_01455_),
    .out0(_01456_));
 b15oai013as1n08x5 _27359_ (.a(_01448_),
    .b(_01452_),
    .c(_01456_),
    .d(net874),
    .o1(_01457_));
 b15and003ah1n04x5 _27360_ (.a(_01437_),
    .b(_01445_),
    .c(_01457_),
    .o(_01458_));
 b15aoi022ar1n02x5 _27361_ (.a(_17446_),
    .b(_15974_),
    .c(_17509_),
    .d(net879),
    .o1(_01459_));
 b15nor002ah1n02x5 _27362_ (.a(net882),
    .b(_01459_),
    .o1(_01460_));
 b15aoi112ah1n02x5 _27363_ (.a(net875),
    .b(_16069_),
    .c(_17487_),
    .d(_16078_),
    .o1(_01461_));
 b15aoi112as1n04x5 _27364_ (.a(net872),
    .b(_01461_),
    .c(_17401_),
    .d(net875),
    .o1(_01462_));
 b15oaoi13ah1n08x5 _27365_ (.a(_01460_),
    .b(net882),
    .c(_16075_),
    .d(_01462_),
    .o1(_01463_));
 b15aoai13an1n03x5 _27366_ (.a(_16096_),
    .b(_17457_),
    .c(_00599_),
    .d(_15943_),
    .o1(_01464_));
 b15aoai13an1n03x5 _27367_ (.a(net885),
    .b(net874),
    .c(_16096_),
    .d(_17457_),
    .o1(_01465_));
 b15aoi112ar1n06x5 _27368_ (.a(\us20.a[2] ),
    .b(_01464_),
    .c(_01465_),
    .d(\us20.a[1] ),
    .o1(_01466_));
 b15oaoi13aq1n04x5 _27369_ (.a(net883),
    .b(_17520_),
    .c(_16134_),
    .d(_16078_),
    .o1(_01467_));
 b15aoi012ar1n04x5 _27370_ (.a(net880),
    .b(_16137_),
    .c(_01025_),
    .o1(_01468_));
 b15oai012al1n12x5 _27371_ (.a(_16045_),
    .b(_01467_),
    .c(_01468_),
    .o1(_01469_));
 b15oab012ar1n02x5 _27372_ (.a(net883),
    .b(_16034_),
    .c(_16047_),
    .out0(_01470_));
 b15aoai13ar1n02x5 _27373_ (.a(_15974_),
    .b(_01470_),
    .c(net880),
    .d(_16034_),
    .o1(_01471_));
 b15nona23as1n04x5 _27374_ (.a(_01466_),
    .b(_16014_),
    .c(_01469_),
    .d(_01471_),
    .out0(_01472_));
 b15oai112aq1n02x5 _27375_ (.a(net872),
    .b(_16129_),
    .c(_16068_),
    .d(_16069_),
    .o1(_01473_));
 b15nor003aq1n06x5 _27376_ (.a(_17463_),
    .b(_16092_),
    .c(_01038_),
    .o1(_01474_));
 b15nand03aq1n03x5 _27377_ (.a(net871),
    .b(net863),
    .c(net877),
    .o1(_01475_));
 b15oai012aq1n08x5 _27378_ (.a(_01475_),
    .b(_01396_),
    .c(net877),
    .o1(_01476_));
 b15oai013aq1n06x5 _27379_ (.a(_00589_),
    .b(_16082_),
    .c(_16080_),
    .d(net877),
    .o1(_01477_));
 b15aoi122ah1n08x5 _27380_ (.a(_17434_),
    .b(_01474_),
    .c(_01476_),
    .d(_01477_),
    .e(_17447_),
    .o1(_01478_));
 b15norp02ar1n03x5 _27381_ (.a(_15993_),
    .b(_16060_),
    .o1(_01479_));
 b15norp03aq1n03x5 _27382_ (.a(_15987_),
    .b(_16021_),
    .c(_15995_),
    .o1(_01480_));
 b15norp02an1n03x5 _27383_ (.a(net873),
    .b(_16060_),
    .o1(_01481_));
 b15oaoi13al1n04x5 _27384_ (.a(_01479_),
    .b(_15959_),
    .c(_01480_),
    .d(_01481_),
    .o1(_01482_));
 b15oai112aq1n08x5 _27385_ (.a(_01473_),
    .b(_01478_),
    .c(_16078_),
    .d(_01482_),
    .o1(_01483_));
 b15aoi012ar1n02x5 _27386_ (.a(_16125_),
    .b(_15947_),
    .c(_16018_),
    .o1(_01484_));
 b15norp03ar1n04x5 _27387_ (.a(_16028_),
    .b(_01454_),
    .c(_01484_),
    .o1(_01485_));
 b15nand03an1n16x5 _27388_ (.a(_16078_),
    .b(_15952_),
    .c(_15955_),
    .o1(_01486_));
 b15aob012aq1n02x5 _27389_ (.a(_16010_),
    .b(_01486_),
    .c(_16031_),
    .out0(_01487_));
 b15oab012aq1n02x5 _27390_ (.a(_16033_),
    .b(_16135_),
    .c(_16077_),
    .out0(_01488_));
 b15oai112an1n12x5 _27391_ (.a(_01485_),
    .b(_01487_),
    .c(_16078_),
    .d(_01488_),
    .o1(_01489_));
 b15norp03an1n02x5 _27392_ (.a(_16018_),
    .b(_15987_),
    .c(_15988_),
    .o1(_01490_));
 b15oaoi13aq1n03x5 _27393_ (.a(net872),
    .b(net880),
    .c(_01490_),
    .d(_16068_),
    .o1(_01491_));
 b15oai022ah1n02x5 _27394_ (.a(_16129_),
    .b(_15988_),
    .c(_17415_),
    .d(net865),
    .o1(_01492_));
 b15aoai13ar1n06x5 _27395_ (.a(_16018_),
    .b(_16047_),
    .c(_01492_),
    .d(_16065_),
    .o1(_01493_));
 b15nandp2ar1n04x5 _27396_ (.a(_16078_),
    .b(_16047_),
    .o1(_01494_));
 b15nano22ah1n03x5 _27397_ (.a(_01494_),
    .b(net883),
    .c(_16084_),
    .out0(_01495_));
 b15nor002al1n06x5 _27398_ (.a(_16078_),
    .b(_16132_),
    .o1(_01496_));
 b15aoi112ah1n03x5 _27399_ (.a(net883),
    .b(_01496_),
    .c(_15963_),
    .d(_17446_),
    .o1(_01497_));
 b15oai112al1n12x5 _27400_ (.a(_01491_),
    .b(_01493_),
    .c(_01495_),
    .d(_01497_),
    .o1(_01498_));
 b15aoi112as1n08x5 _27401_ (.a(_01472_),
    .b(_01483_),
    .c(_01489_),
    .d(_01498_),
    .o1(_01499_));
 b15nandp3as1n24x5 _27402_ (.a(_01458_),
    .b(_01463_),
    .c(_01499_),
    .o1(_01500_));
 b15oaoi13an1n04x5 _27403_ (.a(net759),
    .b(net764),
    .c(net763),
    .d(_01079_),
    .o1(_01501_));
 b15aob012ar1n04x5 _27404_ (.a(net764),
    .b(_16774_),
    .c(_01305_),
    .out0(_01502_));
 b15aoi122as1n06x5 _27405_ (.a(_01501_),
    .b(_01305_),
    .c(_16790_),
    .d(net763),
    .e(_01502_),
    .o1(_01503_));
 b15nandp3ar1n02x5 _27406_ (.a(net763),
    .b(_16898_),
    .c(_16905_),
    .o1(_01504_));
 b15oai112al1n04x5 _27407_ (.a(net755),
    .b(_01504_),
    .c(_16898_),
    .d(_17314_),
    .o1(_01505_));
 b15aoai13ar1n02x5 _27408_ (.a(net766),
    .b(_00735_),
    .c(_16764_),
    .d(net759),
    .o1(_01506_));
 b15oai012ar1n02x5 _27409_ (.a(_16764_),
    .b(_17335_),
    .c(_16786_),
    .o1(_01507_));
 b15aoi012ar1n02x5 _27410_ (.a(_01505_),
    .b(_01506_),
    .c(_01507_),
    .o1(_01508_));
 b15nand02al1n12x5 _27411_ (.a(net766),
    .b(_16915_),
    .o1(_01509_));
 b15nandp2al1n03x5 _27412_ (.a(_16915_),
    .b(_16898_),
    .o1(_01510_));
 b15oai012aq1n04x5 _27413_ (.a(_16760_),
    .b(_16905_),
    .c(_16693_),
    .o1(_01511_));
 b15aoi222al1n08x5 _27414_ (.a(_01509_),
    .b(_00735_),
    .c(_01510_),
    .d(_17373_),
    .e(_16770_),
    .f(_01511_),
    .o1(_01512_));
 b15oab012as1n04x5 _27415_ (.a(_01508_),
    .b(_01512_),
    .c(net755),
    .out0(_01513_));
 b15oai112aq1n02x5 _27416_ (.a(_16785_),
    .b(_16726_),
    .c(_16860_),
    .d(net761),
    .o1(_01514_));
 b15oai112aq1n02x5 _27417_ (.a(_16702_),
    .b(_16708_),
    .c(_16894_),
    .d(net758),
    .o1(_01515_));
 b15mdn022ah1n03x5 _27418_ (.a(_01514_),
    .b(_01515_),
    .o1(_01516_),
    .sa(net754));
 b15nand03an1n02x5 _27419_ (.a(_16783_),
    .b(_16789_),
    .c(_16813_),
    .o1(_01517_));
 b15oai013as1n06x5 _27420_ (.a(_01517_),
    .b(_01308_),
    .c(_16867_),
    .d(_16907_),
    .o1(_01518_));
 b15nand03aq1n03x5 _27421_ (.a(_16873_),
    .b(_16806_),
    .c(_16894_),
    .o1(_01519_));
 b15nand03an1n02x5 _27422_ (.a(_16742_),
    .b(_17390_),
    .c(_00735_),
    .o1(_01520_));
 b15nand02an1n02x5 _27423_ (.a(_16830_),
    .b(_16783_),
    .o1(_01521_));
 b15aoi022ar1n04x5 _27424_ (.a(_16702_),
    .b(_16746_),
    .c(_16831_),
    .d(net754),
    .o1(_01522_));
 b15oai112aq1n08x5 _27425_ (.a(_01519_),
    .b(_01520_),
    .c(_01521_),
    .d(_01522_),
    .o1(_01523_));
 b15norp02aq1n02x5 _27426_ (.a(_17314_),
    .b(_16761_),
    .o1(_01524_));
 b15nor004as1n06x5 _27427_ (.a(_01516_),
    .b(_01518_),
    .c(_01523_),
    .d(_01524_),
    .o1(_01525_));
 b15norp02aq1n03x5 _27428_ (.a(_17389_),
    .b(_16849_),
    .o1(_01526_));
 b15oai112an1n02x5 _27429_ (.a(_16741_),
    .b(_16852_),
    .c(_01526_),
    .d(_17383_),
    .o1(_01527_));
 b15norp03ar1n02x5 _27430_ (.a(_17389_),
    .b(_16849_),
    .c(_16728_),
    .o1(_01528_));
 b15oai012al1n03x5 _27431_ (.a(net760),
    .b(_16851_),
    .c(_01528_),
    .o1(_01529_));
 b15nand02al1n03x5 _27432_ (.a(net748),
    .b(_16852_),
    .o1(_01530_));
 b15nand03aq1n02x5 _27433_ (.a(net750),
    .b(_01127_),
    .c(_16844_),
    .o1(_01531_));
 b15nandp2an1n08x5 _27434_ (.a(_16731_),
    .b(_16798_),
    .o1(_01532_));
 b15oaoi13as1n04x5 _27435_ (.a(_01530_),
    .b(_01531_),
    .c(_17297_),
    .d(_01532_),
    .o1(_01533_));
 b15orn003an1n04x5 _27436_ (.a(_16728_),
    .b(_00789_),
    .c(_01119_),
    .o(_01534_));
 b15nand04as1n06x5 _27437_ (.a(_16907_),
    .b(_16785_),
    .c(_16726_),
    .d(_16861_),
    .o1(_01535_));
 b15oai112as1n16x5 _27438_ (.a(_01534_),
    .b(_01535_),
    .c(_01360_),
    .d(_16908_),
    .o1(_01536_));
 b15nano23an1n08x5 _27439_ (.a(_01527_),
    .b(_01529_),
    .c(_01533_),
    .d(_01536_),
    .out0(_01537_));
 b15aoi022an1n02x5 _27440_ (.a(net761),
    .b(_16798_),
    .c(_16763_),
    .d(net765),
    .o1(_01538_));
 b15oaoi13an1n08x5 _27441_ (.a(_17371_),
    .b(_01538_),
    .c(_16798_),
    .d(_17367_),
    .o1(_01539_));
 b15nandp2aq1n04x5 _27442_ (.a(_16758_),
    .b(_17287_),
    .o1(_01540_));
 b15oaoi13an1n08x5 _27443_ (.a(net754),
    .b(_01540_),
    .c(_00730_),
    .d(_16760_),
    .o1(_01541_));
 b15aoi012ar1n02x5 _27444_ (.a(net761),
    .b(_16728_),
    .c(_16760_),
    .o1(_01542_));
 b15oab012as1n03x5 _27445_ (.a(_16793_),
    .b(_16844_),
    .c(_01542_),
    .out0(_01543_));
 b15nanb02aq1n06x5 _27446_ (.a(net752),
    .b(net757),
    .out0(_01544_));
 b15aoi022al1n02x5 _27447_ (.a(_16710_),
    .b(_16873_),
    .c(_16870_),
    .d(_16726_),
    .o1(_01545_));
 b15nor002ah1n04x5 _27448_ (.a(_01544_),
    .b(_01545_),
    .o1(_01546_));
 b15nor004ah1n12x5 _27449_ (.a(_01539_),
    .b(_01541_),
    .c(_01543_),
    .d(_01546_),
    .o1(_01547_));
 b15nand04as1n16x5 _27450_ (.a(_00736_),
    .b(_01525_),
    .c(_01537_),
    .d(_01547_),
    .o1(_01548_));
 b15nand02ar1n02x5 _27451_ (.a(_16888_),
    .b(_16897_),
    .o1(_01549_));
 b15aoai13ar1n02x5 _27452_ (.a(net763),
    .b(net759),
    .c(_16888_),
    .d(net766),
    .o1(_01550_));
 b15nand04as1n04x5 _27453_ (.a(net755),
    .b(_17367_),
    .c(_01549_),
    .d(_01550_),
    .o1(_01551_));
 b15oai112al1n08x5 _27454_ (.a(_16770_),
    .b(_16856_),
    .c(_16839_),
    .d(_16693_),
    .o1(_01552_));
 b15oai112an1n08x5 _27455_ (.a(_17303_),
    .b(_01552_),
    .c(_16844_),
    .d(_16770_),
    .o1(_01553_));
 b15norp02ar1n03x5 _27456_ (.a(net766),
    .b(_16897_),
    .o1(_01554_));
 b15aoi022as1n08x5 _27457_ (.a(_16768_),
    .b(_00773_),
    .c(_01554_),
    .d(_16798_),
    .o1(_01555_));
 b15oai112al1n16x5 _27458_ (.a(_01551_),
    .b(_01553_),
    .c(_01555_),
    .d(_16770_),
    .o1(_01556_));
 b15nor004as1n12x5 _27459_ (.a(_01503_),
    .b(_01513_),
    .c(_01548_),
    .d(_01556_),
    .o1(_01557_));
 b15xor002ah1n03x5 _27460_ (.a(_01209_),
    .b(_01557_),
    .out0(_01558_));
 b15xor002al1n08x5 _27461_ (.a(_01500_),
    .b(_01558_),
    .out0(_01559_));
 b15aoai13an1n02x5 _27462_ (.a(net604),
    .b(_16473_),
    .c(_16640_),
    .d(_16605_),
    .o1(_01560_));
 b15nonb02ah1n12x5 _27463_ (.a(net599),
    .b(\us13.a[2] ),
    .out0(_01561_));
 b15nand02an1n03x5 _27464_ (.a(_16458_),
    .b(_01561_),
    .o1(_01562_));
 b15aoai13an1n03x5 _27465_ (.a(_16558_),
    .b(net607),
    .c(_01560_),
    .d(_01562_),
    .o1(_01563_));
 b15oai112ar1n12x5 _27466_ (.a(net616),
    .b(_01563_),
    .c(_17077_),
    .d(_16558_),
    .o1(_01564_));
 b15nand03al1n03x5 _27467_ (.a(net612),
    .b(_16577_),
    .c(_16517_),
    .o1(_01565_));
 b15nand02ar1n02x5 _27468_ (.a(_17125_),
    .b(_01565_),
    .o1(_01566_));
 b15nand03ar1n02x5 _27469_ (.a(_16508_),
    .b(_17088_),
    .c(_01566_),
    .o1(_01567_));
 b15oai112al1n04x5 _27470_ (.a(_01564_),
    .b(_01567_),
    .c(_16576_),
    .d(_17088_),
    .o1(_01568_));
 b15oai012ar1n02x5 _27471_ (.a(net608),
    .b(_17085_),
    .c(_16508_),
    .o1(_01569_));
 b15oai022ar1n24x5 _27472_ (.a(net618),
    .b(_16667_),
    .c(_16549_),
    .d(_17574_),
    .o1(_01570_));
 b15aoi013al1n03x5 _27473_ (.a(_01569_),
    .b(_01570_),
    .c(net612),
    .d(_16475_),
    .o1(_01571_));
 b15oaoi13an1n02x5 _27474_ (.a(net620),
    .b(_17085_),
    .c(_17578_),
    .d(_17602_),
    .o1(_01572_));
 b15nandp2ar1n02x5 _27475_ (.a(_16576_),
    .b(_01565_),
    .o1(_01573_));
 b15aoi013al1n03x5 _27476_ (.a(_01572_),
    .b(_01573_),
    .c(_17602_),
    .d(net620),
    .o1(_01574_));
 b15aboi22aq1n08x5 _27477_ (.a(_01568_),
    .b(_16466_),
    .c(_01571_),
    .d(_01574_),
    .out0(_01575_));
 b15aoi022ar1n04x5 _27478_ (.a(net615),
    .b(_16650_),
    .c(_00847_),
    .d(_17562_),
    .o1(_01576_));
 b15and002aq1n02x5 _27479_ (.a(_16659_),
    .b(_17179_),
    .o(_01577_));
 b15aoi012ar1n06x5 _27480_ (.a(_01577_),
    .b(_16446_),
    .c(net606),
    .o1(_01578_));
 b15oai112an1n08x5 _27481_ (.a(_16558_),
    .b(_01576_),
    .c(_01578_),
    .d(_17139_),
    .o1(_01579_));
 b15nand02al1n08x5 _27482_ (.a(_16466_),
    .b(_16577_),
    .o1(_01580_));
 b15oaoi13as1n08x5 _27483_ (.a(_16497_),
    .b(_01580_),
    .c(_16626_),
    .d(_16432_),
    .o1(_01581_));
 b15oai012as1n03x5 _27484_ (.a(_01579_),
    .b(_01581_),
    .c(_16558_),
    .o1(_01582_));
 b15oai122an1n02x5 _27485_ (.a(_16508_),
    .b(net608),
    .c(_17091_),
    .d(_16680_),
    .e(_16498_),
    .o1(_01583_));
 b15aob012an1n03x5 _27486_ (.a(_01583_),
    .b(_16608_),
    .c(net616),
    .out0(_01584_));
 b15aoi013as1n04x5 _27487_ (.a(net612),
    .b(_01277_),
    .c(_01582_),
    .d(_01584_),
    .o1(_01585_));
 b15nand02ar1n02x5 _27488_ (.a(_16518_),
    .b(_16579_),
    .o1(_01586_));
 b15oaoi13al1n02x5 _27489_ (.a(_16518_),
    .b(net601),
    .c(net597),
    .d(_00902_),
    .o1(_01587_));
 b15oai013as1n03x5 _27490_ (.a(_01586_),
    .b(_01587_),
    .c(net612),
    .d(_16538_),
    .o1(_01588_));
 b15aoi022ar1n02x5 _27491_ (.a(_16490_),
    .b(_16519_),
    .c(_16521_),
    .d(_16508_),
    .o1(_01589_));
 b15oai012aq1n03x5 _27492_ (.a(_01588_),
    .b(_01589_),
    .c(net612),
    .o1(_01590_));
 b15nandp3ar1n02x5 _27493_ (.a(net616),
    .b(_16466_),
    .c(_01224_),
    .o1(_01591_));
 b15oai112ar1n04x5 _27494_ (.a(net620),
    .b(_01591_),
    .c(_17131_),
    .d(_17175_),
    .o1(_01592_));
 b15oai022ar1n02x5 _27495_ (.a(_16479_),
    .b(_17183_),
    .c(_17131_),
    .d(_17602_),
    .o1(_01593_));
 b15oai012aq1n04x5 _27496_ (.a(_01592_),
    .b(_01593_),
    .c(net620),
    .o1(_01594_));
 b15oai122as1n02x5 _27497_ (.a(_01277_),
    .b(_00900_),
    .c(_16524_),
    .d(net612),
    .e(_16519_),
    .o1(_01595_));
 b15aoi013an1n04x5 _27498_ (.a(_01595_),
    .b(_16601_),
    .c(_16652_),
    .d(_16475_),
    .o1(_01596_));
 b15oai112an1n12x5 _27499_ (.a(_01590_),
    .b(_01594_),
    .c(_01596_),
    .d(net620),
    .o1(_01597_));
 b15oaoi13ar1n04x5 _27500_ (.a(net610),
    .b(_17119_),
    .c(_16521_),
    .d(net620),
    .o1(_01598_));
 b15oai013as1n03x5 _27501_ (.a(net616),
    .b(_16466_),
    .c(_16516_),
    .d(_17116_),
    .o1(_01599_));
 b15oab012as1n02x5 _27502_ (.a(_16536_),
    .b(_17076_),
    .c(_17117_),
    .out0(_01600_));
 b15oai013ah1n06x5 _27503_ (.a(_16508_),
    .b(net610),
    .c(_17565_),
    .d(_17116_),
    .o1(_01601_));
 b15oai022ah1n08x5 _27504_ (.a(_01598_),
    .b(_01599_),
    .c(_01600_),
    .d(_01601_),
    .o1(_01602_));
 b15nand03aq1n03x5 _27505_ (.a(_16558_),
    .b(_00823_),
    .c(_00851_),
    .o1(_01603_));
 b15oai012ar1n02x5 _27506_ (.a(_01603_),
    .b(_16504_),
    .c(_16498_),
    .o1(_01604_));
 b15aoi022ar1n02x5 _27507_ (.a(_16619_),
    .b(_01581_),
    .c(_01604_),
    .d(_17087_),
    .o1(_01605_));
 b15oai012ar1n02x5 _27508_ (.a(_16674_),
    .b(_16646_),
    .c(_16453_),
    .o1(_01606_));
 b15oaoi13ah1n02x5 _27509_ (.a(_16522_),
    .b(_01606_),
    .c(_00900_),
    .d(_16435_),
    .o1(_01607_));
 b15oai112ah1n16x5 _27510_ (.a(_16597_),
    .b(_01264_),
    .c(_16456_),
    .d(_01215_),
    .o1(_01608_));
 b15nand03an1n04x5 _27511_ (.a(_16475_),
    .b(_16601_),
    .c(_16613_),
    .o1(_01609_));
 b15nand03aq1n04x5 _27512_ (.a(net619),
    .b(_17128_),
    .c(_16524_),
    .o1(_01610_));
 b15nand04an1n12x5 _27513_ (.a(_17536_),
    .b(_01608_),
    .c(_01609_),
    .d(_01610_),
    .o1(_01611_));
 b15nano23al1n05x5 _27514_ (.a(_01602_),
    .b(_01605_),
    .c(_01607_),
    .d(_01611_),
    .out0(_01612_));
 b15aoai13ar1n02x5 _27515_ (.a(_16466_),
    .b(_16643_),
    .c(_16453_),
    .d(net612),
    .o1(_01613_));
 b15aoi022aq1n02x5 _27516_ (.a(_16597_),
    .b(_16481_),
    .c(_16517_),
    .d(_17545_),
    .o1(_01614_));
 b15oai022ar1n02x5 _27517_ (.a(_16558_),
    .b(_16643_),
    .c(_01614_),
    .d(net597),
    .o1(_01615_));
 b15aoi012al1n02x5 _27518_ (.a(_01613_),
    .b(_01615_),
    .c(_16508_),
    .o1(_01616_));
 b15norp03al1n02x5 _27519_ (.a(net612),
    .b(_16439_),
    .c(_01239_),
    .o1(_01617_));
 b15aoi013an1n03x5 _27520_ (.a(_01617_),
    .b(_01224_),
    .c(_16585_),
    .d(net612),
    .o1(_01618_));
 b15aoai13ah1n04x5 _27521_ (.a(_01612_),
    .b(_01616_),
    .c(_01618_),
    .d(net608),
    .o1(_01619_));
 b15nor004as1n12x5 _27522_ (.a(_01575_),
    .b(_01585_),
    .c(_01597_),
    .d(_01619_),
    .o1(_01620_));
 b15norp02ar1n02x5 _27523_ (.a(_16936_),
    .b(_01146_),
    .o1(_01621_));
 b15oai112ar1n02x5 _27524_ (.a(_16258_),
    .b(_16328_),
    .c(_16960_),
    .d(_16390_),
    .o1(_01622_));
 b15oai013aq1n02x5 _27525_ (.a(_01622_),
    .b(_16960_),
    .c(_16282_),
    .d(_16390_),
    .o1(_01623_));
 b15aoai13ah1n03x5 _27526_ (.a(net734),
    .b(_01621_),
    .c(_01623_),
    .d(net732),
    .o1(_01624_));
 b15nand03ah1n04x5 _27527_ (.a(net732),
    .b(_16965_),
    .c(_16315_),
    .o1(_01625_));
 b15xnr002al1n06x5 _27528_ (.a(net722),
    .b(net720),
    .out0(_01626_));
 b15aoai13aq1n02x5 _27529_ (.a(_16289_),
    .b(_16936_),
    .c(_01626_),
    .d(_17055_),
    .o1(_01627_));
 b15aoi022ar1n04x5 _27530_ (.a(net738),
    .b(_17031_),
    .c(_01626_),
    .d(net740),
    .o1(_01628_));
 b15oai022al1n06x5 _27531_ (.a(_16278_),
    .b(_16314_),
    .c(_01628_),
    .d(net716),
    .o1(_01629_));
 b15nanb02aq1n12x5 _27532_ (.a(_01627_),
    .b(_01629_),
    .out0(_01630_));
 b15aoai13al1n08x5 _27533_ (.a(_01624_),
    .b(net734),
    .c(_01625_),
    .d(_01630_),
    .o1(_01631_));
 b15oai022ah1n12x5 _27534_ (.a(net717),
    .b(_16237_),
    .c(_17015_),
    .d(_17022_),
    .o1(_01632_));
 b15nandp3al1n04x5 _27535_ (.a(_16305_),
    .b(_16233_),
    .c(_01632_),
    .o1(_01633_));
 b15aoi012ar1n02x5 _27536_ (.a(net739),
    .b(_16221_),
    .c(_16361_),
    .o1(_01634_));
 b15aoai13ar1n02x5 _27537_ (.a(_16340_),
    .b(_01634_),
    .c(_16957_),
    .d(\us02.a[0] ),
    .o1(_01635_));
 b15oa0022ar1n02x5 _27538_ (.a(net730),
    .b(_16391_),
    .c(_17258_),
    .d(_16347_),
    .o(_01636_));
 b15oai112aq1n04x5 _27539_ (.a(_01633_),
    .b(_01635_),
    .c(_01636_),
    .d(net734),
    .o1(_01637_));
 b15norp02ar1n02x5 _27540_ (.a(_16388_),
    .b(_17258_),
    .o1(_01638_));
 b15oai013ar1n02x5 _27541_ (.a(net742),
    .b(_17206_),
    .c(_00663_),
    .d(_01638_),
    .o1(_01639_));
 b15nand03ar1n03x5 _27542_ (.a(_16367_),
    .b(_16416_),
    .c(_16988_),
    .o1(_01640_));
 b15oai112as1n04x5 _27543_ (.a(_01639_),
    .b(_01640_),
    .c(_16383_),
    .d(_16318_),
    .o1(_01641_));
 b15aoi022ar1n02x5 _27544_ (.a(_16233_),
    .b(_16416_),
    .c(_17008_),
    .d(_16226_),
    .o1(_01642_));
 b15oai022ar1n02x5 _27545_ (.a(_16361_),
    .b(_16389_),
    .c(_01642_),
    .d(\us02.a[0] ),
    .o1(_01643_));
 b15nandp2al1n03x5 _27546_ (.a(net739),
    .b(_01643_),
    .o1(_01644_));
 b15aoi122an1n08x5 _27547_ (.a(net738),
    .b(_16181_),
    .c(_16418_),
    .d(_00927_),
    .e(_16193_),
    .o1(_01645_));
 b15oai112an1n04x5 _27548_ (.a(net716),
    .b(_16224_),
    .c(_17224_),
    .d(_16305_),
    .o1(_01646_));
 b15aoi012al1n04x5 _27549_ (.a(_01645_),
    .b(_01646_),
    .c(net738),
    .o1(_01647_));
 b15nandp3ar1n02x5 _27550_ (.a(net739),
    .b(_16224_),
    .c(_16229_),
    .o1(_01648_));
 b15aoi012an1n02x5 _27551_ (.a(_16221_),
    .b(_16260_),
    .c(_01648_),
    .o1(_01649_));
 b15aoi012ar1n02x5 _27552_ (.a(_16367_),
    .b(_16260_),
    .c(_16231_),
    .o1(_01650_));
 b15oai013an1n06x5 _27553_ (.a(net730),
    .b(_01647_),
    .c(_01649_),
    .d(_01650_),
    .o1(_01651_));
 b15nona23an1n12x5 _27554_ (.a(_01637_),
    .b(_01641_),
    .c(_01644_),
    .d(_01651_),
    .out0(_01652_));
 b15nanb02al1n16x5 _27555_ (.a(_00644_),
    .b(_16419_),
    .out0(_01653_));
 b15aoi012ar1n02x5 _27556_ (.a(net732),
    .b(_16214_),
    .c(_16332_),
    .o1(_01654_));
 b15nandp3ar1n03x5 _27557_ (.a(_16326_),
    .b(_01653_),
    .c(_01654_),
    .o1(_01655_));
 b15oaoi13ar1n02x5 _27558_ (.a(net742),
    .b(_16231_),
    .c(_16383_),
    .d(net734),
    .o1(_01656_));
 b15norp02ar1n02x5 _27559_ (.a(net742),
    .b(_16340_),
    .o1(_01657_));
 b15aoi022ar1n02x5 _27560_ (.a(net742),
    .b(_16383_),
    .c(_01653_),
    .d(_01657_),
    .o1(_01658_));
 b15oai122as1n04x5 _27561_ (.a(net739),
    .b(_01655_),
    .c(_01656_),
    .d(_01658_),
    .e(_16226_),
    .o1(_01659_));
 b15aoi012ar1n02x5 _27562_ (.a(net741),
    .b(net732),
    .c(_16336_),
    .o1(_01660_));
 b15aoi012ar1n02x5 _27563_ (.a(_16958_),
    .b(_16323_),
    .c(net739),
    .o1(_01661_));
 b15oai022as1n02x5 _27564_ (.a(_01149_),
    .b(_17225_),
    .c(_01660_),
    .d(_01661_),
    .o1(_01662_));
 b15norp02ar1n02x5 _27565_ (.a(_16979_),
    .b(_00930_),
    .o1(_01663_));
 b15aoi012ar1n02x5 _27566_ (.a(_01663_),
    .b(_17251_),
    .c(_16997_),
    .o1(_01664_));
 b15orn002ah1n04x5 _27567_ (.a(_16966_),
    .b(_01664_),
    .o(_01665_));
 b15aoai13as1n04x5 _27568_ (.a(_01659_),
    .b(net734),
    .c(_01662_),
    .d(_01665_),
    .o1(_01666_));
 b15xor002al1n03x5 _27569_ (.a(\us02.a[0] ),
    .b(net728),
    .out0(_01667_));
 b15nona23al1n02x5 _27570_ (.a(_16979_),
    .b(_01667_),
    .c(_16405_),
    .d(_16278_),
    .out0(_01668_));
 b15aoi013an1n02x5 _27571_ (.a(net729),
    .b(_16202_),
    .c(_16293_),
    .d(_16960_),
    .o1(_01669_));
 b15aoai13ar1n03x5 _27572_ (.a(_16224_),
    .b(_16223_),
    .c(_16311_),
    .d(_16229_),
    .o1(_01670_));
 b15oai112ah1n04x5 _27573_ (.a(_01668_),
    .b(_01669_),
    .c(net738),
    .d(_01670_),
    .o1(_01671_));
 b15aoai13aq1n06x5 _27574_ (.a(_00942_),
    .b(_00912_),
    .c(_17260_),
    .d(net740),
    .o1(_01672_));
 b15orn003ar1n04x5 _27575_ (.a(net740),
    .b(_16237_),
    .c(_16939_),
    .o(_01673_));
 b15aoi112ar1n08x5 _27576_ (.a(_16248_),
    .b(net716),
    .c(_01672_),
    .d(_01673_),
    .o1(_01674_));
 b15nand02ah1n06x5 _27577_ (.a(net739),
    .b(_16248_),
    .o1(_01675_));
 b15aoai13an1n08x5 _27578_ (.a(\us02.a[3] ),
    .b(_16389_),
    .c(_01675_),
    .d(\us02.a[0] ),
    .o1(_01676_));
 b15nandp3ar1n02x5 _27579_ (.a(net734),
    .b(_16301_),
    .c(_16328_),
    .o1(_01677_));
 b15oaoi13aq1n03x5 _27580_ (.a(net738),
    .b(_01677_),
    .c(_01653_),
    .d(_16283_),
    .o1(_01678_));
 b15oai022ah1n06x5 _27581_ (.a(_01671_),
    .b(_01674_),
    .c(_01676_),
    .d(_01678_),
    .o1(_01679_));
 b15aoi122ar1n06x5 _27582_ (.a(net730),
    .b(_16181_),
    .c(_16418_),
    .d(_16343_),
    .e(net734),
    .o1(_01680_));
 b15aoi112al1n02x5 _27583_ (.a(net720),
    .b(_00696_),
    .c(net734),
    .d(net725),
    .o1(_01681_));
 b15oab012ah1n06x5 _27584_ (.a(_01680_),
    .b(_01681_),
    .c(_16226_),
    .out0(_01682_));
 b15oai012an1n02x5 _27585_ (.a(_16401_),
    .b(_16231_),
    .c(net734),
    .o1(_01683_));
 b15aoi013ah1n03x5 _27586_ (.a(_16283_),
    .b(_16972_),
    .c(_01682_),
    .d(_01683_),
    .o1(_01684_));
 b15nandp3ar1n02x5 _27587_ (.a(_16226_),
    .b(_16230_),
    .c(_16356_),
    .o1(_01685_));
 b15oai012aq1n02x5 _27588_ (.a(_01685_),
    .b(_16237_),
    .c(_16226_),
    .o1(_01686_));
 b15aoi012ar1n04x5 _27589_ (.a(_01682_),
    .b(_01686_),
    .c(_16223_),
    .o1(_01687_));
 b15oai012al1n12x5 _27590_ (.a(_01679_),
    .b(_01684_),
    .c(_01687_),
    .o1(_01688_));
 b15nor004as1n12x5 _27591_ (.a(_01631_),
    .b(_01652_),
    .c(_01666_),
    .d(_01688_),
    .o1(_01689_));
 b15xnr002an1n16x5 _27592_ (.a(_01620_),
    .b(_01689_),
    .out0(_01690_));
 b15xor002as1n03x5 _27593_ (.a(_01559_),
    .b(_01690_),
    .out0(_01691_));
 b15mdn022as1n08x5 _27594_ (.a(_01431_),
    .b(_01691_),
    .o1(_01692_),
    .sa(net540));
 b15xor002as1n16x5 _27595_ (.a(\u0.w[2][5] ),
    .b(_01692_),
    .out0(_00118_));
 b15inv040ah1n02x5 _27596_ (.a(\text_in_r[38] ),
    .o1(_01693_));
 b15nor003aq1n02x5 _27597_ (.a(net750),
    .b(_16839_),
    .c(_01355_),
    .o1(_01694_));
 b15and003ar1n02x5 _27598_ (.a(net753),
    .b(net748),
    .c(_16861_),
    .o(_01695_));
 b15aoai13as1n04x5 _27599_ (.a(_01104_),
    .b(_01694_),
    .c(_01695_),
    .d(net750),
    .o1(_01696_));
 b15aoai13al1n04x5 _27600_ (.a(_16798_),
    .b(_01526_),
    .c(_16902_),
    .d(net767),
    .o1(_01697_));
 b15oai012ah1n04x5 _27601_ (.a(_01696_),
    .b(_01697_),
    .c(net760),
    .o1(_01698_));
 b15nor003ah1n04x5 _27602_ (.a(_17345_),
    .b(_01536_),
    .c(_01698_),
    .o1(_01699_));
 b15aoai13ah1n02x5 _27603_ (.a(net760),
    .b(net756),
    .c(_16774_),
    .d(_17337_),
    .o1(_01700_));
 b15aoi012al1n02x5 _27604_ (.a(_16741_),
    .b(net757),
    .c(_17337_),
    .o1(_01701_));
 b15nor002as1n04x5 _27605_ (.a(net765),
    .b(_00708_),
    .o1(_01702_));
 b15aoai13as1n02x5 _27606_ (.a(_16774_),
    .b(_01702_),
    .c(_01124_),
    .d(net767),
    .o1(_01703_));
 b15aoi012ar1n06x5 _27607_ (.a(_01700_),
    .b(_01701_),
    .c(_01703_),
    .o1(_01704_));
 b15aoi013ar1n02x5 _27608_ (.a(_16851_),
    .b(_17337_),
    .c(_16693_),
    .d(_16844_),
    .o1(_01705_));
 b15norp02al1n04x5 _27609_ (.a(net760),
    .b(_01705_),
    .o1(_01706_));
 b15aob012an1n02x5 _27610_ (.a(_16815_),
    .b(_16832_),
    .c(_17373_),
    .out0(_01707_));
 b15oaoi13ah1n04x5 _27611_ (.a(_00781_),
    .b(_01707_),
    .c(net765),
    .d(_17320_),
    .o1(_01708_));
 b15nor004al1n08x5 _27612_ (.a(_16910_),
    .b(_01704_),
    .c(_01706_),
    .d(_01708_),
    .o1(_01709_));
 b15nandp3ah1n02x5 _27613_ (.a(_16708_),
    .b(_16785_),
    .c(_16894_),
    .o1(_01710_));
 b15nanb02as1n08x5 _27614_ (.a(net767),
    .b(net753),
    .out0(_01711_));
 b15nanb02as1n04x5 _27615_ (.a(_17309_),
    .b(_01711_),
    .out0(_01712_));
 b15nand03ah1n06x5 _27616_ (.a(net760),
    .b(net744),
    .c(_16820_),
    .o1(_01713_));
 b15oaoi13ar1n08x5 _27617_ (.a(_16856_),
    .b(_01710_),
    .c(_01712_),
    .d(_01713_),
    .o1(_01714_));
 b15nand02al1n02x5 _27618_ (.a(net760),
    .b(_16902_),
    .o1(_01715_));
 b15oaoi13al1n04x5 _27619_ (.a(_01324_),
    .b(_01715_),
    .c(net760),
    .d(_17373_),
    .o1(_01716_));
 b15oai012as1n08x5 _27620_ (.a(_00792_),
    .b(_01288_),
    .c(_16780_),
    .o1(_01717_));
 b15and002as1n02x5 _27621_ (.a(_16872_),
    .b(_16824_),
    .o(_01718_));
 b15aoi112ar1n08x5 _27622_ (.a(_01714_),
    .b(_01716_),
    .c(_01717_),
    .d(_01718_),
    .o1(_01719_));
 b15xor002ar1n04x5 _27623_ (.a(net753),
    .b(net744),
    .out0(_01720_));
 b15nand04as1n04x5 _27624_ (.a(_16892_),
    .b(_16788_),
    .c(_16820_),
    .d(_01720_),
    .o1(_01721_));
 b15oai012al1n06x5 _27625_ (.a(_01721_),
    .b(_17371_),
    .c(_17313_),
    .o1(_01722_));
 b15nonb03as1n04x5 _27626_ (.a(net751),
    .b(net744),
    .c(net747),
    .out0(_01723_));
 b15nano22al1n03x5 _27627_ (.a(net760),
    .b(net753),
    .c(net767),
    .out0(_01724_));
 b15oai112al1n12x5 _27628_ (.a(_16798_),
    .b(_01723_),
    .c(_17309_),
    .d(_01724_),
    .o1(_01725_));
 b15aoi022ar1n02x5 _27629_ (.a(net757),
    .b(_16702_),
    .c(_16894_),
    .d(_00802_),
    .o1(_01726_));
 b15oai013an1n04x5 _27630_ (.a(_01725_),
    .b(_01726_),
    .c(_17389_),
    .d(_16741_),
    .o1(_01727_));
 b15nand03aq1n06x5 _27631_ (.a(_16710_),
    .b(_16785_),
    .c(_16836_),
    .o1(_01728_));
 b15aoi013an1n08x5 _27632_ (.a(_01308_),
    .b(_01509_),
    .c(_17380_),
    .d(_01728_),
    .o1(_01729_));
 b15nand03al1n02x5 _27633_ (.a(_16798_),
    .b(_16742_),
    .c(_16894_),
    .o1(_01730_));
 b15mdn022al1n04x5 _27634_ (.a(_16820_),
    .b(_00752_),
    .o1(_01731_),
    .sa(net757));
 b15oai013ar1n06x5 _27635_ (.a(_01730_),
    .b(_01731_),
    .c(_17297_),
    .d(_00719_),
    .o1(_01732_));
 b15nor004ah1n06x5 _27636_ (.a(_01722_),
    .b(_01727_),
    .c(_01729_),
    .d(_01732_),
    .o1(_01733_));
 b15aoai13al1n02x5 _27637_ (.a(_01540_),
    .b(_17382_),
    .c(_16810_),
    .d(_17314_),
    .o1(_01734_));
 b15nandp2as1n04x5 _27638_ (.a(_01051_),
    .b(_01734_),
    .o1(_01735_));
 b15nand04as1n16x5 _27639_ (.a(_00721_),
    .b(_01719_),
    .c(_01733_),
    .d(_01735_),
    .o1(_01736_));
 b15nonb03al1n04x5 _27640_ (.a(net745),
    .b(net746),
    .c(net765),
    .out0(_01737_));
 b15oaoi13aq1n08x5 _27641_ (.a(_16806_),
    .b(_01346_),
    .c(_01737_),
    .d(_16708_),
    .o1(_01738_));
 b15oaoi13aq1n04x5 _27642_ (.a(net758),
    .b(_17352_),
    .c(_01738_),
    .d(_16731_),
    .o1(_01739_));
 b15nand03ah1n03x5 _27643_ (.a(net766),
    .b(net758),
    .c(_16758_),
    .o1(_01740_));
 b15oai112al1n12x5 _27644_ (.a(_16770_),
    .b(_01740_),
    .c(_16810_),
    .d(net766),
    .o1(_01741_));
 b15oai012al1n06x5 _27645_ (.a(net762),
    .b(_16774_),
    .c(_00708_),
    .o1(_01742_));
 b15aoi112as1n08x5 _27646_ (.a(_16741_),
    .b(_01739_),
    .c(_01741_),
    .d(_01742_),
    .o1(_01743_));
 b15oai112aq1n02x5 _27647_ (.a(net759),
    .b(net748),
    .c(_17294_),
    .d(_17292_),
    .o1(_01744_));
 b15aoi012ar1n04x5 _27648_ (.a(_16693_),
    .b(_16786_),
    .c(_01744_),
    .o1(_01745_));
 b15aoai13as1n08x5 _27649_ (.a(net763),
    .b(_01745_),
    .c(_17359_),
    .d(_16896_),
    .o1(_01746_));
 b15oaoi13an1n04x5 _27650_ (.a(net760),
    .b(_16849_),
    .c(_17285_),
    .d(net767),
    .o1(_01747_));
 b15oai112al1n16x5 _27651_ (.a(net757),
    .b(_16710_),
    .c(_00745_),
    .d(_01747_),
    .o1(_01748_));
 b15oab012al1n03x5 _27652_ (.a(_00752_),
    .b(_01711_),
    .c(_00811_),
    .out0(_01749_));
 b15oai013ah1n08x5 _27653_ (.a(_16741_),
    .b(net757),
    .c(_00800_),
    .d(_01749_),
    .o1(_01750_));
 b15oai022aq1n06x5 _27654_ (.a(_17314_),
    .b(_16760_),
    .c(_16775_),
    .d(_16764_),
    .o1(_01751_));
 b15aoi012ar1n06x5 _27655_ (.a(_01750_),
    .b(_01751_),
    .c(_16770_),
    .o1(_01752_));
 b15aoi013aq1n08x5 _27656_ (.a(_01743_),
    .b(_01746_),
    .c(_01748_),
    .d(_01752_),
    .o1(_01753_));
 b15nano23as1n24x5 _27657_ (.a(_01699_),
    .b(_01709_),
    .c(_01736_),
    .d(_01753_),
    .out0(_01754_));
 b15nandp3aq1n02x5 _27658_ (.a(_16018_),
    .b(_01002_),
    .c(_16047_),
    .o1(_01755_));
 b15nor003aq1n06x5 _27659_ (.a(net879),
    .b(_15987_),
    .c(_16021_),
    .o1(_01756_));
 b15oaoi13ar1n04x5 _27660_ (.a(_17424_),
    .b(net882),
    .c(_01756_),
    .d(_01496_),
    .o1(_01757_));
 b15oai112aq1n08x5 _27661_ (.a(_16028_),
    .b(_01755_),
    .c(_01757_),
    .d(_16018_),
    .o1(_01758_));
 b15aoai13aq1n03x5 _27662_ (.a(\us20.a[2] ),
    .b(_16084_),
    .c(_16086_),
    .d(net883),
    .o1(_01759_));
 b15oai012an1n03x5 _27663_ (.a(_17518_),
    .b(_16110_),
    .c(net882),
    .o1(_01760_));
 b15aoi022ar1n08x5 _27664_ (.a(_16066_),
    .b(_17437_),
    .c(_01760_),
    .d(_16047_),
    .o1(_01761_));
 b15nanb02as1n06x5 _27665_ (.a(net865),
    .b(\us20.a[4] ),
    .out0(_01762_));
 b15nand02ar1n04x5 _27666_ (.a(net865),
    .b(\us20.a[2] ),
    .o1(_01763_));
 b15oaoi13al1n04x5 _27667_ (.a(_17479_),
    .b(_01762_),
    .c(_01763_),
    .d(\us20.a[4] ),
    .o1(_01764_));
 b15aoi112al1n04x5 _27668_ (.a(net880),
    .b(_01764_),
    .c(_16058_),
    .d(_16010_),
    .o1(_01765_));
 b15aoi112as1n02x5 _27669_ (.a(_16078_),
    .b(_01454_),
    .c(_00550_),
    .d(net883),
    .o1(_01766_));
 b15oai112ah1n08x5 _27670_ (.a(_01759_),
    .b(_01761_),
    .c(_01765_),
    .d(_01766_),
    .o1(_01767_));
 b15oai012al1n16x5 _27671_ (.a(_01758_),
    .b(_01767_),
    .c(_16028_),
    .o1(_01768_));
 b15aoi012ah1n02x5 _27672_ (.a(_00605_),
    .b(_17487_),
    .c(_16028_),
    .o1(_01769_));
 b15oai122an1n12x5 _27673_ (.a(net876),
    .b(_16031_),
    .c(_16104_),
    .d(_01769_),
    .e(_15959_),
    .o1(_01770_));
 b15nor003an1n04x5 _27674_ (.a(_16092_),
    .b(_01396_),
    .c(_01038_),
    .o1(_01771_));
 b15aoi012ar1n02x5 _27675_ (.a(_01762_),
    .b(_16116_),
    .c(_01038_),
    .o1(_01772_));
 b15oai012aq1n03x5 _27676_ (.a(net869),
    .b(_01771_),
    .c(_01772_),
    .o1(_01773_));
 b15oai022ar1n02x5 _27677_ (.a(_16088_),
    .b(_16021_),
    .c(_00598_),
    .d(_01396_),
    .o1(_01774_));
 b15oai012ar1n02x5 _27678_ (.a(_01385_),
    .b(_15959_),
    .c(net869),
    .o1(_01775_));
 b15aoi022aq1n02x5 _27679_ (.a(net869),
    .b(_01774_),
    .c(_01775_),
    .d(_00545_),
    .o1(_01776_));
 b15oai122ah1n08x5 _27680_ (.a(_01773_),
    .b(_16112_),
    .c(_16135_),
    .d(net880),
    .e(_01776_),
    .o1(_01777_));
 b15oai012ah1n06x5 _27681_ (.a(_01770_),
    .b(_01777_),
    .c(net876),
    .o1(_01778_));
 b15oai022aq1n02x5 _27682_ (.a(_17497_),
    .b(_17455_),
    .c(_00600_),
    .d(net884),
    .o1(_01779_));
 b15aoi122ah1n04x5 _27683_ (.a(net873),
    .b(_17469_),
    .c(_15989_),
    .d(_01779_),
    .e(_17463_),
    .o1(_01780_));
 b15norp02ar1n03x5 _27684_ (.a(_16028_),
    .b(_16034_),
    .o1(_01781_));
 b15aoi112as1n04x5 _27685_ (.a(_16018_),
    .b(_01780_),
    .c(_01781_),
    .d(_00612_),
    .o1(_01782_));
 b15norp02ar1n02x5 _27686_ (.a(net863),
    .b(net877),
    .o1(_01783_));
 b15oai022al1n02x5 _27687_ (.a(_16080_),
    .b(_15995_),
    .c(_00598_),
    .d(_01783_),
    .o1(_01784_));
 b15nandp3ar1n03x5 _27688_ (.a(_16078_),
    .b(_15943_),
    .c(_01784_),
    .o1(_01785_));
 b15nanb03ar1n02x5 _27689_ (.a(net866),
    .b(net881),
    .c(net867),
    .out0(_01786_));
 b15nanb03ar1n02x5 _27690_ (.a(net863),
    .b(net873),
    .c(net871),
    .out0(_01787_));
 b15oaoi13aq1n03x5 _27691_ (.a(_01786_),
    .b(_01787_),
    .c(_17462_),
    .d(_15970_),
    .o1(_01788_));
 b15nor004ar1n04x5 _27692_ (.a(net881),
    .b(_16080_),
    .c(_16113_),
    .d(_15993_),
    .o1(_01789_));
 b15oai012al1n06x5 _27693_ (.a(net884),
    .b(_01788_),
    .c(_01789_),
    .o1(_01790_));
 b15oai013aq1n03x5 _27694_ (.a(_16004_),
    .b(_16021_),
    .c(_00599_),
    .d(_16085_),
    .o1(_01791_));
 b15aoi012al1n02x5 _27695_ (.a(_17420_),
    .b(_16160_),
    .c(net881),
    .o1(_01792_));
 b15oai112al1n08x5 _27696_ (.a(_01025_),
    .b(_01791_),
    .c(_01792_),
    .d(net884),
    .o1(_01793_));
 b15nand04ah1n08x5 _27697_ (.a(_17523_),
    .b(_01785_),
    .c(_01790_),
    .d(_01793_),
    .o1(_01794_));
 b15norp02ar1n03x5 _27698_ (.a(net880),
    .b(_00589_),
    .o1(_01795_));
 b15aoai13ar1n08x5 _27699_ (.a(_00999_),
    .b(_01795_),
    .c(net877),
    .d(_00614_),
    .o1(_01796_));
 b15aoi013al1n06x5 _27700_ (.a(_00540_),
    .b(_00543_),
    .c(_15969_),
    .d(_16025_),
    .o1(_01797_));
 b15orn003ar1n03x5 _27701_ (.a(_16162_),
    .b(_00599_),
    .c(_01797_),
    .o(_01798_));
 b15aoai13ah1n04x5 _27702_ (.a(net883),
    .b(_16042_),
    .c(_00614_),
    .d(_01014_),
    .o1(_01799_));
 b15oai012ah1n02x5 _27703_ (.a(net883),
    .b(_17420_),
    .c(_17447_),
    .o1(_01800_));
 b15nor004ah1n03x5 _27704_ (.a(_16028_),
    .b(_16126_),
    .c(_16082_),
    .d(_16010_),
    .o1(_01801_));
 b15oai012al1n08x5 _27705_ (.a(_01800_),
    .b(_01801_),
    .c(_17490_),
    .o1(_01802_));
 b15nand04ah1n12x5 _27706_ (.a(_01796_),
    .b(_01798_),
    .c(_01799_),
    .d(_01802_),
    .o1(_01803_));
 b15aoai13an1n04x5 _27707_ (.a(_16078_),
    .b(_16042_),
    .c(_00614_),
    .d(_16044_),
    .o1(_01804_));
 b15orn002ar1n02x5 _27708_ (.a(net863),
    .b(net873),
    .o(_01805_));
 b15oai022ar1n02x5 _27709_ (.a(_16011_),
    .b(_01805_),
    .c(_00535_),
    .d(_16116_),
    .o1(_01806_));
 b15nand03aq1n02x5 _27710_ (.a(_16092_),
    .b(_15943_),
    .c(_01806_),
    .o1(_01807_));
 b15nonb03aq1n04x5 _27711_ (.a(net880),
    .b(net884),
    .c(net871),
    .out0(_01808_));
 b15nor004al1n12x5 _27712_ (.a(_01002_),
    .b(_15993_),
    .c(_01416_),
    .d(_01808_),
    .o1(_01809_));
 b15aoi013ah1n02x5 _27713_ (.a(_01809_),
    .b(_00599_),
    .c(_16158_),
    .d(_15989_),
    .o1(_01810_));
 b15nand04ah1n06x5 _27714_ (.a(_16076_),
    .b(_01804_),
    .c(_01807_),
    .d(_01810_),
    .o1(_01811_));
 b15nor004an1n12x5 _27715_ (.a(_01782_),
    .b(_01794_),
    .c(_01803_),
    .d(_01811_),
    .o1(_01812_));
 b15nandp3an1n24x5 _27716_ (.a(_01768_),
    .b(_01778_),
    .c(_01812_),
    .o1(_01813_));
 b15xor002ar1n02x5 _27717_ (.a(_01689_),
    .b(_01813_),
    .out0(_01814_));
 b15xor002aq1n02x5 _27718_ (.a(_01754_),
    .b(_01814_),
    .out0(_01815_));
 b15oai012ar1n02x5 _27719_ (.a(_00650_),
    .b(_16260_),
    .c(_16248_),
    .o1(_01816_));
 b15nand02an1n03x5 _27720_ (.a(_16997_),
    .b(_01816_),
    .o1(_01817_));
 b15aoai13ar1n03x5 _27721_ (.a(_16336_),
    .b(_16282_),
    .c(_16342_),
    .d(_16367_),
    .o1(_01818_));
 b15nandp2al1n04x5 _27722_ (.a(net732),
    .b(_01818_),
    .o1(_01819_));
 b15oai112al1n06x5 _27723_ (.a(_01817_),
    .b(_01819_),
    .c(_16318_),
    .d(_16402_),
    .o1(_01820_));
 b15aoi012ar1n02x5 _27724_ (.a(_16342_),
    .b(_16225_),
    .c(_17005_),
    .o1(_01821_));
 b15aoai13ah1n03x5 _27725_ (.a(net736),
    .b(_01821_),
    .c(_16340_),
    .d(net743),
    .o1(_01822_));
 b15oaoi13aq1n08x5 _27726_ (.a(_16999_),
    .b(_16350_),
    .c(_16416_),
    .d(net741),
    .o1(_01823_));
 b15norp03ah1n04x5 _27727_ (.a(net739),
    .b(_16239_),
    .c(_16367_),
    .o1(_01824_));
 b15oai112an1n16x5 _27728_ (.a(_16226_),
    .b(_01822_),
    .c(_01823_),
    .d(_01824_),
    .o1(_01825_));
 b15nand02ar1n02x5 _27729_ (.a(_16340_),
    .b(_17009_),
    .o1(_01826_));
 b15oai112aq1n04x5 _27730_ (.a(_16414_),
    .b(_01826_),
    .c(_16231_),
    .d(_16311_),
    .o1(_01827_));
 b15aoai13ah1n04x5 _27731_ (.a(_16342_),
    .b(_01820_),
    .c(_01825_),
    .d(_01827_),
    .o1(_01828_));
 b15norp02ar1n02x5 _27732_ (.a(net732),
    .b(_16402_),
    .o1(_01829_));
 b15aoai13as1n02x5 _27733_ (.a(net743),
    .b(_01829_),
    .c(_17062_),
    .d(_16980_),
    .o1(_01830_));
 b15oai112an1n06x5 _27734_ (.a(net732),
    .b(_16379_),
    .c(_16977_),
    .d(_16213_),
    .o1(_01831_));
 b15oai012ar1n06x5 _27735_ (.a(net736),
    .b(_16977_),
    .c(_16283_),
    .o1(_01832_));
 b15aoai13as1n06x5 _27736_ (.a(_01830_),
    .b(_01831_),
    .c(_01832_),
    .d(_16342_),
    .o1(_01833_));
 b15aoi112ar1n04x5 _27737_ (.a(_16226_),
    .b(_16958_),
    .c(_16379_),
    .d(_16311_),
    .o1(_01834_));
 b15oaoi13as1n04x5 _27738_ (.a(_01834_),
    .b(_16320_),
    .c(_17046_),
    .d(_00622_),
    .o1(_01835_));
 b15nor002al1n02x5 _27739_ (.a(net736),
    .b(_17225_),
    .o1(_01836_));
 b15nandp3ar1n02x5 _27740_ (.a(\us02.a[1] ),
    .b(_16995_),
    .c(_16993_),
    .o1(_01837_));
 b15oaoi13as1n02x5 _27741_ (.a(net743),
    .b(_01837_),
    .c(_16993_),
    .d(\us02.a[1] ),
    .o1(_01838_));
 b15nand02ar1n02x5 _27742_ (.a(\us02.a[1] ),
    .b(_16333_),
    .o1(_01839_));
 b15aoi022ar1n02x5 _27743_ (.a(net732),
    .b(_16315_),
    .c(_17225_),
    .d(_01839_),
    .o1(_01840_));
 b15oai013ah1n04x5 _27744_ (.a(_01835_),
    .b(_01836_),
    .c(_01838_),
    .d(_01840_),
    .o1(_01841_));
 b15nand03al1n03x5 _27745_ (.a(net738),
    .b(_16328_),
    .c(_17041_),
    .o1(_01842_));
 b15oaoi13ar1n04x5 _27746_ (.a(_16237_),
    .b(_01842_),
    .c(_00653_),
    .d(net738),
    .o1(_01843_));
 b15oai022an1n04x5 _27747_ (.a(net730),
    .b(_16231_),
    .c(_16396_),
    .d(_16972_),
    .o1(_01844_));
 b15aoi112aq1n06x5 _27748_ (.a(_00969_),
    .b(_01843_),
    .c(_01844_),
    .d(_16214_),
    .o1(_01845_));
 b15aoi022ar1n02x5 _27749_ (.a(net736),
    .b(_16239_),
    .c(_17008_),
    .d(_16283_),
    .o1(_01846_));
 b15oai022al1n02x5 _27750_ (.a(_16225_),
    .b(_01675_),
    .c(_01846_),
    .d(net739),
    .o1(_01847_));
 b15aob012ah1n04x5 _27751_ (.a(_01845_),
    .b(_01847_),
    .c(net732),
    .out0(_01848_));
 b15nor003al1n06x5 _27752_ (.a(_01833_),
    .b(_01841_),
    .c(_01848_),
    .o1(_01849_));
 b15norp03ar1n02x5 _27753_ (.a(net743),
    .b(net736),
    .c(_16260_),
    .o1(_01850_));
 b15aoi112al1n02x5 _27754_ (.a(_16226_),
    .b(_01850_),
    .c(_16403_),
    .d(net743),
    .o1(_01851_));
 b15oai012aq1n04x5 _27755_ (.a(_16402_),
    .b(_16329_),
    .c(net741),
    .o1(_01852_));
 b15aoi222ah1n06x5 _27756_ (.a(net739),
    .b(_16343_),
    .c(_00954_),
    .d(_17223_),
    .e(_01852_),
    .f(net735),
    .o1(_01853_));
 b15aoi012ar1n04x5 _27757_ (.a(_01851_),
    .b(_01853_),
    .c(_16226_),
    .o1(_01854_));
 b15oaoi13an1n08x5 _27758_ (.a(_16325_),
    .b(_16191_),
    .c(_17270_),
    .d(_17271_),
    .o1(_01855_));
 b15nanb02aq1n03x5 _27759_ (.a(_01855_),
    .b(_00954_),
    .out0(_01856_));
 b15norp03an1n02x5 _27760_ (.a(_16283_),
    .b(_16993_),
    .c(_17258_),
    .o1(_01857_));
 b15aoi012ar1n04x5 _27761_ (.a(_01857_),
    .b(_17221_),
    .c(_16365_),
    .o1(_01858_));
 b15oai112al1n12x5 _27762_ (.a(_17050_),
    .b(_01856_),
    .c(_01858_),
    .d(_16342_),
    .o1(_01859_));
 b15oai012ah1n02x5 _27763_ (.a(_16316_),
    .b(_16315_),
    .c(_16321_),
    .o1(_01860_));
 b15oai112as1n06x5 _27764_ (.a(net732),
    .b(_01860_),
    .c(_16414_),
    .d(_16311_),
    .o1(_01861_));
 b15aoi112ah1n06x5 _27765_ (.a(_01854_),
    .b(_01859_),
    .c(_01825_),
    .d(_01861_),
    .o1(_01862_));
 b15oai112ah1n16x5 _27766_ (.a(net740),
    .b(net723),
    .c(_17251_),
    .d(_16419_),
    .o1(_01863_));
 b15oai012ar1n02x5 _27767_ (.a(_01863_),
    .b(_16260_),
    .c(net743),
    .o1(_01864_));
 b15aoi022ar1n02x5 _27768_ (.a(_16390_),
    .b(_16332_),
    .c(_01864_),
    .d(net739),
    .o1(_01865_));
 b15oai112al1n06x5 _27769_ (.a(net736),
    .b(_01819_),
    .c(_01865_),
    .d(net732),
    .o1(_01866_));
 b15nand03as1n12x5 _27770_ (.a(_16181_),
    .b(_16292_),
    .c(_16960_),
    .o1(_01867_));
 b15aoi022aq1n02x5 _27771_ (.a(_16321_),
    .b(_16345_),
    .c(_17008_),
    .d(net732),
    .o1(_01868_));
 b15oai122ah1n08x5 _27772_ (.a(_01867_),
    .b(_01868_),
    .c(net739),
    .d(_16357_),
    .e(_17258_),
    .o1(_01869_));
 b15oai012aq1n08x5 _27773_ (.a(_01866_),
    .b(_01869_),
    .c(\us02.a[2] ),
    .o1(_01870_));
 b15nand04as1n16x5 _27774_ (.a(_01828_),
    .b(_01849_),
    .c(_01862_),
    .d(_01870_),
    .o1(_01871_));
 b15oai112ar1n02x5 _27775_ (.a(_16466_),
    .b(_16482_),
    .c(_00900_),
    .d(net611),
    .o1(_01872_));
 b15oaoi13ar1n02x5 _27776_ (.a(net615),
    .b(_01872_),
    .c(_16629_),
    .d(_16466_),
    .o1(_01873_));
 b15oai012al1n03x5 _27777_ (.a(_16651_),
    .b(_16680_),
    .c(_16524_),
    .o1(_01874_));
 b15aoi022ar1n02x5 _27778_ (.a(_16591_),
    .b(_16650_),
    .c(_01874_),
    .d(net619),
    .o1(_01875_));
 b15aoi012aq1n02x5 _27779_ (.a(_01873_),
    .b(_01875_),
    .c(net615),
    .o1(_01876_));
 b15nandp2ah1n08x5 _27780_ (.a(net603),
    .b(net599),
    .o1(_01877_));
 b15aob012al1n02x5 _27781_ (.a(_16592_),
    .b(_17181_),
    .c(_01877_),
    .out0(_01878_));
 b15oai112al1n06x5 _27782_ (.a(_16604_),
    .b(_01878_),
    .c(_17112_),
    .d(_16453_),
    .o1(_01879_));
 b15aoi012ar1n02x5 _27783_ (.a(_16592_),
    .b(_16577_),
    .c(_16481_),
    .o1(_01880_));
 b15aoi012aq1n02x5 _27784_ (.a(_01879_),
    .b(_01880_),
    .c(_17183_),
    .o1(_01881_));
 b15oai013ar1n02x5 _27785_ (.a(_16519_),
    .b(_17183_),
    .c(net619),
    .d(net608),
    .o1(_01882_));
 b15aoi022ar1n02x5 _27786_ (.a(_16435_),
    .b(_01224_),
    .c(_01882_),
    .d(net615),
    .o1(_01883_));
 b15nor002aq1n02x5 _27787_ (.a(_16460_),
    .b(_01883_),
    .o1(_01884_));
 b15norp03an1n08x5 _27788_ (.a(_01876_),
    .b(_01881_),
    .c(_01884_),
    .o1(_01885_));
 b15nandp2ar1n02x5 _27789_ (.a(_16656_),
    .b(_00823_),
    .o1(_01886_));
 b15oaoi13an1n04x5 _27790_ (.a(net602),
    .b(_01886_),
    .c(_17113_),
    .d(_00823_),
    .o1(_01887_));
 b15nor002ar1n08x5 _27791_ (.a(net596),
    .b(net613),
    .o1(_01888_));
 b15aoai13as1n08x5 _27792_ (.a(_01259_),
    .b(_01887_),
    .c(_16481_),
    .d(_01888_),
    .o1(_01889_));
 b15oaoi13an1n03x5 _27793_ (.a(net608),
    .b(_01889_),
    .c(_01239_),
    .d(_16575_),
    .o1(_01890_));
 b15nand02ar1n02x5 _27794_ (.a(_00902_),
    .b(_17562_),
    .o1(_01891_));
 b15oaoi13ah1n03x5 _27795_ (.a(net612),
    .b(_01891_),
    .c(_17131_),
    .d(_16453_),
    .o1(_01892_));
 b15nor003an1n06x5 _27796_ (.a(_16435_),
    .b(_16490_),
    .c(_16479_),
    .o1(_01893_));
 b15norp02as1n03x5 _27797_ (.a(_16497_),
    .b(_17602_),
    .o1(_01894_));
 b15aoi222as1n12x5 _27798_ (.a(_16670_),
    .b(_16674_),
    .c(_01893_),
    .d(_16672_),
    .e(_01894_),
    .f(_16601_),
    .o1(_01895_));
 b15aoi022aq1n02x5 _27799_ (.a(_16526_),
    .b(_16582_),
    .c(_16650_),
    .d(_16439_),
    .o1(_01896_));
 b15oai012al1n02x5 _27800_ (.a(_01895_),
    .b(_01896_),
    .c(net610),
    .o1(_01897_));
 b15norp02al1n12x5 _27801_ (.a(_16538_),
    .b(_01580_),
    .o1(_01898_));
 b15oai012al1n06x5 _27802_ (.a(_16558_),
    .b(_16614_),
    .c(_01898_),
    .o1(_01899_));
 b15norp02ar1n02x5 _27803_ (.a(_16536_),
    .b(_16581_),
    .o1(_01900_));
 b15oai012as1n03x5 _27804_ (.a(net616),
    .b(_01898_),
    .c(_01900_),
    .o1(_01901_));
 b15nona23an1n12x5 _27805_ (.a(_01892_),
    .b(_01897_),
    .c(_01899_),
    .d(_01901_),
    .out0(_01902_));
 b15norp03an1n02x5 _27806_ (.a(_16522_),
    .b(_16592_),
    .c(_17578_),
    .o1(_01903_));
 b15nor003ar1n02x5 _27807_ (.a(_16643_),
    .b(_17088_),
    .c(_00851_),
    .o1(_01904_));
 b15norp03ar1n02x5 _27808_ (.a(net608),
    .b(_17085_),
    .c(_16582_),
    .o1(_01905_));
 b15norp02ar1n02x5 _27809_ (.a(_16478_),
    .b(_16608_),
    .o1(_01906_));
 b15nor004al1n03x5 _27810_ (.a(_01903_),
    .b(_01904_),
    .c(_01905_),
    .d(_01906_),
    .o1(_01907_));
 b15nand03ar1n02x5 _27811_ (.a(net616),
    .b(_16466_),
    .c(_16650_),
    .o1(_01908_));
 b15aoi112ar1n02x5 _27812_ (.a(_16460_),
    .b(_16490_),
    .c(_17173_),
    .d(_01908_),
    .o1(_01909_));
 b15orn002aq1n03x5 _27813_ (.a(net606),
    .b(net619),
    .o(_01910_));
 b15oai022al1n02x5 _27814_ (.a(_16659_),
    .b(_17088_),
    .c(_01910_),
    .d(net611),
    .o1(_01911_));
 b15oai012ar1n02x5 _27815_ (.a(_00823_),
    .b(_16478_),
    .c(net619),
    .o1(_01912_));
 b15aoi022an1n02x5 _27816_ (.a(_16550_),
    .b(_01911_),
    .c(_01912_),
    .d(_17146_),
    .o1(_01913_));
 b15oab012ar1n02x5 _27817_ (.a(_01909_),
    .b(_01913_),
    .c(_16466_),
    .out0(_01914_));
 b15norp03ar1n02x5 _27818_ (.a(net620),
    .b(net608),
    .c(_16680_),
    .o1(_01915_));
 b15aoi012aq1n02x5 _27819_ (.a(_01915_),
    .b(_17190_),
    .c(_16650_),
    .o1(_01916_));
 b15oai112as1n04x5 _27820_ (.a(_01907_),
    .b(_01914_),
    .c(net612),
    .d(_01916_),
    .o1(_01917_));
 b15nor003ah1n04x5 _27821_ (.a(_01890_),
    .b(_01902_),
    .c(_01917_),
    .o1(_01918_));
 b15nand04al1n06x5 _27822_ (.a(_16458_),
    .b(_16597_),
    .c(\us13.a[2] ),
    .d(_16475_),
    .o1(_01919_));
 b15nanb02al1n06x5 _27823_ (.a(net607),
    .b(net612),
    .out0(_01920_));
 b15oaoi13aq1n03x5 _27824_ (.a(_16458_),
    .b(_01920_),
    .c(_16516_),
    .d(_16659_),
    .o1(_01921_));
 b15aoi012ah1n04x5 _27825_ (.a(_16539_),
    .b(_01921_),
    .c(net604),
    .o1(_01922_));
 b15oaoi13as1n08x5 _27826_ (.a(net617),
    .b(_01919_),
    .c(_01922_),
    .d(_16597_),
    .o1(_01923_));
 b15aoai13ar1n02x5 _27827_ (.a(_16481_),
    .b(_01888_),
    .c(net596),
    .d(net614),
    .o1(_01924_));
 b15oaoi13ar1n02x5 _27828_ (.a(_16616_),
    .b(_01924_),
    .c(_17175_),
    .d(_16665_),
    .o1(_01925_));
 b15oai022ar1n02x5 _27829_ (.a(net614),
    .b(_16482_),
    .c(_16521_),
    .d(net613),
    .o1(_01926_));
 b15and002ar1n02x5 _27830_ (.a(_16558_),
    .b(_01926_),
    .o(_01927_));
 b15orn003as1n02x5 _27831_ (.a(_01923_),
    .b(_01925_),
    .c(_01927_),
    .o(_01928_));
 b15nand04ar1n03x5 _27832_ (.a(_16620_),
    .b(_01877_),
    .c(_16564_),
    .d(_01216_),
    .o1(_01929_));
 b15nandp3ah1n02x5 _27833_ (.a(_16460_),
    .b(\us13.a[3] ),
    .c(_01929_),
    .o1(_01930_));
 b15nandp2ar1n08x5 _27834_ (.a(net599),
    .b(net614),
    .o1(_01931_));
 b15aboi22an1n06x5 _27835_ (.a(_01216_),
    .b(_01931_),
    .c(net603),
    .d(_16561_),
    .out0(_01932_));
 b15oaoi13an1n04x5 _27836_ (.a(net598),
    .b(_17551_),
    .c(_01932_),
    .d(net605),
    .o1(_01933_));
 b15oaoi13as1n08x5 _27837_ (.a(_01928_),
    .b(_01930_),
    .c(_16632_),
    .d(_01933_),
    .o1(_01934_));
 b15oai012ar1n02x5 _27838_ (.a(_16521_),
    .b(_16576_),
    .c(_16508_),
    .o1(_01935_));
 b15nand02al1n02x5 _27839_ (.a(_16619_),
    .b(_01935_),
    .o1(_01936_));
 b15oai112al1n08x5 _27840_ (.a(_16466_),
    .b(_01936_),
    .c(_17125_),
    .d(net616),
    .o1(_01937_));
 b15oaoi13an1n04x5 _27841_ (.a(_16439_),
    .b(_16528_),
    .c(_16576_),
    .d(net616),
    .o1(_01938_));
 b15oaoi13ah1n08x5 _27842_ (.a(_01937_),
    .b(net612),
    .c(_17077_),
    .d(_01938_),
    .o1(_01939_));
 b15oai112as1n16x5 _27843_ (.a(_01885_),
    .b(_01918_),
    .c(_01934_),
    .d(_01939_),
    .o1(_01940_));
 b15xnr002ah1n08x5 _27844_ (.a(_01871_),
    .b(_01940_),
    .out0(_01941_));
 b15xor002ar1n03x5 _27845_ (.a(_01815_),
    .b(_01941_),
    .out0(_01942_));
 b15mdn022ah1n03x5 _27846_ (.a(_01693_),
    .b(_01942_),
    .o1(_01943_),
    .sa(net540));
 b15xor002aq1n06x5 _27847_ (.a(\u0.w[2][6] ),
    .b(_01943_),
    .out0(_00119_));
 b15oai012an1n06x5 _27848_ (.a(net869),
    .b(_00585_),
    .c(_00586_),
    .o1(_01944_));
 b15aoi012al1n02x5 _27849_ (.a(net873),
    .b(_01486_),
    .c(_01944_),
    .o1(_01945_));
 b15aoai13ar1n02x5 _27850_ (.a(_16066_),
    .b(_01945_),
    .c(net873),
    .d(_00550_),
    .o1(_01946_));
 b15nand02aq1n02x5 _27851_ (.a(_16129_),
    .b(_16000_),
    .o1(_01947_));
 b15aoi122al1n04x5 _27852_ (.a(_16028_),
    .b(_16164_),
    .c(_01947_),
    .d(_16033_),
    .e(net875),
    .o1(_01948_));
 b15norp02ar1n02x5 _27853_ (.a(net875),
    .b(_16040_),
    .o1(_01949_));
 b15aoai13as1n03x5 _27854_ (.a(net885),
    .b(_01949_),
    .c(_17427_),
    .d(net875),
    .o1(_01950_));
 b15aoi122al1n04x5 _27855_ (.a(_01756_),
    .b(_16110_),
    .c(_16045_),
    .d(_16145_),
    .e(_00614_),
    .o1(_01951_));
 b15aoi013al1n04x5 _27856_ (.a(net872),
    .b(_01002_),
    .c(_17437_),
    .d(_16018_),
    .o1(_01952_));
 b15aoi013aq1n06x5 _27857_ (.a(_01948_),
    .b(_01950_),
    .c(_01951_),
    .d(_01952_),
    .o1(_01953_));
 b15nand03an1n03x5 _27858_ (.a(net873),
    .b(_16147_),
    .c(_16010_),
    .o1(_01954_));
 b15oai012ar1n08x5 _27859_ (.a(_01954_),
    .b(_01486_),
    .c(_16134_),
    .o1(_01955_));
 b15oai012ar1n02x5 _27860_ (.a(_15959_),
    .b(net873),
    .c(_17420_),
    .o1(_01956_));
 b15aoi012ar1n02x5 _27861_ (.a(_00589_),
    .b(_00599_),
    .c(_01956_),
    .o1(_01957_));
 b15nandp2al1n02x5 _27862_ (.a(net883),
    .b(_00535_),
    .o1(_01958_));
 b15nand03aq1n03x5 _27863_ (.a(_15959_),
    .b(_16000_),
    .c(_17520_),
    .o1(_01959_));
 b15oai112as1n06x5 _27864_ (.a(_01958_),
    .b(_01959_),
    .c(_17490_),
    .d(_17444_),
    .o1(_01960_));
 b15xor002ar1n02x5 _27865_ (.a(_16088_),
    .b(_17469_),
    .out0(_01961_));
 b15nor004al1n02x5 _27866_ (.a(net869),
    .b(net863),
    .c(_16028_),
    .d(_01392_),
    .o1(_01962_));
 b15oai022ar1n02x5 _27867_ (.a(_15959_),
    .b(_16137_),
    .c(_16089_),
    .d(_16028_),
    .o1(_01963_));
 b15aoi022aq1n04x5 _27868_ (.a(_01961_),
    .b(_01962_),
    .c(_01963_),
    .d(_00550_),
    .o1(_01964_));
 b15nona23ar1n12x5 _27869_ (.a(_01955_),
    .b(_01957_),
    .c(_01960_),
    .d(_01964_),
    .out0(_01965_));
 b15nano23aq1n06x5 _27870_ (.a(_17436_),
    .b(_01946_),
    .c(_01953_),
    .d(_01965_),
    .out0(_01966_));
 b15nor004ar1n02x5 _27871_ (.a(_16113_),
    .b(_15955_),
    .c(_16008_),
    .d(_16011_),
    .o1(_01967_));
 b15aoai13an1n02x5 _27872_ (.a(_16028_),
    .b(_01967_),
    .c(_16147_),
    .d(net883),
    .o1(_01968_));
 b15aoi022an1n02x5 _27873_ (.a(_00550_),
    .b(_17469_),
    .c(_17410_),
    .d(_17437_),
    .o1(_01969_));
 b15oai012al1n06x5 _27874_ (.a(_01968_),
    .b(_01969_),
    .c(_16028_),
    .o1(_01970_));
 b15oai012ar1n03x5 _27875_ (.a(_16129_),
    .b(_15997_),
    .c(net869),
    .o1(_01971_));
 b15aoai13as1n04x5 _27876_ (.a(_17480_),
    .b(_01971_),
    .c(net869),
    .d(_15997_),
    .o1(_01972_));
 b15nanb02ar1n06x5 _27877_ (.a(_16122_),
    .b(_17513_),
    .out0(_01973_));
 b15aoi112as1n08x5 _27878_ (.a(\us20.a[7] ),
    .b(_16137_),
    .c(_01972_),
    .d(_01973_),
    .o1(_01974_));
 b15aoi112ar1n02x5 _27879_ (.a(net873),
    .b(_17459_),
    .c(_01486_),
    .d(_16132_),
    .o1(_01975_));
 b15norp03ar1n02x5 _27880_ (.a(net880),
    .b(_15993_),
    .c(_01944_),
    .o1(_01976_));
 b15nor002ar1n02x5 _27881_ (.a(_16028_),
    .b(_16110_),
    .o1(_01977_));
 b15aoi022ar1n06x5 _27882_ (.a(_00550_),
    .b(_16044_),
    .c(_01977_),
    .d(_17446_),
    .o1(_01978_));
 b15norp03aq1n02x5 _27883_ (.a(_16088_),
    .b(_16021_),
    .c(_16112_),
    .o1(_01979_));
 b15oai112ah1n06x5 _27884_ (.a(net869),
    .b(net880),
    .c(_01771_),
    .d(_01979_),
    .o1(_01980_));
 b15nona23ar1n08x5 _27885_ (.a(_01975_),
    .b(_01976_),
    .c(_01978_),
    .d(_01980_),
    .out0(_01981_));
 b15norp03al1n12x5 _27886_ (.a(_01970_),
    .b(_01974_),
    .c(_01981_),
    .o1(_01982_));
 b15oab012ar1n02x5 _27887_ (.a(_00543_),
    .b(_00599_),
    .c(_16040_),
    .out0(_01983_));
 b15aoai13al1n02x5 _27888_ (.a(net879),
    .b(_17437_),
    .c(_16045_),
    .d(net872),
    .o1(_01984_));
 b15aoi013ah1n02x5 _27889_ (.a(_01983_),
    .b(_01984_),
    .c(_17522_),
    .d(_16009_),
    .o1(_01985_));
 b15nor002aq1n02x5 _27890_ (.a(net871),
    .b(_16153_),
    .o1(_01986_));
 b15and003al1n02x5 _27891_ (.a(net871),
    .b(\us20.a[3] ),
    .c(_17415_),
    .o(_01987_));
 b15oai112ah1n08x5 _27892_ (.a(net869),
    .b(_01377_),
    .c(_01986_),
    .d(_01987_),
    .o1(_01988_));
 b15norp02aq1n02x5 _27893_ (.a(_17463_),
    .b(_16100_),
    .o1(_01989_));
 b15norp02ar1n02x5 _27894_ (.a(_16085_),
    .b(_16153_),
    .o1(_01990_));
 b15aoi012aq1n04x5 _27895_ (.a(_01989_),
    .b(_01990_),
    .c(net884),
    .o1(_01991_));
 b15aoi012ar1n06x5 _27896_ (.a(_15943_),
    .b(_17457_),
    .c(\us20.a[0] ),
    .o1(_01992_));
 b15oai122as1n16x5 _27897_ (.a(_01988_),
    .b(_01991_),
    .c(_17503_),
    .d(_17442_),
    .e(_01992_),
    .o1(_01993_));
 b15oai012an1n06x5 _27898_ (.a(_01985_),
    .b(_01993_),
    .c(net876),
    .o1(_01994_));
 b15oaoi13ar1n02x5 _27899_ (.a(_15959_),
    .b(_01494_),
    .c(_17458_),
    .d(_16078_),
    .o1(_01995_));
 b15ao0012al1n03x5 _27900_ (.a(_01995_),
    .b(_17420_),
    .c(_16047_),
    .o(_01996_));
 b15oai012an1n02x5 _27901_ (.a(net879),
    .b(_16047_),
    .c(_16058_),
    .o1(_01997_));
 b15oai112aq1n08x5 _27902_ (.a(net875),
    .b(_01997_),
    .c(_17458_),
    .d(net879),
    .o1(_01998_));
 b15oai112as1n04x5 _27903_ (.a(net882),
    .b(_16078_),
    .c(_16045_),
    .d(_16058_),
    .o1(_01999_));
 b15oai112al1n12x5 _27904_ (.a(_16018_),
    .b(_01999_),
    .c(_16040_),
    .d(_15997_),
    .o1(_02000_));
 b15aoai13ah1n08x5 _27905_ (.a(net874),
    .b(_01996_),
    .c(_01998_),
    .d(_02000_),
    .o1(_02001_));
 b15nand04as1n16x5 _27906_ (.a(_01966_),
    .b(_01982_),
    .c(_01994_),
    .d(_02001_),
    .o1(_02002_));
 b15aoi022ar1n02x5 _27907_ (.a(_16774_),
    .b(_16888_),
    .c(_16772_),
    .d(net763),
    .o1(_02003_));
 b15oai012ar1n02x5 _27908_ (.a(_16832_),
    .b(_16783_),
    .c(_16888_),
    .o1(_02004_));
 b15aoi012aq1n02x5 _27909_ (.a(_16741_),
    .b(_02003_),
    .c(_02004_),
    .o1(_02005_));
 b15nor004an1n03x5 _27910_ (.a(net764),
    .b(net751),
    .c(_00783_),
    .d(_01355_),
    .o1(_02006_));
 b15aoi012an1n02x5 _27911_ (.a(_16748_),
    .b(_16775_),
    .c(net763),
    .o1(_02007_));
 b15nor003ar1n02x5 _27912_ (.a(net759),
    .b(_16888_),
    .c(_16855_),
    .o1(_02008_));
 b15norp03ah1n04x5 _27913_ (.a(_02006_),
    .b(_02007_),
    .c(_02008_),
    .o1(_02009_));
 b15aoi022ar1n02x5 _27914_ (.a(net766),
    .b(_16758_),
    .c(_16846_),
    .d(_16896_),
    .o1(_02010_));
 b15oai022ah1n02x5 _27915_ (.a(_16897_),
    .b(_16855_),
    .c(_02010_),
    .d(_16770_),
    .o1(_02011_));
 b15nandp2ah1n03x5 _27916_ (.a(net759),
    .b(_02011_),
    .o1(_02012_));
 b15aoi013aq1n08x5 _27917_ (.a(_02005_),
    .b(_02009_),
    .c(_02012_),
    .d(_16741_),
    .o1(_02013_));
 b15nano22ar1n02x5 _27918_ (.a(net753),
    .b(net744),
    .c(net757),
    .out0(_02014_));
 b15oai112as1n02x5 _27919_ (.a(_16881_),
    .b(_16872_),
    .c(_01127_),
    .d(_02014_),
    .o1(_02015_));
 b15nandp2ar1n05x5 _27920_ (.a(net767),
    .b(_17337_),
    .o1(_02016_));
 b15oai012al1n03x5 _27921_ (.a(_16693_),
    .b(net757),
    .c(_16742_),
    .o1(_02017_));
 b15aoi013an1n04x5 _27922_ (.a(_02015_),
    .b(_02016_),
    .c(_02017_),
    .d(_16770_),
    .o1(_02018_));
 b15oai012al1n06x5 _27923_ (.a(net757),
    .b(_16907_),
    .c(_17314_),
    .o1(_02019_));
 b15oai112as1n06x5 _27924_ (.a(_16774_),
    .b(_16897_),
    .c(_00730_),
    .d(net765),
    .o1(_02020_));
 b15aoi013al1n08x5 _27925_ (.a(_02018_),
    .b(_02019_),
    .c(_02020_),
    .d(net754),
    .o1(_02021_));
 b15aoi012an1n04x5 _27926_ (.a(_01301_),
    .b(_16788_),
    .c(_17298_),
    .o1(_02022_));
 b15nor003ah1n08x5 _27927_ (.a(_16839_),
    .b(_00751_),
    .c(_02022_),
    .o1(_02023_));
 b15nand02an1n04x5 _27928_ (.a(_16798_),
    .b(_16788_),
    .o1(_02024_));
 b15oai222ah1n12x5 _27929_ (.a(_00722_),
    .b(_17314_),
    .c(_01308_),
    .d(_17373_),
    .e(_02024_),
    .f(_16832_),
    .o1(_02025_));
 b15oai022ah1n06x5 _27930_ (.a(_16713_),
    .b(_16897_),
    .c(_00719_),
    .d(_16903_),
    .o1(_02026_));
 b15aoi112ar1n08x5 _27931_ (.a(_02023_),
    .b(_02025_),
    .c(net765),
    .d(_02026_),
    .o1(_02027_));
 b15aoi012ah1n02x5 _27932_ (.a(net758),
    .b(_01111_),
    .c(_16887_),
    .o1(_02028_));
 b15aoi112ar1n06x5 _27933_ (.a(_16786_),
    .b(_02028_),
    .c(_16834_),
    .d(_16775_),
    .o1(_02029_));
 b15nand02ar1n02x5 _27934_ (.a(net765),
    .b(_16905_),
    .o1(_02030_));
 b15oaoi13ar1n03x5 _27935_ (.a(net754),
    .b(_02030_),
    .c(_17382_),
    .d(_16810_),
    .o1(_02031_));
 b15nor003aq1n06x5 _27936_ (.a(_01518_),
    .b(_02029_),
    .c(_02031_),
    .o1(_02032_));
 b15nand04an1n16x5 _27937_ (.a(_00710_),
    .b(_02021_),
    .c(_02027_),
    .d(_02032_),
    .o1(_02033_));
 b15oai112ar1n02x5 _27938_ (.a(net755),
    .b(_16897_),
    .c(_16898_),
    .d(_00730_),
    .o1(_02034_));
 b15oai012ar1n04x5 _27939_ (.a(_02034_),
    .b(_01702_),
    .c(net755),
    .o1(_02035_));
 b15aoi012aq1n02x5 _27940_ (.a(_16827_),
    .b(_00773_),
    .c(_16693_),
    .o1(_02036_));
 b15oaoi13as1n04x5 _27941_ (.a(net762),
    .b(_02035_),
    .c(_02036_),
    .d(_01532_),
    .o1(_02037_));
 b15aoi013aq1n03x5 _27942_ (.a(_17337_),
    .b(_16726_),
    .c(_16785_),
    .d(net767),
    .o1(_02038_));
 b15oaoi13ah1n04x5 _27943_ (.a(_16774_),
    .b(_02016_),
    .c(_02038_),
    .d(net760),
    .o1(_02039_));
 b15aoi022as1n04x5 _27944_ (.a(_16785_),
    .b(_16726_),
    .c(_17337_),
    .d(net760),
    .o1(_02040_));
 b15aoi013ar1n06x5 _27945_ (.a(_16770_),
    .b(_01723_),
    .c(_01544_),
    .d(_01711_),
    .o1(_02041_));
 b15nand02aq1n04x5 _27946_ (.a(net765),
    .b(net752),
    .o1(_02042_));
 b15aoi013ar1n08x5 _27947_ (.a(net761),
    .b(_16710_),
    .c(_16804_),
    .d(_02042_),
    .o1(_02043_));
 b15oai122an1n16x5 _27948_ (.a(net756),
    .b(_17339_),
    .c(_02040_),
    .d(_02041_),
    .e(_02043_),
    .o1(_02044_));
 b15nand03al1n12x5 _27949_ (.a(_16774_),
    .b(_16785_),
    .c(_16726_),
    .o1(_02045_));
 b15oai122al1n16x5 _27950_ (.a(_16741_),
    .b(_16898_),
    .c(_16793_),
    .d(_17367_),
    .e(_02045_),
    .o1(_02046_));
 b15oaoi13an1n04x5 _27951_ (.a(_16770_),
    .b(_16903_),
    .c(_02045_),
    .d(_16693_),
    .o1(_02047_));
 b15oai022ar1n16x5 _27952_ (.a(_02039_),
    .b(_02044_),
    .c(_02046_),
    .d(_02047_),
    .o1(_02048_));
 b15nandp2an1n02x5 _27953_ (.a(_16815_),
    .b(_16806_),
    .o1(_02049_));
 b15nandp3ar1n03x5 _27954_ (.a(net752),
    .b(_01051_),
    .c(_16726_),
    .o1(_02050_));
 b15aoi012as1n04x5 _27955_ (.a(_01119_),
    .b(_02049_),
    .c(_02050_),
    .o1(_02051_));
 b15nand02as1n02x5 _27956_ (.a(_16708_),
    .b(_16768_),
    .o1(_02052_));
 b15oai013an1n12x5 _27957_ (.a(_02052_),
    .b(_00772_),
    .c(_16713_),
    .d(_16731_),
    .o1(_02053_));
 b15aoai13ar1n08x5 _27958_ (.a(_16770_),
    .b(_02051_),
    .c(_02053_),
    .d(net752),
    .o1(_02054_));
 b15oai013ah1n03x5 _27959_ (.a(_01290_),
    .b(_16908_),
    .c(_00730_),
    .d(_16856_),
    .o1(_02055_));
 b15oai122al1n08x5 _27960_ (.a(_16693_),
    .b(_16764_),
    .c(_16713_),
    .d(_16748_),
    .e(_00719_),
    .o1(_02056_));
 b15nand04ar1n04x5 _27961_ (.a(net758),
    .b(_16702_),
    .c(_16708_),
    .d(_16813_),
    .o1(_02057_));
 b15aob012aq1n06x5 _27962_ (.a(_02057_),
    .b(_16912_),
    .c(net754),
    .out0(_02058_));
 b15oaoi13as1n04x5 _27963_ (.a(_02055_),
    .b(_02056_),
    .c(_16693_),
    .d(_02058_),
    .o1(_02059_));
 b15nand04ah1n16x5 _27964_ (.a(_16721_),
    .b(_02048_),
    .c(_02054_),
    .d(_02059_),
    .o1(_02060_));
 b15nor004as1n12x5 _27965_ (.a(_02013_),
    .b(_02033_),
    .c(_02037_),
    .d(_02060_),
    .o1(_02061_));
 b15xor002al1n02x5 _27966_ (.a(_02002_),
    .b(_02061_),
    .out0(_02062_));
 b15xor002ar1n03x5 _27967_ (.a(_01871_),
    .b(_02062_),
    .out0(_02063_));
 b15nonb03ar1n02x5 _27968_ (.a(\us13.a[7] ),
    .b(\us13.a[3] ),
    .c(net604),
    .out0(_02064_));
 b15aoi012ar1n02x5 _27969_ (.a(_02064_),
    .b(_16542_),
    .c(net604),
    .o1(_02065_));
 b15norp03ah1n02x5 _27970_ (.a(_17093_),
    .b(_17088_),
    .c(_02065_),
    .o1(_02066_));
 b15oai112al1n02x5 _27971_ (.a(net603),
    .b(_16494_),
    .c(_16558_),
    .d(net605),
    .o1(_02067_));
 b15aoai13al1n02x5 _27972_ (.a(_16659_),
    .b(\us13.a[3] ),
    .c(_16558_),
    .d(net599),
    .o1(_02068_));
 b15oaoi13as1n03x5 _27973_ (.a(_16458_),
    .b(_02067_),
    .c(_02068_),
    .d(net603),
    .o1(_02069_));
 b15oaoi13an1n04x5 _27974_ (.a(_02066_),
    .b(_16460_),
    .c(_01898_),
    .d(_02069_),
    .o1(_02070_));
 b15nonb03al1n02x5 _27975_ (.a(net605),
    .b(net598),
    .c(net609),
    .out0(_02071_));
 b15oai013ah1n04x5 _27976_ (.a(_02071_),
    .b(_01561_),
    .c(_00894_),
    .d(net603),
    .o1(_02072_));
 b15nand04an1n08x5 _27977_ (.a(net609),
    .b(_16481_),
    .c(_16520_),
    .d(_16478_),
    .o1(_02073_));
 b15and003aq1n03x5 _27978_ (.a(_16456_),
    .b(_02072_),
    .c(_02073_),
    .o(_02074_));
 b15oai012ar1n12x5 _27979_ (.a(_17541_),
    .b(_16528_),
    .c(_16479_),
    .o1(_02075_));
 b15aoi012as1n02x5 _27980_ (.a(_16429_),
    .b(_16517_),
    .c(_16466_),
    .o1(_02076_));
 b15oai112al1n12x5 _27981_ (.a(_02072_),
    .b(_02073_),
    .c(_16667_),
    .d(_02076_),
    .o1(_02077_));
 b15nand02an1n02x5 _27982_ (.a(_16481_),
    .b(_16621_),
    .o1(_02078_));
 b15oai013an1n08x5 _27983_ (.a(_02078_),
    .b(_16538_),
    .c(_01931_),
    .d(\us13.a[3] ),
    .o1(_02079_));
 b15aoi122al1n08x5 _27984_ (.a(_02075_),
    .b(_02077_),
    .c(\us13.a[0] ),
    .d(_02079_),
    .e(net598),
    .o1(_02080_));
 b15oai022aq1n16x5 _27985_ (.a(net617),
    .b(_02070_),
    .c(_02074_),
    .d(_02080_),
    .o1(_02081_));
 b15nor002aq1n02x5 _27986_ (.a(_16516_),
    .b(_17125_),
    .o1(_02082_));
 b15aoi013ar1n06x5 _27987_ (.a(_02082_),
    .b(_01920_),
    .c(_17559_),
    .d(_17097_),
    .o1(_02083_));
 b15nand02an1n02x5 _27988_ (.a(_16585_),
    .b(_00858_),
    .o1(_02084_));
 b15aoi022al1n06x5 _27989_ (.a(_16435_),
    .b(_01561_),
    .c(_02084_),
    .d(net612),
    .o1(_02085_));
 b15oaoi13ah1n04x5 _27990_ (.a(net610),
    .b(_02083_),
    .c(_02085_),
    .d(_00859_),
    .o1(_02086_));
 b15oai012an1n02x5 _27991_ (.a(_16519_),
    .b(_17131_),
    .c(_16456_),
    .o1(_02087_));
 b15nandp2al1n02x5 _27992_ (.a(net606),
    .b(_16677_),
    .o1(_02088_));
 b15oai022aq1n06x5 _27993_ (.a(_16667_),
    .b(_16513_),
    .c(_17139_),
    .d(_02088_),
    .o1(_02089_));
 b15aoai13ah1n03x5 _27994_ (.a(_16460_),
    .b(_02087_),
    .c(_02089_),
    .d(net604),
    .o1(_02090_));
 b15aoi012as1n02x5 _27995_ (.a(_01248_),
    .b(_17176_),
    .c(_17177_),
    .o1(_02091_));
 b15oai022aq1n02x5 _27996_ (.a(_17602_),
    .b(_17116_),
    .c(_17578_),
    .d(_16516_),
    .o1(_02092_));
 b15aoi012al1n06x5 _27997_ (.a(_02091_),
    .b(_02092_),
    .c(_16466_),
    .o1(_02093_));
 b15nand04ah1n12x5 _27998_ (.a(_16468_),
    .b(_01895_),
    .c(_02090_),
    .d(_02093_),
    .o1(_02094_));
 b15norp03ah1n08x5 _27999_ (.a(_16538_),
    .b(_17139_),
    .c(_01561_),
    .o1(_02095_));
 b15nandp2ah1n02x5 _28000_ (.a(_16558_),
    .b(_17166_),
    .o1(_02096_));
 b15aoi012ar1n04x5 _28001_ (.a(_16504_),
    .b(_16521_),
    .c(_16613_),
    .o1(_02097_));
 b15oai112al1n12x5 _28002_ (.a(_02095_),
    .b(_02096_),
    .c(_02097_),
    .d(_16558_),
    .o1(_02098_));
 b15aoai13ar1n02x5 _28003_ (.a(_17152_),
    .b(_17562_),
    .c(_16473_),
    .d(_16475_),
    .o1(_02099_));
 b15oaoi13as1n02x5 _28004_ (.a(net611),
    .b(_02099_),
    .c(_17116_),
    .d(_16498_),
    .o1(_02100_));
 b15oai012ar1n04x5 _28005_ (.a(_16558_),
    .b(net615),
    .c(_16519_),
    .o1(_02101_));
 b15nand02ar1n02x5 _28006_ (.a(_16659_),
    .b(_16473_),
    .o1(_02102_));
 b15mdn022al1n03x5 _28007_ (.a(_16591_),
    .b(_00847_),
    .o1(_02103_),
    .sa(_17099_));
 b15oai012ar1n04x5 _28008_ (.a(_16519_),
    .b(_02102_),
    .c(_02103_),
    .o1(_02104_));
 b15aoi012aq1n06x5 _28009_ (.a(_02100_),
    .b(_02101_),
    .c(_02104_),
    .o1(_02105_));
 b15norp03ar1n02x5 _28010_ (.a(_16466_),
    .b(_16575_),
    .c(_16673_),
    .o1(_02106_));
 b15nand03ar1n03x5 _28011_ (.a(_16667_),
    .b(_16549_),
    .c(_02106_),
    .o1(_02107_));
 b15norp03al1n02x5 _28012_ (.a(_16458_),
    .b(_16439_),
    .c(_16632_),
    .o1(_02108_));
 b15aoai13al1n02x5 _28013_ (.a(_02108_),
    .b(_01577_),
    .c(_17110_),
    .d(_16579_),
    .o1(_02109_));
 b15aoi022ar1n02x5 _28014_ (.a(net610),
    .b(_16481_),
    .c(_16517_),
    .d(_16544_),
    .o1(_02110_));
 b15orn003al1n02x5 _28015_ (.a(_16667_),
    .b(_17602_),
    .c(_02110_),
    .o(_02111_));
 b15and003ah1n04x5 _28016_ (.a(_02107_),
    .b(_02109_),
    .c(_02111_),
    .o(_02112_));
 b15nand03al1n03x5 _28017_ (.a(_16609_),
    .b(_17553_),
    .c(_17545_),
    .o1(_02113_));
 b15oai012an1n06x5 _28018_ (.a(_02113_),
    .b(_16642_),
    .c(_16521_),
    .o1(_02114_));
 b15nand03al1n02x5 _28019_ (.a(_16577_),
    .b(_16517_),
    .c(_01212_),
    .o1(_02115_));
 b15oai013as1n04x5 _28020_ (.a(_02115_),
    .b(_16528_),
    .c(_16592_),
    .d(_16522_),
    .o1(_02116_));
 b15nor002an1n03x5 _28021_ (.a(_01877_),
    .b(_17175_),
    .o1(_02117_));
 b15oai022an1n08x5 _28022_ (.a(net610),
    .b(_16586_),
    .c(_17139_),
    .d(_01910_),
    .o1(_02118_));
 b15aoi112ar1n08x5 _28023_ (.a(_02114_),
    .b(_02116_),
    .c(_02117_),
    .d(_02118_),
    .o1(_02119_));
 b15nand04as1n16x5 _28024_ (.a(_02098_),
    .b(_02105_),
    .c(_02112_),
    .d(_02119_),
    .o1(_02120_));
 b15nor004as1n12x5 _28025_ (.a(_02081_),
    .b(_02086_),
    .c(_02094_),
    .d(_02120_),
    .o1(_02121_));
 b15xor002as1n16x5 _28026_ (.a(_17068_),
    .b(_02121_),
    .out0(_02122_));
 b15xor002ar1n03x5 _28027_ (.a(_02063_),
    .b(_02122_),
    .out0(_02123_));
 b15cmbn22al1n08x5 _28028_ (.clk1(\text_in_r[39] ),
    .clk2(_02123_),
    .clkout(_02124_),
    .s(net539));
 b15xor002as1n16x5 _28029_ (.a(\u0.w[2][7] ),
    .b(_02124_),
    .out0(_00120_));
 b15bfn000as1n02x5 input13 (.a(key[110]),
    .o(net13));
 b15xor002as1n16x5 _28031_ (.a(_16926_),
    .b(_02002_),
    .out0(_02126_));
 b15xor003an1n16x5 _28032_ (.a(_16690_),
    .b(_17396_),
    .c(_02126_),
    .out0(_02127_));
 b15norp02al1n12x5 _28033_ (.a(net539),
    .b(_02127_),
    .o1(_02128_));
 b15inv040ah1n02x5 _28034_ (.a(\text_in_r[40] ),
    .o1(_02129_));
 b15aoi012aq1n04x5 _28035_ (.a(_02128_),
    .b(_02129_),
    .c(net539),
    .o1(_02130_));
 b15xor002ar1n08x5 _28036_ (.a(net529),
    .b(_02130_),
    .out0(_00081_));
 b15inv020ah1n04x5 _28037_ (.a(\text_in_r[41] ),
    .o1(_02131_));
 b15xor002an1n12x5 _28038_ (.a(_17282_),
    .b(_02126_),
    .out0(_02132_));
 b15xor002as1n08x5 _28039_ (.a(_16168_),
    .b(_17396_),
    .out0(_02133_));
 b15xor002as1n08x5 _28040_ (.a(_00818_),
    .b(_02133_),
    .out0(_02134_));
 b15xor002as1n16x5 _28041_ (.a(_02132_),
    .b(_02134_),
    .out0(_02135_));
 b15mdn022ar1n12x5 _28042_ (.a(_02131_),
    .b(_02135_),
    .o1(_02136_),
    .sa(net539));
 b15xor002ar1n02x5 _28043_ (.a(net528),
    .b(_02136_),
    .out0(_00082_));
 b15xor002as1n12x5 _28044_ (.a(_17526_),
    .b(_00818_),
    .out0(_02137_));
 b15xnr002ah1n08x5 _28045_ (.a(_17615_),
    .b(_02137_),
    .out0(_02138_));
 b15xor002ah1n12x5 _28046_ (.a(_01139_),
    .b(_02138_),
    .out0(_02139_));
 b15cmbn22as1n03x5 _28047_ (.clk1(\text_in_r[42] ),
    .clk2(_02139_),
    .clkout(_02140_),
    .s(net539));
 b15xor002ar1n02x5 _28048_ (.a(\u0.w[2][10] ),
    .b(_02140_),
    .out0(_00083_));
 b15inv040ah1n02x5 _28049_ (.a(\text_in_r[43] ),
    .o1(_02141_));
 b15xor002as1n08x5 _28050_ (.a(_00974_),
    .b(_01138_),
    .out0(_02142_));
 b15xor002ah1n04x5 _28051_ (.a(_00618_),
    .b(_01364_),
    .out0(_02143_));
 b15xor002as1n08x5 _28052_ (.a(_02126_),
    .b(_02143_),
    .out0(_02144_));
 b15xor002ah1n16x5 _28053_ (.a(_02142_),
    .b(_02144_),
    .out0(_02145_));
 b15mdn022an1n04x5 _28054_ (.a(_02141_),
    .b(_02145_),
    .o1(_02146_),
    .sa(net539));
 b15xor002ar1n02x5 _28055_ (.a(\u0.w[2][11] ),
    .b(_02146_),
    .out0(_00084_));
 b15xor002ar1n08x5 _28056_ (.a(_01286_),
    .b(_02126_),
    .out0(_02147_));
 b15xor002as1n12x5 _28057_ (.a(_01049_),
    .b(_01364_),
    .out0(_02148_));
 b15xor002ar1n12x5 _28058_ (.a(_01557_),
    .b(_02148_),
    .out0(_02149_));
 b15xor002as1n06x5 _28059_ (.a(_02147_),
    .b(_02149_),
    .out0(_02150_));
 b15cmbn22as1n04x5 _28060_ (.clk1(\text_in_r[44] ),
    .clk2(_02150_),
    .clkout(_02151_),
    .s(net539));
 b15xor002ah1n12x5 _28061_ (.a(\u0.w[2][12] ),
    .b(_02151_),
    .out0(_00085_));
 b15inv020aq1n08x5 _28062_ (.a(\text_in_r[45] ),
    .o1(_02152_));
 b15xnr002aq1n12x5 _28063_ (.a(_01426_),
    .b(_01557_),
    .out0(_02153_));
 b15xor002as1n06x5 _28064_ (.a(_01754_),
    .b(_02153_),
    .out0(_02154_));
 b15xor002an1n12x5 _28065_ (.a(_01690_),
    .b(_02154_),
    .out0(_02155_));
 b15bfn000ah1n03x5 input12 (.a(key[10]),
    .o(net12));
 b15mdn022al1n16x5 _28067_ (.a(_02152_),
    .b(_02155_),
    .o1(_02157_),
    .sa(net539));
 b15xor002ah1n16x5 _28068_ (.a(\u0.w[2][13] ),
    .b(_02157_),
    .out0(_00086_));
 b15nand02al1n04x5 _28069_ (.a(net539),
    .b(\text_in_r[46] ),
    .o1(_02158_));
 b15xor002al1n16x5 _28070_ (.a(_01500_),
    .b(_01754_),
    .out0(_02159_));
 b15xor002an1n08x5 _28071_ (.a(_02061_),
    .b(_02159_),
    .out0(_02160_));
 b15xor002ah1n04x5 _28072_ (.a(_01941_),
    .b(_02160_),
    .out0(_02161_));
 b15oai012ah1n08x5 _28073_ (.a(_02158_),
    .b(_02161_),
    .c(net539),
    .o1(_02162_));
 b15xor002as1n12x5 _28074_ (.a(\u0.w[2][14] ),
    .b(_02162_),
    .out0(_00087_));
 b15inv000as1n04x5 _28075_ (.a(\text_in_r[47] ),
    .o1(_02163_));
 b15xor002an1n12x5 _28076_ (.a(_01813_),
    .b(_02061_),
    .out0(_02164_));
 b15xor002ah1n04x5 _28077_ (.a(_16926_),
    .b(_02164_),
    .out0(_02165_));
 b15xor002as1n08x5 _28078_ (.a(_02122_),
    .b(_02165_),
    .out0(_02166_));
 b15mdn022ar1n16x5 _28079_ (.a(_02163_),
    .b(_02166_),
    .o1(_02167_),
    .sa(net539));
 b15xor002aq1n16x5 _28080_ (.a(\u0.w[2][15] ),
    .b(_02167_),
    .out0(_00088_));
 b15xnr002as1n16x5 _28081_ (.a(_02002_),
    .b(_02121_),
    .out0(_02168_));
 b15xor003ar1n03x5 _28082_ (.a(_16424_),
    .b(_02133_),
    .c(_02168_),
    .out0(_02169_));
 b15norp02aq1n02x5 _28083_ (.a(net540),
    .b(_02169_),
    .o1(_02170_));
 b15inv020as1n06x5 _28084_ (.a(\text_in_r[48] ),
    .o1(_02171_));
 b15bfn000ah1n04x5 input11 (.a(key[109]),
    .o(net11));
 b15aoi012aq1n06x5 _28086_ (.a(_02170_),
    .b(_02171_),
    .c(net540),
    .o1(_02173_));
 b15xor002as1n06x5 _28087_ (.a(net527),
    .b(_02173_),
    .out0(_00049_));
 b15xor003ar1n04x5 _28088_ (.a(_16168_),
    .b(_16689_),
    .c(_17281_),
    .out0(_02174_));
 b15xor002ar1n03x5 _28089_ (.a(_02137_),
    .b(_02174_),
    .out0(_02175_));
 b15xor002al1n02x5 _28090_ (.a(_02168_),
    .b(_02175_),
    .out0(_02176_));
 b15cmbn22ah1n04x5 _28091_ (.clk1(\text_in_r[49] ),
    .clk2(_02176_),
    .clkout(_02177_),
    .s(net540));
 b15xor002an1n12x5 _28092_ (.a(net526),
    .b(_02177_),
    .out0(_00050_));
 b15inv000as1n06x5 _28093_ (.a(\text_in_r[50] ),
    .o1(_02178_));
 b15xor002aq1n02x5 _28094_ (.a(_17526_),
    .b(_00618_),
    .out0(_02179_));
 b15xor002as1n03x5 _28095_ (.a(_17196_),
    .b(_02179_),
    .out0(_02180_));
 b15xor002ah1n06x5 _28096_ (.a(_01139_),
    .b(_02180_),
    .out0(_02181_));
 b15mdn022al1n16x5 _28097_ (.a(_02178_),
    .b(_02181_),
    .o1(_02182_),
    .sa(net539));
 b15xor002as1n08x5 _28098_ (.a(net525),
    .b(_02182_),
    .out0(_00051_));
 b15inv000as1n03x5 _28099_ (.a(\text_in_r[51] ),
    .o1(_02183_));
 b15xnr002ar1n12x5 _28100_ (.a(_00973_),
    .b(_02148_),
    .out0(_02184_));
 b15xor002an1n08x5 _28101_ (.a(_00619_),
    .b(_02168_),
    .out0(_02185_));
 b15xor002ar1n12x5 _28102_ (.a(_02184_),
    .b(_02185_),
    .out0(_02186_));
 b15mdn022al1n12x5 _28103_ (.a(_02183_),
    .b(_02186_),
    .o1(_02187_),
    .sa(net540));
 b15xor002ar1n03x5 _28104_ (.a(net524),
    .b(_02187_),
    .out0(_00052_));
 b15inv000ar1n12x5 _28105_ (.a(\text_in_r[52] ),
    .o1(_02188_));
 b15xor002aq1n06x5 _28106_ (.a(_01209_),
    .b(_02153_),
    .out0(_02189_));
 b15xnr002ar1n12x5 _28107_ (.a(_00905_),
    .b(_01049_),
    .out0(_02190_));
 b15xor003ar1n16x5 _28108_ (.a(_02168_),
    .b(_02189_),
    .c(_02190_),
    .out0(_02191_));
 b15mdn022ah1n12x5 _28109_ (.a(_02188_),
    .b(_02191_),
    .o1(_02192_),
    .sa(net540));
 b15xor002ah1n16x5 _28110_ (.a(\u0.w[2][20] ),
    .b(_02192_),
    .out0(_00053_));
 b15xor003an1n02x5 _28111_ (.a(_01285_),
    .b(_01426_),
    .c(_01689_),
    .out0(_02193_));
 b15xor002al1n02x5 _28112_ (.a(_02159_),
    .b(_02193_),
    .out0(_02194_));
 b15nor002ar1n03x5 _28113_ (.a(net540),
    .b(_02194_),
    .o1(_02195_));
 b15inv040as1n04x5 _28114_ (.a(\text_in_r[53] ),
    .o1(_02196_));
 b15aoi012al1n08x5 _28115_ (.a(_02195_),
    .b(_02196_),
    .c(net540),
    .o1(_02197_));
 b15xor002an1n12x5 _28116_ (.a(\u0.w[2][21] ),
    .b(_02197_),
    .out0(_00054_));
 b15xor002ar1n03x5 _28117_ (.a(_01871_),
    .b(_02164_),
    .out0(_02198_));
 b15xor002ar1n02x5 _28118_ (.a(_01500_),
    .b(_01620_),
    .out0(_02199_));
 b15xor002al1n02x5 _28119_ (.a(_02198_),
    .b(_02199_),
    .out0(_02200_));
 b15bfn000as1n03x5 input10 (.a(key[108]),
    .o(net10));
 b15cmbn22ah1n04x5 _28121_ (.clk1(\text_in_r[54] ),
    .clk2(_02200_),
    .clkout(_02202_),
    .s(net540));
 b15xor002as1n08x5 _28122_ (.a(\u0.w[2][22] ),
    .b(_02202_),
    .out0(_00055_));
 b15inv040aq1n06x5 _28123_ (.a(\text_in_r[55] ),
    .o1(_02203_));
 b15xor002ar1n03x5 _28124_ (.a(_17068_),
    .b(_01813_),
    .out0(_02204_));
 b15xor002aq1n03x5 _28125_ (.a(_01940_),
    .b(_02204_),
    .out0(_02205_));
 b15xor002ah1n03x5 _28126_ (.a(_02126_),
    .b(_02205_),
    .out0(_02206_));
 b15mdn022aq1n12x5 _28127_ (.a(_02203_),
    .b(_02206_),
    .o1(_02207_),
    .sa(net539));
 b15xor002ah1n06x5 _28128_ (.a(\u0.w[2][23] ),
    .b(_02207_),
    .out0(_00056_));
 b15inv000ar1n16x5 _28129_ (.a(\text_in_r[56] ),
    .o1(_02208_));
 b15xor002al1n02x5 _28130_ (.a(_16689_),
    .b(_02133_),
    .out0(_02209_));
 b15xor002an1n02x5 _28131_ (.a(_02122_),
    .b(_02209_),
    .out0(_02210_));
 b15mdn022al1n04x5 _28132_ (.a(_02208_),
    .b(_02210_),
    .o1(_02211_),
    .sa(net540));
 b15xor002ah1n03x5 _28133_ (.a(net523),
    .b(_02211_),
    .out0(_00017_));
 b15inv020as1n05x5 _28134_ (.a(\text_in_r[57] ),
    .o1(_02212_));
 b15xnr002an1n06x5 _28135_ (.a(_17196_),
    .b(_02137_),
    .out0(_02213_));
 b15xor002ah1n03x5 _28136_ (.a(_16690_),
    .b(_02122_),
    .out0(_02214_));
 b15xor002as1n06x5 _28137_ (.a(_02213_),
    .b(_02214_),
    .out0(_02215_));
 b15mdn022aq1n04x5 _28138_ (.a(_02212_),
    .b(_02215_),
    .o1(_02216_),
    .sa(net539));
 b15xor002an1n08x5 _28139_ (.a(net522),
    .b(_02216_),
    .out0(_00018_));
 b15xor002ar1n03x5 _28140_ (.a(_17282_),
    .b(_01138_),
    .out0(_02217_));
 b15xor002as1n02x5 _28141_ (.a(_00619_),
    .b(_02217_),
    .out0(_02218_));
 b15cmbn22ah1n03x5 _28142_ (.clk1(\text_in_r[58] ),
    .clk2(_02218_),
    .clkout(_02219_),
    .s(net539));
 b15xor002an1n12x5 _28143_ (.a(net521),
    .b(_02219_),
    .out0(_00019_));
 b15xor002ar1n02x5 _28144_ (.a(_00706_),
    .b(_00905_),
    .out0(_02220_));
 b15xor002al1n02x5 _28145_ (.a(_17615_),
    .b(_02220_),
    .out0(_02221_));
 b15xor002an1n02x5 _28146_ (.a(_02122_),
    .b(_02148_),
    .out0(_02222_));
 b15xor002ar1n02x5 _28147_ (.a(_02221_),
    .b(_02222_),
    .out0(_02223_));
 b15cmbn22ar1n02x5 _28148_ (.clk1(\text_in_r[59] ),
    .clk2(_02223_),
    .clkout(_02224_),
    .s(net540));
 b15xor002ar1n03x5 _28149_ (.a(\u0.w[2][27] ),
    .b(_02224_),
    .out0(_00020_));
 b15inv040as1n04x5 _28150_ (.a(\text_in_r[60] ),
    .o1(_02225_));
 b15xor002al1n03x5 _28151_ (.a(_01285_),
    .b(_02153_),
    .out0(_02226_));
 b15xor002al1n02x5 _28152_ (.a(_00974_),
    .b(_02122_),
    .out0(_02227_));
 b15xor002ar1n03x5 _28153_ (.a(_02226_),
    .b(_02227_),
    .out0(_02228_));
 b15mdn022ah1n02x5 _28154_ (.a(_02225_),
    .b(_02228_),
    .o1(_02229_),
    .sa(net539));
 b15xor002ah1n03x5 _28155_ (.a(\u0.w[2][28] ),
    .b(_02229_),
    .out0(_00021_));
 b15xor003ar1n02x5 _28156_ (.a(_01286_),
    .b(_01620_),
    .c(_02159_),
    .out0(_02230_));
 b15norp02ar1n02x5 _28157_ (.a(net539),
    .b(_02230_),
    .o1(_02231_));
 b15inv000an1n04x5 _28158_ (.a(\text_in_r[61] ),
    .o1(_02232_));
 b15aoi012an1n02x5 _28159_ (.a(_02231_),
    .b(_02232_),
    .c(net540),
    .o1(_02233_));
 b15xor002al1n04x5 _28160_ (.a(\u0.w[2][29] ),
    .b(_02233_),
    .out0(_00022_));
 b15xor002ar1n04x5 _28161_ (.a(_01940_),
    .b(_02164_),
    .out0(_02234_));
 b15xor002an1n04x5 _28162_ (.a(_01690_),
    .b(_02234_),
    .out0(_02235_));
 b15cmbn22ar1n02x5 _28163_ (.clk1(\text_in_r[62] ),
    .clk2(_02235_),
    .clkout(_02236_),
    .s(net540));
 b15xor002as1n02x5 _28164_ (.a(\u0.w[2][30] ),
    .b(_02236_),
    .out0(_00023_));
 b15inv040ah1n02x5 _28165_ (.a(\text_in_r[63] ),
    .o1(_02237_));
 b15qgbxo2an1n05x5 _28166_ (.a(_02121_),
    .b(_02126_),
    .out0(_02238_));
 b15xor002an1n03x5 _28167_ (.a(_01941_),
    .b(_02238_),
    .out0(_02239_));
 b15mdn022as1n04x5 _28168_ (.a(_02237_),
    .b(_02239_),
    .o1(_02240_),
    .sa(net539));
 b15xor002ar1n12x5 _28169_ (.a(\u0.w[2][31] ),
    .b(_02240_),
    .out0(_00024_));
 b15bfn000ah1n02x5 input9 (.a(key[107]),
    .o(net9));
 b15inv000as1n48x5 _28171_ (.a(net711),
    .o1(_02242_));
 b15bfm201ah1n02x5 input8 (.a(key[106]),
    .o(net8));
 b15bfn000ah1n02x5 input7 (.a(key[105]),
    .o(net7));
 b15bfn000ar1n02x5 input6 (.a(key[104]),
    .o(net6));
 b15bfn001ah1n12x5 input5 (.a(key[103]),
    .o(net5));
 b15bfn001ah1n08x5 input4 (.a(key[102]),
    .o(net4));
 b15bfn000as1n02x5 input3 (.a(key[101]),
    .o(net3));
 b15bfn000as1n02x5 input2 (.a(key[100]),
    .o(net2));
 b15bfn000aq1n02x5 input1 (.a(key[0]),
    .o(net1));
 b15norp02al1n48x5 _28180_ (.a(net706),
    .b(net701),
    .o1(_02251_));
 b15ztpn00an1n08x5 TAP_780 ();
 b15ztpn00an1n08x5 TAP_779 ();
 b15ztpn00an1n08x5 TAP_778 ();
 b15ztpn00an1n08x5 TAP_777 ();
 b15ztpn00an1n08x5 TAP_776 ();
 b15nandp3as1n04x5 _28186_ (.a(net698),
    .b(net693),
    .c(\us12.a[6] ),
    .o1(_02257_));
 b15ztpn00an1n08x5 TAP_775 ();
 b15orn002as1n32x5 _28188_ (.a(\us12.a[7] ),
    .b(\us12.a[6] ),
    .o(_02259_));
 b15ztpn00an1n08x5 TAP_774 ();
 b15ztpn00an1n08x5 TAP_773 ();
 b15oai012an1n12x5 _28191_ (.a(_02257_),
    .b(_02259_),
    .c(net698),
    .o1(_02262_));
 b15and002al1n02x5 _28192_ (.a(_02251_),
    .b(_02262_),
    .o(_02263_));
 b15ztpn00an1n08x5 TAP_772 ();
 b15ztpn00an1n08x5 TAP_771 ();
 b15ztpn00an1n08x5 TAP_770 ();
 b15ztpn00an1n08x5 TAP_769 ();
 b15ztpn00an1n08x5 TAP_768 ();
 b15ztpn00an1n08x5 TAP_767 ();
 b15ztpn00an1n08x5 TAP_766 ();
 b15ztpn00an1n08x5 TAP_765 ();
 b15ztpn00an1n08x5 TAP_764 ();
 b15qgbna2an1n10x5 _28202_ (.a(net694),
    .b(net714),
    .o1(_02273_));
 b15nand04aq1n12x5 _28203_ (.a(net691),
    .b(net706),
    .c(net702),
    .d(_02273_),
    .o1(_02274_));
 b15nor002ah1n06x5 _28204_ (.a(\us12.a[0] ),
    .b(\us12.a[2] ),
    .o1(_02275_));
 b15inv020ar1n32x5 _28205_ (.a(net693),
    .o1(_02276_));
 b15mdn022ar1n02x5 _28206_ (.a(\us12.a[2] ),
    .b(_02275_),
    .o1(_02277_),
    .sa(_02276_));
 b15ztpn00an1n08x5 TAP_763 ();
 b15nanb02as1n24x5 _28208_ (.a(net701),
    .b(net694),
    .out0(_02279_));
 b15oaoi13an1n02x5 _28209_ (.a(net697),
    .b(_02274_),
    .c(_02277_),
    .d(_02279_),
    .o1(_02280_));
 b15oaoi13ah1n03x5 _28210_ (.a(_02242_),
    .b(net700),
    .c(_02263_),
    .d(_02280_),
    .o1(_02281_));
 b15ztpn00an1n08x5 TAP_762 ();
 b15ztpn00an1n08x5 TAP_761 ();
 b15ztpn00an1n08x5 TAP_760 ();
 b15ztpn00an1n08x5 TAP_759 ();
 b15nonb03aq1n12x5 _28215_ (.a(\us12.a[2] ),
    .b(net705),
    .c(\us12.a[0] ),
    .out0(_02286_));
 b15ztpn00an1n08x5 TAP_758 ();
 b15ztpn00an1n08x5 TAP_757 ();
 b15ztpn00an1n08x5 TAP_756 ();
 b15nona23aq1n32x5 _28219_ (.a(net700),
    .b(net695),
    .c(net692),
    .d(net697),
    .out0(_02290_));
 b15norp02aq1n48x5 _28220_ (.a(net696),
    .b(net699),
    .o1(_02291_));
 b15ztpn00an1n08x5 TAP_755 ();
 b15nonb02as1n16x5 _28222_ (.a(\us12.a[6] ),
    .b(net693),
    .out0(_02293_));
 b15nand02al1n08x5 _28223_ (.a(_02291_),
    .b(_02293_),
    .o1(_02294_));
 b15nandp2an1n08x5 _28224_ (.a(_02290_),
    .b(_02294_),
    .o1(_02295_));
 b15ztpn00an1n08x5 TAP_754 ();
 b15ztpn00an1n08x5 TAP_753 ();
 b15inv000as1n40x5 _28227_ (.a(\us12.a[0] ),
    .o1(_02298_));
 b15nandp3ar1n02x5 _28228_ (.a(net697),
    .b(net692),
    .c(_02298_),
    .o1(_02299_));
 b15nanb02ah1n24x5 _28229_ (.a(\us12.a[2] ),
    .b(\us12.a[0] ),
    .out0(_02300_));
 b15oai013aq1n02x5 _28230_ (.a(_02299_),
    .b(_02300_),
    .c(net692),
    .d(net697),
    .o1(_02301_));
 b15ztpn00an1n08x5 TAP_752 ();
 b15ztpn00an1n08x5 TAP_751 ();
 b15nanb02aq1n04x5 _28233_ (.a(net700),
    .b(net695),
    .out0(_02304_));
 b15nor002al1n02x5 _28234_ (.a(net705),
    .b(_02304_),
    .o1(_02305_));
 b15aoi022an1n06x5 _28235_ (.a(_02286_),
    .b(_02295_),
    .c(_02301_),
    .d(_02305_),
    .o1(_02306_));
 b15ztpn00an1n08x5 TAP_750 ();
 b15ztpn00an1n08x5 TAP_749 ();
 b15nandp2as1n32x5 _28238_ (.a(net692),
    .b(net695),
    .o1(_02309_));
 b15nanb02as1n24x5 _28239_ (.a(net700),
    .b(net697),
    .out0(_02310_));
 b15norp03ar1n16x5 _28240_ (.a(net705),
    .b(_02309_),
    .c(_02310_),
    .o1(_02311_));
 b15ztpn00an1n08x5 TAP_748 ();
 b15nano23ah1n24x5 _28242_ (.a(net697),
    .b(net700),
    .c(net692),
    .d(net695),
    .out0(_02313_));
 b15ztpn00an1n08x5 TAP_747 ();
 b15aoai13an1n04x5 _28244_ (.a(\us12.a[2] ),
    .b(_02311_),
    .c(_02313_),
    .d(net705),
    .o1(_02315_));
 b15aoi013ah1n06x5 _28245_ (.a(_02281_),
    .b(_02306_),
    .c(_02315_),
    .d(_02242_),
    .o1(_02316_));
 b15nanb02as1n24x5 _28246_ (.a(\us12.a[6] ),
    .b(net692),
    .out0(_02317_));
 b15orn002ar1n24x5 _28247_ (.a(net698),
    .b(\us12.a[4] ),
    .o(_02318_));
 b15norp02aq1n32x5 _28248_ (.a(_02317_),
    .b(_02318_),
    .o1(_02319_));
 b15nanb02as1n24x5 _28249_ (.a(net705),
    .b(net709),
    .out0(_02320_));
 b15nonb02as1n16x5 _28250_ (.a(net712),
    .b(net714),
    .out0(_02321_));
 b15ztpn00an1n08x5 TAP_746 ();
 b15norp02al1n02x5 _28252_ (.a(_02320_),
    .b(_02321_),
    .o1(_02323_));
 b15orn002as1n12x5 _28253_ (.a(net708),
    .b(net704),
    .o(_02324_));
 b15orn002an1n32x5 _28254_ (.a(net715),
    .b(\us12.a[1] ),
    .o(_02325_));
 b15nor002al1n16x5 _28255_ (.a(_02324_),
    .b(_02325_),
    .o1(_02326_));
 b15nanb02ah1n24x5 _28256_ (.a(net693),
    .b(\us12.a[6] ),
    .out0(_02327_));
 b15qbfno2bn1n16x5 _28257_ (.a(_02318_),
    .b(_02327_),
    .o1(_02328_));
 b15ao0022an1n04x5 _28258_ (.a(_02319_),
    .b(_02323_),
    .c(_02326_),
    .d(_02328_),
    .o(_02329_));
 b15ztpn00an1n08x5 TAP_745 ();
 b15xor002ar1n02x5 _28260_ (.a(net695),
    .b(net708),
    .out0(_02331_));
 b15nand02ar1n02x5 _28261_ (.a(net692),
    .b(net715),
    .o1(_02332_));
 b15nonb02as1n16x5 _28262_ (.a(net699),
    .b(net696),
    .out0(_02333_));
 b15ztpn00an1n08x5 TAP_744 ();
 b15ztpn00an1n08x5 TAP_743 ();
 b15ztpn00an1n08x5 TAP_742 ();
 b15norp02as1n04x5 _28266_ (.a(net711),
    .b(net704),
    .o1(_02337_));
 b15nona23ah1n02x5 _28267_ (.a(_02331_),
    .b(_02332_),
    .c(_02333_),
    .d(_02337_),
    .out0(_02338_));
 b15ztpn00an1n08x5 TAP_741 ();
 b15xnr002as1n12x5 _28269_ (.a(net715),
    .b(net711),
    .out0(_02340_));
 b15norp02as1n48x5 _28270_ (.a(net693),
    .b(\us12.a[6] ),
    .o1(_02341_));
 b15ztpn00an1n08x5 TAP_740 ();
 b15nonb02as1n16x5 _28272_ (.a(net707),
    .b(net703),
    .out0(_02343_));
 b15ztpn00an1n08x5 TAP_739 ();
 b15ztpn00an1n08x5 TAP_738 ();
 b15nonb02as1n16x5 _28275_ (.a(net698),
    .b(\us12.a[4] ),
    .out0(_02346_));
 b15ztpn00an1n08x5 TAP_737 ();
 b15oai112ar1n04x5 _28277_ (.a(_02341_),
    .b(_02343_),
    .c(_02346_),
    .d(_02333_),
    .o1(_02348_));
 b15oai012aq1n04x5 _28278_ (.a(_02338_),
    .b(_02340_),
    .c(_02348_),
    .o1(_02349_));
 b15nonb02as1n16x5 _28279_ (.a(net711),
    .b(net707),
    .out0(_02350_));
 b15nor004as1n12x5 _28280_ (.a(net696),
    .b(net699),
    .c(net691),
    .d(net694),
    .o1(_02351_));
 b15ztpn00an1n08x5 TAP_736 ();
 b15nand02al1n08x5 _28282_ (.a(_02350_),
    .b(_02351_),
    .o1(_02353_));
 b15nano23as1n24x5 _28283_ (.a(net692),
    .b(net695),
    .c(net697),
    .d(net700),
    .out0(_02354_));
 b15nanb02as1n24x5 _28284_ (.a(net712),
    .b(net714),
    .out0(_02355_));
 b15ztpn00an1n08x5 TAP_735 ();
 b15nanb02as1n24x5 _28286_ (.a(net708),
    .b(net704),
    .out0(_02357_));
 b15norp02as1n03x5 _28287_ (.a(_02355_),
    .b(_02357_),
    .o1(_02358_));
 b15aob012an1n04x5 _28288_ (.a(_02353_),
    .b(_02354_),
    .c(_02358_),
    .out0(_02359_));
 b15ztpn00an1n08x5 TAP_734 ();
 b15nonb03al1n12x5 _28290_ (.a(net708),
    .b(net704),
    .c(net711),
    .out0(_02361_));
 b15nano23ar1n02x5 _28291_ (.a(net700),
    .b(net695),
    .c(net708),
    .d(net692),
    .out0(_02362_));
 b15xor002ar1n02x5 _28292_ (.a(net697),
    .b(net704),
    .out0(_02363_));
 b15aoi022al1n02x5 _28293_ (.a(_02351_),
    .b(_02361_),
    .c(_02362_),
    .d(_02363_),
    .o1(_02364_));
 b15and002aq1n24x5 _28294_ (.a(net691),
    .b(net694),
    .o(_02365_));
 b15nandp2as1n24x5 _28295_ (.a(_02365_),
    .b(_02333_),
    .o1(_02366_));
 b15and002ar1n32x5 _28296_ (.a(net708),
    .b(net704),
    .o(_02367_));
 b15nandp2al1n08x5 _28297_ (.a(_02242_),
    .b(_02367_),
    .o1(_02368_));
 b15oaoi13aq1n03x5 _28298_ (.a(_02298_),
    .b(_02364_),
    .c(_02366_),
    .d(_02368_),
    .o1(_02369_));
 b15nor004ar1n04x5 _28299_ (.a(_02329_),
    .b(_02349_),
    .c(_02359_),
    .d(_02369_),
    .o1(_02370_));
 b15ztpn00an1n08x5 TAP_733 ();
 b15ztpn00an1n08x5 TAP_732 ();
 b15ztpn00an1n08x5 TAP_731 ();
 b15orn003ar1n12x5 _28303_ (.a(net715),
    .b(net711),
    .c(net704),
    .o(_02374_));
 b15norp03as1n24x5 _28304_ (.a(net691),
    .b(net694),
    .c(net707),
    .o1(_02375_));
 b15andc04aq1n16x5 _28305_ (.a(net696),
    .b(net699),
    .c(net691),
    .d(net694),
    .o(_02376_));
 b15ztpn00an1n08x5 TAP_730 ();
 b15aoi022ar1n04x5 _28307_ (.a(_02291_),
    .b(_02375_),
    .c(_02376_),
    .d(net707),
    .o1(_02378_));
 b15aoi012ar1n02x5 _28308_ (.a(_02354_),
    .b(_02351_),
    .c(net713),
    .o1(_02379_));
 b15oa0022al1n03x5 _28309_ (.a(_02374_),
    .b(_02378_),
    .c(_02379_),
    .d(_02368_),
    .o(_02380_));
 b15inv020an1n80x5 _28310_ (.a(net704),
    .o1(_02381_));
 b15ztpn00an1n08x5 TAP_729 ();
 b15ztpn00an1n08x5 TAP_728 ();
 b15ztpn00an1n08x5 TAP_727 ();
 b15nanb02al1n12x5 _28314_ (.a(net705),
    .b(net699),
    .out0(_02385_));
 b15ztpn00an1n08x5 TAP_726 ();
 b15oai022ah1n08x5 _28316_ (.a(_02381_),
    .b(_02310_),
    .c(_02385_),
    .d(net696),
    .o1(_02387_));
 b15norp03as1n04x5 _28317_ (.a(\us12.a[2] ),
    .b(_02327_),
    .c(_02321_),
    .o1(_02388_));
 b15nandp2aq1n32x5 _28318_ (.a(net708),
    .b(net704),
    .o1(_02389_));
 b15nandp2ah1n32x5 _28319_ (.a(\us12.a[0] ),
    .b(\us12.a[1] ),
    .o1(_02390_));
 b15ztpn00an1n08x5 TAP_725 ();
 b15norp02aq1n08x5 _28321_ (.a(_02389_),
    .b(_02390_),
    .o1(_02392_));
 b15aoi222as1n12x5 _28322_ (.a(_02319_),
    .b(_02326_),
    .c(_02387_),
    .d(_02388_),
    .e(_02392_),
    .f(_02313_),
    .o1(_02393_));
 b15nano23ar1n02x5 _28323_ (.a(net692),
    .b(net711),
    .c(net715),
    .d(net697),
    .out0(_02394_));
 b15and002as1n16x5 _28324_ (.a(net714),
    .b(net712),
    .o(_02395_));
 b15ztpn00an1n08x5 TAP_724 ();
 b15aoi013ar1n02x5 _28326_ (.a(_02394_),
    .b(_02395_),
    .c(net695),
    .d(net697),
    .o1(_02397_));
 b15norp03al1n02x5 _28327_ (.a(net700),
    .b(_02324_),
    .c(_02397_),
    .o1(_02398_));
 b15nano22al1n02x5 _28328_ (.a(_02380_),
    .b(_02393_),
    .c(_02398_),
    .out0(_02400_));
 b15ztpn00an1n08x5 TAP_723 ();
 b15nanb02aq1n04x5 _28330_ (.a(net713),
    .b(net699),
    .out0(_02402_));
 b15nano22ar1n12x5 _28331_ (.a(net696),
    .b(net694),
    .c(net691),
    .out0(_02403_));
 b15aoai13al1n06x5 _28332_ (.a(net706),
    .b(net702),
    .c(_02402_),
    .d(_02403_),
    .o1(_02404_));
 b15ztpn00an1n08x5 TAP_722 ();
 b15aoi013ar1n03x5 _28334_ (.a(_02381_),
    .b(_02341_),
    .c(_02346_),
    .d(net710),
    .o1(_02406_));
 b15qbfna2bn1n16x5 _28335_ (.a(_02365_),
    .b(_02346_),
    .o1(_02407_));
 b15oaoi13as1n08x5 _28336_ (.a(_02404_),
    .b(_02406_),
    .c(_02407_),
    .d(_02298_),
    .o1(_02408_));
 b15ztpn00an1n08x5 TAP_721 ();
 b15nonb02as1n16x5 _28338_ (.a(net706),
    .b(net713),
    .out0(_02411_));
 b15nonb02al1n12x5 _28339_ (.a(net714),
    .b(net706),
    .out0(_02412_));
 b15oai112ah1n06x5 _28340_ (.a(net712),
    .b(_02365_),
    .c(_02411_),
    .d(_02412_),
    .o1(_02413_));
 b15ztpn00an1n08x5 TAP_720 ();
 b15nor002ah1n24x5 _28342_ (.a(net712),
    .b(net706),
    .o1(_02415_));
 b15nand03as1n02x5 _28343_ (.a(net714),
    .b(_02341_),
    .c(_02415_),
    .o1(_02416_));
 b15aoi012ar1n06x5 _28344_ (.a(_02318_),
    .b(_02413_),
    .c(_02416_),
    .o1(_02417_));
 b15nanb02ah1n08x5 _28345_ (.a(net709),
    .b(net699),
    .out0(_02418_));
 b15inv040as1n03x5 _28346_ (.a(net698),
    .o1(_02419_));
 b15nandp3ah1n02x5 _28347_ (.a(_02419_),
    .b(_02341_),
    .c(_02395_),
    .o1(_02420_));
 b15aoi012ar1n06x5 _28348_ (.a(_02418_),
    .b(_02420_),
    .c(_02257_),
    .o1(_02422_));
 b15oaoi13as1n08x5 _28349_ (.a(_02408_),
    .b(net705),
    .c(_02417_),
    .d(_02422_),
    .o1(_02423_));
 b15ztpn00an1n08x5 TAP_719 ();
 b15nano23as1n24x5 _28351_ (.a(net697),
    .b(net692),
    .c(net695),
    .d(net700),
    .out0(_02425_));
 b15nonb02as1n12x5 _28352_ (.a(net706),
    .b(net710),
    .out0(_02426_));
 b15nanb02as1n24x5 _28353_ (.a(net708),
    .b(net711),
    .out0(_02427_));
 b15ztpn00an1n08x5 TAP_718 ();
 b15aoai13ar1n03x5 _28355_ (.a(_02425_),
    .b(_02426_),
    .c(_02427_),
    .d(net713),
    .o1(_02429_));
 b15nonb02as1n16x5 _28356_ (.a(net691),
    .b(net694),
    .out0(_02430_));
 b15nandp3al1n08x5 _28357_ (.a(net707),
    .b(_02430_),
    .c(_02291_),
    .o1(_02431_));
 b15norp02ah1n48x5 _28358_ (.a(\us12.a[0] ),
    .b(\us12.a[1] ),
    .o1(_02433_));
 b15ztpn00an1n08x5 TAP_717 ();
 b15oaoi13aq1n08x5 _28360_ (.a(_02381_),
    .b(_02429_),
    .c(_02431_),
    .d(_02433_),
    .o1(_02435_));
 b15nand03al1n03x5 _28361_ (.a(net711),
    .b(_02343_),
    .c(_02351_),
    .o1(_02436_));
 b15and002as1n32x5 _28362_ (.a(net698),
    .b(\us12.a[4] ),
    .o(_02437_));
 b15nandp2ar1n24x5 _28363_ (.a(_02430_),
    .b(_02437_),
    .o1(_02438_));
 b15ztpn00an1n08x5 TAP_716 ();
 b15oai013al1n06x5 _28365_ (.a(_02436_),
    .b(_02438_),
    .c(_02389_),
    .d(_02325_),
    .o1(_02440_));
 b15nano22al1n05x5 _28366_ (.a(net694),
    .b(net702),
    .c(net691),
    .out0(_02441_));
 b15ztpn00an1n08x5 TAP_715 ();
 b15orn002as1n12x5 _28368_ (.a(net710),
    .b(net706),
    .o(_02444_));
 b15aoai13aq1n08x5 _28369_ (.a(_02441_),
    .b(_02291_),
    .c(_02437_),
    .d(_02444_),
    .o1(_02445_));
 b15nand03an1n04x5 _28370_ (.a(net713),
    .b(net710),
    .c(net706),
    .o1(_02446_));
 b15nanb02an1n04x5 _28371_ (.a(net710),
    .b(net696),
    .out0(_02447_));
 b15aoai13ah1n08x5 _28372_ (.a(_02446_),
    .b(net713),
    .c(net706),
    .d(_02447_),
    .o1(_02448_));
 b15nonb02as1n16x5 _28373_ (.a(net714),
    .b(net712),
    .out0(_02449_));
 b15xor002ar1n16x5 _28374_ (.a(net694),
    .b(_02449_),
    .out0(_02450_));
 b15nandp3an1n08x5 _28375_ (.a(net691),
    .b(_02251_),
    .c(_02437_),
    .o1(_02451_));
 b15oai022al1n24x5 _28376_ (.a(_02445_),
    .b(_02448_),
    .c(_02450_),
    .d(_02451_),
    .o1(_02452_));
 b15norp03as1n04x5 _28377_ (.a(_02435_),
    .b(_02440_),
    .c(_02452_),
    .o1(_02453_));
 b15nand04aq1n08x5 _28378_ (.a(_02370_),
    .b(_02400_),
    .c(_02423_),
    .d(_02453_),
    .o1(_02455_));
 b15ztpn00an1n08x5 TAP_714 ();
 b15nanb02aq1n12x5 _28380_ (.a(net712),
    .b(net705),
    .out0(_02457_));
 b15nandp2ah1n03x5 _28381_ (.a(net709),
    .b(_02346_),
    .o1(_02458_));
 b15aoi112ah1n08x5 _28382_ (.a(_02259_),
    .b(_02457_),
    .c(_02458_),
    .d(_02418_),
    .o1(_02459_));
 b15nanb02ah1n12x5 _28383_ (.a(net704),
    .b(net711),
    .out0(_02460_));
 b15inv000ah1n40x5 _28384_ (.a(net708),
    .o1(_02461_));
 b15nano23aq1n24x5 _28385_ (.a(net699),
    .b(net691),
    .c(net694),
    .d(net696),
    .out0(_02462_));
 b15nand02as1n12x5 _28386_ (.a(_02461_),
    .b(_02462_),
    .o1(_02463_));
 b15ztpn00an1n08x5 TAP_713 ();
 b15nona23as1n32x5 _28388_ (.a(net692),
    .b(net695),
    .c(net697),
    .d(net700),
    .out0(_02466_));
 b15oaoi13ar1n02x5 _28389_ (.a(_02460_),
    .b(_02463_),
    .c(_02461_),
    .d(_02466_),
    .o1(_02467_));
 b15nandp3al1n16x5 _28390_ (.a(net711),
    .b(net708),
    .c(net704),
    .o1(_02468_));
 b15nona23as1n32x5 _28391_ (.a(net700),
    .b(net692),
    .c(net695),
    .d(net697),
    .out0(_02469_));
 b15ztpn00an1n08x5 TAP_712 ();
 b15nand04as1n16x5 _28393_ (.a(net698),
    .b(net700),
    .c(net693),
    .d(net695),
    .o1(_02471_));
 b15aoi012ar1n02x5 _28394_ (.a(_02468_),
    .b(_02469_),
    .c(_02471_),
    .o1(_02472_));
 b15nor004an1n03x5 _28395_ (.a(net715),
    .b(_02459_),
    .c(_02467_),
    .d(_02472_),
    .o1(_02473_));
 b15ztpn00an1n08x5 TAP_711 ();
 b15nano23as1n24x5 _28397_ (.a(net699),
    .b(net694),
    .c(net691),
    .d(net696),
    .out0(_02475_));
 b15nanb02al1n02x5 _28398_ (.a(_02468_),
    .b(_02475_),
    .out0(_02477_));
 b15norp03aq1n04x5 _28399_ (.a(net703),
    .b(_02444_),
    .c(_02469_),
    .o1(_02478_));
 b15nano22ar1n03x5 _28400_ (.a(net713),
    .b(_02477_),
    .c(_02478_),
    .out0(_02479_));
 b15nor002ah1n04x5 _28401_ (.a(_02473_),
    .b(_02479_),
    .o1(_02480_));
 b15and003ar1n02x5 _28402_ (.a(net692),
    .b(net695),
    .c(net705),
    .o(_02481_));
 b15oaoi13ar1n02x5 _28403_ (.a(_02481_),
    .b(_02341_),
    .c(_02381_),
    .d(_02325_),
    .o1(_02482_));
 b15aobi12ar1n02x5 _28404_ (.a(\us12.a[0] ),
    .b(\us12.a[1] ),
    .c(net705),
    .out0(_02483_));
 b15oai013ar1n03x5 _28405_ (.a(_02483_),
    .b(_02310_),
    .c(_02259_),
    .d(net712),
    .o1(_02484_));
 b15nona23al1n04x5 _28406_ (.a(\us12.a[2] ),
    .b(_02482_),
    .c(_02346_),
    .d(_02484_),
    .out0(_02485_));
 b15ztpn00an1n08x5 TAP_710 ();
 b15nandp3ah1n03x5 _28408_ (.a(_02321_),
    .b(_02351_),
    .c(_02367_),
    .o1(_02488_));
 b15and002aq1n04x5 _28409_ (.a(_02485_),
    .b(_02488_),
    .o(_02489_));
 b15norp03al1n02x5 _28410_ (.a(net704),
    .b(_02466_),
    .c(_02433_),
    .o1(_02490_));
 b15nonb02al1n12x5 _28411_ (.a(net692),
    .b(net697),
    .out0(_02491_));
 b15qgbna2an1n05x5 _28412_ (.o1(_02492_),
    .a(\us12.a[4] ),
    .b(\us12.a[6] ));
 b15orn002ah1n03x5 _28413_ (.a(net700),
    .b(\us12.a[6] ),
    .o(_02493_));
 b15oai012ar1n16x5 _28414_ (.a(_02492_),
    .b(_02493_),
    .c(_02298_),
    .o1(_02494_));
 b15ztpn00an1n08x5 TAP_709 ();
 b15aoi013al1n03x5 _28416_ (.a(_02490_),
    .b(_02491_),
    .c(_02494_),
    .d(net704),
    .o1(_02496_));
 b15ztpn00an1n08x5 TAP_708 ();
 b15nand03al1n16x5 _28418_ (.a(net709),
    .b(_02430_),
    .c(_02437_),
    .o1(_02499_));
 b15nandp2aq1n24x5 _28419_ (.a(_02293_),
    .b(_02437_),
    .o1(_02500_));
 b15oaoi13al1n02x5 _28420_ (.a(net711),
    .b(_02499_),
    .c(_02500_),
    .d(net707),
    .o1(_02501_));
 b15oab012aq1n04x5 _28421_ (.a(_02501_),
    .b(_02499_),
    .c(_02298_),
    .out0(_02502_));
 b15ztpn00an1n08x5 TAP_707 ();
 b15oai122ah1n08x5 _28423_ (.a(_02489_),
    .b(_02496_),
    .c(net708),
    .d(_02502_),
    .e(net704),
    .o1(_02504_));
 b15nor004an1n08x5 _28424_ (.a(_02316_),
    .b(_02455_),
    .c(_02480_),
    .d(_02504_),
    .o1(_02505_));
 b15ztpn00an1n08x5 TAP_706 ();
 b15nanb02as1n24x5 _28426_ (.a(net831),
    .b(net833),
    .out0(_02507_));
 b15ztpn00an1n08x5 TAP_705 ();
 b15ztpn00an1n08x5 TAP_704 ();
 b15ztpn00an1n08x5 TAP_703 ();
 b15ztpn00an1n08x5 TAP_702 ();
 b15ztpn00an1n08x5 TAP_701 ();
 b15ztpn00an1n08x5 TAP_700 ();
 b15nona23as1n32x5 _28433_ (.a(\us01.a[4] ),
    .b(net823),
    .c(\us01.a[6] ),
    .d(net827),
    .out0(_02515_));
 b15ztpn00an1n08x5 TAP_699 ();
 b15nonb02as1n16x5 _28435_ (.a(\us01.a[4] ),
    .b(net827),
    .out0(_02517_));
 b15ztpn00an1n08x5 TAP_698 ();
 b15ztpn00an1n08x5 TAP_697 ();
 b15ztpn00an1n08x5 TAP_696 ();
 b15ztpn00an1n08x5 TAP_695 ();
 b15ztpn00an1n08x5 TAP_694 ();
 b15nand02ar1n02x5 _28441_ (.a(net825),
    .b(net837),
    .o1(_02524_));
 b15ztpn00an1n08x5 TAP_693 ();
 b15nanb02an1n24x5 _28443_ (.a(net837),
    .b(net840),
    .out0(_02526_));
 b15oaoi13ar1n02x5 _28444_ (.a(net822),
    .b(_02524_),
    .c(_02526_),
    .d(net825),
    .o1(_02527_));
 b15ztpn00an1n08x5 TAP_692 ();
 b15and002ar1n24x5 _28446_ (.a(net823),
    .b(\us01.a[6] ),
    .o(_02529_));
 b15ztpn00an1n08x5 TAP_691 ();
 b15nonb02aq1n12x5 _28448_ (.a(net840),
    .b(net837),
    .out0(_02532_));
 b15aoai13an1n02x5 _28449_ (.a(_02517_),
    .b(_02527_),
    .c(_02529_),
    .d(_02532_),
    .o1(_02533_));
 b15aoi012ar1n04x5 _28450_ (.a(_02507_),
    .b(_02515_),
    .c(_02533_),
    .o1(_02534_));
 b15ztpn00an1n08x5 TAP_690 ();
 b15ztpn00an1n08x5 TAP_689 ();
 b15ztpn00an1n08x5 TAP_688 ();
 b15ztpn00an1n08x5 TAP_687 ();
 b15ztpn00an1n08x5 TAP_686 ();
 b15ztpn00an1n08x5 TAP_685 ();
 b15nor002an1n24x5 _28457_ (.a(net838),
    .b(net835),
    .o1(_02541_));
 b15nand02as1n03x5 _28458_ (.a(net842),
    .b(_02541_),
    .o1(_02543_));
 b15ztpn00an1n08x5 TAP_684 ();
 b15nanb02al1n16x5 _28460_ (.a(net842),
    .b(net835),
    .out0(_02545_));
 b15nanb02as1n24x5 _28461_ (.a(net828),
    .b(net826),
    .out0(_02546_));
 b15nandp2as1n48x5 _28462_ (.a(\us01.a[7] ),
    .b(net824),
    .o1(_02547_));
 b15nor002ar1n32x5 _28463_ (.a(_02546_),
    .b(_02547_),
    .o1(_02548_));
 b15ztpn00an1n08x5 TAP_683 ();
 b15nand04an1n16x5 _28465_ (.a(net832),
    .b(_02543_),
    .c(_02545_),
    .d(_02548_),
    .o1(_02550_));
 b15ztpn00an1n08x5 TAP_682 ();
 b15ztpn00an1n08x5 TAP_681 ();
 b15nandp3an1n24x5 _28468_ (.a(net839),
    .b(\us01.a[2] ),
    .c(\us01.a[3] ),
    .o1(_02554_));
 b15norp03aq1n02x5 _28469_ (.a(net840),
    .b(_02515_),
    .c(_02554_),
    .o1(_02555_));
 b15ztpn00an1n08x5 TAP_680 ();
 b15nanb02as1n24x5 _28471_ (.a(\us01.a[5] ),
    .b(net829),
    .out0(_02557_));
 b15ztpn00an1n08x5 TAP_679 ();
 b15mdn022an1n04x5 _28473_ (.a(_02546_),
    .b(_02557_),
    .o1(_02559_),
    .sa(net831));
 b15ztpn00an1n08x5 TAP_678 ();
 b15ztpn00an1n08x5 TAP_677 ();
 b15nonb02aq1n12x5 _28476_ (.a(net839),
    .b(net840),
    .out0(_02562_));
 b15norp02aq1n03x5 _28477_ (.a(net834),
    .b(_02562_),
    .o1(_02563_));
 b15ztpn00an1n08x5 TAP_676 ();
 b15nonb02aq1n16x5 _28479_ (.a(\us01.a[6] ),
    .b(net823),
    .out0(_02566_));
 b15aoi013ah1n03x5 _28480_ (.a(_02555_),
    .b(_02559_),
    .c(_02563_),
    .d(_02566_),
    .o1(_02567_));
 b15ztpn00an1n08x5 TAP_675 ();
 b15inv000as1n40x5 _28482_ (.a(net835),
    .o1(_02569_));
 b15ztpn00an1n08x5 TAP_674 ();
 b15ztpn00an1n08x5 TAP_673 ();
 b15ztpn00an1n08x5 TAP_672 ();
 b15inv040as1n40x5 _28486_ (.a(net838),
    .o1(_02573_));
 b15ztpn00an1n08x5 TAP_671 ();
 b15nand02ar1n02x5 _28488_ (.a(net827),
    .b(_02573_),
    .o1(_02576_));
 b15norp02as1n08x5 _28489_ (.a(net828),
    .b(net831),
    .o1(_02577_));
 b15ztpn00an1n08x5 TAP_670 ();
 b15and002aq1n12x5 _28491_ (.a(net828),
    .b(net831),
    .o(_02579_));
 b15norp02aq1n16x5 _28492_ (.a(net823),
    .b(\us01.a[6] ),
    .o1(_02580_));
 b15aoi022ar1n02x5 _28493_ (.a(_02529_),
    .b(_02577_),
    .c(_02579_),
    .d(_02580_),
    .o1(_02581_));
 b15ztpn00an1n08x5 TAP_669 ();
 b15nona23as1n32x5 _28495_ (.a(net822),
    .b(net825),
    .c(net826),
    .d(net828),
    .out0(_02583_));
 b15ztpn00an1n08x5 TAP_668 ();
 b15nand02as1n16x5 _28497_ (.a(net840),
    .b(\us01.a[3] ),
    .o1(_02585_));
 b15oa0022aq1n03x5 _28498_ (.a(_02576_),
    .b(_02581_),
    .c(_02583_),
    .d(_02585_),
    .o(_02587_));
 b15oai112al1n16x5 _28499_ (.a(_02550_),
    .b(_02567_),
    .c(_02569_),
    .d(_02587_),
    .o1(_02588_));
 b15ztpn00an1n08x5 TAP_667 ();
 b15ztpn00an1n08x5 TAP_666 ();
 b15ztpn00an1n08x5 TAP_665 ();
 b15ztpn00an1n08x5 TAP_664 ();
 b15nona23as1n32x5 _28504_ (.a(\us01.a[4] ),
    .b(\us01.a[6] ),
    .c(net823),
    .d(net827),
    .out0(_02593_));
 b15nand02ar1n02x5 _28505_ (.a(net831),
    .b(_02593_),
    .o1(_02594_));
 b15nandp2aq1n48x5 _28506_ (.a(\us01.a[5] ),
    .b(net829),
    .o1(_02595_));
 b15nanb02as1n24x5 _28507_ (.a(net824),
    .b(\us01.a[7] ),
    .out0(_02596_));
 b15norp02as1n24x5 _28508_ (.a(_02595_),
    .b(_02596_),
    .o1(_02598_));
 b15ztpn00an1n08x5 TAP_663 ();
 b15oai012al1n02x5 _28510_ (.a(_02594_),
    .b(_02598_),
    .c(net831),
    .o1(_02600_));
 b15ztpn00an1n08x5 TAP_662 ();
 b15nandp2as1n32x5 _28512_ (.a(net837),
    .b(\us01.a[2] ),
    .o1(_02602_));
 b15ztpn00an1n08x5 TAP_661 ();
 b15nanb02ah1n24x5 _28514_ (.a(net834),
    .b(net832),
    .out0(_02604_));
 b15aoi012ar1n02x5 _28515_ (.a(net840),
    .b(_02602_),
    .c(_02604_),
    .o1(_02605_));
 b15ztpn00an1n08x5 TAP_660 ();
 b15ztpn00an1n08x5 TAP_659 ();
 b15nand02ar1n24x5 _28518_ (.a(net837),
    .b(net831),
    .o1(_02609_));
 b15orn002al1n12x5 _28519_ (.a(net836),
    .b(net830),
    .o(_02610_));
 b15inv020an1n80x5 _28520_ (.a(net842),
    .o1(_02611_));
 b15ztpn00an1n08x5 TAP_658 ();
 b15oaoi13an1n03x5 _28522_ (.a(net833),
    .b(_02609_),
    .c(_02610_),
    .d(_02611_),
    .o1(_02613_));
 b15qgbno3an1n05x5 _28523_ (.o1(_02614_),
    .a(_02600_),
    .b(_02605_),
    .c(_02613_));
 b15inv020an1n16x5 _28524_ (.a(net826),
    .o1(_02615_));
 b15nanb02as1n24x5 _28525_ (.a(net840),
    .b(net837),
    .out0(_02616_));
 b15ztpn00an1n08x5 TAP_657 ();
 b15nor002aq1n08x5 _28527_ (.a(net824),
    .b(net833),
    .o1(_02618_));
 b15norp02al1n24x5 _28528_ (.a(net828),
    .b(net822),
    .o1(_02620_));
 b15ztpn00an1n08x5 TAP_656 ();
 b15nand03ah1n06x5 _28530_ (.a(net822),
    .b(net824),
    .c(net830),
    .o1(_02622_));
 b15orn002aq1n32x5 _28531_ (.a(net822),
    .b(net824),
    .o(_02623_));
 b15ztpn00an1n08x5 TAP_655 ();
 b15oai012al1n02x5 _28533_ (.a(_02622_),
    .b(_02623_),
    .c(net830),
    .o1(_02625_));
 b15ztpn00an1n08x5 TAP_654 ();
 b15aoi022as1n02x5 _28535_ (.a(_02618_),
    .b(_02620_),
    .c(_02625_),
    .d(net828),
    .o1(_02627_));
 b15nor003as1n08x5 _28536_ (.a(_02615_),
    .b(_02616_),
    .c(_02627_),
    .o1(_02628_));
 b15nor004al1n08x5 _28537_ (.a(_02534_),
    .b(_02588_),
    .c(_02614_),
    .d(_02628_),
    .o1(_02629_));
 b15inv040al1n40x5 _28538_ (.a(net832),
    .o1(_02631_));
 b15ztpn00an1n08x5 TAP_653 ();
 b15ztpn00an1n08x5 TAP_652 ();
 b15xor002ah1n16x5 _28541_ (.a(net841),
    .b(net836),
    .out0(_02634_));
 b15nano23as1n24x5 _28542_ (.a(net829),
    .b(\us01.a[7] ),
    .c(net824),
    .d(net827),
    .out0(_02635_));
 b15ztpn00an1n08x5 TAP_651 ();
 b15andc04aq1n12x5 _28544_ (.a(net827),
    .b(\us01.a[4] ),
    .c(\us01.a[7] ),
    .d(\us01.a[6] ),
    .o(_02637_));
 b15ztpn00an1n08x5 TAP_650 ();
 b15aoi022ar1n02x5 _28546_ (.a(_02634_),
    .b(_02635_),
    .c(_02637_),
    .d(net836),
    .o1(_02639_));
 b15nandp2ar1n04x5 _28547_ (.a(_02631_),
    .b(_02639_),
    .o1(_02640_));
 b15nandp2aq1n16x5 _28548_ (.a(_02517_),
    .b(_02529_),
    .o1(_02642_));
 b15orn002as1n32x5 _28549_ (.a(\us01.a[5] ),
    .b(net829),
    .o(_02643_));
 b15ztpn00an1n08x5 TAP_649 ();
 b15orn002an1n08x5 _28551_ (.a(net841),
    .b(net834),
    .o(_02645_));
 b15nandp2ar1n05x5 _28552_ (.a(net825),
    .b(_02645_),
    .o1(_02646_));
 b15oai112aq1n08x5 _28553_ (.a(net830),
    .b(_02642_),
    .c(_02643_),
    .d(_02646_),
    .o1(_02647_));
 b15nand02al1n08x5 _28554_ (.a(net824),
    .b(net830),
    .o1(_02648_));
 b15and002ah1n24x5 _28555_ (.a(net840),
    .b(net839),
    .o(_02649_));
 b15oai013aq1n06x5 _28556_ (.a(net834),
    .b(_02648_),
    .c(_02643_),
    .d(_02649_),
    .o1(_02650_));
 b15nandp3ar1n12x5 _28557_ (.o1(_02651_),
    .a(_02640_),
    .b(_02647_),
    .c(_02650_));
 b15oab012ar1n02x5 _28558_ (.a(net840),
    .b(net837),
    .c(net822),
    .out0(_02653_));
 b15orn002ah1n32x5 _28559_ (.a(net833),
    .b(net831),
    .o(_02654_));
 b15ztpn00an1n08x5 TAP_648 ();
 b15nandp3ah1n16x5 _28561_ (.a(net826),
    .b(net828),
    .c(net824),
    .o1(_02656_));
 b15orn003ar1n02x5 _28562_ (.a(_02653_),
    .b(_02654_),
    .c(_02656_),
    .o(_02657_));
 b15nandp2an1n03x5 _28563_ (.a(net826),
    .b(_02529_),
    .o1(_02658_));
 b15aoi012ar1n02x5 _28564_ (.a(_02579_),
    .b(_02649_),
    .c(_02577_),
    .o1(_02659_));
 b15ztpn00an1n08x5 TAP_647 ();
 b15oai013ar1n02x5 _28566_ (.a(_02657_),
    .b(_02658_),
    .c(_02659_),
    .d(net833),
    .o1(_02661_));
 b15and002ar1n12x5 _28567_ (.a(net826),
    .b(net828),
    .o(_02662_));
 b15and002aq1n12x5 _28568_ (.a(net835),
    .b(net832),
    .o(_02664_));
 b15norp02ar1n48x5 _28569_ (.a(net841),
    .b(net836),
    .o1(_02665_));
 b15nonb02ah1n16x5 _28570_ (.a(net823),
    .b(\us01.a[6] ),
    .out0(_02666_));
 b15nand04al1n12x5 _28571_ (.a(_02662_),
    .b(_02664_),
    .c(_02665_),
    .d(_02666_),
    .o1(_02667_));
 b15norp02an1n24x5 _28572_ (.a(net834),
    .b(net830),
    .o1(_02668_));
 b15nandp2as1n12x5 _28573_ (.a(net836),
    .b(_02668_),
    .o1(_02669_));
 b15nanb02ah1n24x5 _28574_ (.a(net826),
    .b(net822),
    .out0(_02670_));
 b15nanb02an1n12x5 _28575_ (.a(net842),
    .b(net824),
    .out0(_02671_));
 b15oai013an1n04x5 _28576_ (.a(_02667_),
    .b(_02669_),
    .c(_02670_),
    .d(_02671_),
    .o1(_02672_));
 b15ztpn00an1n08x5 TAP_646 ();
 b15ztpn00an1n08x5 TAP_645 ();
 b15nandp2an1n08x5 _28579_ (.a(net840),
    .b(net833),
    .o1(_02676_));
 b15norp03ar1n08x5 _28580_ (.a(net826),
    .b(net822),
    .c(net824),
    .o1(_02677_));
 b15nand02aq1n04x5 _28581_ (.a(_02676_),
    .b(_02677_),
    .o1(_02678_));
 b15nor004ar1n02x5 _28582_ (.a(net828),
    .b(_02573_),
    .c(_02631_),
    .d(_02678_),
    .o1(_02679_));
 b15nanb02as1n24x5 _28583_ (.a(\us01.a[7] ),
    .b(net824),
    .out0(_02680_));
 b15nand03al1n24x5 _28584_ (.a(\us01.a[5] ),
    .b(\us01.a[7] ),
    .c(net834),
    .o1(_02681_));
 b15ztpn00an1n08x5 TAP_644 ();
 b15oai022ar1n02x5 _28586_ (.a(net826),
    .b(_02680_),
    .c(_02681_),
    .d(net825),
    .o1(_02683_));
 b15and002aq1n16x5 _28587_ (.a(net841),
    .b(net834),
    .o(_02684_));
 b15norp03ar1n02x5 _28588_ (.a(net828),
    .b(_02610_),
    .c(_02684_),
    .o1(_02686_));
 b15oaoi13ar1n02x5 _28589_ (.a(_02546_),
    .b(_02623_),
    .c(_02547_),
    .d(net839),
    .o1(_02687_));
 b15norp02ar1n02x5 _28590_ (.a(net840),
    .b(_02654_),
    .o1(_02688_));
 b15ao0022al1n02x5 _28591_ (.a(_02683_),
    .b(_02686_),
    .c(_02687_),
    .d(_02688_),
    .o(_02689_));
 b15nor004an1n03x5 _28592_ (.a(_02661_),
    .b(_02672_),
    .c(_02679_),
    .d(_02689_),
    .o1(_02690_));
 b15ztpn00an1n08x5 TAP_643 ();
 b15ornc04ah1n24x5 _28594_ (.a(net826),
    .b(net828),
    .c(net822),
    .d(net825),
    .o(_02692_));
 b15ztpn00an1n08x5 TAP_642 ();
 b15nonb02as1n06x5 _28596_ (.a(net826),
    .b(net822),
    .out0(_02694_));
 b15nanb02aq1n16x5 _28597_ (.a(net831),
    .b(net837),
    .out0(_02695_));
 b15oai112al1n02x5 _28598_ (.a(_02618_),
    .b(_02694_),
    .c(_02695_),
    .d(net828),
    .o1(_02697_));
 b15oai022ar1n02x5 _28599_ (.a(_02507_),
    .b(_02692_),
    .c(_02697_),
    .d(_02579_),
    .o1(_02698_));
 b15ztpn00an1n08x5 TAP_641 ();
 b15nandp2ar1n32x5 _28601_ (.a(_02517_),
    .b(_02580_),
    .o1(_02700_));
 b15nanb02aq1n24x5 _28602_ (.a(net833),
    .b(net837),
    .out0(_02701_));
 b15oai022ar1n02x5 _28603_ (.a(net837),
    .b(_02692_),
    .c(_02700_),
    .d(_02701_),
    .o1(_02702_));
 b15ztpn00an1n08x5 TAP_640 ();
 b15ztpn00an1n08x5 TAP_639 ();
 b15aoai13al1n02x5 _28606_ (.a(net840),
    .b(_02698_),
    .c(_02702_),
    .d(net831),
    .o1(_02705_));
 b15ztpn00an1n08x5 TAP_638 ();
 b15ztpn00an1n08x5 TAP_637 ();
 b15nonb02as1n16x5 _28609_ (.a(\us01.a[3] ),
    .b(\us01.a[2] ),
    .out0(_02709_));
 b15ztpn00an1n08x5 TAP_636 ();
 b15and003aq1n04x5 _28611_ (.a(net826),
    .b(net825),
    .c(net840),
    .o(_02711_));
 b15norp03ar1n02x5 _28612_ (.a(net826),
    .b(net825),
    .c(net831),
    .o1(_02712_));
 b15aoi022ar1n02x5 _28613_ (.a(_02709_),
    .b(_02711_),
    .c(_02712_),
    .d(_02676_),
    .o1(_02713_));
 b15norp02ar1n02x5 _28614_ (.a(net822),
    .b(_02713_),
    .o1(_02714_));
 b15ztpn00an1n08x5 TAP_635 ();
 b15nand02an1n48x5 _28616_ (.a(\us01.a[2] ),
    .b(\us01.a[3] ),
    .o1(_02716_));
 b15ztpn00an1n08x5 TAP_634 ();
 b15norp03al1n02x5 _28618_ (.a(net825),
    .b(_02716_),
    .c(_02670_),
    .o1(_02719_));
 b15oai112an1n04x5 _28619_ (.a(net828),
    .b(net837),
    .c(_02714_),
    .d(_02719_),
    .o1(_02720_));
 b15andc04ah1n04x5 _28620_ (.a(_02651_),
    .b(_02690_),
    .c(_02705_),
    .d(_02720_),
    .o(_02721_));
 b15ztpn00an1n08x5 TAP_633 ();
 b15nor002as1n08x5 _28622_ (.a(_02546_),
    .b(_02623_),
    .o1(_02723_));
 b15nor002an1n24x5 _28623_ (.a(net836),
    .b(net830),
    .o1(_02724_));
 b15oai012ar1n02x5 _28624_ (.a(_02609_),
    .b(_02724_),
    .c(net840),
    .o1(_02725_));
 b15nand02ar1n02x5 _28625_ (.a(_02723_),
    .b(_02725_),
    .o1(_02726_));
 b15norp02as1n16x5 _28626_ (.a(net827),
    .b(\us01.a[4] ),
    .o1(_02727_));
 b15nandp2as1n12x5 _28627_ (.a(_02666_),
    .b(_02727_),
    .o1(_02728_));
 b15ztpn00an1n08x5 TAP_632 ();
 b15oai013al1n04x5 _28629_ (.a(_02726_),
    .b(_02728_),
    .c(_02631_),
    .d(_02573_),
    .o1(_02731_));
 b15nor003an1n06x5 _28630_ (.a(net831),
    .b(_02546_),
    .c(_02623_),
    .o1(_02732_));
 b15ztpn00an1n08x5 TAP_631 ();
 b15aob012as1n03x5 _28632_ (.a(_02728_),
    .b(_02732_),
    .c(_02573_),
    .out0(_02734_));
 b15ztpn00an1n08x5 TAP_630 ();
 b15aoai13ar1n08x5 _28634_ (.a(net833),
    .b(_02731_),
    .c(_02734_),
    .d(net840),
    .o1(_02736_));
 b15nandp2al1n02x5 _28635_ (.a(net828),
    .b(net825),
    .o1(_02737_));
 b15nanb03aq1n16x5 _28636_ (.a(net822),
    .b(net833),
    .c(net826),
    .out0(_02738_));
 b15aoi122ar1n04x5 _28637_ (.a(_02737_),
    .b(_02670_),
    .c(_02738_),
    .d(_02616_),
    .e(_02526_),
    .o1(_02739_));
 b15ztpn00an1n08x5 TAP_629 ();
 b15nonb02al1n16x5 _28639_ (.a(net833),
    .b(net839),
    .out0(_02742_));
 b15nona23as1n32x5 _28640_ (.a(\us01.a[5] ),
    .b(\us01.a[7] ),
    .c(net824),
    .d(net829),
    .out0(_02743_));
 b15norp03al1n03x5 _28641_ (.a(_02611_),
    .b(_02742_),
    .c(_02743_),
    .o1(_02744_));
 b15orn002aq1n24x5 _28642_ (.a(net840),
    .b(net837),
    .o(_02745_));
 b15norp03ar1n02x5 _28643_ (.a(net833),
    .b(_02583_),
    .c(_02745_),
    .o1(_02746_));
 b15oai013ar1n02x5 _28644_ (.a(net831),
    .b(_02739_),
    .c(_02744_),
    .d(_02746_),
    .o1(_02747_));
 b15nor004as1n12x5 _28645_ (.a(net826),
    .b(net828),
    .c(net822),
    .d(net825),
    .o1(_02748_));
 b15ztpn00an1n08x5 TAP_628 ();
 b15ztpn00an1n08x5 TAP_627 ();
 b15norp03as1n16x5 _28648_ (.a(net841),
    .b(_02596_),
    .c(_02643_),
    .o1(_02752_));
 b15aoi022ar1n02x5 _28649_ (.a(net839),
    .b(_02748_),
    .c(_02752_),
    .d(_02602_),
    .o1(_02753_));
 b15oai012ar1n04x5 _28650_ (.a(_02747_),
    .b(_02753_),
    .c(net831),
    .o1(_02754_));
 b15ztpn00an1n08x5 TAP_626 ();
 b15ztpn00an1n08x5 TAP_625 ();
 b15norp02an1n48x5 _28653_ (.a(_02596_),
    .b(_02643_),
    .o1(_02757_));
 b15nandp3ar1n02x5 _28654_ (.a(_02569_),
    .b(net831),
    .c(_02757_),
    .o1(_02758_));
 b15nano23as1n24x5 _28655_ (.a(net827),
    .b(\us01.a[6] ),
    .c(net823),
    .d(\us01.a[4] ),
    .out0(_02759_));
 b15ztpn00an1n08x5 TAP_624 ();
 b15nor003ar1n12x5 _28657_ (.a(_02569_),
    .b(_02680_),
    .c(_02595_),
    .o1(_02761_));
 b15oai012ar1n02x5 _28658_ (.a(_02631_),
    .b(_02759_),
    .c(_02761_),
    .o1(_02763_));
 b15aoi012al1n02x5 _28659_ (.a(_02611_),
    .b(_02758_),
    .c(_02763_),
    .o1(_02764_));
 b15norp02ar1n02x5 _28660_ (.a(net826),
    .b(net825),
    .o1(_02765_));
 b15nor002aq1n03x5 _28661_ (.a(net822),
    .b(net833),
    .o1(_02766_));
 b15oai112al1n06x5 _28662_ (.a(_02765_),
    .b(_02766_),
    .c(_02577_),
    .d(_02579_),
    .o1(_02767_));
 b15nand04as1n16x5 _28663_ (.a(net827),
    .b(\us01.a[4] ),
    .c(net823),
    .d(\us01.a[6] ),
    .o1(_02768_));
 b15oaoi13al1n02x5 _28664_ (.a(_02745_),
    .b(_02767_),
    .c(_02768_),
    .d(_02507_),
    .o1(_02769_));
 b15norp03as1n04x5 _28665_ (.a(_02754_),
    .b(_02764_),
    .c(_02769_),
    .o1(_02770_));
 b15nand04as1n16x5 _28666_ (.a(_02629_),
    .b(_02721_),
    .c(_02736_),
    .d(_02770_),
    .o1(_02771_));
 b15xnr002as1n16x5 _28667_ (.a(net401),
    .b(_02771_),
    .out0(_02772_));
 b15ztpn00an1n08x5 TAP_623 ();
 b15ztpn00an1n08x5 TAP_622 ();
 b15ztpn00an1n08x5 TAP_621 ();
 b15ztpn00an1n08x5 TAP_620 ();
 b15ztpn00an1n08x5 TAP_619 ();
 b15norp02aq1n48x5 _28673_ (.a(net846),
    .b(net849),
    .o1(_02779_));
 b15ztpn00an1n08x5 TAP_618 ();
 b15nonb02as1n16x5 _28675_ (.a(net843),
    .b(\us30.a[6] ),
    .out0(_02781_));
 b15and002aq1n16x5 _28676_ (.a(_02779_),
    .b(_02781_),
    .o(_02782_));
 b15ztpn00an1n08x5 TAP_617 ();
 b15ztpn00an1n08x5 TAP_616 ();
 b15ztpn00an1n08x5 TAP_615 ();
 b15orn002ar1n24x5 _28680_ (.a(net851),
    .b(net853),
    .o(_02787_));
 b15qgbno2an1n10x5 _28681_ (.a(net860),
    .b(_02787_),
    .o1(_02788_));
 b15ztpn00an1n08x5 TAP_614 ();
 b15ztpn00an1n08x5 TAP_613 ();
 b15nonb02as1n16x5 _28684_ (.a(net856),
    .b(net852),
    .out0(_02791_));
 b15ztpn00an1n08x5 TAP_612 ();
 b15ztpn00an1n08x5 TAP_611 ();
 b15nanb02ah1n16x5 _28687_ (.a(net843),
    .b(\us30.a[6] ),
    .out0(_02794_));
 b15ztpn00an1n08x5 TAP_610 ();
 b15ztpn00an1n08x5 TAP_609 ();
 b15nandp2al1n16x5 _28690_ (.a(net846),
    .b(net849),
    .o1(_02798_));
 b15nor002as1n06x5 _28691_ (.a(_02794_),
    .b(_02798_),
    .o1(_02799_));
 b15ztpn00an1n08x5 TAP_608 ();
 b15ztpn00an1n08x5 TAP_607 ();
 b15ztpn00an1n08x5 TAP_606 ();
 b15ztpn00an1n08x5 TAP_605 ();
 b15ztpn00an1n08x5 TAP_604 ();
 b15ztpn00an1n08x5 TAP_603 ();
 b15nona23al1n04x5 _28698_ (.a(net852),
    .b(\us30.a[6] ),
    .c(net849),
    .d(net846),
    .out0(_02807_));
 b15nanb02ah1n16x5 _28699_ (.a(net846),
    .b(\us30.a[6] ),
    .out0(_02808_));
 b15ztpn00an1n08x5 TAP_602 ();
 b15qgbxo2an1n05x5 _28701_ (.a(net856),
    .b(net849),
    .out0(_02810_));
 b15inv020as1n80x5 _28702_ (.a(net850),
    .o1(_02811_));
 b15oai013ar1n12x5 _28703_ (.a(_02807_),
    .b(_02808_),
    .c(_02810_),
    .d(_02811_),
    .o1(_02812_));
 b15aoi222ar1n02x5 _28704_ (.a(_02782_),
    .b(_02788_),
    .c(_02791_),
    .d(_02799_),
    .e(\us30.a[7] ),
    .f(_02812_),
    .o1(_02813_));
 b15orn002aq1n02x5 _28705_ (.a(net857),
    .b(_02813_),
    .o(_02814_));
 b15ztpn00an1n08x5 TAP_601 ();
 b15ztpn00an1n08x5 TAP_600 ();
 b15nonb03ar1n02x5 _28708_ (.a(net861),
    .b(net848),
    .c(\us30.a[6] ),
    .out0(_02818_));
 b15and002aq1n04x5 _28709_ (.a(\us30.a[4] ),
    .b(net844),
    .o(_02819_));
 b15inv000ah1n64x5 _28710_ (.a(net861),
    .o1(_02820_));
 b15ztpn00an1n08x5 TAP_599 ();
 b15aoi012ah1n02x5 _28712_ (.a(_02818_),
    .b(_02819_),
    .c(_02820_),
    .o1(_02822_));
 b15ztpn00an1n08x5 TAP_598 ();
 b15inv000an1n08x5 _28714_ (.a(net847),
    .o1(_02824_));
 b15inv020as1n10x5 _28715_ (.a(net843),
    .o1(_02825_));
 b15ztpn00an1n08x5 TAP_597 ();
 b15nonb02ar1n06x5 _28717_ (.a(net859),
    .b(net852),
    .out0(_02827_));
 b15nand04as1n04x5 _28718_ (.a(net856),
    .b(_02824_),
    .c(_02825_),
    .d(_02827_),
    .o1(_02829_));
 b15ztpn00an1n08x5 TAP_596 ();
 b15norp02aq1n48x5 _28720_ (.a(\us30.a[7] ),
    .b(net844),
    .o1(_02831_));
 b15ztpn00an1n08x5 TAP_595 ();
 b15nonb02as1n16x5 _28722_ (.a(\us30.a[5] ),
    .b(\us30.a[4] ),
    .out0(_02833_));
 b15nand03ah1n16x5 _28723_ (.a(net853),
    .b(_02831_),
    .c(_02833_),
    .o1(_02834_));
 b15ztpn00an1n08x5 TAP_594 ();
 b15ztpn00an1n08x5 TAP_593 ();
 b15nonb02aq1n12x5 _28726_ (.a(net860),
    .b(net858),
    .out0(_02837_));
 b15qgbna2an1n10x5 _28727_ (.a(\us30.a[3] ),
    .b(_02837_),
    .o1(_02838_));
 b15oai022ar1n06x5 _28728_ (.a(_02822_),
    .b(_02829_),
    .c(_02834_),
    .d(_02838_),
    .o1(_02840_));
 b15ztpn00an1n08x5 TAP_592 ();
 b15ztpn00an1n08x5 TAP_591 ();
 b15and002ar1n04x5 _28731_ (.a(net847),
    .b(\us30.a[7] ),
    .o(_02843_));
 b15nor002ah1n24x5 _28732_ (.a(\us30.a[1] ),
    .b(net852),
    .o1(_02844_));
 b15ztpn00an1n08x5 TAP_590 ();
 b15ztpn00an1n08x5 TAP_589 ();
 b15and003ar1n02x5 _28735_ (.a(net856),
    .b(net849),
    .c(net844),
    .o(_02847_));
 b15nor004an1n03x5 _28736_ (.a(\us30.a[0] ),
    .b(net856),
    .c(net849),
    .d(net844),
    .o1(_02848_));
 b15oai112al1n08x5 _28737_ (.a(_02843_),
    .b(_02844_),
    .c(_02847_),
    .d(_02848_),
    .o1(_02849_));
 b15nanb02ar1n02x5 _28738_ (.a(\us30.a[6] ),
    .b(net846),
    .out0(_02851_));
 b15ztpn00an1n08x5 TAP_588 ();
 b15oai012al1n06x5 _28740_ (.a(_02851_),
    .b(_02808_),
    .c(\us30.a[1] ),
    .o1(_02853_));
 b15inv000an1n80x5 _28741_ (.a(net854),
    .o1(_02854_));
 b15ztpn00an1n08x5 TAP_587 ();
 b15nanb02aq1n08x5 _28743_ (.a(\us30.a[7] ),
    .b(net849),
    .out0(_02856_));
 b15ztpn00an1n08x5 TAP_586 ();
 b15nanb02as1n24x5 _28745_ (.a(\us30.a[3] ),
    .b(\us30.a[0] ),
    .out0(_02858_));
 b15norp03ar1n02x5 _28746_ (.a(_02854_),
    .b(_02856_),
    .c(_02858_),
    .o1(_02859_));
 b15aob012aq1n06x5 _28747_ (.a(_02849_),
    .b(_02853_),
    .c(_02859_),
    .out0(_02860_));
 b15ornc04as1n24x5 _28748_ (.a(net846),
    .b(net849),
    .c(net843),
    .d(net845),
    .o(_02862_));
 b15ztpn00an1n08x5 TAP_585 ();
 b15nandp2ar1n48x5 _28750_ (.a(net851),
    .b(net853),
    .o1(_02864_));
 b15ztpn00an1n08x5 TAP_584 ();
 b15ztpn00an1n08x5 TAP_583 ();
 b15nanb02as1n24x5 _28753_ (.a(net862),
    .b(net852),
    .out0(_02867_));
 b15oai112ah1n04x5 _28754_ (.a(_02831_),
    .b(_02833_),
    .c(_02867_),
    .d(net858),
    .o1(_02868_));
 b15ztpn00an1n08x5 TAP_582 ();
 b15oai022ah1n06x5 _28756_ (.a(_02862_),
    .b(_02864_),
    .c(_02868_),
    .d(net855),
    .o1(_02870_));
 b15nandp2ah1n32x5 _28757_ (.a(net859),
    .b(net862),
    .o1(_02871_));
 b15nanb02as1n24x5 _28758_ (.a(net854),
    .b(net850),
    .out0(_02873_));
 b15nanb02as1n02x5 _28759_ (.a(_02871_),
    .b(_02873_),
    .out0(_02874_));
 b15aoi112ar1n06x5 _28760_ (.a(_02840_),
    .b(_02860_),
    .c(_02870_),
    .d(_02874_),
    .o1(_02875_));
 b15nona23as1n32x5 _28761_ (.a(\us30.a[7] ),
    .b(net844),
    .c(\us30.a[5] ),
    .d(\us30.a[4] ),
    .out0(_02876_));
 b15nonb02as1n16x5 _28762_ (.a(net859),
    .b(net862),
    .out0(_02877_));
 b15aoi013ar1n02x5 _28763_ (.a(_02811_),
    .b(net856),
    .c(_02876_),
    .d(_02877_),
    .o1(_02878_));
 b15nanb02ah1n16x5 _28764_ (.a(net849),
    .b(net846),
    .out0(_02879_));
 b15nandp2ah1n32x5 _28765_ (.a(net843),
    .b(\us30.a[6] ),
    .o1(_02880_));
 b15nor002as1n04x5 _28766_ (.a(_02879_),
    .b(_02880_),
    .o1(_02881_));
 b15nandp2as1n48x5 _28767_ (.a(net861),
    .b(net854),
    .o1(_02882_));
 b15ztpn00an1n08x5 TAP_581 ();
 b15nano23an1n16x5 _28769_ (.a(net846),
    .b(net848),
    .c(net843),
    .d(net845),
    .out0(_02885_));
 b15aoai13an1n02x5 _28770_ (.a(_02878_),
    .b(_02881_),
    .c(_02882_),
    .d(_02885_),
    .o1(_02886_));
 b15ztpn00an1n08x5 TAP_580 ();
 b15ztpn00an1n08x5 TAP_579 ();
 b15ztpn00an1n08x5 TAP_578 ();
 b15ztpn00an1n08x5 TAP_577 ();
 b15oaoi13ar1n02x5 _28775_ (.a(net857),
    .b(_02820_),
    .c(net856),
    .d(_02881_),
    .o1(_02891_));
 b15nandp2as1n16x5 _28776_ (.a(net857),
    .b(net850),
    .o1(_02892_));
 b15nona23ar1n02x5 _28777_ (.a(net862),
    .b(net845),
    .c(net849),
    .d(net846),
    .out0(_02893_));
 b15nanb02ar1n02x5 _28778_ (.a(net849),
    .b(net856),
    .out0(_02895_));
 b15oaoi13an1n03x5 _28779_ (.a(_02825_),
    .b(_02893_),
    .c(_02895_),
    .d(_02808_),
    .o1(_02896_));
 b15orn002al1n12x5 _28780_ (.a(net846),
    .b(net849),
    .o(_02897_));
 b15norp02as1n08x5 _28781_ (.a(_02794_),
    .b(_02897_),
    .o1(_02898_));
 b15and002as1n32x5 _28782_ (.a(net846),
    .b(net849),
    .o(_02899_));
 b15and002ar1n12x5 _28783_ (.a(_02899_),
    .b(_02781_),
    .o(_02900_));
 b15oaoi13ar1n02x5 _28784_ (.a(_02896_),
    .b(_02854_),
    .c(_02898_),
    .d(_02900_),
    .o1(_02901_));
 b15oa0022ar1n06x5 _28785_ (.a(_02886_),
    .b(_02891_),
    .c(_02892_),
    .d(_02901_),
    .o(_02902_));
 b15ztpn00an1n08x5 TAP_576 ();
 b15nonb02as1n16x5 _28787_ (.a(net844),
    .b(net843),
    .out0(_02904_));
 b15ztpn00an1n08x5 TAP_575 ();
 b15and003ar1n03x5 _28789_ (.a(net854),
    .b(net846),
    .c(net848),
    .o(_02907_));
 b15nano23an1n24x5 _28790_ (.a(net846),
    .b(net843),
    .c(net845),
    .d(net848),
    .out0(_02908_));
 b15aoi022aq1n04x5 _28791_ (.a(_02904_),
    .b(_02907_),
    .c(_02871_),
    .d(_02908_),
    .o1(_02909_));
 b15ztpn00an1n08x5 TAP_574 ();
 b15norp02an1n08x5 _28793_ (.a(net858),
    .b(net860),
    .o1(_02911_));
 b15ztpn00an1n08x5 TAP_573 ();
 b15nandp2ar1n48x5 _28795_ (.a(_02781_),
    .b(_02833_),
    .o1(_02913_));
 b15aoi112as1n04x5 _28796_ (.a(_02811_),
    .b(_02909_),
    .c(_02911_),
    .d(_02913_),
    .o1(_02914_));
 b15nonb02as1n16x5 _28797_ (.a(\us30.a[4] ),
    .b(\us30.a[5] ),
    .out0(_02915_));
 b15ztpn00an1n08x5 TAP_572 ();
 b15nandp2ah1n16x5 _28799_ (.a(_02904_),
    .b(_02915_),
    .o1(_02918_));
 b15nanb02as1n24x5 _28800_ (.a(net855),
    .b(net860),
    .out0(_02919_));
 b15and002aq1n32x5 _28801_ (.a(net843),
    .b(net844),
    .o(_02920_));
 b15nandp2aq1n48x5 _28802_ (.a(_02920_),
    .b(_02915_),
    .o1(_02921_));
 b15ztpn00an1n08x5 TAP_571 ();
 b15nanb02as1n24x5 _28804_ (.a(net862),
    .b(net859),
    .out0(_02923_));
 b15oai022ar1n02x5 _28805_ (.a(_02918_),
    .b(_02919_),
    .c(_02921_),
    .d(_02923_),
    .o1(_02924_));
 b15ztpn00an1n08x5 TAP_570 ();
 b15aoi012aq1n04x5 _28807_ (.a(_02914_),
    .b(_02924_),
    .c(_02811_),
    .o1(_02926_));
 b15nand04ah1n12x5 _28808_ (.a(_02814_),
    .b(_02875_),
    .c(_02902_),
    .d(_02926_),
    .o1(_02928_));
 b15nandp2as1n32x5 _28809_ (.a(_02831_),
    .b(_02915_),
    .o1(_02929_));
 b15ztpn00an1n08x5 TAP_569 ();
 b15ztpn00an1n08x5 TAP_568 ();
 b15nano23as1n24x5 _28812_ (.a(\us30.a[4] ),
    .b(net844),
    .c(\us30.a[7] ),
    .d(\us30.a[5] ),
    .out0(_02932_));
 b15nanb02al1n12x5 _28813_ (.a(net859),
    .b(net853),
    .out0(_02933_));
 b15nand03ah1n02x5 _28814_ (.a(net850),
    .b(_02932_),
    .c(_02933_),
    .o1(_02934_));
 b15nand02ah1n24x5 _28815_ (.a(net859),
    .b(net856),
    .o1(_02935_));
 b15aoai13ar1n02x5 _28816_ (.a(_02935_),
    .b(net859),
    .c(_02831_),
    .d(_02915_),
    .o1(_02936_));
 b15ztpn00an1n08x5 TAP_567 ();
 b15aoi022ar1n04x5 _28818_ (.a(_02929_),
    .b(_02934_),
    .c(_02936_),
    .d(_02820_),
    .o1(_02939_));
 b15nanb02as1n24x5 _28819_ (.a(net851),
    .b(net853),
    .out0(_02940_));
 b15norp02ar1n03x5 _28820_ (.a(net859),
    .b(_02940_),
    .o1(_02941_));
 b15nandp3ah1n24x5 _28821_ (.a(net852),
    .b(_02831_),
    .c(_02915_),
    .o1(_02942_));
 b15nonb02aq1n16x5 _28822_ (.a(net859),
    .b(net853),
    .out0(_02943_));
 b15aoi012ar1n02x5 _28823_ (.a(_02941_),
    .b(_02942_),
    .c(_02943_),
    .o1(_02944_));
 b15ztpn00an1n08x5 TAP_566 ();
 b15oai012aq1n03x5 _28825_ (.a(_02939_),
    .b(_02944_),
    .c(_02820_),
    .o1(_02946_));
 b15nonb02as1n16x5 _28826_ (.a(\us30.a[0] ),
    .b(net852),
    .out0(_02947_));
 b15nandp2ah1n05x5 _28827_ (.a(_02854_),
    .b(_02947_),
    .o1(_02948_));
 b15nandp2aq1n32x5 _28828_ (.a(_02779_),
    .b(_02781_),
    .o1(_02950_));
 b15inv040as1n60x5 _28829_ (.a(net857),
    .o1(_02951_));
 b15ztpn00an1n08x5 TAP_565 ();
 b15oaoi13an1n03x5 _28831_ (.a(_02948_),
    .b(_02876_),
    .c(_02950_),
    .d(_02951_),
    .o1(_02953_));
 b15nandp2as1n24x5 _28832_ (.a(_02831_),
    .b(_02833_),
    .o1(_02954_));
 b15ztpn00an1n08x5 TAP_564 ();
 b15nanb02as1n24x5 _28834_ (.a(net850),
    .b(net857),
    .out0(_02956_));
 b15orn002as1n12x5 _28835_ (.a(net858),
    .b(net860),
    .o(_02957_));
 b15oai022as1n02x5 _28836_ (.a(_02954_),
    .b(_02956_),
    .c(_02957_),
    .d(_02862_),
    .o1(_02958_));
 b15ztpn00an1n08x5 TAP_563 ();
 b15aoi012an1n08x5 _28838_ (.a(_02953_),
    .b(_02958_),
    .c(net855),
    .o1(_02961_));
 b15ztpn00an1n08x5 TAP_562 ();
 b15ztpn00an1n08x5 TAP_561 ();
 b15nandp2aq1n32x5 _28841_ (.a(_02899_),
    .b(_02781_),
    .o1(_02964_));
 b15nor002ah1n03x5 _28842_ (.a(_02940_),
    .b(_02964_),
    .o1(_02965_));
 b15orn003ar1n02x5 _28843_ (.a(net852),
    .b(_02824_),
    .c(_02856_),
    .o(_02966_));
 b15xor002al1n04x5 _28844_ (.a(\us30.a[1] ),
    .b(net849),
    .out0(_02967_));
 b15nand02an1n06x5 _28845_ (.a(net852),
    .b(\us30.a[7] ),
    .o1(_02968_));
 b15ztpn00an1n08x5 TAP_560 ();
 b15oai013ar1n08x5 _28847_ (.a(_02966_),
    .b(_02967_),
    .c(_02968_),
    .d(net847),
    .o1(_02970_));
 b15ztpn00an1n08x5 TAP_559 ();
 b15aoai13ah1n03x5 _28849_ (.a(net862),
    .b(_02965_),
    .c(_02970_),
    .d(\us30.a[6] ),
    .o1(_02973_));
 b15nano23as1n24x5 _28850_ (.a(net849),
    .b(net843),
    .c(net844),
    .d(net847),
    .out0(_02974_));
 b15ztpn00an1n08x5 TAP_558 ();
 b15oai112al1n06x5 _28852_ (.a(_02951_),
    .b(_02919_),
    .c(_02864_),
    .d(net862),
    .o1(_02976_));
 b15nonb02ah1n12x5 _28853_ (.a(net850),
    .b(net855),
    .out0(_02977_));
 b15aoi012ar1n02x5 _28854_ (.a(_02791_),
    .b(_02977_),
    .c(_02820_),
    .o1(_02978_));
 b15oai112an1n02x5 _28855_ (.a(net859),
    .b(_02978_),
    .c(_02977_),
    .d(_02820_),
    .o1(_02979_));
 b15nandp3al1n04x5 _28856_ (.a(_02974_),
    .b(_02976_),
    .c(_02979_),
    .o1(_02980_));
 b15nand04aq1n12x5 _28857_ (.a(_02946_),
    .b(_02961_),
    .c(_02973_),
    .d(_02980_),
    .o1(_02981_));
 b15ztpn00an1n08x5 TAP_557 ();
 b15nandp2ah1n32x5 _28859_ (.a(_02904_),
    .b(_02779_),
    .o1(_02984_));
 b15nand02as1n12x5 _28860_ (.a(_02854_),
    .b(_02871_),
    .o1(_02985_));
 b15nand02aq1n32x5 _28861_ (.a(_02904_),
    .b(_02899_),
    .o1(_02986_));
 b15ztpn00an1n08x5 TAP_556 ();
 b15oai022ar1n02x5 _28863_ (.a(_02882_),
    .b(_02984_),
    .c(_02985_),
    .d(_02986_),
    .o1(_02988_));
 b15nor002ah1n24x5 _28864_ (.a(net859),
    .b(net855),
    .o1(_02989_));
 b15aoai13ar1n03x5 _28865_ (.a(net850),
    .b(_02988_),
    .c(_02989_),
    .d(_02782_),
    .o1(_02990_));
 b15ztpn00an1n08x5 TAP_555 ();
 b15nandp2as1n16x5 _28867_ (.a(_02833_),
    .b(_02920_),
    .o1(_02992_));
 b15oai013as1n06x5 _28868_ (.a(_02990_),
    .b(_02985_),
    .c(_02992_),
    .d(net850),
    .o1(_02994_));
 b15nand02ar1n24x5 _28869_ (.a(_02951_),
    .b(_02854_),
    .o1(_02995_));
 b15nandp3as1n04x5 _28870_ (.a(net862),
    .b(_02904_),
    .c(_02779_),
    .o1(_02996_));
 b15nona23as1n32x5 _28871_ (.a(net846),
    .b(net849),
    .c(net843),
    .d(net845),
    .out0(_02997_));
 b15oaoi13as1n02x5 _28872_ (.a(_02995_),
    .b(_02996_),
    .c(_02997_),
    .d(net862),
    .o1(_02998_));
 b15ztpn00an1n08x5 TAP_554 ();
 b15nonb02as1n08x5 _28874_ (.a(net846),
    .b(net856),
    .out0(_03000_));
 b15norp03ar1n02x5 _28875_ (.a(net846),
    .b(net848),
    .c(\us30.a[6] ),
    .o1(_03001_));
 b15and002ah1n16x5 _28876_ (.a(net861),
    .b(net854),
    .o(_03002_));
 b15aoi022ar1n02x5 _28877_ (.a(_02819_),
    .b(_03000_),
    .c(_03001_),
    .d(_03002_),
    .o1(_03003_));
 b15nor003aq1n02x5 _28878_ (.a(net857),
    .b(_02825_),
    .c(_03003_),
    .o1(_03005_));
 b15nand03al1n03x5 _28879_ (.a(net859),
    .b(\us30.a[6] ),
    .c(_02833_),
    .o1(_03006_));
 b15nand02ar1n02x5 _28880_ (.a(net856),
    .b(\us30.a[7] ),
    .o1(_03007_));
 b15oaoi13ar1n04x5 _28881_ (.a(_03006_),
    .b(_03007_),
    .c(_02820_),
    .d(\us30.a[7] ),
    .o1(_03008_));
 b15ztpn00an1n08x5 TAP_553 ();
 b15nor002ah1n06x5 _28883_ (.a(net848),
    .b(net843),
    .o1(_03010_));
 b15nandp2al1n16x5 _28884_ (.a(\us30.a[4] ),
    .b(\us30.a[7] ),
    .o1(_03011_));
 b15oab012an1n02x5 _28885_ (.a(_03010_),
    .b(_03011_),
    .c(net861),
    .out0(_03012_));
 b15nand02an1n02x5 _28886_ (.a(net845),
    .b(_03000_),
    .o1(_03013_));
 b15oai122as1n08x5 _28887_ (.a(_02811_),
    .b(_02992_),
    .c(_02882_),
    .d(_03012_),
    .e(_03013_),
    .o1(_03014_));
 b15nor004ar1n06x5 _28888_ (.a(_02998_),
    .b(_03005_),
    .c(_03008_),
    .d(_03014_),
    .o1(_03016_));
 b15aoi012ar1n02x5 _28889_ (.a(_02951_),
    .b(_02996_),
    .c(_02997_),
    .o1(_03017_));
 b15nano23as1n24x5 _28890_ (.a(\us30.a[7] ),
    .b(net844),
    .c(\us30.a[5] ),
    .d(\us30.a[4] ),
    .out0(_03018_));
 b15aoai13ar1n04x5 _28891_ (.a(net855),
    .b(_03017_),
    .c(_03018_),
    .d(net862),
    .o1(_03019_));
 b15nanb02as1n24x5 _28892_ (.a(net858),
    .b(net860),
    .out0(_03020_));
 b15qgbno2an1n10x5 _28893_ (.a(net854),
    .b(_03020_),
    .o1(_03021_));
 b15ztpn00an1n08x5 TAP_552 ();
 b15norp02aq1n16x5 _28895_ (.a(_02798_),
    .b(_02880_),
    .o1(_03023_));
 b15nano23as1n24x5 _28896_ (.a(net846),
    .b(net845),
    .c(net843),
    .d(net849),
    .out0(_03024_));
 b15ztpn00an1n08x5 TAP_551 ();
 b15oaoi13ar1n04x5 _28898_ (.a(_02811_),
    .b(_03021_),
    .c(_03023_),
    .d(_03024_),
    .o1(_03027_));
 b15nand02ah1n12x5 _28899_ (.a(_02904_),
    .b(_02833_),
    .o1(_03028_));
 b15nand04as1n16x5 _28900_ (.a(\us30.a[5] ),
    .b(\us30.a[4] ),
    .c(\us30.a[7] ),
    .d(net844),
    .o1(_03029_));
 b15ztpn00an1n08x5 TAP_550 ();
 b15oai022ar1n02x5 _28902_ (.a(_02951_),
    .b(_03028_),
    .c(_03029_),
    .d(net862),
    .o1(_03031_));
 b15nand02al1n04x5 _28903_ (.a(net855),
    .b(_03031_),
    .o1(_03032_));
 b15aoi022an1n08x5 _28904_ (.a(_03016_),
    .b(_03019_),
    .c(_03027_),
    .d(_03032_),
    .o1(_03033_));
 b15nor004as1n12x5 _28905_ (.a(_02928_),
    .b(_02981_),
    .c(_02994_),
    .d(_03033_),
    .o1(_03034_));
 b15ztpn00an1n08x5 TAP_549 ();
 b15inv020an1n80x5 _28907_ (.a(net581),
    .o1(_03036_));
 b15ztpn00an1n08x5 TAP_548 ();
 b15ztpn00an1n08x5 TAP_547 ();
 b15ztpn00an1n08x5 TAP_546 ();
 b15ztpn00an1n08x5 TAP_545 ();
 b15ztpn00an1n08x5 TAP_544 ();
 b15ztpn00an1n08x5 TAP_543 ();
 b15nona23aq1n24x5 _28914_ (.a(net576),
    .b(net572),
    .c(net570),
    .d(net578),
    .out0(_03044_));
 b15ztpn00an1n08x5 TAP_542 ();
 b15nandp2aq1n48x5 _28916_ (.a(net589),
    .b(net586),
    .o1(_03046_));
 b15norp02ar1n08x5 _28917_ (.a(_03044_),
    .b(_03046_),
    .o1(_03047_));
 b15ztpn00an1n08x5 TAP_541 ();
 b15orn002aq1n24x5 _28919_ (.a(net576),
    .b(net578),
    .o(_03050_));
 b15ztpn00an1n08x5 TAP_540 ();
 b15ztpn00an1n08x5 TAP_539 ();
 b15orn002aq1n32x5 _28922_ (.a(net568),
    .b(net571),
    .o(_03053_));
 b15ztpn00an1n08x5 TAP_538 ();
 b15ztpn00an1n08x5 TAP_537 ();
 b15ztpn00an1n08x5 TAP_536 ();
 b15norp02an1n32x5 _28926_ (.a(net593),
    .b(net589),
    .o1(_03057_));
 b15ztpn00an1n08x5 TAP_535 ();
 b15ztpn00an1n08x5 TAP_534 ();
 b15and003al1n12x5 _28929_ (.a(net593),
    .b(net589),
    .c(net585),
    .o(_03061_));
 b15nor004ar1n02x5 _28930_ (.a(_03050_),
    .b(_03053_),
    .c(_03057_),
    .d(_03061_),
    .o1(_03062_));
 b15orn003ar1n02x5 _28931_ (.a(_03036_),
    .b(_03047_),
    .c(_03062_),
    .o(_03063_));
 b15ztpn00an1n08x5 TAP_533 ();
 b15ztpn00an1n08x5 TAP_532 ();
 b15ztpn00an1n08x5 TAP_531 ();
 b15inv040ah1n36x5 _28935_ (.a(net586),
    .o1(_03067_));
 b15nanb02as1n24x5 _28936_ (.a(net577),
    .b(net574),
    .out0(_03068_));
 b15ztpn00an1n08x5 TAP_530 ();
 b15nandp2ah1n32x5 _28938_ (.a(net568),
    .b(net571),
    .o1(_03071_));
 b15ztpn00an1n08x5 TAP_529 ();
 b15nor003ah1n08x5 _28940_ (.a(_03067_),
    .b(_03068_),
    .c(_03071_),
    .o1(_03073_));
 b15nanb02ah1n12x5 _28941_ (.a(net585),
    .b(net572),
    .out0(_03074_));
 b15nandp2ah1n24x5 _28942_ (.a(net593),
    .b(net586),
    .o1(_03075_));
 b15ztpn00an1n08x5 TAP_528 ();
 b15oai012ar1n02x5 _28944_ (.a(_03074_),
    .b(_03075_),
    .c(net572),
    .o1(_03077_));
 b15ztpn00an1n08x5 TAP_527 ();
 b15nanb02as1n24x5 _28946_ (.a(net576),
    .b(net578),
    .out0(_03079_));
 b15ztpn00an1n08x5 TAP_526 ();
 b15norp02ar1n02x5 _28948_ (.a(net569),
    .b(_03079_),
    .o1(_03082_));
 b15aoi112al1n02x5 _28949_ (.a(net587),
    .b(_03073_),
    .c(_03077_),
    .d(_03082_),
    .o1(_03083_));
 b15ztpn00an1n08x5 TAP_525 ();
 b15ztpn00an1n08x5 TAP_524 ();
 b15nanb02as1n24x5 _28952_ (.a(net572),
    .b(net569),
    .out0(_03086_));
 b15nandp2aq1n32x5 _28953_ (.a(net576),
    .b(net578),
    .o1(_03087_));
 b15norp02ah1n24x5 _28954_ (.a(_03086_),
    .b(_03087_),
    .o1(_03088_));
 b15nor002ah1n12x5 _28955_ (.a(_03079_),
    .b(_03053_),
    .o1(_03089_));
 b15aoi022ar1n02x5 _28956_ (.a(net591),
    .b(_03088_),
    .c(_03089_),
    .d(_03075_),
    .o1(_03090_));
 b15ztpn00an1n08x5 TAP_523 ();
 b15ztpn00an1n08x5 TAP_522 ();
 b15ztpn00an1n08x5 TAP_521 ();
 b15aoi012as1n02x5 _28960_ (.a(_03083_),
    .b(_03090_),
    .c(net587),
    .o1(_03095_));
 b15ztpn00an1n08x5 TAP_520 ();
 b15inv000ah1n20x5 _28962_ (.a(net571),
    .o1(_03097_));
 b15ztpn00an1n08x5 TAP_519 ();
 b15norp03ar1n02x5 _28964_ (.a(net569),
    .b(_03079_),
    .c(_03046_),
    .o1(_03099_));
 b15inv020aq1n32x5 _28965_ (.a(net575),
    .o1(_03100_));
 b15ztpn00an1n08x5 TAP_518 ();
 b15inv000al1n80x5 _28967_ (.a(net591),
    .o1(_03102_));
 b15ztpn00an1n08x5 TAP_517 ();
 b15ztpn00an1n08x5 TAP_516 ();
 b15nonb02ah1n12x5 _28970_ (.a(net579),
    .b(net568),
    .out0(_03106_));
 b15nonb02aq1n16x5 _28971_ (.a(net588),
    .b(net584),
    .out0(_03107_));
 b15nonb02as1n08x5 _28972_ (.a(net568),
    .b(net579),
    .out0(_03108_));
 b15aoi022ar1n02x5 _28973_ (.a(net584),
    .b(_03106_),
    .c(_03107_),
    .d(_03108_),
    .o1(_03109_));
 b15nor003ar1n02x5 _28974_ (.a(_03100_),
    .b(_03102_),
    .c(_03109_),
    .o1(_03110_));
 b15oab012al1n03x5 _28975_ (.a(_03097_),
    .b(_03099_),
    .c(_03110_),
    .out0(_03111_));
 b15ztpn00an1n08x5 TAP_515 ();
 b15ztpn00an1n08x5 TAP_514 ();
 b15ztpn00an1n08x5 TAP_513 ();
 b15oai013as1n04x5 _28979_ (.a(_03063_),
    .b(_03095_),
    .c(_03111_),
    .d(net580),
    .o1(_03116_));
 b15ztpn00an1n08x5 TAP_512 ();
 b15ztpn00an1n08x5 TAP_511 ();
 b15ztpn00an1n08x5 TAP_510 ();
 b15ztpn00an1n08x5 TAP_509 ();
 b15nona23aq1n16x5 _28984_ (.a(net577),
    .b(net568),
    .c(net571),
    .d(net574),
    .out0(_03121_));
 b15nor002aq1n08x5 _28985_ (.a(net580),
    .b(_03121_),
    .o1(_03122_));
 b15nanb02as1n24x5 _28986_ (.a(net593),
    .b(net589),
    .out0(_03123_));
 b15ztpn00an1n08x5 TAP_508 ();
 b15nanb03ah1n08x5 _28988_ (.a(net569),
    .b(net572),
    .c(net580),
    .out0(_03126_));
 b15oaoi13ar1n02x5 _28989_ (.a(_03123_),
    .b(_03121_),
    .c(_03126_),
    .d(_03087_),
    .o1(_03127_));
 b15norp02aq1n08x5 _28990_ (.a(_03087_),
    .b(_03126_),
    .o1(_03128_));
 b15nonb02as1n16x5 _28991_ (.a(net592),
    .b(net588),
    .out0(_03129_));
 b15aoi112an1n02x5 _28992_ (.a(_03122_),
    .b(_03127_),
    .c(_03128_),
    .d(_03129_),
    .o1(_03130_));
 b15ztpn00an1n08x5 TAP_507 ();
 b15nano23as1n24x5 _28994_ (.a(net576),
    .b(\us23.a[6] ),
    .c(net570),
    .d(net578),
    .out0(_03132_));
 b15ztpn00an1n08x5 TAP_506 ();
 b15and002as1n08x5 _28996_ (.a(net587),
    .b(net580),
    .o(_03134_));
 b15nanb02as1n24x5 _28997_ (.a(net568),
    .b(net571),
    .out0(_03135_));
 b15norp02ar1n48x5 _28998_ (.a(_03087_),
    .b(_03135_),
    .o1(_03137_));
 b15aoai13ar1n02x5 _28999_ (.a(net591),
    .b(_03132_),
    .c(_03134_),
    .d(_03137_),
    .o1(_03138_));
 b15ztpn00an1n08x5 TAP_505 ();
 b15qgbno2an1n10x5 _29001_ (.a(net589),
    .b(_03036_),
    .o1(_03140_));
 b15aoi012ar1n02x5 _29002_ (.a(net585),
    .b(_03132_),
    .c(_03140_),
    .o1(_03141_));
 b15aoi022an1n04x5 _29003_ (.a(net585),
    .b(_03130_),
    .c(_03138_),
    .d(_03141_),
    .o1(_03142_));
 b15and002aq1n32x5 _29004_ (.a(net568),
    .b(net573),
    .o(_03143_));
 b15nanb02ah1n12x5 _29005_ (.a(net589),
    .b(net594),
    .out0(_03144_));
 b15nand02ar1n02x5 _29006_ (.a(net585),
    .b(_03144_),
    .o1(_03145_));
 b15oai012ar1n02x5 _29007_ (.a(_03079_),
    .b(_03068_),
    .c(_03129_),
    .o1(_03146_));
 b15aoi013ar1n02x5 _29008_ (.a(_03036_),
    .b(_03143_),
    .c(_03145_),
    .d(_03146_),
    .o1(_03148_));
 b15nor002al1n16x5 _29009_ (.a(_03053_),
    .b(_03068_),
    .o1(_03149_));
 b15nor002aq1n12x5 _29010_ (.a(_03079_),
    .b(_03071_),
    .o1(_03150_));
 b15ztpn00an1n08x5 TAP_504 ();
 b15aoi022ar1n02x5 _29012_ (.a(net585),
    .b(_03149_),
    .c(_03150_),
    .d(net587),
    .o1(_03152_));
 b15ztpn00an1n08x5 TAP_503 ();
 b15ztpn00an1n08x5 TAP_502 ();
 b15oai012al1n02x5 _29015_ (.a(_03148_),
    .b(_03152_),
    .c(net593),
    .o1(_03155_));
 b15ztpn00an1n08x5 TAP_501 ();
 b15andc04as1n16x5 _29017_ (.a(net575),
    .b(net579),
    .c(\us23.a[7] ),
    .d(\us23.a[6] ),
    .o(_03157_));
 b15oab012al1n08x5 _29018_ (.c(net594),
    .a(net586),
    .b(net589),
    .out0(_03159_));
 b15aoi012al1n04x5 _29019_ (.a(net581),
    .b(_03157_),
    .c(_03159_),
    .o1(_03160_));
 b15ztpn00an1n08x5 TAP_500 ();
 b15nonb02as1n16x5 _29021_ (.a(net568),
    .b(net573),
    .out0(_03162_));
 b15inv000as1n40x5 _29022_ (.a(net589),
    .o1(_03163_));
 b15nandp2as1n04x5 _29023_ (.a(_03100_),
    .b(_03163_),
    .o1(_03164_));
 b15nor002al1n16x5 _29024_ (.a(net593),
    .b(net586),
    .o1(_03165_));
 b15nand04ar1n03x5 _29025_ (.a(net577),
    .b(_03162_),
    .c(_03164_),
    .d(_03165_),
    .o1(_03166_));
 b15nand04as1n16x5 _29026_ (.a(net576),
    .b(net578),
    .c(net570),
    .d(\us23.a[6] ),
    .o1(_03167_));
 b15nanb02as1n08x5 _29027_ (.a(net589),
    .b(net586),
    .out0(_03168_));
 b15nor002aq1n08x5 _29028_ (.a(_03167_),
    .b(_03168_),
    .o1(_03170_));
 b15nano23aq1n24x5 _29029_ (.a(net568),
    .b(net571),
    .c(net574),
    .d(net577),
    .out0(_03171_));
 b15aoi012ar1n02x5 _29030_ (.a(_03170_),
    .b(_03171_),
    .c(_03107_),
    .o1(_03172_));
 b15oai112ar1n04x5 _29031_ (.a(_03160_),
    .b(_03166_),
    .c(net591),
    .d(_03172_),
    .o1(_03173_));
 b15ztpn00an1n08x5 TAP_499 ();
 b15nandp2as1n08x5 _29033_ (.a(net577),
    .b(net568),
    .o1(_03175_));
 b15ztpn00an1n08x5 TAP_498 ();
 b15nonb02al1n04x5 _29035_ (.a(net592),
    .b(net571),
    .out0(_03177_));
 b15nanb02al1n02x5 _29036_ (.a(_03175_),
    .b(_03177_),
    .out0(_03178_));
 b15nandp2aq1n05x5 _29037_ (.a(net574),
    .b(net584),
    .o1(_03179_));
 b15orn002al1n32x5 _29038_ (.a(net589),
    .b(net586),
    .o(_03181_));
 b15ztpn00an1n08x5 TAP_497 ();
 b15ztpn00an1n08x5 TAP_496 ();
 b15oaoi13ar1n04x5 _29041_ (.a(_03178_),
    .b(_03179_),
    .c(_03181_),
    .d(net574),
    .o1(_03184_));
 b15oaoi13al1n02x5 _29042_ (.a(_03142_),
    .b(_03155_),
    .c(_03173_),
    .d(_03184_),
    .o1(_03185_));
 b15nonb02as1n16x5 _29043_ (.a(net584),
    .b(net595),
    .out0(_03186_));
 b15nona23as1n32x5 _29044_ (.a(net575),
    .b(net579),
    .c(\us23.a[7] ),
    .d(\us23.a[6] ),
    .out0(_03187_));
 b15ztpn00an1n08x5 TAP_495 ();
 b15norp02al1n12x5 _29046_ (.a(_03036_),
    .b(_03187_),
    .o1(_03189_));
 b15ztpn00an1n08x5 TAP_494 ();
 b15norp03ar1n16x5 _29048_ (.a(net587),
    .b(_03086_),
    .c(_03087_),
    .o1(_03192_));
 b15nanb02ar1n24x5 _29049_ (.a(net582),
    .b(net590),
    .out0(_03193_));
 b15norp03ar1n03x5 _29050_ (.a(_03100_),
    .b(_03053_),
    .c(_03193_),
    .o1(_03194_));
 b15oai013an1n03x5 _29051_ (.a(_03186_),
    .b(_03189_),
    .c(_03192_),
    .d(_03194_),
    .o1(_03195_));
 b15nonb02as1n16x5 _29052_ (.a(net595),
    .b(net584),
    .out0(_03196_));
 b15ztpn00an1n08x5 TAP_493 ();
 b15ztpn00an1n08x5 TAP_492 ();
 b15nano23as1n24x5 _29055_ (.a(net576),
    .b(net578),
    .c(net570),
    .d(\us23.a[6] ),
    .out0(_03199_));
 b15nandp2ar1n03x5 _29056_ (.a(net583),
    .b(_03199_),
    .o1(_03200_));
 b15orn002al1n08x5 _29057_ (.a(net588),
    .b(net582),
    .o(_03201_));
 b15norp02ar1n48x5 _29058_ (.a(\us23.a[7] ),
    .b(net573),
    .o1(_03203_));
 b15nonb02as1n16x5 _29059_ (.a(net575),
    .b(net579),
    .out0(_03204_));
 b15nandp2ah1n24x5 _29060_ (.a(_03203_),
    .b(_03204_),
    .o1(_03205_));
 b15oai012ar1n02x5 _29061_ (.a(_03200_),
    .b(_03201_),
    .c(_03205_),
    .o1(_03206_));
 b15and002an1n16x5 _29062_ (.a(net593),
    .b(net586),
    .o(_03207_));
 b15aoi022an1n02x5 _29063_ (.a(_03189_),
    .b(_03196_),
    .c(_03206_),
    .d(_03207_),
    .o1(_03208_));
 b15ztpn00an1n08x5 TAP_491 ();
 b15orn002ar1n24x5 _29065_ (.a(net594),
    .b(net590),
    .o(_03210_));
 b15nandp3ar1n02x5 _29066_ (.a(_03036_),
    .b(_03210_),
    .c(_03199_),
    .o1(_03211_));
 b15nand02ah1n06x5 _29067_ (.a(net594),
    .b(net583),
    .o1(_03212_));
 b15oaoi13an1n02x5 _29068_ (.a(net586),
    .b(_03211_),
    .c(_03212_),
    .d(_03205_),
    .o1(_03214_));
 b15norp02as1n12x5 _29069_ (.a(_03086_),
    .b(_03050_),
    .o1(_03215_));
 b15norp02ar1n03x5 _29070_ (.a(net592),
    .b(_03201_),
    .o1(_03216_));
 b15orn002al1n32x5 _29071_ (.a(net585),
    .b(net580),
    .o(_03217_));
 b15ztpn00an1n08x5 TAP_490 ();
 b15and002an1n24x5 _29073_ (.a(net586),
    .b(net582),
    .o(_03219_));
 b15aoi022ar1n02x5 _29074_ (.a(net593),
    .b(_03217_),
    .c(_03219_),
    .d(net588),
    .o1(_03220_));
 b15nanb02ar1n02x5 _29075_ (.a(_03216_),
    .b(_03220_),
    .out0(_03221_));
 b15aoi012ah1n02x5 _29076_ (.a(_03214_),
    .b(_03215_),
    .c(_03221_),
    .o1(_03222_));
 b15inv020ar1n32x5 _29077_ (.a(net577),
    .o1(_03223_));
 b15ztpn00an1n08x5 TAP_489 ();
 b15oai022ar1n02x5 _29079_ (.a(net574),
    .b(_03135_),
    .c(_03179_),
    .d(_03086_),
    .o1(_03226_));
 b15and002ah1n03x5 _29080_ (.a(_03223_),
    .b(_03226_),
    .o(_03227_));
 b15and002an1n32x5 _29081_ (.a(net575),
    .b(net579),
    .o(_03228_));
 b15ztpn00an1n08x5 TAP_488 ();
 b15ztpn00an1n08x5 TAP_487 ();
 b15nonb02as1n08x5 _29084_ (.a(net571),
    .b(net568),
    .out0(_03231_));
 b15nandp3ar1n02x5 _29085_ (.a(net592),
    .b(_03228_),
    .c(_03231_),
    .o1(_03232_));
 b15nor002ah1n32x5 _29086_ (.a(net575),
    .b(net579),
    .o1(_03233_));
 b15nand02aq1n16x5 _29087_ (.a(_03162_),
    .b(_03233_),
    .o1(_03234_));
 b15oai012ar1n03x5 _29088_ (.a(_03232_),
    .b(_03234_),
    .c(net592),
    .o1(_03236_));
 b15nor002aq1n32x5 _29089_ (.a(\us23.a[2] ),
    .b(net583),
    .o1(_03237_));
 b15aoi022an1n02x5 _29090_ (.a(_03216_),
    .b(_03227_),
    .c(_03236_),
    .d(_03237_),
    .o1(_03238_));
 b15nand04al1n08x5 _29091_ (.a(_03195_),
    .b(_03208_),
    .c(_03222_),
    .d(_03238_),
    .o1(_03239_));
 b15nor004as1n12x5 _29092_ (.a(net575),
    .b(net579),
    .c(net570),
    .d(\us23.a[6] ),
    .o1(_03240_));
 b15nandp3as1n04x5 _29093_ (.a(_03240_),
    .b(_03057_),
    .c(_03237_),
    .o1(_03241_));
 b15orn002ar1n08x5 _29094_ (.a(net592),
    .b(net584),
    .o(_03242_));
 b15qgbna2an1n05x5 _29095_ (.o1(_03243_),
    .a(_03233_),
    .b(_03242_));
 b15oai013as1n12x5 _29096_ (.a(_03241_),
    .b(_03243_),
    .c(_03061_),
    .d(_03126_),
    .o1(_03244_));
 b15nand02ar1n02x5 _29097_ (.a(_03134_),
    .b(_03157_),
    .o1(_03245_));
 b15nandp2ar1n24x5 _29098_ (.a(_03204_),
    .b(_03143_),
    .o1(_03247_));
 b15oaoi13ar1n02x5 _29099_ (.a(net592),
    .b(_03245_),
    .c(_03201_),
    .d(_03247_),
    .o1(_03248_));
 b15nanb02as1n24x5 _29100_ (.a(net584),
    .b(net580),
    .out0(_03249_));
 b15ztpn00an1n08x5 TAP_486 ();
 b15nonb02as1n16x5 _29102_ (.a(net579),
    .b(net575),
    .out0(_03251_));
 b15nandp2ah1n16x5 _29103_ (.a(_03251_),
    .b(_03203_),
    .o1(_03252_));
 b15xor002as1n16x5 _29104_ (.a(net591),
    .b(net588),
    .out0(_03253_));
 b15oaoi13ah1n02x5 _29105_ (.a(_03249_),
    .b(_03167_),
    .c(_03252_),
    .d(_03253_),
    .o1(_03254_));
 b15nonb02as1n16x5 _29106_ (.a(net585),
    .b(net589),
    .out0(_03255_));
 b15nandp3ar1n02x5 _29107_ (.a(net583),
    .b(_03255_),
    .c(_03171_),
    .o1(_03256_));
 b15oai012ar1n02x5 _29108_ (.a(_03256_),
    .b(_03200_),
    .c(_03210_),
    .o1(_03258_));
 b15nor004aq1n02x5 _29109_ (.a(_03244_),
    .b(_03248_),
    .c(_03254_),
    .d(_03258_),
    .o1(_03259_));
 b15ztpn00an1n08x5 TAP_485 ();
 b15nor003as1n16x5 _29111_ (.a(net579),
    .b(net568),
    .c(net573),
    .o1(_03261_));
 b15ztpn00an1n08x5 TAP_484 ();
 b15aoi112ar1n02x5 _29113_ (.a(net574),
    .b(net580),
    .c(_03075_),
    .d(_03163_),
    .o1(_03263_));
 b15ztpn00an1n08x5 TAP_483 ();
 b15ztpn00an1n08x5 TAP_482 ();
 b15ztpn00an1n08x5 TAP_481 ();
 b15aoai13al1n02x5 _29117_ (.a(_03261_),
    .b(_03263_),
    .c(net574),
    .d(_03134_),
    .o1(_03267_));
 b15ztpn00an1n08x5 TAP_480 ();
 b15nano23as1n24x5 _29119_ (.a(net578),
    .b(\us23.a[6] ),
    .c(net570),
    .d(net576),
    .out0(_03270_));
 b15nand02ar1n02x5 _29120_ (.a(net594),
    .b(_03270_),
    .o1(_03271_));
 b15nand02an1n48x5 _29121_ (.a(_03251_),
    .b(_03143_),
    .o1(_03272_));
 b15oai013al1n04x5 _29122_ (.a(_03271_),
    .b(_03217_),
    .c(_03272_),
    .d(net594),
    .o1(_03273_));
 b15nor002ar1n24x5 _29123_ (.a(net587),
    .b(net581),
    .o1(_03274_));
 b15nand04ah1n02x5 _29124_ (.a(net585),
    .b(_03251_),
    .c(_03143_),
    .d(_03274_),
    .o1(_03275_));
 b15nona23ah1n16x5 _29125_ (.a(net576),
    .b(net569),
    .c(net572),
    .d(net578),
    .out0(_03276_));
 b15oai012an1n03x5 _29126_ (.a(_03275_),
    .b(_03276_),
    .c(net586),
    .o1(_03277_));
 b15ztpn00an1n08x5 TAP_479 ();
 b15aoi022an1n08x5 _29128_ (.a(net589),
    .b(_03273_),
    .c(_03277_),
    .d(net594),
    .o1(_03280_));
 b15nandp2as1n24x5 _29129_ (.a(net591),
    .b(net588),
    .o1(_03281_));
 b15nandp2an1n05x5 _29130_ (.a(_03281_),
    .b(_03237_),
    .o1(_03282_));
 b15nanb02as1n24x5 _29131_ (.a(net584),
    .b(net590),
    .out0(_03283_));
 b15oai012aq1n08x5 _29132_ (.a(_03283_),
    .b(_03255_),
    .c(net591),
    .o1(_03284_));
 b15nano23as1n24x5 _29133_ (.a(net576),
    .b(net570),
    .c(\us23.a[6] ),
    .d(net578),
    .out0(_03285_));
 b15nand02al1n12x5 _29134_ (.a(net580),
    .b(_03285_),
    .o1(_03286_));
 b15nanb03an1n08x5 _29135_ (.a(net578),
    .b(net580),
    .c(net576),
    .out0(_03287_));
 b15orn002ar1n16x5 _29136_ (.a(_03071_),
    .b(_03287_),
    .o(_03288_));
 b15oai222as1n16x5 _29137_ (.a(_03205_),
    .b(_03282_),
    .c(_03284_),
    .d(_03286_),
    .e(_03288_),
    .f(_03075_),
    .o1(_03289_));
 b15nor002ah1n03x5 _29138_ (.a(net588),
    .b(_03217_),
    .o1(_03291_));
 b15oaoi13aq1n03x5 _29139_ (.a(_03289_),
    .b(_03291_),
    .c(_03227_),
    .d(_03137_),
    .o1(_03292_));
 b15nand04an1n06x5 _29140_ (.a(_03259_),
    .b(_03267_),
    .c(_03280_),
    .d(_03292_),
    .o1(_03293_));
 b15nano23al1n06x5 _29141_ (.a(_03116_),
    .b(_03185_),
    .c(_03239_),
    .d(_03293_),
    .out0(_03294_));
 b15nor004al1n04x5 _29142_ (.a(_02546_),
    .b(_02547_),
    .c(_02716_),
    .d(_02745_),
    .o1(_03295_));
 b15nor003ah1n04x5 _29143_ (.a(_02546_),
    .b(_02547_),
    .c(_02554_),
    .o1(_03296_));
 b15nor003an1n08x5 _29144_ (.a(net822),
    .b(_02654_),
    .c(_02656_),
    .o1(_03297_));
 b15oaoi13as1n04x5 _29145_ (.a(_03295_),
    .b(net840),
    .c(_03296_),
    .d(_03297_),
    .o1(_03298_));
 b15nona23aq1n24x5 _29146_ (.a(net827),
    .b(\us01.a[6] ),
    .c(net823),
    .d(\us01.a[4] ),
    .out0(_03299_));
 b15nanb02al1n08x5 _29147_ (.a(net839),
    .b(\us01.a[3] ),
    .out0(_03300_));
 b15nonb02ah1n06x5 _29148_ (.a(net827),
    .b(\us01.a[4] ),
    .out0(_03302_));
 b15nandp3al1n04x5 _29149_ (.a(net840),
    .b(_03302_),
    .c(_02580_),
    .o1(_03303_));
 b15oai022aq1n02x5 _29150_ (.a(_03299_),
    .b(_02695_),
    .c(_03300_),
    .d(_03303_),
    .o1(_03304_));
 b15inv020aq1n08x5 _29151_ (.a(net828),
    .o1(_03305_));
 b15obai22ar1n04x5 _29152_ (.a(_02577_),
    .b(net839),
    .c(_03305_),
    .d(_02609_),
    .out0(_03306_));
 b15nanb02an1n03x5 _29153_ (.a(\us01.a[6] ),
    .b(net840),
    .out0(_03307_));
 b15nonb03al1n04x5 _29154_ (.a(_03306_),
    .b(_03307_),
    .c(_02670_),
    .out0(_03308_));
 b15nonb02as1n08x5 _29155_ (.a(net831),
    .b(net839),
    .out0(_03309_));
 b15nand04an1n03x5 _29156_ (.a(net823),
    .b(_02517_),
    .c(_03309_),
    .d(_03307_),
    .o1(_03310_));
 b15norp03an1n16x5 _29157_ (.a(_02611_),
    .b(_02680_),
    .c(_02643_),
    .o1(_03311_));
 b15nonb02ar1n03x5 _29158_ (.a(net839),
    .b(net831),
    .out0(_03313_));
 b15aob012ar1n03x5 _29159_ (.a(_03310_),
    .b(_03311_),
    .c(_03313_),
    .out0(_03314_));
 b15oai013al1n06x5 _29160_ (.a(net834),
    .b(_03304_),
    .c(_03308_),
    .d(_03314_),
    .o1(_03315_));
 b15nor002aq1n02x5 _29161_ (.a(_02507_),
    .b(_02634_),
    .o1(_03316_));
 b15nand02aq1n12x5 _29162_ (.a(\us01.a[5] ),
    .b(net830),
    .o1(_03317_));
 b15oai012ar1n02x5 _29163_ (.a(_03317_),
    .b(_02610_),
    .c(net826),
    .o1(_03318_));
 b15nanb02al1n12x5 _29164_ (.a(net828),
    .b(net822),
    .out0(_03319_));
 b15norp03ar1n02x5 _29165_ (.a(net833),
    .b(_02671_),
    .c(_03319_),
    .o1(_03320_));
 b15aoi022as1n02x5 _29166_ (.a(_02677_),
    .b(_03316_),
    .c(_03318_),
    .d(_03320_),
    .o1(_03321_));
 b15nanb02as1n02x5 _29167_ (.a(net830),
    .b(net824),
    .out0(_03322_));
 b15norp02ar1n02x5 _29168_ (.a(\us01.a[5] ),
    .b(_03322_),
    .o1(_03324_));
 b15nonb02aq1n12x5 _29169_ (.a(net830),
    .b(net824),
    .out0(_03325_));
 b15ztpn00an1n08x5 TAP_478 ();
 b15aoi012an1n04x5 _29171_ (.a(_03324_),
    .b(_03325_),
    .c(\us01.a[5] ),
    .o1(_03327_));
 b15nandp2al1n08x5 _29172_ (.a(net829),
    .b(net822),
    .o1(_03328_));
 b15oai013aq1n12x5 _29173_ (.a(_03321_),
    .b(_03327_),
    .c(_03328_),
    .d(_02616_),
    .o1(_03329_));
 b15nanb02ah1n16x5 _29174_ (.a(net832),
    .b(net842),
    .out0(_03330_));
 b15oai022ar1n02x5 _29175_ (.a(_02515_),
    .b(_02654_),
    .c(_03330_),
    .d(_02583_),
    .o1(_03331_));
 b15nand02al1n12x5 _29176_ (.a(_02623_),
    .b(_02622_),
    .o1(_03332_));
 b15aoi112al1n03x5 _29177_ (.a(net834),
    .b(_02546_),
    .c(_03313_),
    .d(net840),
    .o1(_03333_));
 b15nonb02as1n06x5 _29178_ (.a(net832),
    .b(net842),
    .out0(_03335_));
 b15oai013ar1n02x5 _29179_ (.a(_02573_),
    .b(_02546_),
    .c(_02623_),
    .d(_03335_),
    .o1(_03336_));
 b15aoi013aq1n02x5 _29180_ (.a(_03331_),
    .b(_03332_),
    .c(_03333_),
    .d(_03336_),
    .o1(_03337_));
 b15oaoi13al1n03x5 _29181_ (.a(net838),
    .b(net832),
    .c(net835),
    .d(_02611_),
    .o1(_03338_));
 b15aoai13aq1n08x5 _29182_ (.a(_03338_),
    .b(_02637_),
    .c(_02635_),
    .d(net832),
    .o1(_03339_));
 b15nor002ah1n06x5 _29183_ (.a(net834),
    .b(_03299_),
    .o1(_03340_));
 b15nano23as1n24x5 _29184_ (.a(net822),
    .b(net825),
    .c(net826),
    .d(net828),
    .out0(_03341_));
 b15aoi012ar1n02x5 _29185_ (.a(_03340_),
    .b(_03341_),
    .c(net834),
    .o1(_03342_));
 b15oai112an1n06x5 _29186_ (.a(_03337_),
    .b(_03339_),
    .c(_03342_),
    .d(_03330_),
    .o1(_03343_));
 b15nano23ar1n08x5 _29187_ (.a(_03298_),
    .b(_03315_),
    .c(_03329_),
    .d(_03343_),
    .out0(_03344_));
 b15norp02aq1n04x5 _29188_ (.a(_02654_),
    .b(_02743_),
    .o1(_03346_));
 b15aoi012an1n02x5 _29189_ (.a(_02507_),
    .b(_02573_),
    .c(_03305_),
    .o1(_03347_));
 b15aoi013al1n04x5 _29190_ (.a(_03346_),
    .b(_03347_),
    .c(_02694_),
    .d(\us01.a[6] ),
    .o1(_03348_));
 b15nandp2al1n08x5 _29191_ (.a(net832),
    .b(_02541_),
    .o1(_03349_));
 b15oai112as1n02x5 _29192_ (.a(net842),
    .b(_03348_),
    .c(_03349_),
    .d(_02515_),
    .o1(_03350_));
 b15norp03ah1n08x5 _29193_ (.a(net832),
    .b(_02596_),
    .c(_02643_),
    .o1(_03351_));
 b15aob012as1n03x5 _29194_ (.a(_02611_),
    .b(_02541_),
    .c(_03351_),
    .out0(_03352_));
 b15nand02ar1n02x5 _29195_ (.a(net833),
    .b(_02620_),
    .o1(_03353_));
 b15oai112an1n04x5 _29196_ (.a(_02615_),
    .b(_03353_),
    .c(_02701_),
    .d(_03328_),
    .o1(_03354_));
 b15nanb02ah1n12x5 _29197_ (.a(net822),
    .b(net828),
    .out0(_03355_));
 b15oai112aq1n02x5 _29198_ (.a(net826),
    .b(_03319_),
    .c(_03355_),
    .d(_02569_),
    .o1(_03357_));
 b15and002ar1n08x5 _29199_ (.a(_03354_),
    .b(_03357_),
    .o(_03358_));
 b15aoai13ar1n08x5 _29200_ (.a(_03350_),
    .b(_03352_),
    .c(_03358_),
    .d(_03325_),
    .o1(_03359_));
 b15oai112al1n06x5 _29201_ (.a(_02631_),
    .b(_02768_),
    .c(_02593_),
    .d(net838),
    .o1(_03360_));
 b15ztpn00an1n08x5 TAP_477 ();
 b15nandp2ah1n16x5 _29203_ (.a(_02566_),
    .b(_02662_),
    .o1(_03362_));
 b15aoi012al1n02x5 _29204_ (.a(net842),
    .b(_02709_),
    .c(_03362_),
    .o1(_03363_));
 b15oai012ar1n04x5 _29205_ (.a(net835),
    .b(_02631_),
    .c(_02768_),
    .o1(_03364_));
 b15nand03ah1n06x5 _29206_ (.a(_03360_),
    .b(_03363_),
    .c(_03364_),
    .o1(_03365_));
 b15orn002ah1n16x5 _29207_ (.a(net838),
    .b(net835),
    .o(_03366_));
 b15oai012al1n04x5 _29208_ (.a(_03362_),
    .b(_02728_),
    .c(_03366_),
    .o1(_03368_));
 b15oai112ah1n08x5 _29209_ (.a(net830),
    .b(_03368_),
    .c(_02684_),
    .d(_02541_),
    .o1(_03369_));
 b15nor002aq1n32x5 _29210_ (.a(_02557_),
    .b(_02623_),
    .o1(_03370_));
 b15ztpn00an1n08x5 TAP_476 ();
 b15oai122ah1n12x5 _29212_ (.a(net832),
    .b(_02745_),
    .c(_03370_),
    .d(_02602_),
    .e(net842),
    .o1(_03372_));
 b15nor002ah1n16x5 _29213_ (.a(_02680_),
    .b(_02643_),
    .o1(_03373_));
 b15aoi012al1n04x5 _29214_ (.a(_03370_),
    .b(_03373_),
    .c(_03366_),
    .o1(_03374_));
 b15oai112as1n16x5 _29215_ (.a(_03365_),
    .b(_03369_),
    .c(_03372_),
    .d(_03374_),
    .o1(_03375_));
 b15xnr002as1n16x5 _29216_ (.a(net839),
    .b(net835),
    .out0(_03376_));
 b15oai012an1n02x5 _29217_ (.a(_03341_),
    .b(_03376_),
    .c(_02532_),
    .o1(_03377_));
 b15nand02ar1n24x5 _29218_ (.a(net841),
    .b(net836),
    .o1(_03379_));
 b15oai112aq1n04x5 _29219_ (.a(net832),
    .b(_03377_),
    .c(_03379_),
    .d(_02642_),
    .o1(_03380_));
 b15nanb03ar1n02x5 _29220_ (.a(\us01.a[6] ),
    .b(net841),
    .c(net829),
    .out0(_03381_));
 b15nanb02aq1n16x5 _29221_ (.a(net829),
    .b(net824),
    .out0(_03382_));
 b15oaoi13aq1n03x5 _29222_ (.a(_02681_),
    .b(_03381_),
    .c(_03382_),
    .d(_02665_),
    .o1(_03383_));
 b15norp03aq1n04x5 _29223_ (.a(net838),
    .b(_02595_),
    .c(_02596_),
    .o1(_03384_));
 b15oai013al1n02x5 _29224_ (.a(_02631_),
    .b(_02546_),
    .c(_02623_),
    .d(_02602_),
    .o1(_03385_));
 b15nor003ah1n03x5 _29225_ (.a(_03383_),
    .b(_03384_),
    .c(_03385_),
    .o1(_03386_));
 b15nor002ah1n04x5 _29226_ (.a(net834),
    .b(_02649_),
    .o1(_03387_));
 b15oai013ar1n02x5 _29227_ (.a(_03387_),
    .b(_03311_),
    .c(_03370_),
    .d(_02548_),
    .o1(_03388_));
 b15aob012ar1n08x5 _29228_ (.a(_03380_),
    .b(_03386_),
    .c(_03388_),
    .out0(_03390_));
 b15nonb02as1n16x5 _29229_ (.a(net834),
    .b(net830),
    .out0(_03391_));
 b15oai012ar1n02x5 _29230_ (.a(_02634_),
    .b(_02709_),
    .c(_03391_),
    .o1(_03392_));
 b15oaoi13al1n03x5 _29231_ (.a(_02743_),
    .b(_03392_),
    .c(_02716_),
    .d(_03379_),
    .o1(_03393_));
 b15ztpn00an1n08x5 TAP_475 ();
 b15nona23ah1n32x5 _29233_ (.a(\us01.a[5] ),
    .b(net829),
    .c(\us01.a[7] ),
    .d(net825),
    .out0(_03395_));
 b15norp02ah1n02x5 _29234_ (.a(_02507_),
    .b(_03395_),
    .o1(_03396_));
 b15nonb02an1n16x5 _29235_ (.a(net842),
    .b(net832),
    .out0(_03397_));
 b15aoi022aq1n02x5 _29236_ (.a(net826),
    .b(_02579_),
    .c(_02727_),
    .d(_03397_),
    .o1(_03398_));
 b15norp03ah1n03x5 _29237_ (.a(net834),
    .b(_02596_),
    .c(_03398_),
    .o1(_03399_));
 b15oaoi13an1n04x5 _29238_ (.a(_03393_),
    .b(net836),
    .c(_03396_),
    .d(_03399_),
    .o1(_03401_));
 b15nor002as1n04x5 _29239_ (.a(net824),
    .b(net839),
    .o1(_03402_));
 b15nanb02aq1n02x5 _29240_ (.a(_03319_),
    .b(_03402_),
    .out0(_03403_));
 b15nanb02an1n06x5 _29241_ (.a(net822),
    .b(net839),
    .out0(_03404_));
 b15and002ar1n02x5 _29242_ (.a(net824),
    .b(net833),
    .o(_03405_));
 b15aoi012ar1n06x5 _29243_ (.a(_03405_),
    .b(_02618_),
    .c(net828),
    .o1(_03406_));
 b15oaoi13as1n08x5 _29244_ (.a(_02615_),
    .b(_03403_),
    .c(_03404_),
    .d(_03406_),
    .o1(_03407_));
 b15aoai13ah1n08x5 _29245_ (.a(net831),
    .b(_03407_),
    .c(_02742_),
    .d(_02748_),
    .o1(_03408_));
 b15norp02ah1n12x5 _29246_ (.a(_02680_),
    .b(_02595_),
    .o1(_03409_));
 b15nandp3ar1n08x5 _29247_ (.a(_02631_),
    .b(_02742_),
    .c(_03409_),
    .o1(_03410_));
 b15nand04ah1n16x5 _29248_ (.a(_03390_),
    .b(_03401_),
    .c(_03408_),
    .d(_03410_),
    .o1(_03412_));
 b15nano23as1n24x5 _29249_ (.a(_03344_),
    .b(_03359_),
    .c(_03375_),
    .d(_03412_),
    .out0(_03413_));
 b15xnr002ar1n02x5 _29250_ (.a(net400),
    .b(_03413_),
    .out0(_03414_));
 b15xor002ar1n02x5 _29251_ (.a(_03034_),
    .b(_03414_),
    .out0(_03415_));
 b15xor002al1n02x5 _29252_ (.a(_02772_),
    .b(_03415_),
    .out0(_03416_));
 b15cmbn22aq1n02x5 _29253_ (.clk1(\text_in_r[64] ),
    .clk2(_03416_),
    .clkout(_03417_),
    .s(net538));
 b15xor002ar1n06x5 _29254_ (.a(\u0.w[1][0] ),
    .b(_03417_),
    .out0(_00105_));
 b15inv020ah1n04x5 _29255_ (.a(\text_in_r[65] ),
    .o1(_03418_));
 b15ztpn00an1n08x5 TAP_474 ();
 b15ztpn00an1n08x5 TAP_473 ();
 b15oai122ar1n04x5 _29258_ (.a(_02951_),
    .b(_02986_),
    .c(_02787_),
    .d(_02862_),
    .e(_02882_),
    .o1(_03422_));
 b15ztpn00an1n08x5 TAP_472 ();
 b15nona23as1n12x5 _29260_ (.a(\us30.a[5] ),
    .b(net844),
    .c(\us30.a[7] ),
    .d(\us30.a[4] ),
    .out0(_03424_));
 b15oai122ah1n04x5 _29261_ (.a(net858),
    .b(_02787_),
    .c(_02929_),
    .d(_03424_),
    .e(_02864_),
    .o1(_03425_));
 b15ztpn00an1n08x5 TAP_471 ();
 b15nand03al1n24x5 _29263_ (.a(_02854_),
    .b(_02899_),
    .c(_02781_),
    .o1(_03427_));
 b15oai022ar1n02x5 _29264_ (.a(_02854_),
    .b(_03028_),
    .c(_03427_),
    .d(_02837_),
    .o1(_03428_));
 b15aoi022ar1n02x5 _29265_ (.a(_03422_),
    .b(_03425_),
    .c(_03428_),
    .d(_02811_),
    .o1(_03429_));
 b15aoai13ar1n02x5 _29266_ (.a(net856),
    .b(_02811_),
    .c(_03018_),
    .d(_02877_),
    .o1(_03430_));
 b15norp02an1n02x5 _29267_ (.a(\us30.a[1] ),
    .b(\us30.a[4] ),
    .o1(_03431_));
 b15aoi013aq1n02x5 _29268_ (.a(net852),
    .b(\us30.a[5] ),
    .c(_02920_),
    .d(_03431_),
    .o1(_03433_));
 b15nandp3ar1n02x5 _29269_ (.a(_02897_),
    .b(_02831_),
    .c(_02877_),
    .o1(_03434_));
 b15aoi012an1n02x5 _29270_ (.a(_03430_),
    .b(_03433_),
    .c(_03434_),
    .o1(_03435_));
 b15ztpn00an1n08x5 TAP_470 ();
 b15ztpn00an1n08x5 TAP_469 ();
 b15ztpn00an1n08x5 TAP_468 ();
 b15aoai13ar1n03x5 _29274_ (.a(_02964_),
    .b(net862),
    .c(_02984_),
    .d(_03029_),
    .o1(_03439_));
 b15aoi013an1n04x5 _29275_ (.a(_03435_),
    .b(_03439_),
    .c(_02791_),
    .d(_02923_),
    .o1(_03440_));
 b15nand03an1n04x5 _29276_ (.a(_02811_),
    .b(_02782_),
    .c(_02911_),
    .o1(_03441_));
 b15nand04aq1n04x5 _29277_ (.a(net858),
    .b(_02867_),
    .c(_02858_),
    .d(_03018_),
    .o1(_03442_));
 b15xnr002ah1n06x5 _29278_ (.a(net858),
    .b(net860),
    .out0(_03444_));
 b15nanb02al1n04x5 _29279_ (.a(_02942_),
    .b(_03444_),
    .out0(_03445_));
 b15aoi013aq1n06x5 _29280_ (.a(net855),
    .b(_03441_),
    .c(_03442_),
    .d(_03445_),
    .o1(_03446_));
 b15orn002al1n08x5 _29281_ (.a(net860),
    .b(net851),
    .o(_03447_));
 b15nandp2ar1n03x5 _29282_ (.a(_02943_),
    .b(_02974_),
    .o1(_03448_));
 b15oaoi13ah1n02x5 _29283_ (.a(_03447_),
    .b(_03448_),
    .c(_02913_),
    .d(_02933_),
    .o1(_03449_));
 b15nano23an1n05x5 _29284_ (.a(_03429_),
    .b(_03440_),
    .c(_03446_),
    .d(_03449_),
    .out0(_03450_));
 b15oaoi13ar1n02x5 _29285_ (.a(net858),
    .b(_02997_),
    .c(_02964_),
    .d(net860),
    .o1(_03451_));
 b15nor004as1n12x5 _29286_ (.a(net846),
    .b(net848),
    .c(net843),
    .d(\us30.a[6] ),
    .o1(_03452_));
 b15nandp2al1n02x5 _29287_ (.a(net858),
    .b(_03452_),
    .o1(_03453_));
 b15aoi012ar1n02x5 _29288_ (.a(net860),
    .b(_02984_),
    .c(_03453_),
    .o1(_03455_));
 b15oab012aq1n04x5 _29289_ (.a(_02864_),
    .b(_03451_),
    .c(_03455_),
    .out0(_03456_));
 b15nand02an1n04x5 _29290_ (.a(net858),
    .b(_02882_),
    .o1(_03457_));
 b15oai122as1n04x5 _29291_ (.a(_02782_),
    .b(_02788_),
    .c(_03457_),
    .d(_02791_),
    .e(net858),
    .o1(_03458_));
 b15nor003ah1n02x5 _29292_ (.a(_02879_),
    .b(_02880_),
    .c(_02882_),
    .o1(_03459_));
 b15norp02ah1n32x5 _29293_ (.a(net861),
    .b(net854),
    .o1(_03460_));
 b15oai012ah1n08x5 _29294_ (.a(_02882_),
    .b(_03460_),
    .c(net857),
    .o1(_03461_));
 b15aoai13aq1n08x5 _29295_ (.a(net850),
    .b(_03459_),
    .c(_03461_),
    .d(_02908_),
    .o1(_03462_));
 b15nandp2aq1n16x5 _29296_ (.a(net853),
    .b(_02932_),
    .o1(_03463_));
 b15oai112as1n06x5 _29297_ (.a(_03458_),
    .b(_03462_),
    .c(_03463_),
    .d(_02956_),
    .o1(_03464_));
 b15nor002aq1n03x5 _29298_ (.a(_02811_),
    .b(_03020_),
    .o1(_03466_));
 b15nor003al1n12x5 _29299_ (.a(_02794_),
    .b(_02798_),
    .c(_02882_),
    .o1(_03467_));
 b15aoi022an1n08x5 _29300_ (.a(_03466_),
    .b(_02898_),
    .c(_03467_),
    .d(_02811_),
    .o1(_03468_));
 b15norp02aq1n24x5 _29301_ (.a(net851),
    .b(net853),
    .o1(_03469_));
 b15nor002an1n08x5 _29302_ (.a(net860),
    .b(_02862_),
    .o1(_03470_));
 b15oai112an1n12x5 _29303_ (.a(_03469_),
    .b(_02923_),
    .c(_02932_),
    .d(_03470_),
    .o1(_03471_));
 b15oai022ar1n02x5 _29304_ (.a(_02858_),
    .b(_03424_),
    .c(_03029_),
    .d(_02867_),
    .o1(_03472_));
 b15nandp2ar1n03x5 _29305_ (.a(_02989_),
    .b(_03472_),
    .o1(_03473_));
 b15nand03ar1n04x5 _29306_ (.a(_03468_),
    .b(_03471_),
    .c(_03473_),
    .o1(_03474_));
 b15oaoi13ar1n03x5 _29307_ (.a(_02873_),
    .b(_02862_),
    .c(_02879_),
    .d(_02880_),
    .o1(_03475_));
 b15nandp2al1n03x5 _29308_ (.a(net861),
    .b(_02862_),
    .o1(_03477_));
 b15oai012an1n04x5 _29309_ (.a(_02820_),
    .b(_02879_),
    .c(_02880_),
    .o1(_03478_));
 b15aoai13as1n06x5 _29310_ (.a(_03475_),
    .b(net857),
    .c(_03477_),
    .d(_03478_),
    .o1(_03479_));
 b15ztpn00an1n08x5 TAP_467 ();
 b15aoi012al1n02x5 _29312_ (.a(_02811_),
    .b(net855),
    .c(_03444_),
    .o1(_03481_));
 b15nanb02al1n24x5 _29313_ (.a(net846),
    .b(net849),
    .out0(_03482_));
 b15qgbno2an1n10x5 _29314_ (.a(_02880_),
    .b(_03482_),
    .o1(_03483_));
 b15ztpn00an1n08x5 TAP_466 ();
 b15aoai13ar1n06x5 _29316_ (.a(_03481_),
    .b(_03483_),
    .c(_02782_),
    .d(net855),
    .o1(_03485_));
 b15nand03an1n03x5 _29317_ (.a(_02904_),
    .b(_02947_),
    .c(_03000_),
    .o1(_03486_));
 b15norp03ar1n02x5 _29318_ (.a(_02787_),
    .b(_03020_),
    .c(_03029_),
    .o1(_03488_));
 b15oab012al1n02x5 _29319_ (.a(_03488_),
    .b(_02892_),
    .c(_02954_),
    .out0(_03489_));
 b15nand04an1n08x5 _29320_ (.a(_03479_),
    .b(_03485_),
    .c(_03486_),
    .d(_03489_),
    .o1(_03490_));
 b15nor004as1n06x5 _29321_ (.a(_03456_),
    .b(_03464_),
    .c(_03474_),
    .d(_03490_),
    .o1(_03491_));
 b15ztpn00an1n08x5 TAP_465 ();
 b15norp02ar1n02x5 _29323_ (.a(_02862_),
    .b(_02935_),
    .o1(_03493_));
 b15aoi112aq1n03x5 _29324_ (.a(net852),
    .b(_03493_),
    .c(_02989_),
    .d(_02898_),
    .o1(_03494_));
 b15ztpn00an1n08x5 TAP_464 ();
 b15nor004al1n03x5 _29326_ (.a(_02951_),
    .b(net856),
    .c(_02794_),
    .d(_02798_),
    .o1(_03496_));
 b15norp03an1n02x5 _29327_ (.a(net859),
    .b(net856),
    .c(_02997_),
    .o1(_03497_));
 b15oai012ah1n04x5 _29328_ (.a(net862),
    .b(_03496_),
    .c(_03497_),
    .o1(_03499_));
 b15nand02as1n06x5 _29329_ (.a(net856),
    .b(net846),
    .o1(_03500_));
 b15norp02ar1n02x5 _29330_ (.a(net843),
    .b(_03500_),
    .o1(_03501_));
 b15ztpn00an1n08x5 TAP_463 ();
 b15nandp3ar1n02x5 _29332_ (.a(net862),
    .b(net849),
    .c(net845),
    .o1(_03503_));
 b15orn003ar1n02x5 _29333_ (.a(net862),
    .b(net849),
    .c(net845),
    .o(_03504_));
 b15aoi012ar1n02x5 _29334_ (.a(net859),
    .b(_03503_),
    .c(_03504_),
    .o1(_03505_));
 b15aoai13aq1n04x5 _29335_ (.a(_03501_),
    .b(_03505_),
    .c(_02877_),
    .d(net845),
    .o1(_03506_));
 b15ztpn00an1n08x5 TAP_462 ();
 b15ztpn00an1n08x5 TAP_461 ();
 b15aoi013al1n06x5 _29338_ (.a(_03494_),
    .b(_03499_),
    .c(_03506_),
    .d(net852),
    .o1(_03510_));
 b15nand02an1n02x5 _29339_ (.a(net862),
    .b(net847),
    .o1(_03511_));
 b15nand02ar1n02x5 _29340_ (.a(_02820_),
    .b(net848),
    .o1(_03512_));
 b15aoi112al1n02x5 _29341_ (.a(_02956_),
    .b(_02880_),
    .c(_03511_),
    .d(_03512_),
    .o1(_03513_));
 b15nandp2al1n24x5 _29342_ (.a(\us30.a[0] ),
    .b(net852),
    .o1(_03514_));
 b15oai022ar1n02x5 _29343_ (.a(_02954_),
    .b(_02923_),
    .c(_02984_),
    .d(_03514_),
    .o1(_03515_));
 b15nandp3ar1n08x5 _29344_ (.a(net862),
    .b(net850),
    .c(_03024_),
    .o1(_03516_));
 b15nona22ah1n04x5 _29345_ (.a(_03513_),
    .b(_03515_),
    .c(_03516_),
    .out0(_03517_));
 b15ztpn00an1n08x5 TAP_460 ();
 b15nandp3ar1n24x5 _29347_ (.a(_02811_),
    .b(_02831_),
    .c(_02833_),
    .o1(_03519_));
 b15qbfna2bn1n16x5 _29348_ (.a(net852),
    .b(_03024_),
    .o1(_03521_));
 b15orn002ah1n03x5 _29349_ (.a(net843),
    .b(net845),
    .o(_03522_));
 b15nor002as1n04x5 _29350_ (.a(_03522_),
    .b(_02879_),
    .o1(_03523_));
 b15norp02as1n16x5 _29351_ (.a(net861),
    .b(net850),
    .o1(_03524_));
 b15aoi022aq1n02x5 _29352_ (.a(net861),
    .b(_03523_),
    .c(_02881_),
    .d(_03524_),
    .o1(_03525_));
 b15aoi013as1n03x5 _29353_ (.a(net857),
    .b(_03519_),
    .c(_03521_),
    .d(_03525_),
    .o1(_03526_));
 b15oaoi13as1n08x5 _29354_ (.a(_03510_),
    .b(_02854_),
    .c(_03517_),
    .d(_03526_),
    .o1(_03527_));
 b15aoi112ar1n02x5 _29355_ (.a(_02811_),
    .b(net855),
    .c(_02950_),
    .d(_02918_),
    .o1(_03528_));
 b15oai112ar1n02x5 _29356_ (.a(_02831_),
    .b(_02844_),
    .c(_02915_),
    .d(_02833_),
    .o1(_03529_));
 b15ztpn00an1n08x5 TAP_459 ();
 b15oaoi13ar1n02x5 _29358_ (.a(_02854_),
    .b(_03529_),
    .c(_02892_),
    .d(_02876_),
    .o1(_03532_));
 b15oai012ar1n02x5 _29359_ (.a(net862),
    .b(_03528_),
    .c(_03532_),
    .o1(_03533_));
 b15oai122as1n04x5 _29360_ (.a(_02820_),
    .b(_02876_),
    .c(_02995_),
    .d(_03029_),
    .e(_02951_),
    .o1(_03534_));
 b15qgbno2an1n05x5 _29361_ (.o1(_03535_),
    .a(net853),
    .b(_03029_));
 b15oai112ah1n06x5 _29362_ (.a(\us30.a[3] ),
    .b(_03534_),
    .c(_03535_),
    .d(_02820_),
    .o1(_03536_));
 b15nand03al1n03x5 _29363_ (.a(net858),
    .b(_03469_),
    .c(_03452_),
    .o1(_03537_));
 b15oai013al1n06x5 _29364_ (.a(_03537_),
    .b(_02921_),
    .c(_03020_),
    .d(_02940_),
    .o1(_03538_));
 b15oaoi13ah1n03x5 _29365_ (.a(_02876_),
    .b(_02948_),
    .c(net858),
    .d(_02864_),
    .o1(_03539_));
 b15oai022an1n06x5 _29366_ (.a(_02787_),
    .b(_02876_),
    .c(_03514_),
    .d(_03463_),
    .o1(_03540_));
 b15aoi112aq1n08x5 _29367_ (.a(_03538_),
    .b(_03539_),
    .c(_03540_),
    .d(net858),
    .o1(_03541_));
 b15and003aq1n03x5 _29368_ (.a(_03533_),
    .b(_03536_),
    .c(_03541_),
    .o(_03543_));
 b15nand04as1n16x5 _29369_ (.a(_03450_),
    .b(_03491_),
    .c(_03527_),
    .d(_03543_),
    .o1(_03544_));
 b15norp03ar1n02x5 _29370_ (.a(_02569_),
    .b(_03379_),
    .c(_02743_),
    .o1(_03545_));
 b15aoi013al1n03x5 _29371_ (.a(_03545_),
    .b(_03373_),
    .c(_03397_),
    .d(_02569_),
    .o1(_03546_));
 b15norp02as1n03x5 _29372_ (.a(net834),
    .b(_02593_),
    .o1(_03547_));
 b15oai122as1n16x5 _29373_ (.a(net831),
    .b(_02761_),
    .c(_03547_),
    .d(_03376_),
    .e(net842),
    .o1(_03548_));
 b15nanb02as1n24x5 _29374_ (.a(net838),
    .b(net835),
    .out0(_03549_));
 b15oai022al1n06x5 _29375_ (.a(net841),
    .b(_03549_),
    .c(_03373_),
    .d(_02631_),
    .o1(_03550_));
 b15aob012ar1n02x5 _29376_ (.a(net841),
    .b(net832),
    .c(_02602_),
    .out0(_03551_));
 b15oai012ah1n04x5 _29377_ (.a(_03551_),
    .b(_02598_),
    .c(net832),
    .o1(_03552_));
 b15oai112aq1n12x5 _29378_ (.a(_03546_),
    .b(_03548_),
    .c(_03550_),
    .d(_03552_),
    .o1(_03554_));
 b15ztpn00an1n08x5 TAP_458 ();
 b15oai013ar1n02x5 _29380_ (.a(_03395_),
    .b(_02596_),
    .c(_02665_),
    .d(_02595_),
    .o1(_03556_));
 b15nand03ah1n02x5 _29381_ (.a(net832),
    .b(_02645_),
    .c(_03556_),
    .o1(_03557_));
 b15ztpn00an1n08x5 TAP_457 ();
 b15oai022al1n02x5 _29383_ (.a(net836),
    .b(_02598_),
    .c(_03341_),
    .d(_02602_),
    .o1(_03559_));
 b15aoi012ah1n04x5 _29384_ (.a(_03557_),
    .b(_03559_),
    .c(net841),
    .o1(_03560_));
 b15aoi022ah1n12x5 _29385_ (.a(_02759_),
    .b(_02745_),
    .c(_02748_),
    .d(_02526_),
    .o1(_03561_));
 b15nandp2ah1n08x5 _29386_ (.a(_03391_),
    .b(_03379_),
    .o1(_03562_));
 b15inv040an1n06x5 _29387_ (.a(net825),
    .o1(_03563_));
 b15nandp2ar1n12x5 _29388_ (.a(_03563_),
    .b(_02620_),
    .o1(_03565_));
 b15oai022ar1n32x5 _29389_ (.a(_02654_),
    .b(_03561_),
    .c(_03562_),
    .d(_03565_),
    .o1(_03566_));
 b15norp02ar1n02x5 _29390_ (.a(_02631_),
    .b(_02692_),
    .o1(_03567_));
 b15nona22ar1n02x5 _29391_ (.a(\us01.a[7] ),
    .b(net834),
    .c(\us01.a[5] ),
    .out0(_03568_));
 b15orn002an1n02x5 _29392_ (.a(net824),
    .b(net830),
    .o(_03569_));
 b15nanb02ar1n02x5 _29393_ (.a(net841),
    .b(net829),
    .out0(_03570_));
 b15oaoi13an1n03x5 _29394_ (.a(_03568_),
    .b(_03569_),
    .c(_02648_),
    .d(_03570_),
    .o1(_03571_));
 b15ztpn00an1n08x5 TAP_456 ();
 b15norp03ar1n16x5 _29396_ (.a(_02507_),
    .b(_02557_),
    .c(_02547_),
    .o1(_03573_));
 b15oai013as1n03x5 _29397_ (.a(net836),
    .b(_03567_),
    .c(_03571_),
    .d(_03573_),
    .o1(_03574_));
 b15orn002ar1n04x5 _29398_ (.a(\us01.a[5] ),
    .b(net830),
    .o(_03576_));
 b15nonb02as1n16x5 _29399_ (.a(net838),
    .b(net835),
    .out0(_03577_));
 b15oai012aq1n02x5 _29400_ (.a(net836),
    .b(_02643_),
    .c(_02611_),
    .o1(_03578_));
 b15ztpn00an1n08x5 TAP_455 ();
 b15aoi022al1n06x5 _29402_ (.a(_02611_),
    .b(_03577_),
    .c(_03578_),
    .d(net834),
    .o1(_03580_));
 b15oai013aq1n08x5 _29403_ (.a(_03574_),
    .b(_03576_),
    .c(_03580_),
    .d(_02596_),
    .o1(_03581_));
 b15nor004as1n12x5 _29404_ (.a(_03554_),
    .b(_03560_),
    .c(_03566_),
    .d(_03581_),
    .o1(_03582_));
 b15nand02an1n12x5 _29405_ (.a(_03302_),
    .b(_02580_),
    .o1(_03583_));
 b15oai122al1n02x5 _29406_ (.a(_02611_),
    .b(_02583_),
    .c(_02716_),
    .d(_02654_),
    .e(_03583_),
    .o1(_03584_));
 b15oai022ar1n02x5 _29407_ (.a(net832),
    .b(_02583_),
    .c(_03362_),
    .d(_03349_),
    .o1(_03585_));
 b15oai012al1n02x5 _29408_ (.a(_03584_),
    .b(_03585_),
    .c(_02611_),
    .o1(_03587_));
 b15oai012an1n02x5 _29409_ (.a(_02684_),
    .b(_02768_),
    .c(net838),
    .o1(_03588_));
 b15nor002ar1n02x5 _29410_ (.a(_02768_),
    .b(_03335_),
    .o1(_03589_));
 b15oai112ar1n08x5 _29411_ (.a(_02669_),
    .b(_03588_),
    .c(_03589_),
    .d(_03370_),
    .o1(_03590_));
 b15aoi112ar1n06x5 _29412_ (.a(_03309_),
    .b(_03590_),
    .c(_02541_),
    .d(_02700_),
    .o1(_03591_));
 b15nano23aq1n24x5 _29413_ (.a(\us01.a[4] ),
    .b(\us01.a[6] ),
    .c(net823),
    .d(net827),
    .out0(_03592_));
 b15nand02ar1n02x5 _29414_ (.a(net831),
    .b(_03592_),
    .o1(_03593_));
 b15oaoi13ar1n02x5 _29415_ (.a(_02569_),
    .b(_03593_),
    .c(_03362_),
    .d(net831),
    .o1(_03594_));
 b15oab012ar1n04x5 _29416_ (.a(_02745_),
    .b(_03346_),
    .c(_03594_),
    .out0(_03595_));
 b15nano23ah1n06x5 _29417_ (.a(_03298_),
    .b(_03587_),
    .c(_03591_),
    .d(_03595_),
    .out0(_03596_));
 b15nano23as1n16x5 _29418_ (.a(net827),
    .b(net823),
    .c(\us01.a[6] ),
    .d(\us01.a[4] ),
    .out0(_03598_));
 b15aoi222aq1n02x5 _29419_ (.a(_02517_),
    .b(_02529_),
    .c(_03577_),
    .d(_03341_),
    .e(_03598_),
    .f(_02573_),
    .o1(_03599_));
 b15ztpn00an1n08x5 TAP_454 ();
 b15oai022aq1n04x5 _29421_ (.a(net835),
    .b(_02583_),
    .c(_03599_),
    .d(\us01.a[3] ),
    .o1(_03601_));
 b15nano23as1n24x5 _29422_ (.a(net827),
    .b(\us01.a[4] ),
    .c(net823),
    .d(\us01.a[6] ),
    .out0(_03602_));
 b15oai012ar1n03x5 _29423_ (.a(_02709_),
    .b(_02548_),
    .c(_03602_),
    .o1(_03603_));
 b15nand03al1n03x5 _29424_ (.a(net842),
    .b(_02709_),
    .c(_02757_),
    .o1(_03604_));
 b15nand02as1n16x5 _29425_ (.a(_02566_),
    .b(_02727_),
    .o1(_03605_));
 b15oai112an1n06x5 _29426_ (.a(_03603_),
    .b(_03604_),
    .c(_03330_),
    .d(_03605_),
    .o1(_03606_));
 b15aoi022an1n08x5 _29427_ (.a(net842),
    .b(_03601_),
    .c(_03606_),
    .d(_02573_),
    .o1(_03607_));
 b15norp02ar1n02x5 _29428_ (.a(_02631_),
    .b(_02748_),
    .o1(_03609_));
 b15aoi013ar1n02x5 _29429_ (.a(\us01.a[3] ),
    .b(_03302_),
    .c(_02529_),
    .d(_02562_),
    .o1(_03610_));
 b15nandp3ar1n02x5 _29430_ (.a(_02611_),
    .b(_02566_),
    .c(_02727_),
    .o1(_03611_));
 b15nand02ar1n02x5 _29431_ (.a(net840),
    .b(_03341_),
    .o1(_03612_));
 b15aoi013aq1n02x5 _29432_ (.a(_03609_),
    .b(_03610_),
    .c(_03611_),
    .d(_03612_),
    .o1(_03613_));
 b15nandp3ar1n02x5 _29433_ (.a(_02611_),
    .b(_02759_),
    .c(_03300_),
    .o1(_03614_));
 b15oai112aq1n02x5 _29434_ (.a(net835),
    .b(_03614_),
    .c(_03300_),
    .d(_02583_),
    .o1(_03615_));
 b15aoi122as1n02x5 _29435_ (.a(\us01.a[3] ),
    .b(_02665_),
    .c(_03341_),
    .d(_03598_),
    .e(net838),
    .o1(_03616_));
 b15qgbna2an1n05x5 _29436_ (.o1(_03617_),
    .a(net839),
    .b(_02759_));
 b15nandp3ar1n02x5 _29437_ (.a(_02611_),
    .b(_03302_),
    .c(_02529_),
    .o1(_03618_));
 b15aoi013ar1n02x5 _29438_ (.a(_03616_),
    .b(_03617_),
    .c(_03618_),
    .d(\us01.a[3] ),
    .o1(_03620_));
 b15oa0022ar1n06x5 _29439_ (.a(_03613_),
    .b(_03615_),
    .c(_03620_),
    .d(net835),
    .o(_03621_));
 b15oai013an1n02x5 _29440_ (.a(_03577_),
    .b(_02645_),
    .c(_02547_),
    .d(_02557_),
    .o1(_03622_));
 b15oai112an1n06x5 _29441_ (.a(\us01.a[7] ),
    .b(_03622_),
    .c(_02635_),
    .d(net836),
    .o1(_03623_));
 b15aoi022ah1n06x5 _29442_ (.a(net829),
    .b(_02646_),
    .c(_02684_),
    .d(_03382_),
    .o1(_03624_));
 b15oaoi13as1n08x5 _29443_ (.a(_03623_),
    .b(_02656_),
    .c(net826),
    .d(_03624_),
    .o1(_03625_));
 b15nor002al1n32x5 _29444_ (.a(\us01.a[0] ),
    .b(\us01.a[2] ),
    .o1(_03626_));
 b15aoai13ah1n02x5 _29445_ (.a(_03626_),
    .b(_03592_),
    .c(_02757_),
    .d(net838),
    .o1(_03627_));
 b15nor002an1n03x5 _29446_ (.a(net835),
    .b(_02743_),
    .o1(_03628_));
 b15oab012an1n02x5 _29447_ (.a(_03628_),
    .b(_02545_),
    .c(_02642_),
    .out0(_03629_));
 b15oai012ar1n08x5 _29448_ (.a(_03627_),
    .b(_03629_),
    .c(net838),
    .o1(_03631_));
 b15oaoi13ar1n08x5 _29449_ (.a(_03621_),
    .b(\us01.a[3] ),
    .c(_03625_),
    .d(_03631_),
    .o1(_03632_));
 b15nand04as1n16x5 _29450_ (.a(_03582_),
    .b(_03596_),
    .c(_03607_),
    .d(_03632_),
    .o1(_03633_));
 b15xor002an1n04x5 _29451_ (.a(_03544_),
    .b(_03633_),
    .out0(_03634_));
 b15oai112ar1n02x5 _29452_ (.a(net696),
    .b(_02365_),
    .c(net713),
    .d(net699),
    .o1(_03635_));
 b15nand02al1n16x5 _29453_ (.a(net711),
    .b(net708),
    .o1(_03636_));
 b15oai022ar1n02x5 _29454_ (.a(_02407_),
    .b(_02444_),
    .c(_03635_),
    .d(_03636_),
    .o1(_03637_));
 b15nandp2an1n05x5 _29455_ (.a(net702),
    .b(_03637_),
    .o1(_03638_));
 b15ztpn00an1n08x5 TAP_453 ();
 b15nandp3an1n04x5 _29457_ (.a(net711),
    .b(net707),
    .c(_02376_),
    .o1(_03640_));
 b15nandp3aq1n08x5 _29458_ (.a(net703),
    .b(_02365_),
    .c(_02346_),
    .o1(_03642_));
 b15oaoi13an1n08x5 _29459_ (.a(net713),
    .b(_03640_),
    .c(_03642_),
    .d(net711),
    .o1(_03643_));
 b15xnr002as1n16x5 _29460_ (.a(\us12.a[1] ),
    .b(\us12.a[2] ),
    .out0(_03644_));
 b15and002al1n08x5 _29461_ (.a(net714),
    .b(net701),
    .o(_03645_));
 b15nand04ar1n12x5 _29462_ (.a(_02430_),
    .b(_02291_),
    .c(_03644_),
    .d(_03645_),
    .o1(_03646_));
 b15nand04as1n06x5 _29463_ (.a(_02341_),
    .b(_02343_),
    .c(_02346_),
    .d(_02390_),
    .o1(_03647_));
 b15nanb02as1n24x5 _29464_ (.a(net697),
    .b(net700),
    .out0(_03648_));
 b15nanb03ar1n02x5 _29465_ (.a(net694),
    .b(net712),
    .c(net701),
    .out0(_03649_));
 b15oa0022as1n03x5 _29466_ (.a(_02279_),
    .b(_02310_),
    .c(_03648_),
    .d(_03649_),
    .o(_03650_));
 b15nandp2ah1n16x5 _29467_ (.a(net713),
    .b(net706),
    .o1(_03651_));
 b15nand03as1n04x5 _29468_ (.a(_02276_),
    .b(_02325_),
    .c(_03651_),
    .o1(_03653_));
 b15oai112as1n16x5 _29469_ (.a(_03646_),
    .b(_03647_),
    .c(_03650_),
    .d(_03653_),
    .o1(_03654_));
 b15and002al1n04x5 _29470_ (.a(net713),
    .b(net707),
    .o(_03655_));
 b15nand04an1n08x5 _29471_ (.a(net703),
    .b(_02293_),
    .c(_02437_),
    .d(_03655_),
    .o1(_03656_));
 b15nanb02as1n24x5 _29472_ (.a(\us12.a[0] ),
    .b(\us12.a[1] ),
    .out0(_03657_));
 b15ztpn00an1n08x5 TAP_452 ();
 b15nandp3aq1n08x5 _29474_ (.a(net702),
    .b(_02293_),
    .c(_02437_),
    .o1(_03659_));
 b15nandp3ah1n04x5 _29475_ (.a(_02343_),
    .b(_02430_),
    .c(_02437_),
    .o1(_03660_));
 b15aoai13ah1n06x5 _29476_ (.a(_03656_),
    .b(_03657_),
    .c(_03659_),
    .d(_03660_),
    .o1(_03661_));
 b15nandp2an1n05x5 _29477_ (.a(_02381_),
    .b(_02425_),
    .o1(_03662_));
 b15oaoi13ah1n02x5 _29478_ (.a(_02355_),
    .b(_03662_),
    .c(_02499_),
    .d(_02381_),
    .o1(_03664_));
 b15nor004aq1n06x5 _29479_ (.a(_03643_),
    .b(_03654_),
    .c(_03661_),
    .d(_03664_),
    .o1(_03665_));
 b15nand02an1n32x5 _29480_ (.a(_02341_),
    .b(_02333_),
    .o1(_03666_));
 b15nandp2an1n12x5 _29481_ (.a(net709),
    .b(_02321_),
    .o1(_03667_));
 b15aoi112ah1n02x5 _29482_ (.a(net703),
    .b(_03666_),
    .c(_02444_),
    .d(_03667_),
    .o1(_03668_));
 b15ztpn00an1n08x5 TAP_451 ();
 b15norp03aq1n24x5 _29484_ (.a(net696),
    .b(net699),
    .c(net691),
    .o1(_03670_));
 b15aoi022ar1n02x5 _29485_ (.a(_02242_),
    .b(_03670_),
    .c(_02395_),
    .d(_02475_),
    .o1(_03671_));
 b15nor002aq1n02x5 _29486_ (.a(_02320_),
    .b(_03671_),
    .o1(_03672_));
 b15nona23aq1n24x5 _29487_ (.a(net696),
    .b(net691),
    .c(net694),
    .d(net699),
    .out0(_03673_));
 b15oai022al1n06x5 _29488_ (.a(_03667_),
    .b(_02438_),
    .c(_03673_),
    .d(_02444_),
    .o1(_03675_));
 b15aoi112aq1n06x5 _29489_ (.a(_03668_),
    .b(_03672_),
    .c(net703),
    .d(_03675_),
    .o1(_03676_));
 b15nona23as1n32x5 _29490_ (.a(net697),
    .b(net700),
    .c(net692),
    .d(net695),
    .out0(_03677_));
 b15nand03an1n02x5 _29491_ (.a(_02320_),
    .b(_02433_),
    .c(_02357_),
    .o1(_03678_));
 b15nonb02as1n08x5 _29492_ (.a(net705),
    .b(net709),
    .out0(_03679_));
 b15nor002as1n04x5 _29493_ (.a(_02343_),
    .b(_03679_),
    .o1(_03680_));
 b15oaoi13al1n04x5 _29494_ (.a(_03677_),
    .b(_03678_),
    .c(_03680_),
    .d(_02390_),
    .o1(_03681_));
 b15ztpn00an1n08x5 TAP_450 ();
 b15oai022an1n02x5 _29496_ (.a(_03677_),
    .b(_02389_),
    .c(_03662_),
    .d(net709),
    .o1(_03683_));
 b15ztpn00an1n08x5 TAP_449 ();
 b15aoi012aq1n04x5 _29498_ (.a(_03681_),
    .b(_03683_),
    .c(net710),
    .o1(_03686_));
 b15nand04ah1n16x5 _29499_ (.a(_03638_),
    .b(_03665_),
    .c(_03676_),
    .d(_03686_),
    .o1(_03687_));
 b15norp02ar1n12x5 _29500_ (.a(_02309_),
    .b(_03648_),
    .o1(_03688_));
 b15nor002ah1n06x5 _29501_ (.a(_03657_),
    .b(_02357_),
    .o1(_03689_));
 b15nor004ar1n02x5 _29502_ (.a(net703),
    .b(_02309_),
    .c(_02300_),
    .d(_03648_),
    .o1(_03690_));
 b15oai022ar1n02x5 _29503_ (.a(_02319_),
    .b(_03688_),
    .c(_03689_),
    .d(_03690_),
    .o1(_03691_));
 b15norp02al1n03x5 _29504_ (.a(net695),
    .b(_02324_),
    .o1(_03692_));
 b15aoi022ar1n02x5 _29505_ (.a(_02367_),
    .b(_02403_),
    .c(_02491_),
    .d(_03692_),
    .o1(_03693_));
 b15oai013ar1n02x5 _29506_ (.a(_03691_),
    .b(_03693_),
    .c(_03657_),
    .d(net700),
    .o1(_03694_));
 b15nandp2an1n24x5 _29507_ (.a(net698),
    .b(\us12.a[4] ),
    .o1(_03695_));
 b15norp02ar1n08x5 _29508_ (.a(_02327_),
    .b(_03695_),
    .o1(_03697_));
 b15aoai13an1n02x5 _29509_ (.a(_02323_),
    .b(_02319_),
    .c(_02298_),
    .d(_03697_),
    .o1(_03698_));
 b15nona23as1n32x5 _29510_ (.a(net698),
    .b(\us12.a[6] ),
    .c(net693),
    .d(\us12.a[4] ),
    .out0(_03699_));
 b15ztpn00an1n08x5 TAP_448 ();
 b15nor002aq1n06x5 _29512_ (.a(net701),
    .b(_03699_),
    .o1(_03701_));
 b15oai022ar1n02x5 _29513_ (.a(_02355_),
    .b(_02357_),
    .c(_02389_),
    .d(net710),
    .o1(_03702_));
 b15aoi022as1n04x5 _29514_ (.a(_02426_),
    .b(_03701_),
    .c(_03702_),
    .d(_02313_),
    .o1(_03703_));
 b15norp03al1n03x5 _29515_ (.a(_02320_),
    .b(_02325_),
    .c(_02469_),
    .o1(_03704_));
 b15norp03ah1n03x5 _29516_ (.a(net691),
    .b(_02310_),
    .c(_02427_),
    .o1(_03705_));
 b15nanb02an1n12x5 _29517_ (.a(net694),
    .b(net701),
    .out0(_03706_));
 b15aoi013al1n06x5 _29518_ (.a(_03704_),
    .b(_03705_),
    .c(_03706_),
    .d(_02279_),
    .o1(_03708_));
 b15nor002al1n06x5 _29519_ (.a(_02259_),
    .b(_02310_),
    .o1(_03709_));
 b15norp02ah1n12x5 _29520_ (.a(_02357_),
    .b(_02390_),
    .o1(_03710_));
 b15norp02an1n12x5 _29521_ (.a(_02276_),
    .b(_03695_),
    .o1(_03711_));
 b15nor002al1n02x5 _29522_ (.a(_02461_),
    .b(_03657_),
    .o1(_03712_));
 b15aoi222as1n06x5 _29523_ (.a(_02326_),
    .b(_03709_),
    .c(_03710_),
    .d(_03711_),
    .e(_03712_),
    .f(_02311_),
    .o1(_03713_));
 b15nand04al1n06x5 _29524_ (.a(_03698_),
    .b(_03703_),
    .c(_03708_),
    .d(_03713_),
    .o1(_03714_));
 b15ztpn00an1n08x5 TAP_447 ();
 b15ztpn00an1n08x5 TAP_446 ();
 b15ztpn00an1n08x5 TAP_445 ();
 b15nonb03ar1n02x5 _29528_ (.a(net710),
    .b(net699),
    .c(net696),
    .out0(_03719_));
 b15oai112ah1n02x5 _29529_ (.a(net714),
    .b(_02293_),
    .c(_02437_),
    .d(_03719_),
    .o1(_03720_));
 b15aoai13ar1n02x5 _29530_ (.a(_02355_),
    .b(_02351_),
    .c(_02475_),
    .d(_02242_),
    .o1(_03721_));
 b15aoi013as1n02x5 _29531_ (.a(net706),
    .b(_02381_),
    .c(_03720_),
    .d(_03721_),
    .o1(_03722_));
 b15xor002ar1n08x5 _29532_ (.a(\us12.a[6] ),
    .b(_02321_),
    .out0(_03723_));
 b15nand02as1n06x5 _29533_ (.a(net693),
    .b(_02346_),
    .o1(_03724_));
 b15and002al1n08x5 _29534_ (.a(\us12.a[4] ),
    .b(net693),
    .o(_03725_));
 b15nor002ah1n06x5 _29535_ (.a(\us12.a[4] ),
    .b(net693),
    .o1(_03726_));
 b15nor002al1n06x5 _29536_ (.a(\us12.a[6] ),
    .b(net712),
    .o1(_03727_));
 b15mdn022an1n06x5 _29537_ (.a(_03725_),
    .b(_03726_),
    .o1(_03728_),
    .sa(_03727_));
 b15oai122aq1n16x5 _29538_ (.a(net701),
    .b(_03723_),
    .c(_03724_),
    .d(_03728_),
    .e(net698),
    .o1(_03730_));
 b15nand02as1n08x5 _29539_ (.a(_03722_),
    .b(_03730_),
    .o1(_03731_));
 b15nand02ar1n02x5 _29540_ (.a(_02340_),
    .b(_02475_),
    .o1(_03732_));
 b15oai012al1n03x5 _29541_ (.a(_03732_),
    .b(_02340_),
    .c(_02294_),
    .o1(_03733_));
 b15nor002ar1n02x5 _29542_ (.a(_02325_),
    .b(_02366_),
    .o1(_03734_));
 b15oai013an1n06x5 _29543_ (.a(_02367_),
    .b(_03733_),
    .c(_03734_),
    .d(_02351_),
    .o1(_03735_));
 b15nona23as1n04x5 _29544_ (.a(_03694_),
    .b(_03714_),
    .c(_03731_),
    .d(_03735_),
    .out0(_03736_));
 b15nand02as1n02x5 _29545_ (.a(_02321_),
    .b(_03701_),
    .o1(_03737_));
 b15oai012al1n06x5 _29546_ (.a(_02437_),
    .b(_02293_),
    .c(_02430_),
    .o1(_03738_));
 b15qbfna2bn1n16x5 _29547_ (.a(net702),
    .b(_02449_),
    .o1(_03739_));
 b15oaoi13ah1n08x5 _29548_ (.a(net709),
    .b(_03737_),
    .c(_03738_),
    .d(_03739_),
    .o1(_03741_));
 b15nor002ar1n06x5 _29549_ (.a(_02389_),
    .b(_03699_),
    .o1(_03742_));
 b15aoi022an1n08x5 _29550_ (.a(_03688_),
    .b(_02392_),
    .c(_02475_),
    .d(_03689_),
    .o1(_03743_));
 b15nand03al1n08x5 _29551_ (.a(_02251_),
    .b(_02328_),
    .c(_02449_),
    .o1(_03744_));
 b15nano22aq1n08x5 _29552_ (.a(net714),
    .b(net709),
    .c(net705),
    .out0(_03745_));
 b15aoi112as1n04x5 _29553_ (.a(_03710_),
    .b(_03745_),
    .c(_02321_),
    .d(_02367_),
    .o1(_03746_));
 b15oai112ah1n16x5 _29554_ (.a(_03743_),
    .b(_03744_),
    .c(_02466_),
    .d(_03746_),
    .o1(_03747_));
 b15nor003ah1n08x5 _29555_ (.a(_03741_),
    .b(_03742_),
    .c(_03747_),
    .o1(_03748_));
 b15ztpn00an1n08x5 TAP_444 ();
 b15aoi013ah1n03x5 _29557_ (.a(_02449_),
    .b(_02375_),
    .c(net712),
    .d(_02437_),
    .o1(_03750_));
 b15nonb02an1n12x5 _29558_ (.a(\us12.a[2] ),
    .b(net698),
    .out0(_03752_));
 b15aoi022as1n06x5 _29559_ (.a(net698),
    .b(_02375_),
    .c(_03752_),
    .d(_02365_),
    .o1(_03753_));
 b15norp03aq1n12x5 _29560_ (.a(_02385_),
    .b(_03750_),
    .c(_03753_),
    .o1(_03754_));
 b15norp03al1n08x5 _29561_ (.a(_02242_),
    .b(_02309_),
    .c(_03648_),
    .o1(_03755_));
 b15nor002an1n03x5 _29562_ (.a(\us12.a[1] ),
    .b(_02471_),
    .o1(_03756_));
 b15oai012an1n04x5 _29563_ (.a(net708),
    .b(_03755_),
    .c(_03756_),
    .o1(_03757_));
 b15norp02ah1n12x5 _29564_ (.a(_02317_),
    .b(_03695_),
    .o1(_03758_));
 b15norp02ar1n02x5 _29565_ (.a(_03677_),
    .b(_03644_),
    .o1(_03759_));
 b15aoi022al1n04x5 _29566_ (.a(_02275_),
    .b(_03758_),
    .c(_03759_),
    .d(\us12.a[0] ),
    .o1(_03760_));
 b15aoi012al1n06x5 _29567_ (.a(net705),
    .b(_03757_),
    .c(_03760_),
    .o1(_03761_));
 b15ztpn00an1n08x5 TAP_443 ();
 b15norp02an1n16x5 _29569_ (.a(_02259_),
    .b(_03648_),
    .o1(_03764_));
 b15aoi022an1n02x5 _29570_ (.a(_02343_),
    .b(_03670_),
    .c(_03764_),
    .d(_02361_),
    .o1(_03765_));
 b15nandp3al1n03x5 _29571_ (.a(net703),
    .b(_02313_),
    .c(_02415_),
    .o1(_03766_));
 b15aoi012ar1n06x5 _29572_ (.a(net715),
    .b(_03765_),
    .c(_03766_),
    .o1(_03767_));
 b15norp03ar1n16x5 _29573_ (.a(_03754_),
    .b(_03761_),
    .c(_03767_),
    .o1(_03768_));
 b15nona23as1n32x5 _29574_ (.a(_03687_),
    .b(_03736_),
    .c(_03748_),
    .d(_03768_),
    .out0(_03769_));
 b15xor002ah1n03x5 _29575_ (.a(_03034_),
    .b(_03769_),
    .out0(_03770_));
 b15xor002aq1n08x5 _29576_ (.a(_03634_),
    .b(_03770_),
    .out0(_03771_));
 b15ztpn00an1n08x5 TAP_442 ();
 b15ztpn00an1n08x5 TAP_441 ();
 b15nonb02as1n16x5 _29579_ (.a(net584),
    .b(net582),
    .out0(_03775_));
 b15ztpn00an1n08x5 TAP_440 ();
 b15norp02an1n02x5 _29581_ (.a(_03163_),
    .b(_03249_),
    .o1(_03777_));
 b15ztpn00an1n08x5 TAP_439 ();
 b15aoi022aq1n02x5 _29583_ (.a(_03199_),
    .b(_03775_),
    .c(_03777_),
    .d(_03157_),
    .o1(_03779_));
 b15ztpn00an1n08x5 TAP_438 ();
 b15ztpn00an1n08x5 TAP_437 ();
 b15nanb02al1n08x5 _29586_ (.a(net571),
    .b(net595),
    .out0(_03782_));
 b15nand04ar1n04x5 _29587_ (.a(net568),
    .b(_03228_),
    .c(_03782_),
    .d(_03219_),
    .o1(_03783_));
 b15ztpn00an1n08x5 TAP_436 ();
 b15aoi013ar1n02x5 _29589_ (.a(_03163_),
    .b(net582),
    .c(_03132_),
    .d(_03186_),
    .o1(_03786_));
 b15and002an1n02x5 _29590_ (.a(_03783_),
    .b(_03786_),
    .o(_03787_));
 b15ztpn00an1n08x5 TAP_435 ();
 b15nor004as1n12x5 _29592_ (.a(_03223_),
    .b(net569),
    .c(_03036_),
    .d(_03074_),
    .o1(_03789_));
 b15norp02an1n04x5 _29593_ (.a(net573),
    .b(net582),
    .o1(_03790_));
 b15aoai13al1n02x5 _29594_ (.a(net574),
    .b(_03789_),
    .c(_03790_),
    .d(_03108_),
    .o1(_03791_));
 b15oaoi13an1n03x5 _29595_ (.a(_03102_),
    .b(_03779_),
    .c(_03787_),
    .d(_03791_),
    .o1(_03792_));
 b15ztpn00an1n08x5 TAP_434 ();
 b15nand04ar1n02x5 _29597_ (.a(net595),
    .b(_03162_),
    .c(_03228_),
    .d(_03219_),
    .o1(_03794_));
 b15nand02as1n24x5 _29598_ (.a(_03203_),
    .b(_03228_),
    .o1(_03796_));
 b15oai112ar1n02x5 _29599_ (.a(_03163_),
    .b(_03794_),
    .c(_03249_),
    .d(_03796_),
    .o1(_03797_));
 b15nanb02as1n24x5 _29600_ (.a(net591),
    .b(net584),
    .out0(_03798_));
 b15nor002ar1n06x5 _29601_ (.a(net575),
    .b(_03097_),
    .o1(_03799_));
 b15nanb02ah1n03x5 _29602_ (.a(net571),
    .b(net575),
    .out0(_03800_));
 b15nandp2ar1n02x5 _29603_ (.a(_03106_),
    .b(_03800_),
    .o1(_03801_));
 b15nor004an1n04x5 _29604_ (.a(net582),
    .b(_03798_),
    .c(_03799_),
    .d(_03801_),
    .o1(_03802_));
 b15norp02ar1n02x5 _29605_ (.a(_03797_),
    .b(_03802_),
    .o1(_03803_));
 b15ztpn00an1n08x5 TAP_433 ();
 b15ztpn00an1n08x5 TAP_432 ();
 b15nano23ah1n24x5 _29608_ (.a(net578),
    .b(net570),
    .c(\us23.a[6] ),
    .d(net576),
    .out0(_03807_));
 b15aoai13ah1n06x5 _29609_ (.a(net583),
    .b(_03807_),
    .c(_03171_),
    .d(_03186_),
    .o1(_03808_));
 b15aoi012an1n02x5 _29610_ (.a(_03787_),
    .b(_03803_),
    .c(_03808_),
    .o1(_03809_));
 b15nandp3aq1n03x5 _29611_ (.a(net594),
    .b(_03162_),
    .c(_03233_),
    .o1(_03810_));
 b15aoai13ar1n08x5 _29612_ (.a(_03810_),
    .b(net590),
    .c(_03205_),
    .d(_03234_),
    .o1(_03811_));
 b15nand03ah1n06x5 _29613_ (.a(net584),
    .b(_03203_),
    .c(_03204_),
    .o1(_03812_));
 b15oai012al1n08x5 _29614_ (.a(_03812_),
    .b(_03234_),
    .c(_03283_),
    .o1(_03813_));
 b15nor002ah1n24x5 _29615_ (.a(net595),
    .b(net582),
    .o1(_03814_));
 b15aoi022al1n16x5 _29616_ (.a(_03775_),
    .b(_03811_),
    .c(_03813_),
    .d(_03814_),
    .o1(_03815_));
 b15ztpn00an1n08x5 TAP_431 ();
 b15and002as1n08x5 _29618_ (.a(net590),
    .b(net584),
    .o(_03818_));
 b15and003ar1n02x5 _29619_ (.a(net568),
    .b(_03204_),
    .c(_03814_),
    .o(_03819_));
 b15orn002as1n08x5 _29620_ (.a(net575),
    .b(net568),
    .o(_03820_));
 b15nandp2ah1n04x5 _29621_ (.a(net579),
    .b(net595),
    .o1(_03821_));
 b15ztpn00an1n08x5 TAP_430 ();
 b15nandp2ar1n08x5 _29623_ (.a(_03102_),
    .b(net582),
    .o1(_03823_));
 b15oaoi13ar1n02x5 _29624_ (.a(_03820_),
    .b(_03821_),
    .c(net579),
    .d(_03823_),
    .o1(_03824_));
 b15oai112aq1n02x5 _29625_ (.a(net571),
    .b(_03818_),
    .c(_03819_),
    .d(_03824_),
    .o1(_03825_));
 b15ztpn00an1n08x5 TAP_429 ();
 b15nandp2aq1n24x5 _29627_ (.a(net584),
    .b(net580),
    .o1(_03827_));
 b15nanb02an1n24x5 _29628_ (.a(net590),
    .b(net573),
    .out0(_03829_));
 b15nor004an1n02x5 _29629_ (.a(net592),
    .b(_03827_),
    .c(_03820_),
    .d(_03829_),
    .o1(_03830_));
 b15nor003as1n08x5 _29630_ (.a(net574),
    .b(net569),
    .c(net572),
    .o1(_03831_));
 b15aoai13ah1n03x5 _29631_ (.a(net577),
    .b(_03830_),
    .c(_03831_),
    .d(_03291_),
    .o1(_03832_));
 b15ztpn00an1n08x5 TAP_428 ();
 b15nor004as1n03x5 _29633_ (.a(net577),
    .b(_03827_),
    .c(_03820_),
    .d(_03829_),
    .o1(_03834_));
 b15norp03ar1n16x5 _29634_ (.a(net580),
    .b(_03050_),
    .c(_03135_),
    .o1(_03835_));
 b15norp02ar1n48x5 _29635_ (.a(\us23.a[1] ),
    .b(\us23.a[2] ),
    .o1(_03836_));
 b15aoai13as1n06x5 _29636_ (.a(net592),
    .b(_03834_),
    .c(_03835_),
    .d(_03836_),
    .o1(_03837_));
 b15nand04aq1n06x5 _29637_ (.a(_03815_),
    .b(_03825_),
    .c(_03832_),
    .d(_03837_),
    .o1(_03838_));
 b15norp03ar1n08x5 _29638_ (.a(_03792_),
    .b(_03809_),
    .c(_03838_),
    .o1(_03840_));
 b15nand02ar1n02x5 _29639_ (.a(net571),
    .b(_03836_),
    .o1(_03841_));
 b15oaoi13ar1n02x5 _29640_ (.a(_03820_),
    .b(_03841_),
    .c(net571),
    .d(_03046_),
    .o1(_03842_));
 b15nand02ah1n24x5 _29641_ (.a(net575),
    .b(net568),
    .o1(_03843_));
 b15norp02ar1n02x5 _29642_ (.a(_03046_),
    .b(_03843_),
    .o1(_03844_));
 b15oai112an1n04x5 _29643_ (.a(net577),
    .b(_03814_),
    .c(_03842_),
    .d(_03844_),
    .o1(_03845_));
 b15nonb02aq1n06x5 _29644_ (.a(net588),
    .b(net592),
    .out0(_03846_));
 b15oab012ar1n02x5 _29645_ (.a(_03121_),
    .b(_03196_),
    .c(_03846_),
    .out0(_03847_));
 b15oab012an1n06x5 _29646_ (.a(net583),
    .b(_03170_),
    .c(_03847_),
    .out0(_03848_));
 b15qgbno2an1n10x5 _29647_ (.a(net574),
    .b(net571),
    .o1(_03849_));
 b15nonb03al1n04x5 _29648_ (.a(net584),
    .b(net582),
    .c(net588),
    .out0(_03851_));
 b15nona23al1n04x5 _29649_ (.a(_03106_),
    .b(_03108_),
    .c(_03849_),
    .d(_03851_),
    .out0(_03852_));
 b15nonb02aq1n16x5 _29650_ (.a(net582),
    .b(net586),
    .out0(_03853_));
 b15nandp3an1n03x5 _29651_ (.a(net588),
    .b(_03853_),
    .c(_03831_),
    .o1(_03854_));
 b15nano23an1n03x5 _29652_ (.a(net588),
    .b(net583),
    .c(net569),
    .d(net572),
    .out0(_03855_));
 b15aoi022ah1n06x5 _29653_ (.a(_03240_),
    .b(_03775_),
    .c(_03855_),
    .d(_03251_),
    .o1(_03856_));
 b15oai112an1n12x5 _29654_ (.a(_03852_),
    .b(_03854_),
    .c(net592),
    .d(_03856_),
    .o1(_03857_));
 b15nand03ah1n03x5 _29655_ (.a(_03233_),
    .b(_03231_),
    .c(_03851_),
    .o1(_03858_));
 b15oai013an1n03x5 _29656_ (.a(_03858_),
    .b(_03217_),
    .c(_03205_),
    .d(_03210_),
    .o1(_03859_));
 b15nor003ar1n02x5 _29657_ (.a(_03100_),
    .b(net588),
    .c(_03053_),
    .o1(_03860_));
 b15norp03as1n02x5 _29658_ (.a(net574),
    .b(_03281_),
    .c(_03071_),
    .o1(_03862_));
 b15oai112as1n04x5 _29659_ (.a(net577),
    .b(_03219_),
    .c(_03860_),
    .d(_03862_),
    .o1(_03863_));
 b15nano22ah1n08x5 _29660_ (.a(net575),
    .b(net579),
    .c(net573),
    .out0(_03864_));
 b15nonb02ah1n12x5 _29661_ (.a(net573),
    .b(net582),
    .out0(_03865_));
 b15aoi022ar1n02x5 _29662_ (.a(_03134_),
    .b(_03864_),
    .c(_03865_),
    .d(_03233_),
    .o1(_03866_));
 b15ztpn00an1n08x5 TAP_427 ();
 b15oai013an1n03x5 _29664_ (.a(_03863_),
    .b(_03866_),
    .c(_03798_),
    .d(net569),
    .o1(_03868_));
 b15nor004an1n06x5 _29665_ (.a(_03848_),
    .b(_03857_),
    .c(_03859_),
    .d(_03868_),
    .o1(_03869_));
 b15aoi022ar1n02x5 _29666_ (.a(_03122_),
    .b(_03255_),
    .c(_03270_),
    .d(_03777_),
    .o1(_03870_));
 b15nor002al1n02x5 _29667_ (.a(net595),
    .b(_03870_),
    .o1(_03871_));
 b15ztpn00an1n08x5 TAP_426 ();
 b15norp03ar1n02x5 _29669_ (.a(net582),
    .b(_03057_),
    .c(_03272_),
    .o1(_03874_));
 b15aoai13al1n02x5 _29670_ (.a(net584),
    .b(_03874_),
    .c(_03240_),
    .d(net582),
    .o1(_03875_));
 b15aoi012ar1n02x5 _29671_ (.a(_03079_),
    .b(_03210_),
    .c(net573),
    .o1(_03876_));
 b15nandp3ar1n02x5 _29672_ (.a(net569),
    .b(_03219_),
    .c(_03876_),
    .o1(_03877_));
 b15nanb02as1n04x5 _29673_ (.a(net583),
    .b(net592),
    .out0(_03878_));
 b15oai022al1n12x5 _29674_ (.a(_03086_),
    .b(_03823_),
    .c(_03878_),
    .d(_03135_),
    .o1(_03879_));
 b15aoi022ar1n02x5 _29675_ (.a(_03036_),
    .b(_03240_),
    .c(_03879_),
    .d(_03233_),
    .o1(_03880_));
 b15oai112ar1n04x5 _29676_ (.a(_03875_),
    .b(_03877_),
    .c(_03880_),
    .d(_03283_),
    .o1(_03881_));
 b15nano23ah1n03x5 _29677_ (.a(_03845_),
    .b(_03869_),
    .c(_03871_),
    .d(_03881_),
    .out0(_03882_));
 b15ztpn00an1n08x5 TAP_425 ();
 b15ztpn00an1n08x5 TAP_424 ();
 b15ztpn00an1n08x5 TAP_423 ();
 b15nand02aq1n24x5 _29681_ (.a(\us23.a[1] ),
    .b(net583),
    .o1(_03887_));
 b15oai022aq1n04x5 _29682_ (.a(net582),
    .b(_03187_),
    .c(_03234_),
    .d(_03887_),
    .o1(_03888_));
 b15aoi122ar1n06x5 _29683_ (.a(_03067_),
    .b(_03189_),
    .c(net590),
    .d(_03888_),
    .e(net595),
    .o1(_03889_));
 b15nandp2an1n08x5 _29684_ (.a(_03163_),
    .b(net583),
    .o1(_03890_));
 b15aoi012an1n02x5 _29685_ (.a(_03890_),
    .b(_03810_),
    .c(_03247_),
    .o1(_03891_));
 b15ztpn00an1n08x5 TAP_422 ();
 b15nonb02al1n03x5 _29687_ (.a(net590),
    .b(net579),
    .out0(_03893_));
 b15aoai13ah1n03x5 _29688_ (.a(_03231_),
    .b(_03893_),
    .c(_03100_),
    .d(_03163_),
    .o1(_03895_));
 b15nor002ar1n08x5 _29689_ (.a(_03102_),
    .b(_03163_),
    .o1(_03896_));
 b15ztpn00an1n08x5 TAP_421 ();
 b15aoi022as1n04x5 _29691_ (.a(_03896_),
    .b(_03106_),
    .c(_03108_),
    .d(_03123_),
    .o1(_03898_));
 b15oai112an1n12x5 _29692_ (.a(net582),
    .b(_03895_),
    .c(_03898_),
    .d(_03800_),
    .o1(_03899_));
 b15ztpn00an1n08x5 TAP_420 ();
 b15aoi112al1n02x5 _29694_ (.a(_03100_),
    .b(_03053_),
    .c(_03821_),
    .d(_03163_),
    .o1(_03901_));
 b15norp02al1n08x5 _29695_ (.a(net574),
    .b(_03071_),
    .o1(_03902_));
 b15oai012ar1n02x5 _29696_ (.a(net595),
    .b(net590),
    .c(net579),
    .o1(_03903_));
 b15oai012al1n03x5 _29697_ (.a(_03903_),
    .b(_03210_),
    .c(net579),
    .o1(_03904_));
 b15aoi012an1n04x5 _29698_ (.a(_03901_),
    .b(_03902_),
    .c(_03904_),
    .o1(_03906_));
 b15ztpn00an1n08x5 TAP_419 ();
 b15aoi022ar1n02x5 _29700_ (.a(_03102_),
    .b(_03088_),
    .c(_03285_),
    .d(net590),
    .o1(_03908_));
 b15nandp3ar1n02x5 _29701_ (.a(_03036_),
    .b(_03906_),
    .c(_03908_),
    .o1(_03909_));
 b15aoi012ah1n02x5 _29702_ (.a(_03891_),
    .b(_03899_),
    .c(_03909_),
    .o1(_03910_));
 b15aoi012al1n06x5 _29703_ (.a(_03889_),
    .b(_03910_),
    .c(_03067_),
    .o1(_03911_));
 b15nona22aq1n24x5 _29704_ (.a(net591),
    .b(net587),
    .c(net585),
    .out0(_03912_));
 b15norp03al1n04x5 _29705_ (.a(_03071_),
    .b(_03912_),
    .c(_03287_),
    .o1(_03913_));
 b15nor003ar1n06x5 _29706_ (.a(_03046_),
    .b(_03071_),
    .c(_03287_),
    .o1(_03914_));
 b15nor003ar1n06x5 _29707_ (.a(_03087_),
    .b(_03135_),
    .c(_03217_),
    .o1(_03915_));
 b15oaoi13as1n08x5 _29708_ (.a(_03913_),
    .b(net591),
    .c(_03914_),
    .d(_03915_),
    .o1(_03917_));
 b15nand02an1n03x5 _29709_ (.a(_03123_),
    .b(_03075_),
    .o1(_03918_));
 b15aobi12as1n06x5 _29710_ (.a(_03241_),
    .b(_03918_),
    .c(_03128_),
    .out0(_03919_));
 b15nonb03an1n06x5 _29711_ (.a(net573),
    .b(net579),
    .c(net575),
    .out0(_03920_));
 b15aoi012aq1n02x5 _29712_ (.a(_03864_),
    .b(_03920_),
    .c(net590),
    .o1(_03921_));
 b15nor003an1n04x5 _29713_ (.a(_03102_),
    .b(_03249_),
    .c(_03921_),
    .o1(_03922_));
 b15nandp2as1n16x5 _29714_ (.a(_03102_),
    .b(_03107_),
    .o1(_03923_));
 b15and002ar1n08x5 _29715_ (.a(net573),
    .b(net582),
    .o(_03924_));
 b15nandp2al1n08x5 _29716_ (.a(_03204_),
    .b(_03924_),
    .o1(_03925_));
 b15norp02an1n03x5 _29717_ (.a(_03790_),
    .b(_03924_),
    .o1(_03926_));
 b15oaoi13aq1n04x5 _29718_ (.a(_03923_),
    .b(_03925_),
    .c(_03079_),
    .d(_03926_),
    .o1(_03928_));
 b15oai012aq1n12x5 _29719_ (.a(net569),
    .b(_03922_),
    .c(_03928_),
    .o1(_03929_));
 b15nandp3ar1n16x5 _29720_ (.a(_03917_),
    .b(_03919_),
    .c(_03929_),
    .o1(_03930_));
 b15nano23an1n16x5 _29721_ (.a(_03840_),
    .b(_03882_),
    .c(_03911_),
    .d(_03930_),
    .out0(_03931_));
 b15xor002ar1n03x5 _29722_ (.a(_02771_),
    .b(_03413_),
    .out0(_03932_));
 b15xor002aq1n03x5 _29723_ (.a(net393),
    .b(_03932_),
    .out0(_03933_));
 b15xor002aq1n06x5 _29724_ (.a(_03771_),
    .b(_03933_),
    .out0(_03934_));
 b15ztpn00an1n08x5 TAP_418 ();
 b15mdn022al1n12x5 _29726_ (.a(_03418_),
    .b(_03934_),
    .o1(_03936_),
    .sa(net537));
 b15xor002as1n12x5 _29727_ (.a(\u0.w[1][1] ),
    .b(_03936_),
    .out0(_00106_));
 b15aoai13al1n02x5 _29728_ (.a(net584),
    .b(_03122_),
    .c(_03270_),
    .d(net582),
    .o1(_03938_));
 b15aoi022an1n02x5 _29729_ (.a(_03036_),
    .b(_03251_),
    .c(_03204_),
    .d(_03924_),
    .o1(_03939_));
 b15oai013as1n04x5 _29730_ (.a(_03938_),
    .b(_03939_),
    .c(_03283_),
    .d(net569),
    .o1(_03940_));
 b15nandp3ar1n02x5 _29731_ (.a(\us23.a[2] ),
    .b(_03036_),
    .c(_03270_),
    .o1(_03941_));
 b15aoi022ar1n02x5 _29732_ (.a(_03203_),
    .b(_03237_),
    .c(_03924_),
    .d(net568),
    .o1(_03942_));
 b15nand02ar1n02x5 _29733_ (.a(_03100_),
    .b(_03942_),
    .o1(_03943_));
 b15obai22al1n12x5 _29734_ (.a(_03865_),
    .b(net569),
    .c(_03086_),
    .d(_03827_),
    .out0(_03944_));
 b15oai012ah1n03x5 _29735_ (.a(_03943_),
    .b(_03944_),
    .c(_03100_),
    .o1(_03945_));
 b15oaoi13ah1n03x5 _29736_ (.a(net590),
    .b(_03941_),
    .c(_03945_),
    .d(net579),
    .o1(_03946_));
 b15oai012aq1n12x5 _29737_ (.a(net594),
    .b(_03940_),
    .c(_03946_),
    .o1(_03947_));
 b15norp02al1n02x5 _29738_ (.a(_03123_),
    .b(_03276_),
    .o1(_03949_));
 b15oai112al1n06x5 _29739_ (.a(net581),
    .b(_03046_),
    .c(_03215_),
    .d(_03949_),
    .o1(_03950_));
 b15aoi012ar1n04x5 _29740_ (.a(_03205_),
    .b(_03107_),
    .c(net593),
    .o1(_03951_));
 b15oai112al1n08x5 _29741_ (.a(net581),
    .b(_03798_),
    .c(_03951_),
    .d(_03157_),
    .o1(_03952_));
 b15nand02ar1n02x5 _29742_ (.a(net585),
    .b(_03167_),
    .o1(_03953_));
 b15oaoi13ah1n03x5 _29743_ (.a(net587),
    .b(_03953_),
    .c(_03149_),
    .d(net585),
    .o1(_03954_));
 b15aoi022al1n06x5 _29744_ (.a(_03157_),
    .b(_03274_),
    .c(_03219_),
    .d(_03150_),
    .o1(_03955_));
 b15oai122ar1n12x5 _29745_ (.a(_03950_),
    .b(_03952_),
    .c(_03954_),
    .d(_03955_),
    .e(net593),
    .o1(_03956_));
 b15nona23as1n08x5 _29746_ (.a(net578),
    .b(net572),
    .c(net569),
    .d(net576),
    .out0(_03957_));
 b15norp03ar1n02x5 _29747_ (.a(net581),
    .b(_03057_),
    .c(_03957_),
    .o1(_03958_));
 b15nonb02ar1n12x5 _29748_ (.a(net583),
    .b(net592),
    .out0(_03960_));
 b15aoai13al1n03x5 _29749_ (.a(net585),
    .b(_03958_),
    .c(_03960_),
    .d(_03088_),
    .o1(_03961_));
 b15norp02as1n12x5 _29750_ (.a(_03050_),
    .b(_03135_),
    .o1(_03962_));
 b15oai112al1n06x5 _29751_ (.a(net587),
    .b(_03962_),
    .c(_03219_),
    .d(_03165_),
    .o1(_03963_));
 b15nor002ah1n04x5 _29752_ (.a(net593),
    .b(_03249_),
    .o1(_03964_));
 b15aoi022an1n04x5 _29753_ (.a(_03157_),
    .b(_03775_),
    .c(_03964_),
    .d(_03132_),
    .o1(_03965_));
 b15oai112ah1n06x5 _29754_ (.a(_03961_),
    .b(_03963_),
    .c(_03965_),
    .d(net587),
    .o1(_03966_));
 b15aoi013al1n03x5 _29755_ (.a(_03067_),
    .b(net581),
    .c(_03240_),
    .d(_03123_),
    .o1(_03967_));
 b15ao0022al1n02x5 _29756_ (.a(_03036_),
    .b(_03807_),
    .c(_03240_),
    .d(_03960_),
    .o(_03968_));
 b15aoi022ar1n08x5 _29757_ (.a(_03807_),
    .b(_03140_),
    .c(_03968_),
    .d(net589),
    .o1(_03969_));
 b15aoi012an1n08x5 _29758_ (.a(_03967_),
    .b(_03969_),
    .c(_03067_),
    .o1(_03971_));
 b15nor003ar1n08x5 _29759_ (.a(_03956_),
    .b(_03966_),
    .c(_03971_),
    .o1(_03972_));
 b15nand03aq1n02x5 _29760_ (.a(net575),
    .b(\us23.a[7] ),
    .c(net582),
    .o1(_03973_));
 b15orn002aq1n02x5 _29761_ (.a(\us23.a[7] ),
    .b(net582),
    .o(_03974_));
 b15oai012aq1n06x5 _29762_ (.a(_03973_),
    .b(_03974_),
    .c(net575),
    .o1(_03975_));
 b15norp03as1n04x5 _29763_ (.a(net579),
    .b(net573),
    .c(net595),
    .o1(_03976_));
 b15aoi022ar1n16x5 _29764_ (.a(_03240_),
    .b(_03775_),
    .c(_03975_),
    .d(_03976_),
    .o1(_03977_));
 b15norp02ar1n02x5 _29765_ (.a(net585),
    .b(_03187_),
    .o1(_03978_));
 b15aoi112ar1n02x5 _29766_ (.a(_03036_),
    .b(_03978_),
    .c(_03150_),
    .d(net585),
    .o1(_03979_));
 b15aoi022ar1n02x5 _29767_ (.a(_03089_),
    .b(_03186_),
    .c(_03196_),
    .d(_03157_),
    .o1(_03980_));
 b15aoai13an1n02x5 _29768_ (.a(_03977_),
    .b(_03979_),
    .c(_03980_),
    .d(_03036_),
    .o1(_03982_));
 b15nand02ar1n16x5 _29769_ (.a(_03162_),
    .b(_03228_),
    .o1(_03983_));
 b15aoi012aq1n16x5 _29770_ (.a(_03102_),
    .b(_03046_),
    .c(_03181_),
    .o1(_03984_));
 b15obai22aq1n04x5 _29771_ (.a(_03923_),
    .b(_03234_),
    .c(_03983_),
    .d(_03984_),
    .out0(_03985_));
 b15aoai13ar1n02x5 _29772_ (.a(_03102_),
    .b(_03107_),
    .c(_03255_),
    .d(_03205_),
    .o1(_03986_));
 b15oai012aq1n04x5 _29773_ (.a(_03205_),
    .b(_03796_),
    .c(_03896_),
    .o1(_03987_));
 b15aoi012ar1n02x5 _29774_ (.a(_03985_),
    .b(_03986_),
    .c(_03987_),
    .o1(_03988_));
 b15aoai13ar1n02x5 _29775_ (.a(net594),
    .b(_03137_),
    .c(_03962_),
    .d(_03163_),
    .o1(_03989_));
 b15aoai13al1n02x5 _29776_ (.a(_03988_),
    .b(_03836_),
    .c(_03187_),
    .d(_03989_),
    .o1(_03990_));
 b15aoi022as1n04x5 _29777_ (.a(net587),
    .b(_03982_),
    .c(_03990_),
    .d(_03036_),
    .o1(_03991_));
 b15nandp2ar1n02x5 _29778_ (.a(net577),
    .b(_03067_),
    .o1(_03993_));
 b15nor002aq1n12x5 _29779_ (.a(net573),
    .b(net595),
    .o1(_03994_));
 b15nanb02ar1n02x5 _29780_ (.a(_03843_),
    .b(_03994_),
    .out0(_03995_));
 b15nanb02aq1n04x5 _29781_ (.a(net590),
    .b(net568),
    .out0(_03996_));
 b15aoi022al1n06x5 _29782_ (.a(_03143_),
    .b(_03253_),
    .c(_03996_),
    .d(_03177_),
    .o1(_03997_));
 b15oaoi13an1n04x5 _29783_ (.a(_03993_),
    .b(_03995_),
    .c(_03997_),
    .d(net574),
    .o1(_03998_));
 b15aoi012aq1n04x5 _29784_ (.a(_03247_),
    .b(_03284_),
    .c(_03923_),
    .o1(_03999_));
 b15oai013aq1n03x5 _29785_ (.a(net583),
    .b(_03242_),
    .c(_03796_),
    .d(net588),
    .o1(_04000_));
 b15aoi022ar1n02x5 _29786_ (.a(_03846_),
    .b(_03132_),
    .c(_03199_),
    .d(net592),
    .o1(_04001_));
 b15nor002an1n02x5 _29787_ (.a(_03067_),
    .b(_04001_),
    .o1(_04002_));
 b15nor004ah1n06x5 _29788_ (.a(_03998_),
    .b(_03999_),
    .c(_04000_),
    .d(_04002_),
    .o1(_04004_));
 b15aoi012ar1n02x5 _29789_ (.a(net584),
    .b(_03086_),
    .c(_03135_),
    .o1(_04005_));
 b15nanb02an1n02x5 _29790_ (.a(net584),
    .b(net568),
    .out0(_04006_));
 b15ao0022ar1n02x5 _29791_ (.a(net574),
    .b(_04005_),
    .c(_04006_),
    .d(_03849_),
    .o(_04007_));
 b15nor002an1n04x5 _29792_ (.a(_03100_),
    .b(_03135_),
    .o1(_04008_));
 b15aoi022aq1n04x5 _29793_ (.a(net577),
    .b(_04007_),
    .c(_04008_),
    .d(_03207_),
    .o1(_04009_));
 b15oai012as1n08x5 _29794_ (.a(_04004_),
    .b(_04009_),
    .c(net588),
    .o1(_04010_));
 b15aoi012ar1n02x5 _29795_ (.a(net581),
    .b(_03150_),
    .c(_03196_),
    .o1(_04011_));
 b15oai012al1n02x5 _29796_ (.a(net587),
    .b(_03073_),
    .c(_03150_),
    .o1(_04012_));
 b15aob012ar1n12x5 _29797_ (.a(_04010_),
    .b(_04011_),
    .c(_04012_),
    .out0(_04013_));
 b15nand04aq1n16x5 _29798_ (.a(_03947_),
    .b(_03972_),
    .c(_03991_),
    .d(_04013_),
    .o1(_04015_));
 b15nonb03as1n08x5 _29799_ (.a(net710),
    .b(net707),
    .c(net713),
    .out0(_04016_));
 b15oaoi13aq1n03x5 _29800_ (.a(_02381_),
    .b(_02351_),
    .c(_03655_),
    .d(_04016_),
    .o1(_04017_));
 b15qgbna2an1n05x5 _29801_ (.o1(_04018_),
    .a(net707),
    .b(_02351_));
 b15aoai13aq1n08x5 _29802_ (.a(_04017_),
    .b(net710),
    .c(_02463_),
    .d(_04018_),
    .o1(_04019_));
 b15nandp3ar1n02x5 _29803_ (.a(net711),
    .b(_02341_),
    .c(_02333_),
    .o1(_04020_));
 b15oaoi13ah1n02x5 _29804_ (.a(_02300_),
    .b(_04020_),
    .c(_02366_),
    .d(net711),
    .o1(_04021_));
 b15oai012ar1n02x5 _29805_ (.a(_02381_),
    .b(_03667_),
    .c(_03666_),
    .o1(_04022_));
 b15oai012ar1n02x5 _29806_ (.a(_04019_),
    .b(_04021_),
    .c(_04022_),
    .o1(_04023_));
 b15nano23al1n24x5 _29807_ (.a(net697),
    .b(net695),
    .c(net692),
    .d(net700),
    .out0(_04024_));
 b15nandp2ar1n02x5 _29808_ (.a(net708),
    .b(_04024_),
    .o1(_04026_));
 b15oaoi13ar1n02x5 _29809_ (.a(_02340_),
    .b(_04026_),
    .c(_02366_),
    .d(net708),
    .o1(_04027_));
 b15norp03an1n02x5 _29810_ (.a(net708),
    .b(_02325_),
    .c(_02469_),
    .o1(_04028_));
 b15oai012as1n03x5 _29811_ (.a(net704),
    .b(_04027_),
    .c(_04028_),
    .o1(_04029_));
 b15oai022ar1n02x5 _29812_ (.a(_02427_),
    .b(_02471_),
    .c(_02500_),
    .d(_02368_),
    .o1(_04030_));
 b15nanb02as1n12x5 _29813_ (.a(net706),
    .b(\us12.a[6] ),
    .out0(_04031_));
 b15norp02al1n12x5 _29814_ (.a(net699),
    .b(net701),
    .o1(_04032_));
 b15nonb02an1n04x5 _29815_ (.a(net699),
    .b(net694),
    .out0(_04033_));
 b15aoi022as1n08x5 _29816_ (.a(_04031_),
    .b(_04032_),
    .c(_04033_),
    .d(_02367_),
    .o1(_04034_));
 b15nanb02aq1n16x5 _29817_ (.a(net691),
    .b(net696),
    .out0(_04035_));
 b15nand02al1n24x5 _29818_ (.a(_02430_),
    .b(_02291_),
    .o1(_04037_));
 b15oai122ah1n02x5 _29819_ (.a(_02477_),
    .b(_04034_),
    .c(_04035_),
    .d(_04037_),
    .e(net707),
    .o1(_04038_));
 b15oai013aq1n03x5 _29820_ (.a(net713),
    .b(_02478_),
    .c(_04030_),
    .d(_04038_),
    .o1(_04039_));
 b15nand03as1n02x5 _29821_ (.a(_04023_),
    .b(_04029_),
    .c(_04039_),
    .o1(_04040_));
 b15oai012al1n06x5 _29822_ (.a(_02343_),
    .b(_03755_),
    .c(_03756_),
    .o1(_04041_));
 b15and002ar1n02x5 _29823_ (.a(_02449_),
    .b(_03670_),
    .o(_04042_));
 b15aoai13ar1n03x5 _29824_ (.a(_03692_),
    .b(_04042_),
    .c(_02355_),
    .d(_03711_),
    .o1(_04043_));
 b15norp02an1n24x5 _29825_ (.a(_02309_),
    .b(_02310_),
    .o1(_04044_));
 b15nor002al1n04x5 _29826_ (.a(net711),
    .b(_02389_),
    .o1(_04045_));
 b15aoi222ah1n06x5 _29827_ (.a(_04044_),
    .b(_02358_),
    .c(_04045_),
    .d(_03764_),
    .e(_03710_),
    .f(_02462_),
    .o1(_04046_));
 b15nor003an1n08x5 _29828_ (.a(_02259_),
    .b(_02320_),
    .c(_02310_),
    .o1(_04048_));
 b15nand02as1n08x5 _29829_ (.a(net710),
    .b(net702),
    .o1(_04049_));
 b15aoi112al1n04x5 _29830_ (.a(net709),
    .b(_02471_),
    .c(_04049_),
    .d(_02374_),
    .o1(_04050_));
 b15nor002an1n06x5 _29831_ (.a(_02324_),
    .b(_02390_),
    .o1(_04051_));
 b15inv000ah1n05x5 _29832_ (.a(\us12.a[4] ),
    .o1(_04052_));
 b15norp02as1n03x5 _29833_ (.a(_04052_),
    .b(_02327_),
    .o1(_04053_));
 b15aoi112ah1n03x5 _29834_ (.a(_04048_),
    .b(_04050_),
    .c(_04051_),
    .d(_04053_),
    .o1(_04054_));
 b15nand04an1n08x5 _29835_ (.a(_04041_),
    .b(_04043_),
    .c(_04046_),
    .d(_04054_),
    .o1(_04055_));
 b15nor002ar1n02x5 _29836_ (.a(net696),
    .b(_02457_),
    .o1(_04056_));
 b15norp03aq1n02x5 _29837_ (.a(_02298_),
    .b(_02310_),
    .c(_02460_),
    .o1(_04057_));
 b15oai112as1n06x5 _29838_ (.a(net709),
    .b(_02430_),
    .c(_04056_),
    .d(_04057_),
    .o1(_04059_));
 b15nanb02aq1n12x5 _29839_ (.a(net696),
    .b(net691),
    .out0(_04060_));
 b15norp03al1n02x5 _29840_ (.a(net709),
    .b(_02279_),
    .c(_04060_),
    .o1(_04061_));
 b15aoai13ah1n03x5 _29841_ (.a(net710),
    .b(_04061_),
    .c(_03758_),
    .d(_02411_),
    .o1(_04062_));
 b15aoi022ah1n06x5 _29842_ (.a(_02321_),
    .b(_03670_),
    .c(_03711_),
    .d(net715),
    .o1(_04063_));
 b15nand02ah1n03x5 _29843_ (.a(net694),
    .b(_02367_),
    .o1(_04064_));
 b15oai112ah1n12x5 _29844_ (.a(_04059_),
    .b(_04062_),
    .c(_04063_),
    .d(_04064_),
    .o1(_04065_));
 b15nandp2as1n04x5 _29845_ (.a(net704),
    .b(_02350_),
    .o1(_04066_));
 b15xor002as1n03x5 _29846_ (.a(net694),
    .b(net713),
    .out0(_04067_));
 b15mdn022ar1n02x5 _29847_ (.a(_02333_),
    .b(_02346_),
    .o1(_04068_),
    .sa(_04067_));
 b15norp03an1n03x5 _29848_ (.a(net692),
    .b(_04066_),
    .c(_04068_),
    .o1(_04070_));
 b15nand04al1n02x5 _29849_ (.a(_02298_),
    .b(net703),
    .c(_02365_),
    .d(_02333_),
    .o1(_04071_));
 b15oai012an1n04x5 _29850_ (.a(_04071_),
    .b(_03662_),
    .c(_02298_),
    .o1(_04072_));
 b15aoi012ah1n02x5 _29851_ (.a(_04070_),
    .b(_04072_),
    .c(_02426_),
    .o1(_04073_));
 b15nanb02aq1n12x5 _29852_ (.a(net713),
    .b(net703),
    .out0(_04074_));
 b15norp03ah1n08x5 _29853_ (.a(_02242_),
    .b(_02290_),
    .c(_04074_),
    .o1(_04075_));
 b15nor004as1n04x5 _29854_ (.a(_02242_),
    .b(_02309_),
    .c(_02320_),
    .d(_02310_),
    .o1(_04076_));
 b15aoi112an1n08x5 _29855_ (.a(_04075_),
    .b(_04076_),
    .c(_02328_),
    .d(_03689_),
    .o1(_04077_));
 b15nand03ar1n03x5 _29856_ (.a(_02461_),
    .b(_02319_),
    .c(_02460_),
    .o1(_04078_));
 b15nandp2ah1n03x5 _29857_ (.a(_02321_),
    .b(_03679_),
    .o1(_04079_));
 b15oai022an1n06x5 _29858_ (.a(_02366_),
    .b(_02468_),
    .c(_02438_),
    .d(_04079_),
    .o1(_04081_));
 b15nano23ar1n02x5 _29859_ (.a(_04077_),
    .b(_04078_),
    .c(_04081_),
    .d(_02440_),
    .out0(_04082_));
 b15nona23as1n02x5 _29860_ (.a(_04055_),
    .b(_04065_),
    .c(_04073_),
    .d(_04082_),
    .out0(_04083_));
 b15aoai13ar1n02x5 _29861_ (.a(net696),
    .b(_02365_),
    .c(_02341_),
    .d(net710),
    .o1(_04084_));
 b15nonb02ah1n08x5 _29862_ (.a(net710),
    .b(net696),
    .out0(_04085_));
 b15nand02ar1n02x5 _29863_ (.a(_02293_),
    .b(_04085_),
    .o1(_04086_));
 b15aoi112an1n02x5 _29864_ (.a(net699),
    .b(_02389_),
    .c(_04084_),
    .d(_04086_),
    .o1(_04087_));
 b15nonb02ah1n03x5 _29865_ (.a(net696),
    .b(net694),
    .out0(_04088_));
 b15ztpn00an1n08x5 TAP_417 ();
 b15nonb03ar1n02x5 _29867_ (.a(net699),
    .b(net691),
    .c(net703),
    .out0(_04090_));
 b15nano22ar1n02x5 _29868_ (.a(net691),
    .b(net703),
    .c(net699),
    .out0(_04092_));
 b15oai112al1n02x5 _29869_ (.a(net706),
    .b(_04088_),
    .c(_04090_),
    .d(_04092_),
    .o1(_04093_));
 b15nand04al1n02x5 _29870_ (.a(net691),
    .b(net694),
    .c(net703),
    .d(_02291_),
    .o1(_04094_));
 b15aoi012ah1n02x5 _29871_ (.a(net710),
    .b(_04093_),
    .c(_04094_),
    .o1(_04095_));
 b15oai012al1n06x5 _29872_ (.a(net713),
    .b(_04087_),
    .c(_04095_),
    .o1(_04096_));
 b15nor002al1n03x5 _29873_ (.a(_02276_),
    .b(_02318_),
    .o1(_04097_));
 b15aoi022ah1n08x5 _29874_ (.a(net714),
    .b(_02293_),
    .c(_03727_),
    .d(net693),
    .o1(_04098_));
 b15oai022an1n08x5 _29875_ (.a(_02327_),
    .b(_02355_),
    .c(_04098_),
    .d(_02419_),
    .o1(_04099_));
 b15aoai13as1n08x5 _29876_ (.a(_02343_),
    .b(_04097_),
    .c(_04099_),
    .d(net699),
    .o1(_04100_));
 b15aoi013ar1n02x5 _29877_ (.a(_02381_),
    .b(_02365_),
    .c(_02346_),
    .d(_04016_),
    .o1(_04101_));
 b15and002an1n08x5 _29878_ (.a(net696),
    .b(net694),
    .o(_04103_));
 b15nano22al1n02x5 _29879_ (.a(net691),
    .b(net707),
    .c(net699),
    .out0(_04104_));
 b15norp02aq1n02x5 _29880_ (.a(net691),
    .b(net707),
    .o1(_04105_));
 b15aoai13ah1n04x5 _29881_ (.a(_04103_),
    .b(_04104_),
    .c(net699),
    .d(_04105_),
    .o1(_04106_));
 b15aoi022ar1n02x5 _29882_ (.a(_02333_),
    .b(_02375_),
    .c(_02475_),
    .d(_03655_),
    .o1(_04107_));
 b15aoai13ar1n02x5 _29883_ (.a(_04101_),
    .b(net710),
    .c(_04106_),
    .d(_04107_),
    .o1(_04108_));
 b15nand04aq1n16x5 _29884_ (.a(net706),
    .b(_02291_),
    .c(_02293_),
    .d(_02449_),
    .o1(_04109_));
 b15nand03aq1n16x5 _29885_ (.a(_02461_),
    .b(_02291_),
    .c(_02293_),
    .o1(_04110_));
 b15nand02an1n04x5 _29886_ (.a(net706),
    .b(_02425_),
    .o1(_04111_));
 b15aoai13as1n08x5 _29887_ (.a(_04109_),
    .b(_03657_),
    .c(_04110_),
    .d(_04111_),
    .o1(_04112_));
 b15oai012as1n03x5 _29888_ (.a(_04108_),
    .b(_04112_),
    .c(net703),
    .o1(_04114_));
 b15nand03al1n16x5 _29889_ (.a(_02381_),
    .b(_02341_),
    .c(_02346_),
    .o1(_04115_));
 b15nandp2ar1n03x5 _29890_ (.a(_02437_),
    .b(_02375_),
    .o1(_04116_));
 b15oaoi13an1n04x5 _29891_ (.a(net712),
    .b(_04115_),
    .c(_04116_),
    .d(net714),
    .o1(_04117_));
 b15aoi022as1n08x5 _29892_ (.a(_02286_),
    .b(_02313_),
    .c(_02354_),
    .d(_03679_),
    .o1(_04118_));
 b15nor002aq1n04x5 _29893_ (.a(net698),
    .b(net694),
    .o1(_04119_));
 b15norp03ar1n02x5 _29894_ (.a(\us12.a[4] ),
    .b(net693),
    .c(net714),
    .o1(_04120_));
 b15oai112aq1n04x5 _29895_ (.a(_02251_),
    .b(_04119_),
    .c(_03725_),
    .d(_04120_),
    .o1(_04121_));
 b15aoi012an1n04x5 _29896_ (.a(_02242_),
    .b(_04118_),
    .c(_04121_),
    .o1(_04122_));
 b15aoi013as1n02x5 _29897_ (.a(net701),
    .b(_02341_),
    .c(_02437_),
    .d(net714),
    .o1(_04123_));
 b15inv040ah1n02x5 _29898_ (.a(\us12.a[6] ),
    .o1(_04125_));
 b15nandp2ah1n04x5 _29899_ (.a(net698),
    .b(_04125_),
    .o1(_04126_));
 b15nanb02ah1n04x5 _29900_ (.a(net693),
    .b(\us12.a[4] ),
    .out0(_04127_));
 b15nanb02al1n06x5 _29901_ (.a(\us12.a[4] ),
    .b(net693),
    .out0(_04128_));
 b15nandp2al1n08x5 _29902_ (.a(_04127_),
    .b(_04128_),
    .o1(_04129_));
 b15oaoi13ah1n04x5 _29903_ (.a(_04123_),
    .b(net701),
    .c(_04126_),
    .d(_04129_),
    .o1(_04130_));
 b15aoi112as1n08x5 _29904_ (.a(_04117_),
    .b(_04122_),
    .c(_02415_),
    .d(_04130_),
    .o1(_04131_));
 b15nand04ah1n08x5 _29905_ (.a(_04096_),
    .b(_04100_),
    .c(_04114_),
    .d(_04131_),
    .o1(_04132_));
 b15nor003aq1n06x5 _29906_ (.a(_04040_),
    .b(_04083_),
    .c(_04132_),
    .o1(_04133_));
 b15nona22ar1n02x5 _29907_ (.a(net828),
    .b(net839),
    .c(net822),
    .out0(_04134_));
 b15aoi112an1n03x5 _29908_ (.a(net824),
    .b(_02569_),
    .c(_03404_),
    .d(_04134_),
    .o1(_04136_));
 b15and003ar1n02x5 _29909_ (.a(net825),
    .b(_02620_),
    .c(_03577_),
    .o(_04137_));
 b15nor004al1n08x5 _29910_ (.a(_03305_),
    .b(_02569_),
    .c(_02566_),
    .d(_02666_),
    .o1(_04138_));
 b15oai013aq1n02x5 _29911_ (.a(net826),
    .b(_04136_),
    .c(_04137_),
    .d(_04138_),
    .o1(_04139_));
 b15oai112an1n06x5 _29912_ (.a(net831),
    .b(_04139_),
    .c(_02700_),
    .d(net833),
    .o1(_04140_));
 b15aoi112ar1n02x5 _29913_ (.a(net833),
    .b(_02757_),
    .c(_03370_),
    .d(net839),
    .o1(_04141_));
 b15aoi012ah1n02x5 _29914_ (.a(_04141_),
    .b(_02593_),
    .c(net833),
    .o1(_04142_));
 b15oai112an1n12x5 _29915_ (.a(net840),
    .b(_04140_),
    .c(_04142_),
    .d(net831),
    .o1(_04143_));
 b15oai012ar1n04x5 _29916_ (.a(_03317_),
    .b(_03330_),
    .c(net826),
    .o1(_04144_));
 b15nand03an1n08x5 _29917_ (.a(_02620_),
    .b(_03402_),
    .c(_04144_),
    .o1(_04145_));
 b15aoai13as1n02x5 _29918_ (.a(net838),
    .b(_03341_),
    .c(_03397_),
    .d(_03592_),
    .o1(_04147_));
 b15aoi012al1n06x5 _29919_ (.a(net834),
    .b(_04145_),
    .c(_04147_),
    .o1(_04148_));
 b15aoi012ah1n02x5 _29920_ (.a(_02611_),
    .b(_02573_),
    .c(_02759_),
    .o1(_04149_));
 b15norp02aq1n03x5 _29921_ (.a(net840),
    .b(_02598_),
    .o1(_04150_));
 b15aoi112ah1n06x5 _29922_ (.a(_02716_),
    .b(_04149_),
    .c(_04150_),
    .d(_03617_),
    .o1(_04151_));
 b15norp02ar1n02x5 _29923_ (.a(net831),
    .b(_02515_),
    .o1(_04152_));
 b15aoai13an1n02x5 _29924_ (.a(net840),
    .b(_04152_),
    .c(_03341_),
    .d(net831),
    .o1(_04153_));
 b15inv000al1n02x5 _29925_ (.a(_03355_),
    .o1(_04154_));
 b15oai012ar1n02x5 _29926_ (.a(_02716_),
    .b(net833),
    .c(net828),
    .o1(_04155_));
 b15aoi022as1n04x5 _29927_ (.a(net831),
    .b(_04154_),
    .c(_04155_),
    .d(net822),
    .o1(_04156_));
 b15oai013ar1n08x5 _29928_ (.a(_04153_),
    .b(_04156_),
    .c(net825),
    .d(net826),
    .o1(_04158_));
 b15aoi112an1n06x5 _29929_ (.a(_04148_),
    .b(_04151_),
    .c(_04158_),
    .d(_02573_),
    .o1(_04159_));
 b15ztpn00an1n08x5 TAP_416 ();
 b15aoai13as1n06x5 _29931_ (.a(_03391_),
    .b(_02757_),
    .c(_02562_),
    .d(_03602_),
    .o1(_04161_));
 b15inv000ah1n10x5 _29932_ (.a(\us01.a[7] ),
    .o1(_04162_));
 b15nor003an1n06x5 _29933_ (.a(net824),
    .b(_02616_),
    .c(_02643_),
    .o1(_04163_));
 b15norp02as1n03x5 _29934_ (.a(net839),
    .b(_02656_),
    .o1(_04164_));
 b15oai112as1n16x5 _29935_ (.a(_04162_),
    .b(_02709_),
    .c(_04163_),
    .d(_04164_),
    .o1(_04165_));
 b15aoi022aq1n08x5 _29936_ (.a(net831),
    .b(_02757_),
    .c(_02732_),
    .d(_02616_),
    .o1(_04166_));
 b15oai112as1n16x5 _29937_ (.a(_04161_),
    .b(_04165_),
    .c(_04166_),
    .d(net833),
    .o1(_04167_));
 b15norp02aq1n02x5 _29938_ (.a(net828),
    .b(_02547_),
    .o1(_04169_));
 b15nona23ar1n02x5 _29939_ (.a(net825),
    .b(net840),
    .c(net839),
    .d(net828),
    .out0(_04170_));
 b15oaoi13ah1n02x5 _29940_ (.a(net822),
    .b(_04170_),
    .c(_02526_),
    .d(_03563_),
    .o1(_04171_));
 b15oai112al1n08x5 _29941_ (.a(_02615_),
    .b(_03391_),
    .c(_04169_),
    .d(_04171_),
    .o1(_04172_));
 b15nor003ar1n02x5 _29942_ (.a(_02631_),
    .b(_02562_),
    .c(_02692_),
    .o1(_04173_));
 b15nand02ar1n24x5 _29943_ (.a(net824),
    .b(net840),
    .o1(_04174_));
 b15nor004ar1n08x5 _29944_ (.a(_02615_),
    .b(net822),
    .c(net831),
    .d(_04174_),
    .o1(_04175_));
 b15oai013ah1n02x5 _29945_ (.a(net833),
    .b(_02732_),
    .c(_04173_),
    .d(_04175_),
    .o1(_04176_));
 b15oai012ar1n02x5 _29946_ (.a(net833),
    .b(net831),
    .c(_02649_),
    .o1(_04177_));
 b15nor002al1n12x5 _29947_ (.a(net832),
    .b(_02768_),
    .o1(_04178_));
 b15aoai13ah1n02x5 _29948_ (.a(_04177_),
    .b(_02598_),
    .c(_02616_),
    .d(_04178_),
    .o1(_04180_));
 b15oaoi13al1n03x5 _29949_ (.a(_02611_),
    .b(_02609_),
    .c(_02654_),
    .d(net839),
    .o1(_04181_));
 b15oai112ah1n06x5 _29950_ (.a(_04172_),
    .b(_04176_),
    .c(_04180_),
    .d(_04181_),
    .o1(_04182_));
 b15aoi022ar1n02x5 _29951_ (.a(_03391_),
    .b(_02748_),
    .c(_04175_),
    .d(net828),
    .o1(_04183_));
 b15nandp2ah1n08x5 _29952_ (.a(_02611_),
    .b(net830),
    .o1(_04184_));
 b15aoi022ar1n04x5 _29953_ (.a(_03391_),
    .b(_03598_),
    .c(_04184_),
    .d(_03340_),
    .o1(_04185_));
 b15aoi012ar1n02x5 _29954_ (.a(_02573_),
    .b(_04183_),
    .c(_04185_),
    .o1(_04186_));
 b15norp02aq1n12x5 _29955_ (.a(_02573_),
    .b(_02768_),
    .o1(_04187_));
 b15nor002as1n02x5 _29956_ (.a(\us01.a[0] ),
    .b(_02515_),
    .o1(_04188_));
 b15aoai13as1n02x5 _29957_ (.a(_02709_),
    .b(_04187_),
    .c(_02573_),
    .d(_04188_),
    .o1(_04189_));
 b15nor002ah1n02x5 _29958_ (.a(net831),
    .b(_02623_),
    .o1(_04191_));
 b15oai022ah1n04x5 _29959_ (.a(_02526_),
    .b(_02595_),
    .c(_02616_),
    .d(_02643_),
    .o1(_04192_));
 b15nor002al1n02x5 _29960_ (.a(net826),
    .b(net822),
    .o1(_04193_));
 b15aob012as1n02x5 _29961_ (.a(_02681_),
    .b(_04193_),
    .c(_03626_),
    .out0(_04194_));
 b15nor003ah1n03x5 _29962_ (.a(net828),
    .b(_03563_),
    .c(_02695_),
    .o1(_04195_));
 b15aoi022aq1n12x5 _29963_ (.a(_04191_),
    .b(_04192_),
    .c(_04194_),
    .d(_04195_),
    .o1(_04196_));
 b15aoi012al1n02x5 _29964_ (.a(\us01.a[0] ),
    .b(_03366_),
    .c(_02554_),
    .o1(_04197_));
 b15nand04as1n04x5 _29965_ (.a(_02631_),
    .b(_02517_),
    .c(_02529_),
    .d(_03549_),
    .o1(_04198_));
 b15nanb03aq1n06x5 _29966_ (.a(net835),
    .b(net839),
    .c(\us01.a[0] ),
    .out0(_04199_));
 b15nand04aq1n04x5 _29967_ (.a(\us01.a[3] ),
    .b(_03302_),
    .c(_02529_),
    .d(_04199_),
    .o1(_04200_));
 b15aoi012ar1n06x5 _29968_ (.a(_04197_),
    .b(_04198_),
    .c(_04200_),
    .o1(_04202_));
 b15nand03aq1n03x5 _29969_ (.a(\us01.a[3] ),
    .b(_02517_),
    .c(_02529_),
    .o1(_04203_));
 b15mdn022ah1n02x5 _29970_ (.a(_03366_),
    .b(_03376_),
    .o1(_04204_),
    .sa(_02611_));
 b15mdn022aq1n03x5 _29971_ (.a(_03602_),
    .b(_02635_),
    .o1(_04205_),
    .sa(_02631_));
 b15oai022an1n08x5 _29972_ (.a(_04203_),
    .b(_04204_),
    .c(_04205_),
    .d(_03366_),
    .o1(_04206_));
 b15nano23al1n12x5 _29973_ (.a(_04189_),
    .b(_04196_),
    .c(_04202_),
    .d(_04206_),
    .out0(_04207_));
 b15aoi012ar1n02x5 _29974_ (.a(\us01.a[6] ),
    .b(net839),
    .c(net828),
    .o1(_04208_));
 b15nand03al1n04x5 _29975_ (.a(_03626_),
    .b(_02694_),
    .c(_04208_),
    .o1(_04209_));
 b15qgbna2an1n05x5 _29976_ (.o1(_04210_),
    .a(_02684_),
    .b(_03592_));
 b15oai112al1n08x5 _29977_ (.a(_04209_),
    .b(_04210_),
    .c(_02602_),
    .d(_03605_),
    .o1(_04211_));
 b15aoi013ar1n02x5 _29978_ (.a(_03598_),
    .b(_04193_),
    .c(net825),
    .d(_02569_),
    .o1(_04213_));
 b15oai022ah1n02x5 _29979_ (.a(_02526_),
    .b(_03362_),
    .c(_04213_),
    .d(_02616_),
    .o1(_04214_));
 b15oai012al1n06x5 _29980_ (.a(net831),
    .b(_04211_),
    .c(_04214_),
    .o1(_04215_));
 b15nona23ah1n12x5 _29981_ (.a(_04182_),
    .b(_04186_),
    .c(_04207_),
    .d(_04215_),
    .out0(_04216_));
 b15nano23as1n24x5 _29982_ (.a(_04143_),
    .b(_04159_),
    .c(_04167_),
    .d(_04216_),
    .out0(_04217_));
 b15qgbxo2an1n10x5 _29983_ (.a(net399),
    .b(_04217_),
    .out0(_04218_));
 b15xor002an1n03x5 _29984_ (.a(net392),
    .b(_04218_),
    .out0(_04219_));
 b15nandp2ar1n03x5 _29985_ (.a(net853),
    .b(_02782_),
    .o1(_04220_));
 b15nandp2ar1n32x5 _29986_ (.a(_02854_),
    .b(_03018_),
    .o1(_04221_));
 b15oaoi13ar1n02x5 _29987_ (.a(net859),
    .b(_04220_),
    .c(_04221_),
    .d(net860),
    .o1(_04222_));
 b15norp02ar1n02x5 _29988_ (.a(_02871_),
    .b(_04221_),
    .o1(_04224_));
 b15norp03ah1n03x5 _29989_ (.a(\us30.a[3] ),
    .b(_04222_),
    .c(_04224_),
    .o1(_04225_));
 b15oai022ar1n02x5 _29990_ (.a(net853),
    .b(_02913_),
    .c(_03463_),
    .d(net862),
    .o1(_04226_));
 b15orn002al1n32x5 _29991_ (.a(\us30.a[0] ),
    .b(net856),
    .o(_04227_));
 b15oai122an1n08x5 _29992_ (.a(net843),
    .b(_02879_),
    .c(_02882_),
    .d(_03482_),
    .e(_04227_),
    .o1(_04228_));
 b15oai022as1n02x5 _29993_ (.a(_02854_),
    .b(_02798_),
    .c(_02897_),
    .d(net862),
    .o1(_04229_));
 b15oai112al1n12x5 _29994_ (.a(net859),
    .b(_04228_),
    .c(_04229_),
    .d(net843),
    .o1(_04230_));
 b15ztpn00an1n08x5 TAP_415 ();
 b15aoi022as1n06x5 _29996_ (.a(_02854_),
    .b(_02779_),
    .c(_03002_),
    .d(_02899_),
    .o1(_04232_));
 b15and003ar1n02x5 _29997_ (.a(_02824_),
    .b(_03002_),
    .c(_03010_),
    .o(_04233_));
 b15oai012aq1n03x5 _29998_ (.a(_02879_),
    .b(_03482_),
    .c(_02854_),
    .o1(_04235_));
 b15aoi013ah1n04x5 _29999_ (.a(_04233_),
    .b(_04235_),
    .c(_02882_),
    .d(net843),
    .o1(_04236_));
 b15oai122as1n16x5 _30000_ (.a(_04230_),
    .b(_04232_),
    .c(net843),
    .d(_04236_),
    .e(net859),
    .o1(_04237_));
 b15aoi022an1n02x5 _30001_ (.a(_02923_),
    .b(_04226_),
    .c(_04237_),
    .d(net844),
    .o1(_04238_));
 b15aoi012ar1n06x5 _30002_ (.a(_04225_),
    .b(_04238_),
    .c(\us30.a[3] ),
    .o1(_04239_));
 b15oai022ar1n02x5 _30003_ (.a(_02986_),
    .b(_02867_),
    .c(_02913_),
    .d(net850),
    .o1(_04240_));
 b15aoi022an1n02x5 _30004_ (.a(_02799_),
    .b(_03466_),
    .c(_04240_),
    .d(net857),
    .o1(_04241_));
 b15oai012an1n06x5 _30005_ (.a(_03541_),
    .b(_04241_),
    .c(net854),
    .o1(_04242_));
 b15nanb02ah1n24x5 _30006_ (.a(net860),
    .b(net853),
    .out0(_04243_));
 b15aoi012an1n02x5 _30007_ (.a(_02951_),
    .b(_04243_),
    .c(_03514_),
    .o1(_04244_));
 b15oai012as1n02x5 _30008_ (.a(_03023_),
    .b(_04244_),
    .c(_02941_),
    .o1(_04246_));
 b15nor003ar1n06x5 _30009_ (.a(_02880_),
    .b(_03482_),
    .c(_02935_),
    .o1(_04247_));
 b15nor004ar1n02x5 _30010_ (.a(net846),
    .b(net848),
    .c(_02940_),
    .d(_02880_),
    .o1(_04248_));
 b15oai012ar1n02x5 _30011_ (.a(net862),
    .b(_04247_),
    .c(_04248_),
    .o1(_04249_));
 b15norp02as1n04x5 _30012_ (.a(net856),
    .b(net844),
    .o1(_04250_));
 b15nor004an1n02x5 _30013_ (.a(_02897_),
    .b(_02871_),
    .c(_02968_),
    .d(_04250_),
    .o1(_04251_));
 b15aoi012ar1n02x5 _30014_ (.a(_04251_),
    .b(_04247_),
    .c(_02811_),
    .o1(_04252_));
 b15nanb02an1n03x5 _30015_ (.a(net848),
    .b(\us30.a[7] ),
    .out0(_04253_));
 b15norp02ar1n02x5 _30016_ (.a(_04227_),
    .b(_04253_),
    .o1(_04254_));
 b15nandp3ar1n02x5 _30017_ (.a(net852),
    .b(net847),
    .c(net844),
    .o1(_04255_));
 b15oai013ar1n02x5 _30018_ (.a(_04255_),
    .b(_02956_),
    .c(net844),
    .d(net846),
    .o1(_04257_));
 b15oai012as1n04x5 _30019_ (.a(_02864_),
    .b(_03469_),
    .c(net857),
    .o1(_04258_));
 b15aoi022ar1n02x5 _30020_ (.a(_04254_),
    .b(_04257_),
    .c(_04258_),
    .d(_02974_),
    .o1(_04259_));
 b15andc04ar1n02x5 _30021_ (.a(_04246_),
    .b(_04249_),
    .c(_04252_),
    .d(_04259_),
    .o(_04260_));
 b15nona23aq1n02x5 _30022_ (.a(net856),
    .b(net848),
    .c(_02904_),
    .d(_02947_),
    .out0(_04261_));
 b15nonb02ar1n02x5 _30023_ (.a(net852),
    .b(\us30.a[7] ),
    .out0(_04262_));
 b15nonb02al1n04x5 _30024_ (.a(\us30.a[7] ),
    .b(net852),
    .out0(_04263_));
 b15aoi012as1n02x5 _30025_ (.a(_04262_),
    .b(_04263_),
    .c(_02820_),
    .o1(_04264_));
 b15nanb02as1n12x5 _30026_ (.a(\us30.a[2] ),
    .b(\us30.a[1] ),
    .out0(_04265_));
 b15inv040as1n06x5 _30027_ (.a(net844),
    .o1(_04266_));
 b15nandp2ar1n05x5 _30028_ (.a(net848),
    .b(_04266_),
    .o1(_04268_));
 b15oai013as1n06x5 _30029_ (.a(_04261_),
    .b(_04264_),
    .c(_04265_),
    .d(_04268_),
    .o1(_04269_));
 b15nor003an1n03x5 _30030_ (.a(net847),
    .b(\us30.a[6] ),
    .c(_02995_),
    .o1(_04270_));
 b15oai022aq1n02x5 _30031_ (.a(net852),
    .b(_02856_),
    .c(_04253_),
    .d(_03514_),
    .o1(_04271_));
 b15nandp2ar1n02x5 _30032_ (.a(net847),
    .b(_02791_),
    .o1(_04272_));
 b15oai013al1n04x5 _30033_ (.a(_02942_),
    .b(_04272_),
    .c(net848),
    .d(_02880_),
    .o1(_04273_));
 b15aoi222ah1n06x5 _30034_ (.a(_02824_),
    .b(_04269_),
    .c(_04270_),
    .d(_04271_),
    .e(_04273_),
    .f(_02877_),
    .o1(_04274_));
 b15aoai13ar1n02x5 _30035_ (.a(net852),
    .b(_02989_),
    .c(_02877_),
    .d(net856),
    .o1(_04275_));
 b15oai012ar1n02x5 _30036_ (.a(net861),
    .b(_02791_),
    .c(_02977_),
    .o1(_04276_));
 b15aoi012ar1n02x5 _30037_ (.a(_02876_),
    .b(_04275_),
    .c(_04276_),
    .o1(_04277_));
 b15aoi012ar1n02x5 _30038_ (.a(_02779_),
    .b(_02899_),
    .c(_02820_),
    .o1(_04279_));
 b15oai022ar1n04x5 _30039_ (.a(net862),
    .b(_02897_),
    .c(_04279_),
    .d(net859),
    .o1(_04280_));
 b15aoi013ar1n03x5 _30040_ (.a(_04277_),
    .b(_04280_),
    .c(_02904_),
    .d(_02791_),
    .o1(_04281_));
 b15aoi012ah1n04x5 _30041_ (.a(_03452_),
    .b(_02957_),
    .c(_02854_),
    .o1(_04282_));
 b15oai012ah1n06x5 _30042_ (.a(_02811_),
    .b(_02919_),
    .c(_03024_),
    .o1(_04283_));
 b15oaoi13an1n04x5 _30043_ (.a(_02951_),
    .b(_02882_),
    .c(_03024_),
    .d(net855),
    .o1(_04284_));
 b15nor003as1n12x5 _30044_ (.a(_04282_),
    .b(_04283_),
    .c(_04284_),
    .o1(_04285_));
 b15nand04al1n16x5 _30045_ (.a(net862),
    .b(_02854_),
    .c(_02899_),
    .d(_02781_),
    .o1(_04286_));
 b15and002ar1n02x5 _30046_ (.a(net856),
    .b(net844),
    .o(_04287_));
 b15aoi012ar1n02x5 _30047_ (.a(_04287_),
    .b(_04250_),
    .c(\us30.a[1] ),
    .o1(_04288_));
 b15nand02ar1n02x5 _30048_ (.a(_02820_),
    .b(net843),
    .o1(_04290_));
 b15oai013al1n02x5 _30049_ (.a(_04286_),
    .b(_04288_),
    .c(_04290_),
    .d(_02897_),
    .o1(_04291_));
 b15aoi012al1n02x5 _30050_ (.a(_04285_),
    .b(_04291_),
    .c(net852),
    .o1(_04292_));
 b15nand04an1n06x5 _30051_ (.a(_04260_),
    .b(_04274_),
    .c(_04281_),
    .d(_04292_),
    .o1(_04293_));
 b15orn002as1n04x5 _30052_ (.a(_04242_),
    .b(_04293_),
    .o(_04294_));
 b15nandp3ar1n02x5 _30053_ (.a(_02811_),
    .b(_02932_),
    .c(_02989_),
    .o1(_04295_));
 b15ztpn00an1n08x5 TAP_414 ();
 b15oaoi13al1n02x5 _30055_ (.a(net860),
    .b(_04295_),
    .c(_03521_),
    .d(_02951_),
    .o1(_04297_));
 b15nonb02aq1n04x5 _30056_ (.a(net861),
    .b(net854),
    .out0(_04298_));
 b15nano22ar1n03x5 _30057_ (.a(net849),
    .b(net843),
    .c(net846),
    .out0(_04299_));
 b15and002al1n04x5 _30058_ (.a(_04298_),
    .b(_04299_),
    .o(_04301_));
 b15norp02ar1n32x5 _30059_ (.a(net860),
    .b(_02854_),
    .o1(_04302_));
 b15aoi013ar1n06x5 _30060_ (.a(_04301_),
    .b(_03010_),
    .c(_04302_),
    .d(net847),
    .o1(_04303_));
 b15nor003as1n03x5 _30061_ (.a(net850),
    .b(_04266_),
    .c(_04303_),
    .o1(_04304_));
 b15oaoi13ar1n02x5 _30062_ (.a(_02858_),
    .b(_04220_),
    .c(net853),
    .d(_02986_),
    .o1(_04305_));
 b15aoi012ah1n02x5 _30063_ (.a(_03447_),
    .b(_03427_),
    .c(_02954_),
    .o1(_04306_));
 b15nor004aq1n03x5 _30064_ (.a(_04297_),
    .b(_04304_),
    .c(_04305_),
    .d(_04306_),
    .o1(_04307_));
 b15xor002ar1n02x5 _30065_ (.a(net852),
    .b(net845),
    .out0(_04308_));
 b15nano22an1n05x5 _30066_ (.a(_03010_),
    .b(_03000_),
    .c(_04308_),
    .out0(_04309_));
 b15aoi013ar1n02x5 _30067_ (.a(_04309_),
    .b(_02932_),
    .c(_02947_),
    .d(net853),
    .o1(_04310_));
 b15oai112an1n04x5 _30068_ (.a(net858),
    .b(_04310_),
    .c(_02964_),
    .d(_04243_),
    .o1(_04312_));
 b15oai022ar1n04x5 _30069_ (.a(_02940_),
    .b(_02954_),
    .c(_02964_),
    .d(_03514_),
    .o1(_04313_));
 b15oai012al1n06x5 _30070_ (.a(_04312_),
    .b(_04313_),
    .c(net858),
    .o1(_04314_));
 b15oai122aq1n08x5 _30071_ (.a(net851),
    .b(_02918_),
    .c(_02985_),
    .d(_02989_),
    .e(_02862_),
    .o1(_04315_));
 b15oai022an1n02x5 _30072_ (.a(_03020_),
    .b(_02913_),
    .c(_02929_),
    .d(_04243_),
    .o1(_04316_));
 b15oai012ar1n06x5 _30073_ (.a(_04315_),
    .b(_04316_),
    .c(\us30.a[3] ),
    .o1(_04317_));
 b15nandp3al1n08x5 _30074_ (.a(_04307_),
    .b(_04314_),
    .c(_04317_),
    .o1(_04318_));
 b15orn003al1n24x5 _30075_ (.a(_04239_),
    .b(_04294_),
    .c(_04318_),
    .o(_04319_));
 b15xor002an1n03x5 _30076_ (.a(_03633_),
    .b(_04319_),
    .out0(_04320_));
 b15xor002an1n06x5 _30077_ (.a(_04219_),
    .b(_04320_),
    .out0(_04321_));
 b15cmbn22al1n08x5 _30078_ (.clk1(\text_in_r[66] ),
    .clk2(_04321_),
    .clkout(_04323_),
    .s(net537));
 b15xor002aq1n16x5 _30079_ (.a(\u0.w[1][2] ),
    .b(_04323_),
    .out0(_00107_));
 b15oai122aq1n04x5 _30080_ (.a(net703),
    .b(_02407_),
    .c(_03636_),
    .d(_04106_),
    .e(net713),
    .o1(_04324_));
 b15oaoi13as1n02x5 _30081_ (.a(_03651_),
    .b(_03699_),
    .c(net710),
    .d(_02500_),
    .o1(_04325_));
 b15nandp3ar1n02x5 _30082_ (.a(_02411_),
    .b(_02293_),
    .c(_02437_),
    .o1(_04326_));
 b15aoi013ar1n02x5 _30083_ (.a(_02462_),
    .b(_02437_),
    .c(_02293_),
    .d(net713),
    .o1(_04327_));
 b15oaoi13as1n02x5 _30084_ (.a(_02242_),
    .b(_04326_),
    .c(_04327_),
    .d(net706),
    .o1(_04328_));
 b15oai013an1n06x5 _30085_ (.a(_04324_),
    .b(_04325_),
    .c(_04328_),
    .d(net703),
    .o1(_04329_));
 b15nand02aq1n06x5 _30086_ (.a(_02461_),
    .b(_02354_),
    .o1(_04330_));
 b15oaoi13an1n02x5 _30087_ (.a(net704),
    .b(_04330_),
    .c(_03666_),
    .d(net713),
    .o1(_04331_));
 b15nandp3ah1n08x5 _30088_ (.a(_02341_),
    .b(_02346_),
    .c(_03645_),
    .o1(_04333_));
 b15oai122al1n04x5 _30089_ (.a(_04333_),
    .b(_04074_),
    .c(_02466_),
    .d(net703),
    .e(_03666_),
    .o1(_04334_));
 b15aoai13an1n02x5 _30090_ (.a(_02242_),
    .b(_04331_),
    .c(_04334_),
    .d(net707),
    .o1(_04335_));
 b15and002ar1n24x5 _30091_ (.a(net711),
    .b(net708),
    .o(_04336_));
 b15oai013an1n06x5 _30092_ (.a(_02469_),
    .b(_02427_),
    .c(_03648_),
    .d(_02259_),
    .o1(_04337_));
 b15aoi222ah1n12x5 _30093_ (.a(_04336_),
    .b(_04024_),
    .c(_03764_),
    .d(_02433_),
    .e(\us12.a[0] ),
    .f(_04337_),
    .o1(_04338_));
 b15norp02ar1n02x5 _30094_ (.a(net711),
    .b(_02469_),
    .o1(_04339_));
 b15aoai13ar1n04x5 _30095_ (.a(net715),
    .b(_04339_),
    .c(_02319_),
    .d(_02461_),
    .o1(_04340_));
 b15aoi122ar1n06x5 _30096_ (.a(net704),
    .b(_02319_),
    .c(_02433_),
    .d(_02350_),
    .e(_04024_),
    .o1(_04341_));
 b15aoi022as1n08x5 _30097_ (.a(net704),
    .b(_04338_),
    .c(_04340_),
    .d(_04341_),
    .o1(_04342_));
 b15oai013ar1n08x5 _30098_ (.a(_03677_),
    .b(_03695_),
    .c(_02317_),
    .d(_02381_),
    .o1(_04344_));
 b15aoi112ah1n06x5 _30099_ (.a(_02298_),
    .b(_04048_),
    .c(_04344_),
    .d(_02350_),
    .o1(_04345_));
 b15norp03ar1n02x5 _30100_ (.a(net711),
    .b(net708),
    .c(_02471_),
    .o1(_04346_));
 b15aoai13aq1n03x5 _30101_ (.a(net704),
    .b(_04346_),
    .c(_04336_),
    .d(_02425_),
    .o1(_04347_));
 b15nandp3al1n03x5 _30102_ (.a(net711),
    .b(net704),
    .c(_02319_),
    .o1(_04348_));
 b15aoi012aq1n02x5 _30103_ (.a(net715),
    .b(_02425_),
    .c(_02361_),
    .o1(_04349_));
 b15aoi022aq1n08x5 _30104_ (.a(_04345_),
    .b(_04347_),
    .c(_04348_),
    .d(_04349_),
    .o1(_04350_));
 b15nano23ar1n05x5 _30105_ (.a(_04329_),
    .b(_04335_),
    .c(_04342_),
    .d(_04350_),
    .out0(_04351_));
 b15norp02ar1n02x5 _30106_ (.a(_03706_),
    .b(_04128_),
    .o1(_04352_));
 b15oaoi13ar1n02x5 _30107_ (.a(_04127_),
    .b(_02273_),
    .c(net701),
    .d(net694),
    .o1(_04353_));
 b15oai012as1n03x5 _30108_ (.a(_04085_),
    .b(_04352_),
    .c(_04353_),
    .o1(_04355_));
 b15aoi022ah1n04x5 _30109_ (.a(net701),
    .b(_04044_),
    .c(_02351_),
    .d(net710),
    .o1(_04356_));
 b15oaoi13as1n08x5 _30110_ (.a(net706),
    .b(_04355_),
    .c(_04356_),
    .d(_02321_),
    .o1(_04357_));
 b15aoi013ar1n02x5 _30111_ (.a(net710),
    .b(_02343_),
    .c(_02291_),
    .d(_02293_),
    .o1(_04358_));
 b15nandp2ar1n12x5 _30112_ (.a(net713),
    .b(net702),
    .o1(_04359_));
 b15aoai13ar1n02x5 _30113_ (.a(_04358_),
    .b(_04359_),
    .c(_03699_),
    .d(_04110_),
    .o1(_04360_));
 b15oaoi13ar1n02x5 _30114_ (.a(net703),
    .b(_04110_),
    .c(_03651_),
    .d(_02366_),
    .o1(_04361_));
 b15oai012ar1n02x5 _30115_ (.a(net710),
    .b(_03699_),
    .c(_04074_),
    .o1(_04362_));
 b15oa0012al1n03x5 _30116_ (.a(_04360_),
    .b(_04361_),
    .c(_04362_),
    .o(_04363_));
 b15nor002an1n06x5 _30117_ (.a(_02381_),
    .b(_03673_),
    .o1(_04364_));
 b15oai022ar1n02x5 _30118_ (.a(_02242_),
    .b(_02324_),
    .c(_03657_),
    .d(_02357_),
    .o1(_04366_));
 b15aoi112aq1n02x5 _30119_ (.a(_04364_),
    .b(_03742_),
    .c(_04366_),
    .d(_02425_),
    .o1(_04367_));
 b15oai022ar1n02x5 _30120_ (.a(_04037_),
    .b(_02368_),
    .c(_02460_),
    .d(_02290_),
    .o1(_04368_));
 b15aob012aq1n02x5 _30121_ (.a(_04367_),
    .b(_04368_),
    .c(net715),
    .out0(_04369_));
 b15oaoi13ar1n02x5 _30122_ (.a(_02367_),
    .b(_02242_),
    .c(net703),
    .d(_02411_),
    .o1(_04370_));
 b15aoi022ar1n02x5 _30123_ (.a(net711),
    .b(_02367_),
    .c(_03680_),
    .d(net713),
    .o1(_04371_));
 b15oai022ar1n02x5 _30124_ (.a(_03677_),
    .b(_04370_),
    .c(_04371_),
    .d(_02438_),
    .o1(_04372_));
 b15nor004aq1n03x5 _30125_ (.a(_04357_),
    .b(_04363_),
    .c(_04369_),
    .d(_04372_),
    .o1(_04373_));
 b15nandp3ar1n02x5 _30126_ (.a(net711),
    .b(net704),
    .c(_02376_),
    .o1(_04374_));
 b15nand02aq1n03x5 _30127_ (.a(_02242_),
    .b(_02381_),
    .o1(_04375_));
 b15oaoi13an1n03x5 _30128_ (.a(net713),
    .b(_04374_),
    .c(_02366_),
    .d(_04375_),
    .o1(_04377_));
 b15and002as1n04x5 _30129_ (.a(net711),
    .b(net704),
    .o(_04378_));
 b15aoai13ar1n02x5 _30130_ (.a(net707),
    .b(_04377_),
    .c(_04378_),
    .d(_03688_),
    .o1(_04379_));
 b15norp03ar1n12x5 _30131_ (.a(_02381_),
    .b(_02317_),
    .c(_03695_),
    .o1(_04380_));
 b15norp03ah1n03x5 _30132_ (.a(_04052_),
    .b(_02276_),
    .c(_02279_),
    .o1(_04381_));
 b15nandp2aq1n03x5 _30133_ (.a(net698),
    .b(net712),
    .o1(_04382_));
 b15oai012ar1n08x5 _30134_ (.a(_04382_),
    .b(_02355_),
    .c(net698),
    .o1(_04383_));
 b15aoi022an1n12x5 _30135_ (.a(_02433_),
    .b(_04380_),
    .c(_04381_),
    .d(_04383_),
    .o1(_04384_));
 b15oa0012an1n02x5 _30136_ (.a(_04379_),
    .b(_04384_),
    .c(net707),
    .o(_04385_));
 b15nand02al1n04x5 _30137_ (.a(_02343_),
    .b(_04044_),
    .o1(_04386_));
 b15oai012al1n02x5 _30138_ (.a(_02471_),
    .b(_02327_),
    .c(_02318_),
    .o1(_04388_));
 b15aoi022as1n04x5 _30139_ (.a(_02367_),
    .b(_03670_),
    .c(_04388_),
    .d(_02251_),
    .o1(_04389_));
 b15aoai13as1n03x5 _30140_ (.a(net712),
    .b(_02311_),
    .c(_02351_),
    .d(net708),
    .o1(_04390_));
 b15aoi013ah1n06x5 _30141_ (.a(net715),
    .b(_04386_),
    .c(_04389_),
    .d(_04390_),
    .o1(_04391_));
 b15nandp3ar1n02x5 _30142_ (.a(_02461_),
    .b(net702),
    .c(_02376_),
    .o1(_04392_));
 b15aob012an1n04x5 _30143_ (.a(net710),
    .b(_03660_),
    .c(_04392_),
    .out0(_04393_));
 b15oai112al1n02x5 _30144_ (.a(_02343_),
    .b(_02340_),
    .c(_02376_),
    .d(_02313_),
    .o1(_04394_));
 b15nandp3ar1n02x5 _30145_ (.a(_02262_),
    .b(_02449_),
    .c(_04032_),
    .o1(_04395_));
 b15oai012al1n02x5 _30146_ (.a(_02286_),
    .b(_02328_),
    .c(_03758_),
    .o1(_04396_));
 b15nand04aq1n04x5 _30147_ (.a(_04393_),
    .b(_04394_),
    .c(_04395_),
    .d(_04396_),
    .o1(_04397_));
 b15oai022ar1n02x5 _30148_ (.a(_02366_),
    .b(_04049_),
    .c(_04115_),
    .d(net710),
    .o1(_04399_));
 b15and002an1n02x5 _30149_ (.a(net714),
    .b(_04399_),
    .o(_04400_));
 b15nand02an1n02x5 _30150_ (.a(net714),
    .b(_02475_),
    .o1(_04401_));
 b15oaoi13an1n08x5 _30151_ (.a(_02461_),
    .b(_04401_),
    .c(_03659_),
    .d(_02355_),
    .o1(_04402_));
 b15nor004aq1n08x5 _30152_ (.a(_04391_),
    .b(_04397_),
    .c(_04400_),
    .d(_04402_),
    .o1(_04403_));
 b15nand04ah1n08x5 _30153_ (.a(_04351_),
    .b(_04373_),
    .c(_04385_),
    .d(_04403_),
    .o1(_04404_));
 b15norp03ar1n02x5 _30154_ (.a(_02546_),
    .b(_02547_),
    .c(_02585_),
    .o1(_04405_));
 b15aoi012an1n02x5 _30155_ (.a(_04405_),
    .b(_02757_),
    .c(_02724_),
    .o1(_04406_));
 b15aoi112aq1n03x5 _30156_ (.a(_03341_),
    .b(_03573_),
    .c(_02664_),
    .d(_03370_),
    .o1(_04407_));
 b15oai022al1n08x5 _30157_ (.a(net835),
    .b(_04406_),
    .c(_04407_),
    .d(_02745_),
    .o1(_04408_));
 b15oai022ah1n08x5 _30158_ (.a(_03299_),
    .b(_02669_),
    .c(_04210_),
    .d(net831),
    .o1(_04410_));
 b15norp02ah1n04x5 _30159_ (.a(_02557_),
    .b(_02547_),
    .o1(_04411_));
 b15aoi022as1n04x5 _30160_ (.a(net836),
    .b(_04411_),
    .c(_02723_),
    .d(_02532_),
    .o1(_04412_));
 b15oabi12ar1n08x5 _30161_ (.a(_04410_),
    .b(_04412_),
    .c(_02716_),
    .out0(_04413_));
 b15aoai13ar1n02x5 _30162_ (.a(net839),
    .b(_03626_),
    .c(_02604_),
    .d(net840),
    .o1(_04414_));
 b15oaoi13ar1n02x5 _30163_ (.a(_02593_),
    .b(_04414_),
    .c(_02507_),
    .d(_02745_),
    .o1(_04415_));
 b15oai012ar1n02x5 _30164_ (.a(_02664_),
    .b(_02635_),
    .c(_03341_),
    .o1(_04416_));
 b15aoi022ar1n02x5 _30165_ (.a(_03391_),
    .b(_02665_),
    .c(_02709_),
    .d(net838),
    .o1(_04417_));
 b15oai012ar1n03x5 _30166_ (.a(_04416_),
    .b(_04417_),
    .c(_02728_),
    .o1(_04418_));
 b15oab012an1n02x5 _30167_ (.a(_03296_),
    .b(_03303_),
    .c(_02507_),
    .out0(_04419_));
 b15nona22an1n08x5 _30168_ (.a(_04415_),
    .b(_04418_),
    .c(_04419_),
    .out0(_04421_));
 b15oai022ar1n02x5 _30169_ (.a(_02595_),
    .b(_02541_),
    .c(_02643_),
    .d(_03549_),
    .o1(_04422_));
 b15aoi022al1n04x5 _30170_ (.a(_02541_),
    .b(_02635_),
    .c(_04422_),
    .d(_02666_),
    .o1(_04423_));
 b15norp03an1n02x5 _30171_ (.a(net835),
    .b(_02631_),
    .c(_02768_),
    .o1(_04424_));
 b15aoi012al1n04x5 _30172_ (.a(_04424_),
    .b(_02635_),
    .c(net835),
    .o1(_04425_));
 b15oai022ah1n06x5 _30173_ (.a(_02585_),
    .b(_04423_),
    .c(_04425_),
    .d(_02611_),
    .o1(_04426_));
 b15nor004al1n12x5 _30174_ (.a(_04408_),
    .b(_04413_),
    .c(_04421_),
    .d(_04426_),
    .o1(_04427_));
 b15aoi022ar1n02x5 _30175_ (.a(net838),
    .b(_02598_),
    .c(_04187_),
    .d(_03397_),
    .o1(_04428_));
 b15aoi012ar1n02x5 _30176_ (.a(_02598_),
    .b(_02637_),
    .c(_02573_),
    .o1(_04429_));
 b15oai013aq1n02x5 _30177_ (.a(_04428_),
    .b(_04429_),
    .c(net832),
    .d(net842),
    .o1(_04430_));
 b15nand02ar1n08x5 _30178_ (.a(net835),
    .b(_04430_),
    .o1(_04432_));
 b15oaoi13as1n02x5 _30179_ (.a(_03330_),
    .b(_03583_),
    .c(_02642_),
    .d(net835),
    .o1(_04433_));
 b15nand02ar1n02x5 _30180_ (.a(_02611_),
    .b(_03602_),
    .o1(_04434_));
 b15oaoi13ar1n02x5 _30181_ (.a(_02569_),
    .b(_04434_),
    .c(_03605_),
    .d(net832),
    .o1(_04435_));
 b15oab012an1n03x5 _30182_ (.a(net838),
    .b(_04433_),
    .c(_04435_),
    .out0(_04436_));
 b15oai012aq1n03x5 _30183_ (.a(_02569_),
    .b(_03341_),
    .c(_03351_),
    .o1(_04437_));
 b15oai013ar1n02x5 _30184_ (.a(net841),
    .b(net832),
    .c(_02515_),
    .d(_03549_),
    .o1(_04438_));
 b15aoi013an1n03x5 _30185_ (.a(_04438_),
    .b(_03409_),
    .c(_02664_),
    .d(_02573_),
    .o1(_04439_));
 b15nand02aq1n08x5 _30186_ (.a(_02709_),
    .b(_03409_),
    .o1(_04440_));
 b15aoi012al1n02x5 _30187_ (.a(net841),
    .b(_03391_),
    .c(_03373_),
    .o1(_04441_));
 b15aoi022ah1n06x5 _30188_ (.a(_04437_),
    .b(_04439_),
    .c(_04440_),
    .d(_04441_),
    .o1(_04443_));
 b15nor003aq1n04x5 _30189_ (.a(_02611_),
    .b(_02515_),
    .c(_02604_),
    .o1(_04444_));
 b15aoi013ah1n08x5 _30190_ (.a(_04444_),
    .b(_03370_),
    .c(_03391_),
    .d(_02573_),
    .o1(_04445_));
 b15aoai13ar1n02x5 _30191_ (.a(_03335_),
    .b(_04187_),
    .c(_02548_),
    .d(net835),
    .o1(_04446_));
 b15and003al1n04x5 _30192_ (.a(net840),
    .b(_02602_),
    .c(_03300_),
    .o(_04447_));
 b15norp02ar1n02x5 _30193_ (.a(_02545_),
    .b(_02724_),
    .o1(_04448_));
 b15nor004al1n02x5 _30194_ (.a(net832),
    .b(_02680_),
    .c(_02595_),
    .d(_02541_),
    .o1(_04449_));
 b15oai022ar1n04x5 _30195_ (.a(_04447_),
    .b(_04448_),
    .c(_04449_),
    .d(_02748_),
    .o1(_04450_));
 b15oai012ar1n02x5 _30196_ (.a(_02649_),
    .b(_03573_),
    .c(_03628_),
    .o1(_04451_));
 b15nand04as1n03x5 _30197_ (.a(_04445_),
    .b(_04446_),
    .c(_04450_),
    .d(_04451_),
    .o1(_04452_));
 b15aoai13ar1n02x5 _30198_ (.a(_02668_),
    .b(_04187_),
    .c(_02598_),
    .d(net842),
    .o1(_04454_));
 b15norp02ar1n02x5 _30199_ (.a(net841),
    .b(_02604_),
    .o1(_04455_));
 b15aoai13ah1n04x5 _30200_ (.a(_04455_),
    .b(_03384_),
    .c(_02635_),
    .d(net838),
    .o1(_04456_));
 b15norp02ar1n02x5 _30201_ (.a(_02548_),
    .b(_03311_),
    .o1(_04457_));
 b15oai112ah1n02x5 _30202_ (.a(_04454_),
    .b(_04456_),
    .c(_03349_),
    .d(_04457_),
    .o1(_04458_));
 b15nor004aq1n06x5 _30203_ (.a(_04436_),
    .b(_04443_),
    .c(_04452_),
    .d(_04458_),
    .o1(_04459_));
 b15orn003ar1n04x5 _30204_ (.a(\us01.a[7] ),
    .b(net825),
    .c(net834),
    .o(_04460_));
 b15oai022as1n06x5 _30205_ (.a(_02547_),
    .b(_03379_),
    .c(_04460_),
    .d(_02634_),
    .o1(_04461_));
 b15nand02ar1n02x5 _30206_ (.a(_02517_),
    .b(_04461_),
    .o1(_04462_));
 b15oab012ar1n02x5 _30207_ (.a(_03592_),
    .b(_03605_),
    .c(_02545_),
    .out0(_04463_));
 b15norp02ah1n02x5 _30208_ (.a(_02569_),
    .b(_02665_),
    .o1(_04465_));
 b15aoi022ah1n08x5 _30209_ (.a(_02562_),
    .b(_02757_),
    .c(_04465_),
    .d(_02759_),
    .o1(_04466_));
 b15nand04aq1n03x5 _30210_ (.a(net832),
    .b(_04462_),
    .c(_04463_),
    .d(_04466_),
    .o1(_04467_));
 b15norp03ar1n02x5 _30211_ (.a(net842),
    .b(_02546_),
    .c(_02547_),
    .o1(_04468_));
 b15oai122ah1n02x5 _30212_ (.a(_02515_),
    .b(_02557_),
    .c(_02623_),
    .d(_02643_),
    .e(_02680_),
    .o1(_04469_));
 b15aoai13an1n02x5 _30213_ (.a(net838),
    .b(_04468_),
    .c(_04469_),
    .d(_02569_),
    .o1(_04470_));
 b15oai022ar1n02x5 _30214_ (.a(net835),
    .b(_02515_),
    .c(_02583_),
    .d(_02602_),
    .o1(_04471_));
 b15aoi112ar1n02x5 _30215_ (.a(_02611_),
    .b(_04471_),
    .c(_02548_),
    .d(_02573_),
    .o1(_04472_));
 b15oai013al1n02x5 _30216_ (.a(_02569_),
    .b(_02637_),
    .c(_03370_),
    .d(_03373_),
    .o1(_04473_));
 b15aoi012ar1n02x5 _30217_ (.a(net842),
    .b(net835),
    .c(_02548_),
    .o1(_04474_));
 b15aoai13as1n02x5 _30218_ (.a(_04470_),
    .b(_04472_),
    .c(_04473_),
    .d(_04474_),
    .o1(_04476_));
 b15oai012an1n06x5 _30219_ (.a(_04467_),
    .b(_04476_),
    .c(net832),
    .o1(_04477_));
 b15nand04as1n16x5 _30220_ (.a(_04427_),
    .b(_04432_),
    .c(_04459_),
    .d(_04477_),
    .o1(_04478_));
 b15xor002aq1n06x5 _30221_ (.a(net398),
    .b(_04478_),
    .out0(_04479_));
 b15norp02as1n03x5 _30222_ (.a(_03020_),
    .b(_02997_),
    .o1(_04480_));
 b15oai012ah1n04x5 _30223_ (.a(_04221_),
    .b(_03028_),
    .c(_04243_),
    .o1(_04481_));
 b15aoai13al1n08x5 _30224_ (.a(net851),
    .b(_04480_),
    .c(_04481_),
    .d(net858),
    .o1(_04482_));
 b15nandp3ar1n02x5 _30225_ (.a(_02951_),
    .b(net851),
    .c(_03024_),
    .o1(_04483_));
 b15oaoi13ar1n03x5 _30226_ (.a(net853),
    .b(_04483_),
    .c(_02984_),
    .d(_02951_),
    .o1(_04484_));
 b15oaoi13aq1n02x5 _30227_ (.a(net851),
    .b(_02964_),
    .c(_02929_),
    .d(_02935_),
    .o1(_04485_));
 b15oai012an1n06x5 _30228_ (.a(_02820_),
    .b(_04484_),
    .c(_04485_),
    .o1(_04487_));
 b15aoi012as1n02x5 _30229_ (.a(_03020_),
    .b(_02876_),
    .c(_03463_),
    .o1(_04488_));
 b15oaoi13al1n03x5 _30230_ (.a(_02876_),
    .b(_02995_),
    .c(_02923_),
    .d(_02854_),
    .o1(_04489_));
 b15nor003ah1n06x5 _30231_ (.a(\us30.a[3] ),
    .b(_04488_),
    .c(_04489_),
    .o1(_04490_));
 b15aoi022al1n02x5 _30232_ (.a(_04302_),
    .b(_02900_),
    .c(_03021_),
    .d(_02881_),
    .o1(_04491_));
 b15nandp3ar1n02x5 _30233_ (.a(net861),
    .b(net854),
    .c(_02908_),
    .o1(_04492_));
 b15aoi012ah1n02x5 _30234_ (.a(net857),
    .b(_03427_),
    .c(_04492_),
    .o1(_04493_));
 b15nand02ah1n02x5 _30235_ (.a(net857),
    .b(_02908_),
    .o1(_04494_));
 b15aoi012aq1n02x5 _30236_ (.a(net861),
    .b(_03427_),
    .c(_04494_),
    .o1(_04495_));
 b15nano23ah1n06x5 _30237_ (.a(net850),
    .b(_04491_),
    .c(_04493_),
    .d(_04495_),
    .out0(_04496_));
 b15oai112aq1n16x5 _30238_ (.a(_04482_),
    .b(_04487_),
    .c(_04490_),
    .d(_04496_),
    .o1(_04498_));
 b15oai022an1n02x5 _30239_ (.a(_04227_),
    .b(_02876_),
    .c(_02882_),
    .d(_03028_),
    .o1(_04499_));
 b15aoi112ah1n02x5 _30240_ (.a(net859),
    .b(_02965_),
    .c(_04499_),
    .d(net852),
    .o1(_04500_));
 b15nandp2ar1n02x5 _30241_ (.a(_02899_),
    .b(_04250_),
    .o1(_04501_));
 b15oai012ah1n03x5 _30242_ (.a(net856),
    .b(_02833_),
    .c(_02915_),
    .o1(_04502_));
 b15oai012an1n04x5 _30243_ (.a(_04501_),
    .b(_04502_),
    .c(_04266_),
    .o1(_04503_));
 b15oai022ar1n02x5 _30244_ (.a(_02854_),
    .b(_02984_),
    .c(_02921_),
    .d(_04227_),
    .o1(_04504_));
 b15aoi022ar1n04x5 _30245_ (.a(_04263_),
    .b(_04503_),
    .c(_04504_),
    .d(net852),
    .o1(_04505_));
 b15aoi012aq1n06x5 _30246_ (.a(_04500_),
    .b(_04505_),
    .c(net859),
    .o1(_04506_));
 b15oai013as1n02x5 _30247_ (.a(_02950_),
    .b(_02858_),
    .c(_02989_),
    .d(_02986_),
    .o1(_04507_));
 b15aoai13ar1n04x5 _30248_ (.a(net858),
    .b(_02788_),
    .c(net853),
    .d(\us30.a[3] ),
    .o1(_04509_));
 b15ztpn00an1n08x5 TAP_413 ();
 b15oai022al1n06x5 _30250_ (.a(_02954_),
    .b(_03460_),
    .c(_02989_),
    .d(_02997_),
    .o1(_04511_));
 b15aoi022ah1n06x5 _30251_ (.a(_04507_),
    .b(_04509_),
    .c(_04511_),
    .d(_02811_),
    .o1(_04512_));
 b15aoi012ar1n02x5 _30252_ (.a(net858),
    .b(_02942_),
    .c(_03519_),
    .o1(_04513_));
 b15oai022ar1n02x5 _30253_ (.a(_02986_),
    .b(_02838_),
    .c(_03448_),
    .d(\us30.a[3] ),
    .o1(_04514_));
 b15norp02al1n04x5 _30254_ (.a(_04513_),
    .b(_04514_),
    .o1(_04515_));
 b15oai112ar1n06x5 _30255_ (.a(\us30.a[3] ),
    .b(_03463_),
    .c(_02995_),
    .d(_02921_),
    .o1(_04516_));
 b15nand02aq1n02x5 _30256_ (.a(_02819_),
    .b(_02943_),
    .o1(_04517_));
 b15oai022al1n02x5 _30257_ (.a(_02854_),
    .b(_02913_),
    .c(_04517_),
    .d(_02825_),
    .o1(_04518_));
 b15oai112an1n06x5 _30258_ (.a(net860),
    .b(_04516_),
    .c(_04518_),
    .d(\us30.a[3] ),
    .o1(_04520_));
 b15nand04ah1n03x5 _30259_ (.a(net855),
    .b(_02833_),
    .c(_02923_),
    .d(_02920_),
    .o1(_04521_));
 b15xor002ah1n03x5 _30260_ (.a(_02854_),
    .b(_02877_),
    .out0(_04522_));
 b15oaoi13as1n08x5 _30261_ (.a(_02811_),
    .b(_04521_),
    .c(_04522_),
    .d(_02862_),
    .o1(_04523_));
 b15aoi112ar1n02x5 _30262_ (.a(net853),
    .b(_02871_),
    .c(_02929_),
    .d(_03521_),
    .o1(_04524_));
 b15oab012ar1n02x5 _30263_ (.a(_04263_),
    .b(_02867_),
    .c(\us30.a[7] ),
    .out0(_04525_));
 b15norp03ar1n03x5 _30264_ (.a(\us30.a[5] ),
    .b(_04517_),
    .c(_04525_),
    .o1(_04526_));
 b15nor003as1n02x5 _30265_ (.a(_04523_),
    .b(_04524_),
    .c(_04526_),
    .o1(_04527_));
 b15nand04ah1n08x5 _30266_ (.a(_04512_),
    .b(_04515_),
    .c(_04520_),
    .d(_04527_),
    .o1(_04528_));
 b15nand02as1n02x5 _30267_ (.a(_02933_),
    .b(_04265_),
    .o1(_04529_));
 b15nandp3an1n03x5 _30268_ (.a(net853),
    .b(_02920_),
    .c(_02915_),
    .o1(_04531_));
 b15aoi222aq1n08x5 _30269_ (.a(net860),
    .b(_04529_),
    .c(_04531_),
    .d(_02954_),
    .e(_04302_),
    .f(_02921_),
    .o1(_04532_));
 b15norp03ar1n02x5 _30270_ (.a(net859),
    .b(\us30.a[5] ),
    .c(net844),
    .o1(_04533_));
 b15aoi013ar1n02x5 _30271_ (.a(_04533_),
    .b(_02943_),
    .c(net844),
    .d(\us30.a[5] ),
    .o1(_04534_));
 b15nor002aq1n02x5 _30272_ (.a(_03011_),
    .b(_04534_),
    .o1(_04535_));
 b15orn002ar1n08x5 _30273_ (.a(_02854_),
    .b(_03029_),
    .o(_04536_));
 b15oaoi13an1n04x5 _30274_ (.a(_02820_),
    .b(_04536_),
    .c(_03424_),
    .d(net853),
    .o1(_04537_));
 b15oai013aq1n08x5 _30275_ (.a(\us30.a[3] ),
    .b(_04532_),
    .c(_04535_),
    .d(_04537_),
    .o1(_04538_));
 b15nandp2al1n16x5 _30276_ (.a(_02951_),
    .b(net851),
    .o1(_04539_));
 b15oai022aq1n06x5 _30277_ (.a(_02858_),
    .b(_02921_),
    .c(_04539_),
    .d(_02986_),
    .o1(_04540_));
 b15nandp2al1n08x5 _30278_ (.a(_02811_),
    .b(_02932_),
    .o1(_04542_));
 b15oai022aq1n06x5 _30279_ (.a(_02867_),
    .b(_02992_),
    .c(_04542_),
    .d(_02820_),
    .o1(_04543_));
 b15aoi112as1n08x5 _30280_ (.a(net853),
    .b(_04540_),
    .c(_04543_),
    .d(net858),
    .o1(_04544_));
 b15oai122ah1n02x5 _30281_ (.a(net855),
    .b(_02956_),
    .c(_02913_),
    .d(_03514_),
    .e(_02876_),
    .o1(_04545_));
 b15inv040as1n02x5 _30282_ (.a(_04545_),
    .o1(_04546_));
 b15oai112al1n06x5 _30283_ (.a(net858),
    .b(_02862_),
    .c(_03028_),
    .d(_02820_),
    .o1(_04547_));
 b15oai012an1n02x5 _30284_ (.a(net862),
    .b(_02854_),
    .c(_03024_),
    .o1(_04548_));
 b15nand04al1n06x5 _30285_ (.a(_02951_),
    .b(_02996_),
    .c(_03029_),
    .d(_04548_),
    .o1(_04549_));
 b15aoi012aq1n02x5 _30286_ (.a(net858),
    .b(_02862_),
    .c(_03028_),
    .o1(_04550_));
 b15oai112ah1n08x5 _30287_ (.a(_04547_),
    .b(_04549_),
    .c(_04550_),
    .d(_02919_),
    .o1(_04551_));
 b15oai122al1n16x5 _30288_ (.a(_04538_),
    .b(_04544_),
    .c(_04546_),
    .d(_04551_),
    .e(net851),
    .o1(_04553_));
 b15nor004as1n12x5 _30289_ (.a(_04498_),
    .b(_04506_),
    .c(_04528_),
    .d(_04553_),
    .o1(_04554_));
 b15xor002an1n08x5 _30290_ (.a(_03034_),
    .b(_04554_),
    .out0(_04555_));
 b15xor002al1n12x5 _30291_ (.a(_04479_),
    .b(_04555_),
    .out0(_04556_));
 b15norp02aq1n02x5 _30292_ (.a(_03281_),
    .b(_03957_),
    .o1(_04557_));
 b15aoi013ar1n06x5 _30293_ (.a(_04557_),
    .b(_03962_),
    .c(_03181_),
    .d(_03046_),
    .o1(_04558_));
 b15oaoi13ar1n02x5 _30294_ (.a(net583),
    .b(_04558_),
    .c(_03912_),
    .d(_03167_),
    .o1(_04559_));
 b15nor002ah1n06x5 _30295_ (.a(net579),
    .b(net568),
    .o1(_04560_));
 b15nand02an1n03x5 _30296_ (.a(_03097_),
    .b(net590),
    .o1(_04561_));
 b15nand04ah1n08x5 _30297_ (.a(net575),
    .b(net595),
    .c(_04560_),
    .d(_04561_),
    .o1(_04562_));
 b15nanb02ar1n02x5 _30298_ (.a(net571),
    .b(net579),
    .out0(_04564_));
 b15nanb02aq1n24x5 _30299_ (.a(net577),
    .b(net571),
    .out0(_04565_));
 b15aoi012ar1n02x5 _30300_ (.a(net575),
    .b(_04564_),
    .c(_04565_),
    .o1(_04566_));
 b15nor003ar1n03x5 _30301_ (.a(net571),
    .b(_03281_),
    .c(_03068_),
    .o1(_04567_));
 b15oai012aq1n04x5 _30302_ (.a(net568),
    .b(_04566_),
    .c(_04567_),
    .o1(_04568_));
 b15aoi012aq1n06x5 _30303_ (.a(_03827_),
    .b(_04562_),
    .c(_04568_),
    .o1(_04569_));
 b15nandp3ar1n02x5 _30304_ (.a(_03036_),
    .b(_03144_),
    .c(_03157_),
    .o1(_04570_));
 b15oaoi13an1n02x5 _30305_ (.a(net586),
    .b(_04570_),
    .c(_03212_),
    .d(_03247_),
    .o1(_04571_));
 b15oaoi13ar1n02x5 _30306_ (.a(_03798_),
    .b(_03288_),
    .c(_03796_),
    .d(net588),
    .o1(_04572_));
 b15nor004ar1n03x5 _30307_ (.a(_04559_),
    .b(_04569_),
    .c(_04571_),
    .d(_04572_),
    .o1(_04573_));
 b15nandp2al1n04x5 _30308_ (.a(net569),
    .b(net580),
    .o1(_04575_));
 b15xor002an1n02x5 _30309_ (.a(net572),
    .b(net587),
    .out0(_04576_));
 b15oai013an1n06x5 _30310_ (.a(net591),
    .b(_03079_),
    .c(_04575_),
    .d(_04576_),
    .o1(_04577_));
 b15oai013an1n08x5 _30311_ (.a(_03102_),
    .b(_03163_),
    .c(_03249_),
    .d(_03957_),
    .o1(_04578_));
 b15nor003ar1n08x5 _30312_ (.a(net587),
    .b(net581),
    .c(_03187_),
    .o1(_04579_));
 b15oai012as1n04x5 _30313_ (.a(_04577_),
    .b(_04578_),
    .c(_04579_),
    .o1(_04580_));
 b15nor004aq1n03x5 _30314_ (.a(net580),
    .b(_03053_),
    .c(_03068_),
    .d(_03107_),
    .o1(_04581_));
 b15nanb02ah1n12x5 _30315_ (.a(net580),
    .b(net584),
    .out0(_04582_));
 b15aoai13an1n06x5 _30316_ (.a(net591),
    .b(_04581_),
    .c(_04582_),
    .d(_03171_),
    .o1(_04583_));
 b15norp02ar1n02x5 _30317_ (.a(net593),
    .b(_03044_),
    .o1(_04584_));
 b15aoai13as1n02x5 _30318_ (.a(_03134_),
    .b(_04584_),
    .c(_03196_),
    .d(_03089_),
    .o1(_04586_));
 b15nandp2as1n12x5 _30319_ (.a(net590),
    .b(_03237_),
    .o1(_04587_));
 b15oai012ar1n02x5 _30320_ (.a(net593),
    .b(_03067_),
    .c(_03274_),
    .o1(_04588_));
 b15aob012an1n02x5 _30321_ (.a(_03132_),
    .b(_04587_),
    .c(_04588_),
    .out0(_04589_));
 b15nand04as1n06x5 _30322_ (.a(_04580_),
    .b(_04583_),
    .c(_04586_),
    .d(_04589_),
    .o1(_04590_));
 b15norp02an1n08x5 _30323_ (.a(_03068_),
    .b(_03071_),
    .o1(_04591_));
 b15aobi12aq1n08x5 _30324_ (.a(net585),
    .b(net589),
    .c(net593),
    .out0(_04592_));
 b15nand02al1n03x5 _30325_ (.a(_04591_),
    .b(_04592_),
    .o1(_04593_));
 b15aoai13as1n02x5 _30326_ (.a(_03150_),
    .b(_03984_),
    .c(_03102_),
    .d(_03255_),
    .o1(_04594_));
 b15nor002aq1n03x5 _30327_ (.a(net572),
    .b(_03050_),
    .o1(_04595_));
 b15qgbno2an1n10x5 _30328_ (.a(net569),
    .b(net587),
    .o1(_04597_));
 b15oai122al1n16x5 _30329_ (.a(_04595_),
    .b(_04578_),
    .c(_04579_),
    .d(_03067_),
    .e(_04597_),
    .o1(_04598_));
 b15aoi013al1n04x5 _30330_ (.a(net581),
    .b(_04593_),
    .c(_04594_),
    .d(_04598_),
    .o1(_04599_));
 b15nor002an1n04x5 _30331_ (.a(net585),
    .b(_03044_),
    .o1(_04600_));
 b15oaoi13aq1n02x5 _30332_ (.a(net581),
    .b(_03181_),
    .c(_04600_),
    .d(net593),
    .o1(_04601_));
 b15oaoi13an1n04x5 _30333_ (.a(_04601_),
    .b(_03276_),
    .c(_03044_),
    .d(net581),
    .o1(_04602_));
 b15nor003ah1n02x5 _30334_ (.a(net580),
    .b(_03086_),
    .c(_03087_),
    .o1(_04603_));
 b15aoi012ah1n02x5 _30335_ (.a(_03165_),
    .b(_03255_),
    .c(net591),
    .o1(_04604_));
 b15mdn022al1n06x5 _30336_ (.a(_04603_),
    .b(_03128_),
    .o1(_04605_),
    .sa(_04604_));
 b15norp03ar1n03x5 _30337_ (.a(_03067_),
    .b(_03086_),
    .c(_03050_),
    .o1(_04606_));
 b15nor003an1n03x5 _30338_ (.a(net585),
    .b(_03050_),
    .c(_03135_),
    .o1(_04608_));
 b15oai112as1n06x5 _30339_ (.a(net580),
    .b(_03129_),
    .c(_04606_),
    .d(_04608_),
    .o1(_04609_));
 b15aoai13an1n06x5 _30340_ (.a(_03102_),
    .b(_03835_),
    .c(_03140_),
    .d(_03089_),
    .o1(_04610_));
 b15norp03ar1n04x5 _30341_ (.a(_03068_),
    .b(_03071_),
    .c(_03249_),
    .o1(_04611_));
 b15aoai13ar1n08x5 _30342_ (.a(_03163_),
    .b(_04611_),
    .c(_03814_),
    .d(_03215_),
    .o1(_04612_));
 b15nand04al1n12x5 _30343_ (.a(_04605_),
    .b(_04609_),
    .c(_04610_),
    .d(_04612_),
    .o1(_04613_));
 b15nor004as1n08x5 _30344_ (.a(_04590_),
    .b(_04599_),
    .c(_04602_),
    .d(_04613_),
    .o1(_04614_));
 b15aoi013ah1n02x5 _30345_ (.a(net575),
    .b(net579),
    .c(net582),
    .d(_03143_),
    .o1(_04615_));
 b15nandp2aq1n02x5 _30346_ (.a(_04560_),
    .b(_03994_),
    .o1(_04616_));
 b15oai012ah1n06x5 _30347_ (.a(_04615_),
    .b(_04616_),
    .c(net582),
    .o1(_04617_));
 b15oai012as1n03x5 _30348_ (.a(net575),
    .b(_03036_),
    .c(_04565_),
    .o1(_04619_));
 b15nor004ar1n08x5 _30349_ (.a(net582),
    .b(_03162_),
    .c(_03231_),
    .d(_03821_),
    .o1(_04620_));
 b15oai112an1n12x5 _30350_ (.a(_03818_),
    .b(_04617_),
    .c(_04619_),
    .d(_04620_),
    .o1(_04621_));
 b15aoi013aq1n02x5 _30351_ (.a(_03189_),
    .b(_03285_),
    .c(_03036_),
    .d(_03186_),
    .o1(_04622_));
 b15oai012aq1n06x5 _30352_ (.a(_04621_),
    .b(_04622_),
    .c(net590),
    .o1(_04623_));
 b15oai022aq1n08x5 _30353_ (.a(_03050_),
    .b(_03053_),
    .c(_03175_),
    .d(_03100_),
    .o1(_04624_));
 b15oaoi13ar1n02x5 _30354_ (.a(net594),
    .b(net590),
    .c(net586),
    .d(_03157_),
    .o1(_04625_));
 b15norp02ar1n02x5 _30355_ (.a(_03067_),
    .b(_03240_),
    .o1(_04626_));
 b15aoi012ah1n04x5 _30356_ (.a(net586),
    .b(_03162_),
    .c(_03228_),
    .o1(_04627_));
 b15oai013as1n02x5 _30357_ (.a(_04625_),
    .b(_04626_),
    .c(_04627_),
    .d(net590),
    .o1(_04628_));
 b15aoi022ar1n04x5 _30358_ (.a(net586),
    .b(_03983_),
    .c(_03167_),
    .d(_03836_),
    .o1(_04630_));
 b15oai112al1n08x5 _30359_ (.a(_04624_),
    .b(_04628_),
    .c(_04630_),
    .d(_03102_),
    .o1(_04631_));
 b15aoi022ar1n02x5 _30360_ (.a(net587),
    .b(_03215_),
    .c(_03962_),
    .d(net585),
    .o1(_04632_));
 b15oab012al1n02x5 _30361_ (.a(_03036_),
    .b(_03207_),
    .c(_04632_),
    .out0(_04633_));
 b15oai013an1n02x5 _30362_ (.a(_03252_),
    .b(_03843_),
    .c(_03057_),
    .d(net579),
    .o1(_04634_));
 b15oai012ar1n03x5 _30363_ (.a(net586),
    .b(_03252_),
    .c(net590),
    .o1(_04635_));
 b15aoi012ar1n02x5 _30364_ (.a(_03285_),
    .b(_03203_),
    .c(_03251_),
    .o1(_04636_));
 b15aoi022al1n02x5 _30365_ (.a(_03247_),
    .b(_03836_),
    .c(_04636_),
    .d(net590),
    .o1(_04637_));
 b15oai112al1n06x5 _30366_ (.a(_04634_),
    .b(_04635_),
    .c(_03102_),
    .d(_04637_),
    .o1(_04638_));
 b15oai112as1n08x5 _30367_ (.a(_03228_),
    .b(_03231_),
    .c(net594),
    .d(_03818_),
    .o1(_04639_));
 b15oab012ar1n02x5 _30368_ (.a(net583),
    .b(_03984_),
    .c(_04639_),
    .out0(_04641_));
 b15aoi022aq1n02x5 _30369_ (.a(_04631_),
    .b(_04633_),
    .c(_04638_),
    .d(_04641_),
    .o1(_04642_));
 b15nano23al1n06x5 _30370_ (.a(_04573_),
    .b(_04614_),
    .c(_04623_),
    .d(_04642_),
    .out0(_04643_));
 b15xnr002ar1n02x5 _30371_ (.a(_04217_),
    .b(net397),
    .out0(_04644_));
 b15xor002ar1n02x5 _30372_ (.a(_03413_),
    .b(_04644_),
    .out0(_04645_));
 b15xor002al1n02x5 _30373_ (.a(_04556_),
    .b(_04645_),
    .out0(_04646_));
 b15cmbn22ar1n08x5 _30374_ (.clk1(\text_in_r[67] ),
    .clk2(_04646_),
    .clkout(_04647_),
    .s(net538));
 b15xor002ar1n16x5 _30375_ (.a(\u0.w[1][3] ),
    .b(_04647_),
    .out0(_00108_));
 b15inv040aq1n04x5 _30376_ (.a(\text_in_r[68] ),
    .o1(_04648_));
 b15nand02ar1n02x5 _30377_ (.a(net702),
    .b(_02376_),
    .o1(_04649_));
 b15nonb03ar1n02x5 _30378_ (.a(net691),
    .b(net714),
    .c(net699),
    .out0(_04651_));
 b15aoi013ah1n02x5 _30379_ (.a(_04651_),
    .b(_02325_),
    .c(_02276_),
    .d(net699),
    .o1(_04652_));
 b15oai013al1n04x5 _30380_ (.a(_04649_),
    .b(_04652_),
    .c(net696),
    .d(_02279_),
    .o1(_04653_));
 b15nand02al1n08x5 _30381_ (.a(net709),
    .b(_04653_),
    .o1(_04654_));
 b15nand04ar1n02x5 _30382_ (.a(_02381_),
    .b(_02293_),
    .c(_02437_),
    .d(_02433_),
    .o1(_04655_));
 b15oai012an1n04x5 _30383_ (.a(_04655_),
    .b(_04110_),
    .c(_02381_),
    .o1(_04656_));
 b15nanb02al1n12x5 _30384_ (.a(\us12.a[1] ),
    .b(\us12.a[2] ),
    .out0(_04657_));
 b15oaoi13as1n08x5 _30385_ (.a(net714),
    .b(_04115_),
    .c(_02471_),
    .d(_04657_),
    .o1(_04658_));
 b15oaoi13ar1n04x5 _30386_ (.a(_04359_),
    .b(_04018_),
    .c(_02444_),
    .d(_03666_),
    .o1(_04659_));
 b15nand02ah1n06x5 _30387_ (.a(_02242_),
    .b(_02343_),
    .o1(_04660_));
 b15ornc04al1n16x5 _30388_ (.a(net698),
    .b(\us12.a[4] ),
    .c(net693),
    .d(\us12.a[6] ),
    .o(_04662_));
 b15oaoi13aq1n08x5 _30389_ (.a(_04660_),
    .b(_03666_),
    .c(net714),
    .d(_04662_),
    .o1(_04663_));
 b15nor004aq1n06x5 _30390_ (.a(_04656_),
    .b(_04658_),
    .c(_04659_),
    .d(_04663_),
    .o1(_04664_));
 b15aoai13ar1n02x5 _30391_ (.a(net713),
    .b(_04336_),
    .c(_02415_),
    .d(net703),
    .o1(_04665_));
 b15oai012ar1n08x5 _30392_ (.a(net707),
    .b(_02337_),
    .c(_04378_),
    .o1(_04666_));
 b15aoi012al1n02x5 _30393_ (.a(_02466_),
    .b(_04665_),
    .c(_04666_),
    .o1(_04667_));
 b15aoai13al1n03x5 _30394_ (.a(net706),
    .b(net702),
    .c(_02293_),
    .d(_02437_),
    .o1(_04668_));
 b15oa0022ar1n03x5 _30395_ (.a(net696),
    .b(_02402_),
    .c(_04085_),
    .d(net699),
    .o(_04669_));
 b15oaoi13ah1n04x5 _30396_ (.a(_04668_),
    .b(net702),
    .c(_02259_),
    .d(_04669_),
    .o1(_04670_));
 b15oai012ar1n04x5 _30397_ (.a(net704),
    .b(net711),
    .c(net715),
    .o1(_04671_));
 b15nand04as1n06x5 _30398_ (.a(_02461_),
    .b(_02351_),
    .c(_02374_),
    .d(_04671_),
    .o1(_04673_));
 b15nand02aq1n16x5 _30399_ (.a(_02251_),
    .b(_02395_),
    .o1(_04674_));
 b15oai122as1n16x5 _30400_ (.a(_04673_),
    .b(_04674_),
    .c(_03666_),
    .d(_04037_),
    .e(_04066_),
    .o1(_04675_));
 b15nor004aq1n06x5 _30401_ (.a(_02435_),
    .b(_04667_),
    .c(_04670_),
    .d(_04675_),
    .o1(_04676_));
 b15and003ar1n02x5 _30402_ (.a(net700),
    .b(net695),
    .c(net704),
    .o(_04677_));
 b15nor004ar1n04x5 _30403_ (.a(net700),
    .b(net695),
    .c(net715),
    .d(net704),
    .o1(_04678_));
 b15oai112aq1n08x5 _30404_ (.a(_02350_),
    .b(_02491_),
    .c(_04677_),
    .d(_04678_),
    .o1(_04679_));
 b15aoai13ar1n04x5 _30405_ (.a(_04679_),
    .b(_04375_),
    .c(_02431_),
    .d(_04330_),
    .o1(_04680_));
 b15nor002an1n06x5 _30406_ (.a(_04081_),
    .b(_04680_),
    .o1(_04681_));
 b15nand04as1n16x5 _30407_ (.a(_04654_),
    .b(_04664_),
    .c(_04676_),
    .d(_04681_),
    .o1(_04682_));
 b15oai012as1n06x5 _30408_ (.a(_02390_),
    .b(_04024_),
    .c(\us12.a[0] ),
    .o1(_04684_));
 b15nandp2aq1n04x5 _30409_ (.a(\us12.a[1] ),
    .b(_02354_),
    .o1(_04685_));
 b15aoi222as1n12x5 _30410_ (.a(net708),
    .b(_04684_),
    .c(_04685_),
    .d(_02275_),
    .e(_03677_),
    .f(_02469_),
    .o1(_04686_));
 b15nand03aq1n03x5 _30411_ (.a(net710),
    .b(_02475_),
    .c(_03651_),
    .o1(_04687_));
 b15oai112ah1n06x5 _30412_ (.a(net702),
    .b(_04687_),
    .c(_03651_),
    .d(_02407_),
    .o1(_04688_));
 b15nor002an1n03x5 _30413_ (.a(_04686_),
    .b(_04688_),
    .o1(_04689_));
 b15nand03ar1n08x5 _30414_ (.a(net713),
    .b(_02425_),
    .c(_04336_),
    .o1(_04690_));
 b15oaoi13ah1n03x5 _30415_ (.a(_03699_),
    .b(_03667_),
    .c(_02390_),
    .d(net709),
    .o1(_04691_));
 b15nand03al1n02x5 _30416_ (.a(net694),
    .b(net709),
    .c(_03670_),
    .o1(_04692_));
 b15nanb03ah1n06x5 _30417_ (.a(net694),
    .b(net691),
    .c(net696),
    .out0(_04693_));
 b15oaoi13ar1n04x5 _30418_ (.a(net713),
    .b(_04692_),
    .c(_04693_),
    .d(_02427_),
    .o1(_04695_));
 b15oaoi13aq1n04x5 _30419_ (.a(_02355_),
    .b(_02499_),
    .c(net709),
    .d(_02290_),
    .o1(_04696_));
 b15nonb02al1n08x5 _30420_ (.a(net712),
    .b(net699),
    .out0(_04697_));
 b15nano22ar1n02x5 _30421_ (.a(net696),
    .b(net706),
    .c(net714),
    .out0(_04698_));
 b15oai112al1n06x5 _30422_ (.a(_02293_),
    .b(_04697_),
    .c(_04698_),
    .d(_02412_),
    .o1(_04699_));
 b15xor002ar1n06x5 _30423_ (.a(_02276_),
    .b(_02433_),
    .out0(_04700_));
 b15oai013an1n08x5 _30424_ (.a(_04699_),
    .b(_04700_),
    .c(_04031_),
    .d(_02310_),
    .o1(_04701_));
 b15nor004al1n08x5 _30425_ (.a(_04691_),
    .b(_04695_),
    .c(_04696_),
    .d(_04701_),
    .o1(_04702_));
 b15aoi013as1n08x5 _30426_ (.a(_04689_),
    .b(_04690_),
    .c(_04702_),
    .d(_02381_),
    .o1(_04703_));
 b15aoai13ah1n03x5 _30427_ (.a(_02343_),
    .b(_04044_),
    .c(_04129_),
    .d(_04119_),
    .o1(_04704_));
 b15nandp3ar1n03x5 _30428_ (.a(\us12.a[4] ),
    .b(net693),
    .c(\us12.a[6] ),
    .o1(_04706_));
 b15nona23ar1n04x5 _30429_ (.a(_03752_),
    .b(_04706_),
    .c(_04382_),
    .d(net705),
    .out0(_04707_));
 b15aob012ar1n03x5 _30430_ (.a(net714),
    .b(_04704_),
    .c(_04707_),
    .out0(_04708_));
 b15nand02as1n02x5 _30431_ (.a(_02298_),
    .b(_02381_),
    .o1(_04709_));
 b15oai112aq1n08x5 _30432_ (.a(net710),
    .b(_04333_),
    .c(_04709_),
    .d(_02366_),
    .o1(_04710_));
 b15mdn022al1n02x5 _30433_ (.a(_03725_),
    .b(_03726_),
    .o1(_04711_),
    .sa(_03645_));
 b15nonb03ah1n08x5 _30434_ (.a(\us12.a[4] ),
    .b(net701),
    .c(net698),
    .out0(_04712_));
 b15aoi013ar1n02x5 _30435_ (.a(_04712_),
    .b(_02346_),
    .c(net701),
    .d(net693),
    .o1(_04713_));
 b15oai022ar1n02x5 _30436_ (.a(_04126_),
    .b(_04711_),
    .c(_04713_),
    .d(_04031_),
    .o1(_04714_));
 b15oai012ah1n02x5 _30437_ (.a(_04710_),
    .b(_04714_),
    .c(net712),
    .o1(_04715_));
 b15oai012ar1n02x5 _30438_ (.a(_02500_),
    .b(_03699_),
    .c(_02415_),
    .o1(_04717_));
 b15aoi022ar1n02x5 _30439_ (.a(_02412_),
    .b(_03699_),
    .c(_02500_),
    .d(_02411_),
    .o1(_04718_));
 b15oai112ah1n04x5 _30440_ (.a(net701),
    .b(_04717_),
    .c(_04718_),
    .d(_02242_),
    .o1(_04719_));
 b15nandp3aq1n08x5 _30441_ (.a(_04708_),
    .b(_04715_),
    .c(_04719_),
    .o1(_04720_));
 b15norp03as1n24x5 _30442_ (.a(_04682_),
    .b(_04703_),
    .c(_04720_),
    .o1(_04721_));
 b15norp03aq1n12x5 _30443_ (.a(_03036_),
    .b(_03053_),
    .c(_03068_),
    .o1(_04722_));
 b15norp03aq1n03x5 _30444_ (.a(_03068_),
    .b(_03071_),
    .c(_03878_),
    .o1(_04723_));
 b15aoi112aq1n06x5 _30445_ (.a(_04722_),
    .b(_04723_),
    .c(_03814_),
    .d(_03171_),
    .o1(_04724_));
 b15oai012an1n06x5 _30446_ (.a(net584),
    .b(_03887_),
    .c(_03796_),
    .o1(_04725_));
 b15nanb02an1n12x5 _30447_ (.a(net569),
    .b(net580),
    .out0(_04726_));
 b15oa0022an1n03x5 _30448_ (.a(_03843_),
    .b(_03193_),
    .c(_04726_),
    .d(net574),
    .o(_04728_));
 b15oa0012an1n06x5 _30449_ (.a(_03996_),
    .b(_03102_),
    .c(net568),
    .o(_04729_));
 b15oai222ah1n16x5 _30450_ (.a(_03272_),
    .b(_03201_),
    .c(_04565_),
    .d(_04728_),
    .e(_04729_),
    .f(_03925_),
    .o1(_04730_));
 b15obai22ar1n16x5 _30451_ (.a(_04724_),
    .b(_04725_),
    .c(_04730_),
    .d(net584),
    .out0(_04731_));
 b15oai022an1n02x5 _30452_ (.a(_03167_),
    .b(_03212_),
    .c(_03217_),
    .d(_03187_),
    .o1(_04732_));
 b15aoi013al1n02x5 _30453_ (.a(_03163_),
    .b(_03036_),
    .c(_03207_),
    .d(_03285_),
    .o1(_04733_));
 b15oai012ar1n06x5 _30454_ (.a(_04733_),
    .b(_03276_),
    .c(_03249_),
    .o1(_04734_));
 b15aoi022ar1n02x5 _30455_ (.a(net586),
    .b(_03270_),
    .c(_03285_),
    .d(_03237_),
    .o1(_04735_));
 b15nor002al1n02x5 _30456_ (.a(net594),
    .b(_04735_),
    .o1(_04736_));
 b15oai022al1n06x5 _30457_ (.a(net589),
    .b(_04732_),
    .c(_04734_),
    .d(_04736_),
    .o1(_04737_));
 b15aoi022ar1n02x5 _30458_ (.a(net586),
    .b(_03270_),
    .c(_03285_),
    .d(_03836_),
    .o1(_04739_));
 b15oai222al1n06x5 _30459_ (.a(_03983_),
    .b(_03890_),
    .c(_03217_),
    .d(_03247_),
    .e(net583),
    .f(_04739_),
    .o1(_04740_));
 b15nand02an1n03x5 _30460_ (.a(net594),
    .b(_04740_),
    .o1(_04741_));
 b15oai012as1n02x5 _30461_ (.a(\us23.a[1] ),
    .b(net582),
    .c(_03272_),
    .o1(_04742_));
 b15nand02an1n02x5 _30462_ (.a(net582),
    .b(_03261_),
    .o1(_04743_));
 b15nand03aq1n08x5 _30463_ (.a(net575),
    .b(net573),
    .c(\us23.a[2] ),
    .o1(_04744_));
 b15nand02ah1n02x5 _30464_ (.a(net579),
    .b(_03974_),
    .o1(_04745_));
 b15oai012ar1n08x5 _30465_ (.a(_04743_),
    .b(_04744_),
    .c(_04745_),
    .o1(_04746_));
 b15oai112aq1n12x5 _30466_ (.a(_03102_),
    .b(_04742_),
    .c(_04746_),
    .d(net590),
    .o1(_04747_));
 b15nand04ah1n08x5 _30467_ (.a(_04731_),
    .b(_04737_),
    .c(_04741_),
    .d(_04747_),
    .o1(_04748_));
 b15norp02ar1n02x5 _30468_ (.a(_03223_),
    .b(_03036_),
    .o1(_04750_));
 b15aoai13as1n02x5 _30469_ (.a(_04750_),
    .b(_04008_),
    .c(_03100_),
    .d(_03162_),
    .o1(_04751_));
 b15norp02al1n02x5 _30470_ (.a(net588),
    .b(_03044_),
    .o1(_04752_));
 b15aoi112al1n03x5 _30471_ (.a(_03798_),
    .b(_04752_),
    .c(net588),
    .d(_03137_),
    .o1(_04753_));
 b15oai022an1n02x5 _30472_ (.a(_03807_),
    .b(_03281_),
    .c(_03137_),
    .d(net588),
    .o1(_04754_));
 b15aoi112aq1n04x5 _30473_ (.a(_04751_),
    .b(_04753_),
    .c(_03067_),
    .d(_04754_),
    .o1(_04755_));
 b15oai112an1n02x5 _30474_ (.a(_03274_),
    .b(_03831_),
    .c(net577),
    .d(_03102_),
    .o1(_04756_));
 b15nanb02as1n06x5 _30475_ (.a(net568),
    .b(net576),
    .out0(_04757_));
 b15orn003ah1n04x5 _30476_ (.a(net571),
    .b(_03281_),
    .c(_04757_),
    .o(_04758_));
 b15oaoi13al1n03x5 _30477_ (.a(_03067_),
    .b(_04756_),
    .c(_04758_),
    .d(_03223_),
    .o1(_04759_));
 b15nandp2aq1n02x5 _30478_ (.a(_03036_),
    .b(_03240_),
    .o1(_04761_));
 b15oai012an1n04x5 _30479_ (.a(_04761_),
    .b(_03890_),
    .c(_03252_),
    .o1(_04762_));
 b15nandp2as1n08x5 _30480_ (.a(_03159_),
    .b(_04762_),
    .o1(_04763_));
 b15nand02ar1n02x5 _30481_ (.a(net584),
    .b(_03106_),
    .o1(_04764_));
 b15aoi022ar1n02x5 _30482_ (.a(_03960_),
    .b(_03849_),
    .c(_03865_),
    .d(net574),
    .o1(_04765_));
 b15nor002al1n03x5 _30483_ (.a(_04764_),
    .b(_04765_),
    .o1(_04766_));
 b15nandp2as1n04x5 _30484_ (.a(net584),
    .b(_03281_),
    .o1(_04767_));
 b15norp02ah1n02x5 _30485_ (.a(net588),
    .b(_03196_),
    .o1(_04768_));
 b15oai222as1n08x5 _30486_ (.a(_03121_),
    .b(_04767_),
    .c(_04768_),
    .d(_03272_),
    .e(_04758_),
    .f(net577),
    .o1(_04769_));
 b15aoi112an1n06x5 _30487_ (.a(_03289_),
    .b(_04766_),
    .c(_04769_),
    .d(net583),
    .o1(_04770_));
 b15nona23as1n16x5 _30488_ (.a(_04755_),
    .b(_04759_),
    .c(_04763_),
    .d(_04770_),
    .out0(_04772_));
 b15nand03al1n08x5 _30489_ (.a(_03067_),
    .b(_03162_),
    .c(_03228_),
    .o1(_04773_));
 b15aoi022ar1n16x5 _30490_ (.a(_03088_),
    .b(_03255_),
    .c(_04600_),
    .d(net589),
    .o1(_04774_));
 b15oai022ar1n06x5 _30491_ (.a(_03123_),
    .b(_04773_),
    .c(_04774_),
    .d(_03102_),
    .o1(_04775_));
 b15aob012al1n06x5 _30492_ (.a(_03815_),
    .b(_04775_),
    .c(_03036_),
    .out0(_04776_));
 b15oai112ar1n04x5 _30493_ (.a(net569),
    .b(_03233_),
    .c(_03046_),
    .d(_03097_),
    .o1(_04777_));
 b15oai122aq1n04x5 _30494_ (.a(_04777_),
    .b(_03923_),
    .c(_03983_),
    .d(_03067_),
    .e(_03167_),
    .o1(_04778_));
 b15aoi012ar1n02x5 _30495_ (.a(net594),
    .b(\us23.a[2] ),
    .c(_03157_),
    .o1(_04779_));
 b15aoi012ah1n02x5 _30496_ (.a(_04779_),
    .b(_03187_),
    .c(_03067_),
    .o1(_04780_));
 b15oai112al1n08x5 _30497_ (.a(net582),
    .b(_04778_),
    .c(_04780_),
    .d(net590),
    .o1(_04781_));
 b15nand02an1n06x5 _30498_ (.a(_04560_),
    .b(_03865_),
    .o1(_04783_));
 b15nand02as1n04x5 _30499_ (.a(net574),
    .b(_03836_),
    .o1(_04784_));
 b15oai012ah1n02x5 _30500_ (.a(net584),
    .b(net590),
    .c(_03100_),
    .o1(_04785_));
 b15aoi112an1n04x5 _30501_ (.a(net595),
    .b(_04783_),
    .c(_04784_),
    .d(_04785_),
    .o1(_04786_));
 b15nand04an1n03x5 _30502_ (.a(net590),
    .b(_03036_),
    .c(_03251_),
    .d(_03203_),
    .o1(_04787_));
 b15aoi022an1n02x5 _30503_ (.a(net584),
    .b(_03233_),
    .c(_03228_),
    .d(_03836_),
    .o1(_04788_));
 b15nand02al1n03x5 _30504_ (.a(net582),
    .b(_03203_),
    .o1(_04789_));
 b15oai122al1n08x5 _30505_ (.a(_04787_),
    .b(_04788_),
    .c(_04789_),
    .d(_04783_),
    .e(_03283_),
    .o1(_04790_));
 b15aoi012as1n06x5 _30506_ (.a(_04786_),
    .b(_04790_),
    .c(net595),
    .o1(_04791_));
 b15nanb02al1n16x5 _30507_ (.a(net576),
    .b(net569),
    .out0(_04792_));
 b15orn003al1n02x5 _30508_ (.a(net571),
    .b(_03046_),
    .c(_04792_),
    .o(_04794_));
 b15oaoi13an1n08x5 _30509_ (.a(net591),
    .b(_04794_),
    .c(_04757_),
    .d(_03829_),
    .o1(_04795_));
 b15nand03aq1n02x5 _30510_ (.a(net576),
    .b(_03097_),
    .c(net585),
    .o1(_04796_));
 b15oai012al1n06x5 _30511_ (.a(_04796_),
    .b(_03074_),
    .c(net576),
    .o1(_04797_));
 b15aoai13as1n08x5 _30512_ (.a(net578),
    .b(_04795_),
    .c(_04797_),
    .d(_04597_),
    .o1(_04798_));
 b15oai112aq1n16x5 _30513_ (.a(_04781_),
    .b(_04791_),
    .c(net582),
    .d(_04798_),
    .o1(_04799_));
 b15nor004as1n12x5 _30514_ (.a(_04748_),
    .b(_04772_),
    .c(_04776_),
    .d(_04799_),
    .o1(_04800_));
 b15xor002aq1n06x5 _30515_ (.a(_04721_),
    .b(_04800_),
    .out0(_04801_));
 b15xor002ah1n03x5 _30516_ (.a(_03413_),
    .b(_04478_),
    .out0(_04802_));
 b15xor002aq1n06x5 _30517_ (.a(_04801_),
    .b(_04802_),
    .out0(_04803_));
 b15nand02ar1n02x5 _30518_ (.a(net844),
    .b(_03431_),
    .o1(_04805_));
 b15oai012aq1n03x5 _30519_ (.a(_04805_),
    .b(_04268_),
    .c(\us30.a[0] ),
    .o1(_04806_));
 b15aoi013as1n04x5 _30520_ (.a(net852),
    .b(_02843_),
    .c(_04227_),
    .d(_04806_),
    .o1(_04807_));
 b15nand03as1n12x5 _30521_ (.a(net862),
    .b(_02854_),
    .c(_03452_),
    .o1(_04808_));
 b15nand02al1n02x5 _30522_ (.a(_02820_),
    .b(_02899_),
    .o1(_04809_));
 b15aoai13as1n03x5 _30523_ (.a(_04808_),
    .b(_02880_),
    .c(_04809_),
    .d(_04502_),
    .o1(_04810_));
 b15aob012as1n06x5 _30524_ (.a(_02794_),
    .b(_02781_),
    .c(net856),
    .out0(_04811_));
 b15aoi022an1n12x5 _30525_ (.a(\us30.a[1] ),
    .b(_04810_),
    .c(_04811_),
    .d(_02915_),
    .o1(_04812_));
 b15aoi012al1n16x5 _30526_ (.a(_04807_),
    .b(_04812_),
    .c(net852),
    .o1(_04813_));
 b15aoai13ar1n03x5 _30527_ (.a(net857),
    .b(_03460_),
    .c(_02873_),
    .d(net861),
    .o1(_04814_));
 b15oaoi13an1n04x5 _30528_ (.a(_02913_),
    .b(_04814_),
    .c(_02957_),
    .d(_02940_),
    .o1(_04816_));
 b15aoai13an1n04x5 _30529_ (.a(_02904_),
    .b(_02779_),
    .c(_04227_),
    .d(_02899_),
    .o1(_04817_));
 b15oai012ah1n04x5 _30530_ (.a(_02811_),
    .b(_02882_),
    .c(_02951_),
    .o1(_04818_));
 b15aoai13aq1n04x5 _30531_ (.a(_02919_),
    .b(net860),
    .c(_02904_),
    .d(_02779_),
    .o1(_04819_));
 b15aoi112ar1n08x5 _30532_ (.a(_04817_),
    .b(_04818_),
    .c(_04819_),
    .d(_02951_),
    .o1(_04820_));
 b15nandp2ah1n02x5 _30533_ (.a(_04298_),
    .b(_03024_),
    .o1(_04821_));
 b15qgbxo2an1n05x5 _30534_ (.a(_02951_),
    .b(_03002_),
    .out0(_04822_));
 b15oaoi13as1n08x5 _30535_ (.a(_02811_),
    .b(_04821_),
    .c(_04822_),
    .d(_02950_),
    .o1(_04823_));
 b15aoai13an1n02x5 _30536_ (.a(_03469_),
    .b(_03452_),
    .c(_02899_),
    .d(_02781_),
    .o1(_04824_));
 b15oaoi13an1n04x5 _30537_ (.a(_02820_),
    .b(_04824_),
    .c(_02964_),
    .d(_02864_),
    .o1(_04825_));
 b15nor004as1n08x5 _30538_ (.a(_04816_),
    .b(_04820_),
    .c(_04823_),
    .d(_04825_),
    .o1(_04827_));
 b15nand02al1n12x5 _30539_ (.a(net854),
    .b(_02957_),
    .o1(_04828_));
 b15nand03aq1n03x5 _30540_ (.a(_02811_),
    .b(_03452_),
    .c(_02871_),
    .o1(_04829_));
 b15aoi012an1n06x5 _30541_ (.a(_04828_),
    .b(_04829_),
    .c(_03521_),
    .o1(_04830_));
 b15aoi012ah1n02x5 _30542_ (.a(_03452_),
    .b(_02833_),
    .c(_02920_),
    .o1(_04831_));
 b15aoi013ar1n04x5 _30543_ (.a(net855),
    .b(_02833_),
    .c(_02923_),
    .d(_02920_),
    .o1(_04832_));
 b15nor004an1n08x5 _30544_ (.a(_02811_),
    .b(_03002_),
    .c(_04831_),
    .d(_04832_),
    .o1(_04833_));
 b15nanb02al1n02x5 _30545_ (.a(net856),
    .b(net849),
    .out0(_04834_));
 b15xor002ar1n04x5 _30546_ (.a(net862),
    .b(_04834_),
    .out0(_04835_));
 b15nano23al1n08x5 _30547_ (.a(_04835_),
    .b(_02844_),
    .c(_02808_),
    .d(_02825_),
    .out0(_04836_));
 b15nonb03ar1n12x5 _30548_ (.a(net849),
    .b(net844),
    .c(net847),
    .out0(_04838_));
 b15aoi012ar1n08x5 _30549_ (.a(net852),
    .b(net856),
    .c(\us30.a[1] ),
    .o1(_04839_));
 b15aoi022al1n24x5 _30550_ (.a(_02947_),
    .b(_02974_),
    .c(_04838_),
    .d(_04839_),
    .o1(_04840_));
 b15oaoi13ar1n08x5 _30551_ (.a(_04840_),
    .b(_02882_),
    .c(net861),
    .d(_02929_),
    .o1(_04841_));
 b15nor004ah1n12x5 _30552_ (.a(_04830_),
    .b(_04833_),
    .c(_04836_),
    .d(_04841_),
    .o1(_04842_));
 b15nand03an1n04x5 _30553_ (.a(_02904_),
    .b(_02899_),
    .c(_03460_),
    .o1(_04843_));
 b15oaoi13ar1n04x5 _30554_ (.a(_02811_),
    .b(_04843_),
    .c(_02997_),
    .d(_03460_),
    .o1(_04844_));
 b15oab012ar1n03x5 _30555_ (.a(_04539_),
    .b(_03467_),
    .c(_03018_),
    .out0(_04845_));
 b15oaoi13aq1n03x5 _30556_ (.a(_02820_),
    .b(_04221_),
    .c(_02935_),
    .d(_02921_),
    .o1(_04846_));
 b15aoi112an1n06x5 _30557_ (.a(_04844_),
    .b(_04845_),
    .c(_02811_),
    .d(_04846_),
    .o1(_04847_));
 b15nano23ar1n02x5 _30558_ (.a(net854),
    .b(net846),
    .c(net843),
    .d(net845),
    .out0(_04849_));
 b15nanb02ar1n02x5 _30559_ (.a(net857),
    .b(net848),
    .out0(_04850_));
 b15aoi022ar1n02x5 _30560_ (.a(_02951_),
    .b(_03024_),
    .c(_04849_),
    .d(_04850_),
    .o1(_04851_));
 b15norp02ah1n04x5 _30561_ (.a(_02820_),
    .b(_04851_),
    .o1(_04852_));
 b15aoai13ah1n06x5 _30562_ (.a(_02811_),
    .b(_04852_),
    .c(_03024_),
    .d(_02943_),
    .o1(_04853_));
 b15nand04ah1n16x5 _30563_ (.a(_04827_),
    .b(_04842_),
    .c(_04847_),
    .d(_04853_),
    .o1(_04854_));
 b15oaoi13ar1n02x5 _30564_ (.a(_02871_),
    .b(_02921_),
    .c(_02929_),
    .d(net853),
    .o1(_04855_));
 b15oai122an1n04x5 _30565_ (.a(net851),
    .b(_04243_),
    .c(_02984_),
    .d(_02957_),
    .e(_02929_),
    .o1(_04856_));
 b15aoi013ar1n02x5 _30566_ (.a(_02951_),
    .b(net860),
    .c(\us30.a[7] ),
    .d(_02899_),
    .o1(_04857_));
 b15aoi012aq1n02x5 _30567_ (.a(_04857_),
    .b(_02964_),
    .c(_02820_),
    .o1(_04858_));
 b15aoi013ar1n02x5 _30568_ (.a(net853),
    .b(_02837_),
    .c(_02984_),
    .d(_03029_),
    .o1(_04860_));
 b15aoi112as1n02x5 _30569_ (.a(_04855_),
    .b(_04856_),
    .c(_04858_),
    .d(_04860_),
    .o1(_04861_));
 b15aoai13ar1n02x5 _30570_ (.a(_02811_),
    .b(_02957_),
    .c(_04536_),
    .d(_02950_),
    .o1(_04862_));
 b15oai022ar1n02x5 _30571_ (.a(net853),
    .b(_02950_),
    .c(_04536_),
    .d(_02951_),
    .o1(_04863_));
 b15aoi012ar1n02x5 _30572_ (.a(_04862_),
    .b(_04863_),
    .c(net860),
    .o1(_04864_));
 b15nor002aq1n04x5 _30573_ (.a(_04861_),
    .b(_04864_),
    .o1(_04865_));
 b15oaoi13an1n02x5 _30574_ (.a(_02838_),
    .b(_02834_),
    .c(net853),
    .d(_03424_),
    .o1(_04866_));
 b15nor002ah1n02x5 _30575_ (.a(net853),
    .b(_03424_),
    .o1(_04867_));
 b15aoi013an1n03x5 _30576_ (.a(_04866_),
    .b(_04867_),
    .c(_02877_),
    .d(\us30.a[3] ),
    .o1(_04868_));
 b15nand03an1n06x5 _30577_ (.a(_02833_),
    .b(_02920_),
    .c(_03524_),
    .o1(_04869_));
 b15orn003al1n08x5 _30578_ (.a(net845),
    .b(_03500_),
    .c(_03011_),
    .o(_04871_));
 b15aoi013an1n08x5 _30579_ (.a(_02951_),
    .b(_04869_),
    .c(_04840_),
    .d(_04871_),
    .o1(_04872_));
 b15oai022ar1n02x5 _30580_ (.a(_02954_),
    .b(_02858_),
    .c(_02876_),
    .d(_04243_),
    .o1(_04873_));
 b15aoi012aq1n02x5 _30581_ (.a(_04872_),
    .b(_04873_),
    .c(_02951_),
    .o1(_04874_));
 b15nand02ar1n02x5 _30582_ (.a(_02837_),
    .b(_03463_),
    .o1(_04875_));
 b15aoai13as1n03x5 _30583_ (.a(_04875_),
    .b(_03535_),
    .c(_02932_),
    .d(net860),
    .o1(_04876_));
 b15oai112al1n12x5 _30584_ (.a(_04868_),
    .b(_04874_),
    .c(_04876_),
    .d(\us30.a[3] ),
    .o1(_04877_));
 b15nor004as1n12x5 _30585_ (.a(_04813_),
    .b(_04854_),
    .c(_04865_),
    .d(_04877_),
    .o1(_04878_));
 b15nandp3al1n03x5 _30586_ (.a(net824),
    .b(_02620_),
    .c(_02668_),
    .o1(_04879_));
 b15nanb02an1n03x5 _30587_ (.a(_03328_),
    .b(_03325_),
    .out0(_04880_));
 b15aoi112ah1n04x5 _30588_ (.a(\us01.a[5] ),
    .b(_02611_),
    .c(_04879_),
    .d(_04880_),
    .o1(_04882_));
 b15oai012ar1n02x5 _30589_ (.a(_02738_),
    .b(_02670_),
    .c(net833),
    .o1(_04883_));
 b15nand04as1n03x5 _30590_ (.a(net828),
    .b(_03563_),
    .c(net830),
    .d(_04883_),
    .o1(_04884_));
 b15aoi012ar1n02x5 _30591_ (.a(_02573_),
    .b(_02668_),
    .c(_02752_),
    .o1(_04885_));
 b15nand02an1n02x5 _30592_ (.a(_04884_),
    .b(_04885_),
    .o1(_04886_));
 b15oai022ar1n16x5 _30593_ (.a(net832),
    .b(_03583_),
    .c(_03395_),
    .d(_02585_),
    .o1(_04887_));
 b15oai022as1n06x5 _30594_ (.a(_04882_),
    .b(_04886_),
    .c(_04887_),
    .d(net836),
    .o1(_04888_));
 b15nor003aq1n06x5 _30595_ (.a(net836),
    .b(_02557_),
    .c(_02547_),
    .o1(_04889_));
 b15oaoi13ar1n02x5 _30596_ (.a(net830),
    .b(_02692_),
    .c(_02547_),
    .d(_02546_),
    .o1(_04890_));
 b15oai012ar1n02x5 _30597_ (.a(net841),
    .b(_04889_),
    .c(_04890_),
    .o1(_04891_));
 b15oaoi13al1n02x5 _30598_ (.a(_04889_),
    .b(net836),
    .c(_02548_),
    .d(_02748_),
    .o1(_04893_));
 b15oaoi13as1n03x5 _30599_ (.a(net834),
    .b(_04891_),
    .c(_04893_),
    .d(net830),
    .o1(_04894_));
 b15oai012as1n02x5 _30600_ (.a(net831),
    .b(_02680_),
    .c(_02595_),
    .o1(_04895_));
 b15aoi112aq1n06x5 _30601_ (.a(_02593_),
    .b(_02742_),
    .c(_02701_),
    .d(_02611_),
    .o1(_04896_));
 b15oai112ah1n08x5 _30602_ (.a(_04199_),
    .b(_04895_),
    .c(_04896_),
    .d(net831),
    .o1(_04897_));
 b15aoi022ah1n06x5 _30603_ (.a(_02649_),
    .b(_03340_),
    .c(_03376_),
    .d(_04188_),
    .o1(_04898_));
 b15aoi022as1n06x5 _30604_ (.a(_03602_),
    .b(_03397_),
    .c(_03335_),
    .d(_02759_),
    .o1(_04899_));
 b15oai122as1n16x5 _30605_ (.a(_04897_),
    .b(_04898_),
    .c(\us01.a[3] ),
    .d(_04899_),
    .e(_02569_),
    .o1(_04900_));
 b15aoi122al1n04x5 _30606_ (.a(net841),
    .b(_03391_),
    .c(_03341_),
    .d(_03309_),
    .e(_02748_),
    .o1(_04901_));
 b15nand03an1n08x5 _30607_ (.a(_02664_),
    .b(_02666_),
    .c(_02727_),
    .o1(_04902_));
 b15nandp3aq1n03x5 _30608_ (.a(net836),
    .b(_02759_),
    .c(_02668_),
    .o1(_04904_));
 b15aoi013al1n06x5 _30609_ (.a(_04901_),
    .b(_04902_),
    .c(_04904_),
    .d(net841),
    .o1(_04905_));
 b15oai012an1n03x5 _30610_ (.a(_02579_),
    .b(_02532_),
    .c(net833),
    .o1(_04906_));
 b15aoi012ah1n04x5 _30611_ (.a(_04906_),
    .b(_02678_),
    .c(_02658_),
    .o1(_04907_));
 b15aoi112ar1n02x5 _30612_ (.a(_02546_),
    .b(_02547_),
    .c(_03366_),
    .d(_02676_),
    .o1(_04908_));
 b15oai022ar1n02x5 _30613_ (.a(_02557_),
    .b(_02547_),
    .c(_02596_),
    .d(_02643_),
    .o1(_04909_));
 b15aoai13ah1n02x5 _30614_ (.a(net830),
    .b(_04908_),
    .c(_04909_),
    .d(net836),
    .o1(_04910_));
 b15nona23ar1n05x5 _30615_ (.a(_04905_),
    .b(_04907_),
    .c(_04910_),
    .d(_04445_),
    .out0(_04911_));
 b15norp03as1n02x5 _30616_ (.a(_02631_),
    .b(_02583_),
    .c(_03366_),
    .o1(_04912_));
 b15aoai13an1n06x5 _30617_ (.a(net841),
    .b(_04912_),
    .c(_02757_),
    .d(_03391_),
    .o1(_04913_));
 b15oai012an1n02x5 _30618_ (.a(_02573_),
    .b(_02654_),
    .c(_02743_),
    .o1(_04915_));
 b15oai022ar1n04x5 _30619_ (.a(_02596_),
    .b(_03317_),
    .c(_03576_),
    .d(_02680_),
    .o1(_04916_));
 b15aoi013an1n04x5 _30620_ (.a(_04915_),
    .b(_04916_),
    .c(net841),
    .d(net829),
    .o1(_04917_));
 b15nor004an1n03x5 _30621_ (.a(net841),
    .b(net830),
    .c(_02557_),
    .d(_02547_),
    .o1(_04918_));
 b15oai022ar1n04x5 _30622_ (.a(_02507_),
    .b(_02743_),
    .c(_03395_),
    .d(_02604_),
    .o1(_04919_));
 b15nor004ar1n04x5 _30623_ (.a(_02631_),
    .b(_02595_),
    .c(_02596_),
    .d(_02645_),
    .o1(_04920_));
 b15nor004aq1n06x5 _30624_ (.a(_02573_),
    .b(_04918_),
    .c(_04919_),
    .d(_04920_),
    .o1(_04921_));
 b15nandp3ar1n02x5 _30625_ (.a(net824),
    .b(net836),
    .c(net830),
    .o1(_04922_));
 b15oai022al1n02x5 _30626_ (.a(_02546_),
    .b(_03569_),
    .c(_04922_),
    .d(_02557_),
    .o1(_04923_));
 b15nandp2al1n05x5 _30627_ (.a(_04162_),
    .b(_04923_),
    .o1(_04924_));
 b15oai122an1n16x5 _30628_ (.a(_04913_),
    .b(_04917_),
    .c(_04921_),
    .d(net841),
    .e(_04924_),
    .o1(_04926_));
 b15nor004al1n08x5 _30629_ (.a(_04894_),
    .b(_04900_),
    .c(_04911_),
    .d(_04926_),
    .o1(_04927_));
 b15nor003al1n04x5 _30630_ (.a(net829),
    .b(\us01.a[7] ),
    .c(_02648_),
    .o1(_04928_));
 b15oai022as1n02x5 _30631_ (.a(net830),
    .b(_02623_),
    .c(_02671_),
    .d(_04162_),
    .o1(_04929_));
 b15aoai13as1n06x5 _30632_ (.a(\us01.a[5] ),
    .b(_04928_),
    .c(_04929_),
    .d(net829),
    .o1(_04930_));
 b15oaoi13aq1n03x5 _30633_ (.a(_03549_),
    .b(_04930_),
    .c(net830),
    .d(_02728_),
    .o1(_04931_));
 b15xor002ar1n02x5 _30634_ (.a(\us01.a[5] ),
    .b(net833),
    .out0(_04932_));
 b15nanb02al1n06x5 _30635_ (.a(net824),
    .b(net836),
    .out0(_04933_));
 b15nano23aq1n03x5 _30636_ (.a(_02611_),
    .b(_04932_),
    .c(_04933_),
    .d(_03328_),
    .out0(_04934_));
 b15oaoi13ar1n02x5 _30637_ (.a(_04934_),
    .b(_03409_),
    .c(_02665_),
    .d(net834),
    .o1(_04935_));
 b15oaoi13aq1n03x5 _30638_ (.a(net830),
    .b(_04935_),
    .c(_02700_),
    .d(_03379_),
    .o1(_04937_));
 b15norp02ar1n02x5 _30639_ (.a(net834),
    .b(_02532_),
    .o1(_04938_));
 b15oai022al1n02x5 _30640_ (.a(_02701_),
    .b(_02723_),
    .c(_04938_),
    .d(_03598_),
    .o1(_04939_));
 b15oai012ar1n02x5 _30641_ (.a(_02573_),
    .b(net834),
    .c(_02723_),
    .o1(_04940_));
 b15aoi012aq1n02x5 _30642_ (.a(_04939_),
    .b(_04940_),
    .c(_02611_),
    .o1(_04941_));
 b15aoi112an1n06x5 _30643_ (.a(_04931_),
    .b(_04937_),
    .c(_04941_),
    .d(net830),
    .o1(_04942_));
 b15aoai13al1n04x5 _30644_ (.a(net830),
    .b(_03373_),
    .c(_03592_),
    .d(net836),
    .o1(_04943_));
 b15oai112ar1n08x5 _30645_ (.a(_02569_),
    .b(_04943_),
    .c(_03395_),
    .d(_02610_),
    .o1(_04944_));
 b15oai012ar1n02x5 _30646_ (.a(_03325_),
    .b(net842),
    .c(\us01.a[5] ),
    .o1(_04945_));
 b15oai013ar1n02x5 _30647_ (.a(_04945_),
    .b(_03322_),
    .c(net842),
    .d(\us01.a[5] ),
    .o1(_04946_));
 b15aob012al1n06x5 _30648_ (.a(net833),
    .b(_02620_),
    .c(_04946_),
    .out0(_04948_));
 b15aoi012ar1n02x5 _30649_ (.a(_02631_),
    .b(_02635_),
    .c(_02573_),
    .o1(_04949_));
 b15aoi012ar1n02x5 _30650_ (.a(net830),
    .b(_02665_),
    .c(_02748_),
    .o1(_04950_));
 b15aob012ar1n02x5 _30651_ (.a(_03382_),
    .b(_03402_),
    .c(net828),
    .out0(_04951_));
 b15nand04al1n02x5 _30652_ (.a(\us01.a[5] ),
    .b(net822),
    .c(net842),
    .d(_04951_),
    .o1(_04952_));
 b15aoi012aq1n02x5 _30653_ (.a(_04949_),
    .b(_04950_),
    .c(_04952_),
    .o1(_04953_));
 b15oai012ah1n06x5 _30654_ (.a(_04944_),
    .b(_04948_),
    .c(_04953_),
    .o1(_04954_));
 b15nand04as1n16x5 _30655_ (.a(_04888_),
    .b(_04927_),
    .c(_04942_),
    .d(_04954_),
    .o1(_04955_));
 b15xor002al1n08x5 _30656_ (.a(_04878_),
    .b(_04955_),
    .out0(_04956_));
 b15xor002ah1n02x5 _30657_ (.a(_03034_),
    .b(_04956_),
    .out0(_04957_));
 b15xor002ah1n03x5 _30658_ (.a(_04803_),
    .b(_04957_),
    .out0(_04959_));
 b15mdn022al1n03x5 _30659_ (.a(_04648_),
    .b(_04959_),
    .o1(_04960_),
    .sa(net542));
 b15xor002ar1n03x5 _30660_ (.a(\u0.w[1][4] ),
    .b(_04960_),
    .out0(_00109_));
 b15nand02ar1n02x5 _30661_ (.a(net574),
    .b(_03162_),
    .o1(_04961_));
 b15oaoi13an1n03x5 _30662_ (.a(_03129_),
    .b(_04961_),
    .c(net574),
    .d(_03135_),
    .o1(_04962_));
 b15oai022aq1n06x5 _30663_ (.a(_03123_),
    .b(_03799_),
    .c(_03994_),
    .d(_03164_),
    .o1(_04963_));
 b15aoai13an1n08x5 _30664_ (.a(net577),
    .b(_04962_),
    .c(_04963_),
    .d(net568),
    .o1(_04964_));
 b15norp03as1n04x5 _30665_ (.a(net568),
    .b(net571),
    .c(net588),
    .o1(_04965_));
 b15nor002aq1n03x5 _30666_ (.a(net577),
    .b(_03071_),
    .o1(_04966_));
 b15oai112al1n16x5 _30667_ (.a(_03100_),
    .b(_03102_),
    .c(_04965_),
    .d(_04966_),
    .o1(_04967_));
 b15aoi012an1n16x5 _30668_ (.a(_03249_),
    .b(_04964_),
    .c(_04967_),
    .o1(_04969_));
 b15nandp3aq1n02x5 _30669_ (.a(_03251_),
    .b(_03143_),
    .c(_03853_),
    .o1(_04970_));
 b15aoi022aq1n08x5 _30670_ (.a(_03853_),
    .b(_03864_),
    .c(_03920_),
    .d(_03775_),
    .o1(_04971_));
 b15oaoi13ar1n08x5 _30671_ (.a(_03102_),
    .b(_04970_),
    .c(_04971_),
    .d(\us23.a[7] ),
    .o1(_04972_));
 b15aoai13ar1n06x5 _30672_ (.a(net588),
    .b(_04972_),
    .c(_03775_),
    .d(_03137_),
    .o1(_04973_));
 b15oa0022al1n03x5 _30673_ (.a(_03175_),
    .b(_03193_),
    .c(_04726_),
    .d(net577),
    .o(_04974_));
 b15oai122ah1n02x5 _30674_ (.a(net594),
    .b(_03252_),
    .c(_04587_),
    .d(_04744_),
    .e(_04974_),
    .o1(_04975_));
 b15nor003as1n04x5 _30675_ (.a(_03053_),
    .b(_03068_),
    .c(_04582_),
    .o1(_04976_));
 b15oai022an1n12x5 _30676_ (.a(_03843_),
    .b(_03827_),
    .c(_03820_),
    .d(_03217_),
    .o1(_04977_));
 b15norp02ar1n08x5 _30677_ (.a(net578),
    .b(_03097_),
    .o1(_04978_));
 b15aoi013ah1n06x5 _30678_ (.a(_04976_),
    .b(_04977_),
    .c(net587),
    .d(_04978_),
    .o1(_04980_));
 b15aob012al1n04x5 _30679_ (.a(_04975_),
    .b(_04980_),
    .c(_03102_),
    .out0(_04981_));
 b15oaoi13an1n03x5 _30680_ (.a(net594),
    .b(_04773_),
    .c(_03272_),
    .d(_03046_),
    .o1(_04982_));
 b15oai122ah1n08x5 _30681_ (.a(_03163_),
    .b(net586),
    .c(_03247_),
    .d(_03252_),
    .e(_03798_),
    .o1(_04983_));
 b15oai112al1n08x5 _30682_ (.a(net589),
    .b(_04773_),
    .c(_03252_),
    .d(_03075_),
    .o1(_04984_));
 b15aoai13as1n06x5 _30683_ (.a(_03036_),
    .b(_04982_),
    .c(_04983_),
    .d(_04984_),
    .o1(_04985_));
 b15norp03ar1n04x5 _30684_ (.a(_03102_),
    .b(_03983_),
    .c(_03193_),
    .o1(_04986_));
 b15oaoi13as1n02x5 _30685_ (.a(_03036_),
    .b(_03796_),
    .c(_03167_),
    .d(net594),
    .o1(_04987_));
 b15oai012al1n08x5 _30686_ (.a(net586),
    .b(_04986_),
    .c(_04987_),
    .o1(_04988_));
 b15nand04as1n12x5 _30687_ (.a(_04973_),
    .b(_04981_),
    .c(_04985_),
    .d(_04988_),
    .o1(_04989_));
 b15nandp3ar1n02x5 _30688_ (.a(net574),
    .b(_03123_),
    .c(_03261_),
    .o1(_04991_));
 b15aoi012ar1n02x5 _30689_ (.a(net572),
    .b(_03057_),
    .c(net577),
    .o1(_04992_));
 b15oaoi13ah1n03x5 _30690_ (.a(_03217_),
    .b(_04991_),
    .c(_04992_),
    .d(_04792_),
    .o1(_04993_));
 b15nor003ar1n08x5 _30691_ (.a(_03848_),
    .b(_03857_),
    .c(_04993_),
    .o1(_04994_));
 b15nand03ah1n02x5 _30692_ (.a(net568),
    .b(_03204_),
    .c(_03994_),
    .o1(_04995_));
 b15nandp2ar1n16x5 _30693_ (.a(_03196_),
    .b(_03270_),
    .o1(_04996_));
 b15aoi012al1n04x5 _30694_ (.a(_03193_),
    .b(_04995_),
    .c(_04996_),
    .o1(_04997_));
 b15aoai13aq1n03x5 _30695_ (.a(net582),
    .b(_03255_),
    .c(_03196_),
    .d(_03132_),
    .o1(_04998_));
 b15aoai13al1n04x5 _30696_ (.a(\us23.a[7] ),
    .b(_03864_),
    .c(_03920_),
    .d(net595),
    .o1(_04999_));
 b15nand02ah1n03x5 _30697_ (.a(net575),
    .b(_04560_),
    .o1(_05000_));
 b15aoi012ah1n02x5 _30698_ (.a(_03994_),
    .b(_03196_),
    .c(net573),
    .o1(_05002_));
 b15oaoi13aq1n04x5 _30699_ (.a(_04998_),
    .b(_04999_),
    .c(_05000_),
    .d(_05002_),
    .o1(_05003_));
 b15oai112as1n02x5 _30700_ (.a(net574),
    .b(_03162_),
    .c(_03186_),
    .d(_03223_),
    .o1(_05004_));
 b15aoi022aq1n02x5 _30701_ (.a(_03108_),
    .b(_03790_),
    .c(_03924_),
    .d(_03106_),
    .o1(_05005_));
 b15oai022as1n06x5 _30702_ (.a(_03887_),
    .b(_05004_),
    .c(_05005_),
    .d(_04784_),
    .o1(_05006_));
 b15nor004an1n12x5 _30703_ (.a(_03244_),
    .b(_04997_),
    .c(_05003_),
    .d(_05006_),
    .o1(_05007_));
 b15aoi013aq1n02x5 _30704_ (.a(_03855_),
    .b(_03253_),
    .c(_03143_),
    .d(_03036_),
    .o1(_05008_));
 b15nor003as1n03x5 _30705_ (.a(_03067_),
    .b(_03050_),
    .c(_05008_),
    .o1(_05009_));
 b15oaoi13ar1n02x5 _30706_ (.a(_03102_),
    .b(_03249_),
    .c(_03775_),
    .d(_03163_),
    .o1(_05010_));
 b15aoi012ar1n02x5 _30707_ (.a(_03036_),
    .b(_03283_),
    .c(_03912_),
    .o1(_05011_));
 b15oab012an1n03x5 _30708_ (.a(_03234_),
    .b(_05010_),
    .c(_05011_),
    .out0(_05013_));
 b15aob012aq1n04x5 _30709_ (.a(_03812_),
    .b(_03196_),
    .c(_03137_),
    .out0(_05014_));
 b15aoi112ar1n08x5 _30710_ (.a(_05009_),
    .b(_05013_),
    .c(_03274_),
    .d(_05014_),
    .o1(_05015_));
 b15nand04an1n03x5 _30711_ (.a(_03251_),
    .b(_03203_),
    .c(_03129_),
    .d(_03219_),
    .o1(_05016_));
 b15nand03ah1n06x5 _30712_ (.a(_03846_),
    .b(_03199_),
    .c(_03237_),
    .o1(_05017_));
 b15oai112aq1n06x5 _30713_ (.a(_05016_),
    .b(_05017_),
    .c(_03205_),
    .d(_03249_),
    .o1(_05018_));
 b15aoi122ah1n06x5 _30714_ (.a(net581),
    .b(_03240_),
    .c(_03159_),
    .d(_03270_),
    .e(_04592_),
    .o1(_05019_));
 b15oaoi13an1n08x5 _30715_ (.a(_05019_),
    .b(net583),
    .c(_03984_),
    .d(_04639_),
    .o1(_05020_));
 b15nandp3ar1n04x5 _30716_ (.a(net582),
    .b(_03186_),
    .c(_03261_),
    .o1(_05021_));
 b15xor002an1n04x5 _30717_ (.a(net575),
    .b(net590),
    .out0(_05022_));
 b15mdn022an1n04x5 _30718_ (.a(_03186_),
    .b(_03196_),
    .o1(_05024_),
    .sa(_03223_));
 b15orn003ar1n03x5 _30719_ (.a(net582),
    .b(_03843_),
    .c(_03829_),
    .o(_05025_));
 b15oai022ah1n08x5 _30720_ (.a(_05021_),
    .b(_05022_),
    .c(_05024_),
    .d(_05025_),
    .o1(_05026_));
 b15oaoi13aq1n03x5 _30721_ (.a(_03102_),
    .b(_03858_),
    .c(_03288_),
    .d(_03283_),
    .o1(_05027_));
 b15nor004ah1n06x5 _30722_ (.a(_05018_),
    .b(_05020_),
    .c(_05026_),
    .d(_05027_),
    .o1(_05028_));
 b15nand04ah1n16x5 _30723_ (.a(_04994_),
    .b(_05007_),
    .c(_05015_),
    .d(_05028_),
    .o1(_05029_));
 b15norp03as1n24x5 _30724_ (.a(_04969_),
    .b(_04989_),
    .c(_05029_),
    .o1(_05030_));
 b15xor002ah1n03x5 _30725_ (.a(net711),
    .b(_04067_),
    .out0(_05031_));
 b15nand03ah1n03x5 _30726_ (.a(_02276_),
    .b(_02343_),
    .c(_02333_),
    .o1(_05032_));
 b15aoi022an1n04x5 _30727_ (.a(net707),
    .b(_02376_),
    .c(_02462_),
    .d(_02350_),
    .o1(_05033_));
 b15oai022as1n08x5 _30728_ (.a(_05031_),
    .b(_05032_),
    .c(_05033_),
    .d(_04074_),
    .o1(_05035_));
 b15mdn022an1n06x5 _30729_ (.a(_02350_),
    .b(_02426_),
    .o1(_05036_),
    .sa(net699));
 b15nor004aq1n12x5 _30730_ (.a(_02381_),
    .b(_02273_),
    .c(_04060_),
    .d(_05036_),
    .o1(_05037_));
 b15nandp2al1n04x5 _30731_ (.a(_02251_),
    .b(_02433_),
    .o1(_05038_));
 b15nandp2aq1n04x5 _30732_ (.a(_04378_),
    .b(_03651_),
    .o1(_05039_));
 b15oai222as1n16x5 _30733_ (.a(_02290_),
    .b(_05038_),
    .c(_02463_),
    .d(_03739_),
    .e(_05039_),
    .f(_02438_),
    .o1(_05040_));
 b15nand04aq1n03x5 _30734_ (.a(_02343_),
    .b(_02291_),
    .c(_02293_),
    .d(_02395_),
    .o1(_05041_));
 b15oai013an1n08x5 _30735_ (.a(_05041_),
    .b(_02444_),
    .c(_02407_),
    .d(net702),
    .o1(_05042_));
 b15nor004as1n12x5 _30736_ (.a(_05035_),
    .b(_05037_),
    .c(_05040_),
    .d(_05042_),
    .o1(_05043_));
 b15nor003ar1n02x5 _30737_ (.a(_03657_),
    .b(_02385_),
    .c(_03753_),
    .o1(_05044_));
 b15norp02as1n03x5 _30738_ (.a(\us12.a[6] ),
    .b(net705),
    .o1(_05046_));
 b15nonb02aq1n03x5 _30739_ (.a(net698),
    .b(net706),
    .out0(_05047_));
 b15oai112as1n12x5 _30740_ (.a(_05046_),
    .b(_03726_),
    .c(_05047_),
    .d(_03752_),
    .o1(_05048_));
 b15oai022al1n02x5 _30741_ (.a(_02460_),
    .b(_02500_),
    .c(_05048_),
    .d(net714),
    .o1(_05049_));
 b15aoi012an1n04x5 _30742_ (.a(_05044_),
    .b(_05049_),
    .c(net709),
    .o1(_05050_));
 b15nanb02an1n02x5 _30743_ (.a(_04380_),
    .b(net709),
    .out0(_05051_));
 b15nand03aq1n24x5 _30744_ (.a(net704),
    .b(_02341_),
    .c(_02333_),
    .o1(_05052_));
 b15nandp2al1n02x5 _30745_ (.a(net714),
    .b(_02381_),
    .o1(_05053_));
 b15oai022al1n06x5 _30746_ (.a(net714),
    .b(_05052_),
    .c(_05053_),
    .d(_02500_),
    .o1(_05054_));
 b15oai112ah1n08x5 _30747_ (.a(_02242_),
    .b(_05051_),
    .c(_05054_),
    .d(net709),
    .o1(_05055_));
 b15oai112al1n04x5 _30748_ (.a(_04052_),
    .b(net705),
    .c(_02411_),
    .d(_04125_),
    .o1(_05057_));
 b15aoi013ar1n02x5 _30749_ (.a(_03745_),
    .b(_03679_),
    .c(_02298_),
    .d(\us12.a[6] ),
    .o1(_05058_));
 b15oai012as1n03x5 _30750_ (.a(_05057_),
    .b(_05058_),
    .c(_04052_),
    .o1(_05059_));
 b15nand04an1n12x5 _30751_ (.a(net698),
    .b(net693),
    .c(net712),
    .d(_05059_),
    .o1(_05060_));
 b15nand04ah1n16x5 _30752_ (.a(_05043_),
    .b(_05050_),
    .c(_05055_),
    .d(_05060_),
    .o1(_05061_));
 b15and002ar1n03x5 _30753_ (.a(net699),
    .b(net702),
    .o(_05062_));
 b15nona22ar1n02x5 _30754_ (.a(net696),
    .b(net691),
    .c(net694),
    .out0(_05063_));
 b15oai022ar1n02x5 _30755_ (.a(_02325_),
    .b(_04693_),
    .c(_05063_),
    .d(_02449_),
    .o1(_05064_));
 b15oai022ah1n02x5 _30756_ (.a(_02290_),
    .b(_03657_),
    .c(_03648_),
    .d(_02309_),
    .o1(_05065_));
 b15ao0022an1n03x5 _30757_ (.a(_05062_),
    .b(_05064_),
    .c(_05065_),
    .d(_04049_),
    .o(_05066_));
 b15aoi022ar1n16x5 _30758_ (.a(_02381_),
    .b(_04112_),
    .c(_05066_),
    .d(_02461_),
    .o1(_05068_));
 b15oai012ar1n02x5 _30759_ (.a(net701),
    .b(_02500_),
    .c(net712),
    .o1(_05069_));
 b15oai112al1n02x5 _30760_ (.a(_02381_),
    .b(_03677_),
    .c(_03699_),
    .d(_02325_),
    .o1(_05070_));
 b15nand03as1n04x5 _30761_ (.a(_02461_),
    .b(_05069_),
    .c(_05070_),
    .o1(_05071_));
 b15nand02an1n06x5 _30762_ (.a(\us12.a[6] ),
    .b(_02298_),
    .o1(_05072_));
 b15oa0022ar1n02x5 _30763_ (.a(_04660_),
    .b(_04127_),
    .c(_04128_),
    .d(net706),
    .o(_05073_));
 b15oa0022ar1n04x5 _30764_ (.a(_04660_),
    .b(_03724_),
    .c(_05073_),
    .d(net698),
    .o(_05074_));
 b15oai112as1n16x5 _30765_ (.a(_05068_),
    .b(_05071_),
    .c(_05072_),
    .d(_05074_),
    .o1(_05075_));
 b15nandp3aq1n02x5 _30766_ (.a(_02343_),
    .b(_02321_),
    .c(_02354_),
    .o1(_05076_));
 b15norp02an1n02x5 _30767_ (.a(_02242_),
    .b(_02412_),
    .o1(_05077_));
 b15oai122aq1n08x5 _30768_ (.a(_05076_),
    .b(_05077_),
    .c(_05048_),
    .d(_03673_),
    .e(_04674_),
    .o1(_05079_));
 b15nonb02an1n02x5 _30769_ (.a(net694),
    .b(net699),
    .out0(_05080_));
 b15aoi022al1n02x5 _30770_ (.a(_02412_),
    .b(_05080_),
    .c(_04033_),
    .d(net706),
    .o1(_05081_));
 b15oai012aq1n04x5 _30771_ (.a(_02353_),
    .b(_04035_),
    .c(_05081_),
    .o1(_05082_));
 b15aoi012ar1n08x5 _30772_ (.a(_05079_),
    .b(_05082_),
    .c(net702),
    .o1(_05083_));
 b15norp03as1n04x5 _30773_ (.a(_02466_),
    .b(_02357_),
    .c(_02390_),
    .o1(_05084_));
 b15aoi122as1n08x5 _30774_ (.a(_05084_),
    .b(_02351_),
    .c(_02326_),
    .d(_02319_),
    .e(_04051_),
    .o1(_05085_));
 b15oai022ar1n02x5 _30775_ (.a(net696),
    .b(net706),
    .c(_03651_),
    .d(_04085_),
    .o1(_05086_));
 b15nor004as1n03x5 _30776_ (.a(net699),
    .b(net691),
    .c(_03706_),
    .d(_05086_),
    .o1(_05087_));
 b15nonb02al1n04x5 _30777_ (.a(_05085_),
    .b(_05087_),
    .out0(_05088_));
 b15aoi012al1n02x5 _30778_ (.a(_02461_),
    .b(_02346_),
    .c(_02441_),
    .o1(_05090_));
 b15aoi022ar1n04x5 _30779_ (.a(_02365_),
    .b(_04032_),
    .c(_05062_),
    .d(_02341_),
    .o1(_05091_));
 b15oai013an1n06x5 _30780_ (.a(_05090_),
    .b(_05091_),
    .c(net710),
    .d(net696),
    .o1(_05092_));
 b15nand03an1n04x5 _30781_ (.a(_02242_),
    .b(_02381_),
    .c(_02425_),
    .o1(_05093_));
 b15oai012aq1n12x5 _30782_ (.a(_05093_),
    .b(_03642_),
    .c(_02242_),
    .o1(_05094_));
 b15oai112al1n16x5 _30783_ (.a(net714),
    .b(_05092_),
    .c(_05094_),
    .d(net706),
    .o1(_05095_));
 b15nand04as1n02x5 _30784_ (.a(net701),
    .b(_02411_),
    .c(_02430_),
    .d(_02291_),
    .o1(_05096_));
 b15oai112ar1n08x5 _30785_ (.a(_02343_),
    .b(_03725_),
    .c(_04103_),
    .d(_04119_),
    .o1(_05097_));
 b15aoi012aq1n06x5 _30786_ (.a(net710),
    .b(_05096_),
    .c(_05097_),
    .o1(_05098_));
 b15nor004as1n08x5 _30787_ (.a(_02452_),
    .b(_03654_),
    .c(_04675_),
    .d(_05098_),
    .o1(_05099_));
 b15nand04ah1n16x5 _30788_ (.a(_05083_),
    .b(_05088_),
    .c(_05095_),
    .d(_05099_),
    .o1(_05101_));
 b15norp03as1n24x5 _30789_ (.a(_05061_),
    .b(_05075_),
    .c(_05101_),
    .o1(_05102_));
 b15xnr002ah1n08x5 _30790_ (.a(_05030_),
    .b(_05102_),
    .out0(_05103_));
 b15xor002an1n12x5 _30791_ (.a(_04955_),
    .b(_05103_),
    .out0(_05104_));
 b15oai012ar1n02x5 _30792_ (.a(net854),
    .b(_02974_),
    .c(_03024_),
    .o1(_05105_));
 b15oaoi13al1n02x5 _30793_ (.a(_02811_),
    .b(_05105_),
    .c(_02964_),
    .d(_02820_),
    .o1(_05106_));
 b15oai013ar1n03x5 _30794_ (.a(_03519_),
    .b(_03524_),
    .c(net854),
    .d(_02992_),
    .o1(_05107_));
 b15nor003as1n03x5 _30795_ (.a(net857),
    .b(_05106_),
    .c(_05107_),
    .o1(_05108_));
 b15oai012ar1n04x5 _30796_ (.a(net856),
    .b(_03024_),
    .c(_04299_),
    .o1(_05109_));
 b15aoi012al1n02x5 _30797_ (.a(net861),
    .b(_03427_),
    .c(_05109_),
    .o1(_05110_));
 b15norp02aq1n02x5 _30798_ (.a(net848),
    .b(_02880_),
    .o1(_05112_));
 b15aoi112aq1n04x5 _30799_ (.a(_02956_),
    .b(_05110_),
    .c(_05112_),
    .d(_03000_),
    .o1(_05113_));
 b15aoi112aq1n03x5 _30800_ (.a(_02892_),
    .b(_03483_),
    .c(net861),
    .d(_03523_),
    .o1(_05114_));
 b15norp03an1n12x5 _30801_ (.a(_05108_),
    .b(_05113_),
    .c(_05114_),
    .o1(_05115_));
 b15aoi012ar1n02x5 _30802_ (.a(_02951_),
    .b(_04227_),
    .c(_02882_),
    .o1(_05116_));
 b15oai012an1n06x5 _30803_ (.a(_02908_),
    .b(_03021_),
    .c(_05116_),
    .o1(_05117_));
 b15oai022an1n08x5 _30804_ (.a(net853),
    .b(_02862_),
    .c(_02929_),
    .d(_02820_),
    .o1(_05118_));
 b15nandp2al1n08x5 _30805_ (.a(net853),
    .b(_03018_),
    .o1(_05119_));
 b15oai012al1n08x5 _30806_ (.a(_05119_),
    .b(_02921_),
    .c(net853),
    .o1(_05120_));
 b15oai022aq1n06x5 _30807_ (.a(net860),
    .b(_02984_),
    .c(_02929_),
    .d(net858),
    .o1(_05121_));
 b15aoi222as1n12x5 _30808_ (.a(net858),
    .b(_05118_),
    .c(_05120_),
    .d(_02820_),
    .e(_05121_),
    .f(net853),
    .o1(_05123_));
 b15aoi013al1n06x5 _30809_ (.a(net851),
    .b(_04808_),
    .c(_05117_),
    .d(_05123_),
    .o1(_05124_));
 b15oai012an1n02x5 _30810_ (.a(net851),
    .b(net853),
    .c(_02871_),
    .o1(_05125_));
 b15nandp2ar1n05x5 _30811_ (.a(_03452_),
    .b(_02919_),
    .o1(_05126_));
 b15oaoi13al1n04x5 _30812_ (.a(_05125_),
    .b(_02986_),
    .c(_02877_),
    .d(_05126_),
    .o1(_05127_));
 b15oai012ar1n08x5 _30813_ (.a(_03519_),
    .b(_02942_),
    .c(_02854_),
    .o1(_05128_));
 b15oai022al1n08x5 _30814_ (.a(_04302_),
    .b(_04542_),
    .c(_04536_),
    .d(net860),
    .o1(_05129_));
 b15aoi122ar1n08x5 _30815_ (.a(_05127_),
    .b(_05128_),
    .c(_02820_),
    .d(_05129_),
    .e(_02951_),
    .o1(_05130_));
 b15aoi012al1n06x5 _30816_ (.a(_02856_),
    .b(_04266_),
    .c(\us30.a[1] ),
    .o1(_05131_));
 b15oaoi13an1n04x5 _30817_ (.a(_02820_),
    .b(_02856_),
    .c(_02880_),
    .d(net848),
    .o1(_05132_));
 b15oai112ah1n16x5 _30818_ (.a(net847),
    .b(_02791_),
    .c(_05131_),
    .d(_05132_),
    .o1(_05133_));
 b15norp02ar1n02x5 _30819_ (.a(_02876_),
    .b(_02892_),
    .o1(_05134_));
 b15aoai13ah1n02x5 _30820_ (.a(net855),
    .b(_05134_),
    .c(_03470_),
    .d(_02844_),
    .o1(_05135_));
 b15nor003aq1n03x5 _30821_ (.a(net845),
    .b(_02892_),
    .c(_03011_),
    .o1(_05136_));
 b15norp02as1n03x5 _30822_ (.a(_02820_),
    .b(net847),
    .o1(_05137_));
 b15norp02ar1n02x5 _30823_ (.a(net855),
    .b(_02837_),
    .o1(_05138_));
 b15oai022ah1n02x5 _30824_ (.a(_03029_),
    .b(_05138_),
    .c(_03457_),
    .d(_02918_),
    .o1(_05139_));
 b15aoi122ar1n04x5 _30825_ (.a(_04823_),
    .b(_05136_),
    .c(_05137_),
    .d(_05139_),
    .e(net851),
    .o1(_05140_));
 b15nand04aq1n08x5 _30826_ (.a(_05130_),
    .b(_05133_),
    .c(_05135_),
    .d(_05140_),
    .o1(_05141_));
 b15nandp3ar1n02x5 _30827_ (.a(net860),
    .b(_02977_),
    .c(_02885_),
    .o1(_05142_));
 b15nand03aq1n12x5 _30828_ (.a(net850),
    .b(_02831_),
    .c(_02833_),
    .o1(_05144_));
 b15nandp3ar1n02x5 _30829_ (.a(_02811_),
    .b(_02904_),
    .c(_02899_),
    .o1(_05145_));
 b15aoai13an1n02x5 _30830_ (.a(_05142_),
    .b(net860),
    .c(_05144_),
    .d(_05145_),
    .o1(_05146_));
 b15aoi012ar1n02x5 _30831_ (.a(_02951_),
    .b(net860),
    .c(_03024_),
    .o1(_05147_));
 b15nand02al1n03x5 _30832_ (.a(_02820_),
    .b(_03024_),
    .o1(_05148_));
 b15aoi013ar1n02x5 _30833_ (.a(_05147_),
    .b(_05148_),
    .c(_02921_),
    .d(_02951_),
    .o1(_05149_));
 b15ao0022ah1n03x5 _30834_ (.a(_02951_),
    .b(_05146_),
    .c(_05149_),
    .d(_03469_),
    .o(_05150_));
 b15nand02ar1n02x5 _30835_ (.a(_02811_),
    .b(_02837_),
    .o1(_05151_));
 b15oai112aq1n02x5 _30836_ (.a(net855),
    .b(_05144_),
    .c(_05151_),
    .d(_02964_),
    .o1(_05152_));
 b15nona23ah1n02x5 _30837_ (.a(_02892_),
    .b(_03011_),
    .c(_03511_),
    .d(_04266_),
    .out0(_05153_));
 b15nand02ar1n02x5 _30838_ (.a(_02844_),
    .b(_03018_),
    .o1(_05155_));
 b15aoi013ar1n02x5 _30839_ (.a(net854),
    .b(_02904_),
    .c(_02779_),
    .d(net850),
    .o1(_05156_));
 b15nandp3al1n02x5 _30840_ (.a(_05153_),
    .b(_05155_),
    .c(_05156_),
    .o1(_05157_));
 b15norp03ar1n02x5 _30841_ (.a(net857),
    .b(net843),
    .c(net845),
    .o1(_05158_));
 b15oai112aq1n04x5 _30842_ (.a(net852),
    .b(net848),
    .c(_02920_),
    .d(_05158_),
    .o1(_05159_));
 b15aoi022an1n02x5 _30843_ (.a(net848),
    .b(_02781_),
    .c(_03010_),
    .d(net845),
    .o1(_05160_));
 b15oai012an1n08x5 _30844_ (.a(_05159_),
    .b(_05160_),
    .c(_02951_),
    .o1(_05161_));
 b15aoai13ar1n04x5 _30845_ (.a(_05152_),
    .b(_05157_),
    .c(_05161_),
    .d(_05137_),
    .o1(_05162_));
 b15nona23as1n04x5 _30846_ (.a(_03464_),
    .b(_05150_),
    .c(_05162_),
    .d(_04482_),
    .out0(_05163_));
 b15nor004as1n12x5 _30847_ (.a(_05115_),
    .b(_05124_),
    .c(_05141_),
    .d(_05163_),
    .o1(_05164_));
 b15oaoi13an1n02x5 _30848_ (.a(_02616_),
    .b(_02642_),
    .c(_03382_),
    .d(_02738_),
    .o1(_05166_));
 b15aoi012ar1n02x5 _30849_ (.a(_02742_),
    .b(_02701_),
    .c(net842),
    .o1(_05167_));
 b15oai022as1n02x5 _30850_ (.a(_03299_),
    .b(_03549_),
    .c(_05167_),
    .d(_02768_),
    .o1(_05168_));
 b15oaoi13ar1n02x5 _30851_ (.a(net834),
    .b(_02642_),
    .c(_02583_),
    .d(_02616_),
    .o1(_05169_));
 b15nor003as1n03x5 _30852_ (.a(_05166_),
    .b(_05168_),
    .c(_05169_),
    .o1(_05170_));
 b15nor002aq1n03x5 _30853_ (.a(net834),
    .b(_02623_),
    .o1(_05171_));
 b15oai012ah1n02x5 _30854_ (.a(_04460_),
    .b(_02684_),
    .c(_02547_),
    .o1(_05172_));
 b15aoi022ar1n08x5 _30855_ (.a(net841),
    .b(_05171_),
    .c(_05172_),
    .d(_02573_),
    .o1(_05173_));
 b15oaoi13al1n04x5 _30856_ (.a(net830),
    .b(_05170_),
    .c(_05173_),
    .d(_02546_),
    .o1(_05174_));
 b15nanb02ar1n02x5 _30857_ (.a(_04174_),
    .b(_04162_),
    .out0(_05175_));
 b15oaoi13al1n03x5 _30858_ (.a(net829),
    .b(_05175_),
    .c(_04933_),
    .d(_04162_),
    .o1(_05177_));
 b15norp03ar1n02x5 _30859_ (.a(_04162_),
    .b(_02541_),
    .c(_02671_),
    .o1(_05178_));
 b15norp02ar1n02x5 _30860_ (.a(_02623_),
    .b(_03387_),
    .o1(_05179_));
 b15oaoi13ah1n02x5 _30861_ (.a(_05177_),
    .b(net829),
    .c(_05178_),
    .d(_05179_),
    .o1(_05180_));
 b15nor002as1n04x5 _30862_ (.a(_03317_),
    .b(_05180_),
    .o1(_05181_));
 b15nor002aq1n02x5 _30863_ (.a(_02716_),
    .b(_02596_),
    .o1(_05182_));
 b15oai022al1n06x5 _30864_ (.a(_02634_),
    .b(_02643_),
    .c(_02649_),
    .d(_02595_),
    .o1(_05183_));
 b15norp03al1n02x5 _30865_ (.a(_02611_),
    .b(_03391_),
    .c(_03309_),
    .o1(_05184_));
 b15aoi013an1n03x5 _30866_ (.a(_05184_),
    .b(_02669_),
    .c(_02716_),
    .d(_02611_),
    .o1(_05185_));
 b15oai022an1n02x5 _30867_ (.a(_02695_),
    .b(_02700_),
    .c(_03362_),
    .d(_02604_),
    .o1(_05186_));
 b15aoi222as1n06x5 _30868_ (.a(_05182_),
    .b(_05183_),
    .c(_05185_),
    .d(_03373_),
    .e(net842),
    .f(_05186_),
    .o1(_05188_));
 b15aoi022ar1n02x5 _30869_ (.a(_02569_),
    .b(_03598_),
    .c(_03341_),
    .d(_02745_),
    .o1(_05189_));
 b15norp03aq1n02x5 _30870_ (.a(net830),
    .b(_02649_),
    .c(_05189_),
    .o1(_05190_));
 b15oai112ar1n02x5 _30871_ (.a(_02620_),
    .b(_03325_),
    .c(_02615_),
    .d(net833),
    .o1(_05191_));
 b15oaoi13an1n03x5 _30872_ (.a(_05191_),
    .b(net842),
    .c(_02573_),
    .d(_02692_),
    .o1(_05192_));
 b15oaoi13ar1n02x5 _30873_ (.a(_03562_),
    .b(_02743_),
    .c(_02593_),
    .d(_02573_),
    .o1(_05193_));
 b15nand02ar1n02x5 _30874_ (.a(_02579_),
    .b(_02634_),
    .o1(_05194_));
 b15nand03an1n03x5 _30875_ (.a(_02615_),
    .b(net822),
    .c(_02618_),
    .o1(_05195_));
 b15oaoi13ar1n03x5 _30876_ (.a(_05194_),
    .b(_05195_),
    .c(_03563_),
    .d(_02738_),
    .o1(_05196_));
 b15nor004ah1n03x5 _30877_ (.a(_05190_),
    .b(_05192_),
    .c(_05193_),
    .d(_05196_),
    .o1(_05197_));
 b15nandp3an1n03x5 _30878_ (.a(_02611_),
    .b(_03391_),
    .c(_03370_),
    .o1(_05199_));
 b15aoi012ah1n06x5 _30879_ (.a(net836),
    .b(_04440_),
    .c(_05199_),
    .o1(_05200_));
 b15aoi022al1n02x5 _30880_ (.a(_02724_),
    .b(_02635_),
    .c(_03341_),
    .d(_02709_),
    .o1(_05201_));
 b15nand04al1n06x5 _30881_ (.a(net826),
    .b(net825),
    .c(net836),
    .d(net833),
    .o1(_05202_));
 b15oa0022ar1n03x5 _30882_ (.a(_04184_),
    .b(_03319_),
    .c(_03355_),
    .d(net830),
    .o(_05203_));
 b15oai022as1n06x5 _30883_ (.a(net842),
    .b(_05201_),
    .c(_05202_),
    .d(_05203_),
    .o1(_05204_));
 b15nano23ah1n08x5 _30884_ (.a(_05188_),
    .b(_05197_),
    .c(_05200_),
    .d(_05204_),
    .out0(_05205_));
 b15nor002aq1n02x5 _30885_ (.a(_02643_),
    .b(_03322_),
    .o1(_05206_));
 b15norp02al1n04x5 _30886_ (.a(_02595_),
    .b(_04933_),
    .o1(_05207_));
 b15aoai13ar1n08x5 _30887_ (.a(net822),
    .b(_05206_),
    .c(_05207_),
    .d(net830),
    .o1(_05208_));
 b15oai022aq1n12x5 _30888_ (.a(_02557_),
    .b(_02547_),
    .c(_02643_),
    .d(_02680_),
    .o1(_05210_));
 b15aoai13as1n06x5 _30889_ (.a(net830),
    .b(_04889_),
    .c(_05210_),
    .d(net841),
    .o1(_05211_));
 b15norp02as1n04x5 _30890_ (.a(net831),
    .b(_02743_),
    .o1(_05212_));
 b15oai022as1n06x5 _30891_ (.a(_02609_),
    .b(_03319_),
    .c(_03355_),
    .d(_02610_),
    .o1(_05213_));
 b15oai012al1n06x5 _30892_ (.a(_02609_),
    .b(_02724_),
    .c(_02611_),
    .o1(_05214_));
 b15aoi222as1n12x5 _30893_ (.a(_02649_),
    .b(_05212_),
    .c(_05213_),
    .d(_02711_),
    .e(_05214_),
    .f(_02757_),
    .o1(_05215_));
 b15aoi013al1n08x5 _30894_ (.a(net833),
    .b(_05208_),
    .c(_05211_),
    .d(_05215_),
    .o1(_05216_));
 b15oai022ar1n02x5 _30895_ (.a(net825),
    .b(_02546_),
    .c(_02557_),
    .d(_02532_),
    .o1(_05217_));
 b15aoi022an1n04x5 _30896_ (.a(_02598_),
    .b(_03626_),
    .c(_02766_),
    .d(_05217_),
    .o1(_05218_));
 b15nor002ar1n08x5 _30897_ (.a(_02631_),
    .b(_05218_),
    .o1(_05219_));
 b15nandp2ah1n03x5 _30898_ (.a(_02668_),
    .b(_02748_),
    .o1(_05221_));
 b15oai013an1n02x5 _30899_ (.a(net842),
    .b(_02595_),
    .c(_02596_),
    .d(_02695_),
    .o1(_05222_));
 b15nor002ar1n02x5 _30900_ (.a(net838),
    .b(_02716_),
    .o1(_05223_));
 b15oaoi13al1n04x5 _30901_ (.a(_05222_),
    .b(_05223_),
    .c(_03341_),
    .d(_03370_),
    .o1(_05224_));
 b15qgbna2an1n05x5 _30902_ (.o1(_05225_),
    .a(_02662_),
    .b(_02666_));
 b15oa0022ar1n06x5 _30903_ (.a(_05225_),
    .b(_02654_),
    .c(_02700_),
    .d(_02554_),
    .o(_05226_));
 b15aoi022as1n08x5 _30904_ (.a(_05221_),
    .b(_05224_),
    .c(_05226_),
    .d(_02611_),
    .o1(_05227_));
 b15nor004as1n12x5 _30905_ (.a(_03566_),
    .b(_05216_),
    .c(_05219_),
    .d(_05227_),
    .o1(_05228_));
 b15nona23an1n32x5 _30906_ (.a(_05174_),
    .b(_05181_),
    .c(_05205_),
    .d(_05228_),
    .out0(_05229_));
 b15qgbxo2an1n10x5 _30907_ (.a(_05164_),
    .b(_05229_),
    .out0(_05230_));
 b15xor002ar1n12x5 _30908_ (.a(_05104_),
    .b(_05230_),
    .out0(_05232_));
 b15cmbn22ar1n02x5 _30909_ (.clk1(\text_in_r[69] ),
    .clk2(_05232_),
    .clkout(_05233_),
    .s(net542));
 b15xor002ar1n02x5 _30910_ (.a(\u0.w[1][5] ),
    .b(_05233_),
    .out0(_00110_));
 b15oai012al1n06x5 _30911_ (.a(_03286_),
    .b(_03217_),
    .c(_03272_),
    .o1(_05234_));
 b15nandp2al1n04x5 _30912_ (.a(_03129_),
    .b(_03286_),
    .o1(_05235_));
 b15nand04aq1n16x5 _30913_ (.a(_03168_),
    .b(_03923_),
    .c(_05234_),
    .d(_05235_),
    .o1(_05236_));
 b15norp03as1n04x5 _30914_ (.a(_03050_),
    .b(_03135_),
    .c(_03144_),
    .o1(_05237_));
 b15aoai13al1n03x5 _30915_ (.a(net581),
    .b(_05237_),
    .c(_03089_),
    .d(net587),
    .o1(_05238_));
 b15aoai13as1n02x5 _30916_ (.a(_03814_),
    .b(_03215_),
    .c(net587),
    .d(_03962_),
    .o1(_05239_));
 b15aoi012ar1n06x5 _30917_ (.a(_03067_),
    .b(_05238_),
    .c(_05239_),
    .o1(_05240_));
 b15nanb02ar1n02x5 _30918_ (.a(net579),
    .b(net568),
    .out0(_05242_));
 b15nor002an1n03x5 _30919_ (.a(_05242_),
    .b(_03829_),
    .o1(_05243_));
 b15nor002ar1n04x5 _30920_ (.a(_03053_),
    .b(_03893_),
    .o1(_05244_));
 b15aoai13as1n08x5 _30921_ (.a(net575),
    .b(_05243_),
    .c(_05244_),
    .d(_03196_),
    .o1(_05245_));
 b15aoai13an1n06x5 _30922_ (.a(net585),
    .b(_05237_),
    .c(_03149_),
    .d(net587),
    .o1(_05246_));
 b15nandp3al1n04x5 _30923_ (.a(net585),
    .b(_03210_),
    .c(_03157_),
    .o1(_05247_));
 b15aoi013al1n06x5 _30924_ (.a(net581),
    .b(_05245_),
    .c(_05246_),
    .d(_05247_),
    .o1(_05248_));
 b15aoi013al1n03x5 _30925_ (.a(_04722_),
    .b(_03088_),
    .c(_03036_),
    .d(net594),
    .o1(_05249_));
 b15norp02ar1n02x5 _30926_ (.a(net581),
    .b(_03798_),
    .o1(_05250_));
 b15aoi022al1n02x5 _30927_ (.a(_03149_),
    .b(_03853_),
    .c(_05250_),
    .d(_03088_),
    .o1(_05251_));
 b15oai022an1n06x5 _30928_ (.a(_03168_),
    .b(_05249_),
    .c(_05251_),
    .d(_03163_),
    .o1(_05253_));
 b15nor004as1n08x5 _30929_ (.a(_03971_),
    .b(_05240_),
    .c(_05248_),
    .d(_05253_),
    .o1(_05254_));
 b15aoi012ar1n02x5 _30930_ (.a(net594),
    .b(_03887_),
    .c(_03181_),
    .o1(_05255_));
 b15nandp3ar1n02x5 _30931_ (.a(net581),
    .b(_03144_),
    .c(_03199_),
    .o1(_05256_));
 b15aoi012aq1n02x5 _30932_ (.a(_05255_),
    .b(_05256_),
    .c(_04761_),
    .o1(_05257_));
 b15aoai13aq1n03x5 _30933_ (.a(net583),
    .b(_03270_),
    .c(_03228_),
    .d(_03162_),
    .o1(_05258_));
 b15norp02al1n04x5 _30934_ (.a(_03067_),
    .b(_03270_),
    .o1(_05259_));
 b15oaoi13as1n08x5 _30935_ (.a(_05258_),
    .b(\us23.a[1] ),
    .c(_04627_),
    .d(_05259_),
    .o1(_05260_));
 b15oai112ar1n04x5 _30936_ (.a(_03036_),
    .b(_03285_),
    .c(_03061_),
    .d(_03057_),
    .o1(_05261_));
 b15nandp3ar1n02x5 _30937_ (.a(_03807_),
    .b(_03057_),
    .c(_03237_),
    .o1(_05262_));
 b15oai112ar1n02x5 _30938_ (.a(net581),
    .b(_03123_),
    .c(_03132_),
    .d(net586),
    .o1(_05264_));
 b15aoi022ar1n02x5 _30939_ (.a(_03162_),
    .b(_03233_),
    .c(_03075_),
    .d(_03132_),
    .o1(_05265_));
 b15oai112ar1n02x5 _30940_ (.a(_05261_),
    .b(_05262_),
    .c(_05264_),
    .d(_05265_),
    .o1(_05266_));
 b15and002al1n08x5 _30941_ (.a(net578),
    .b(net572),
    .o(_05267_));
 b15nonb03ar1n02x5 _30942_ (.a(net576),
    .b(net570),
    .c(net581),
    .out0(_05268_));
 b15nano22ar1n02x5 _30943_ (.a(net570),
    .b(net581),
    .c(net576),
    .out0(_05269_));
 b15oai112as1n02x5 _30944_ (.a(_03165_),
    .b(_05267_),
    .c(_05268_),
    .d(_05269_),
    .o1(_05270_));
 b15nano23al1n02x5 _30945_ (.a(net576),
    .b(net589),
    .c(net581),
    .d(net570),
    .out0(_05271_));
 b15nano23aq1n03x5 _30946_ (.a(net570),
    .b(net581),
    .c(net589),
    .d(net576),
    .out0(_05272_));
 b15oai112as1n04x5 _30947_ (.a(_03207_),
    .b(_05267_),
    .c(_05271_),
    .d(_05272_),
    .o1(_05273_));
 b15aoi012ar1n06x5 _30948_ (.a(_03228_),
    .b(_03144_),
    .c(_03233_),
    .o1(_05275_));
 b15nandp3ar1n02x5 _30949_ (.a(_03162_),
    .b(_03123_),
    .c(_03237_),
    .o1(_05276_));
 b15oai112aq1n04x5 _30950_ (.a(_05270_),
    .b(_05273_),
    .c(_05275_),
    .d(_05276_),
    .o1(_05277_));
 b15nor004aq1n03x5 _30951_ (.a(_05257_),
    .b(_05260_),
    .c(_05266_),
    .d(_05277_),
    .o1(_05278_));
 b15nand02ar1n02x5 _30952_ (.a(net586),
    .b(_03807_),
    .o1(_05279_));
 b15oaoi13ar1n02x5 _30953_ (.a(_03102_),
    .b(_05279_),
    .c(_03252_),
    .d(_03181_),
    .o1(_05280_));
 b15norp02ar1n02x5 _30954_ (.a(net589),
    .b(_05279_),
    .o1(_05281_));
 b15oai012an1n04x5 _30955_ (.a(net581),
    .b(_05280_),
    .c(_05281_),
    .o1(_05282_));
 b15oaoi13as1n02x5 _30956_ (.a(_03181_),
    .b(_03276_),
    .c(_03102_),
    .d(_03187_),
    .o1(_05283_));
 b15oaoi13ar1n03x5 _30957_ (.a(_03102_),
    .b(_03276_),
    .c(_03187_),
    .d(_03046_),
    .o1(_05284_));
 b15nor003al1n06x5 _30958_ (.a(net581),
    .b(_05283_),
    .c(_05284_),
    .o1(_05286_));
 b15oaoi13ah1n03x5 _30959_ (.a(_03187_),
    .b(_03181_),
    .c(net593),
    .d(_03818_),
    .o1(_05287_));
 b15aoi112ah1n02x5 _30960_ (.a(_03050_),
    .b(_03242_),
    .c(_03135_),
    .d(_03086_),
    .o1(_05288_));
 b15nor003ah1n06x5 _30961_ (.a(_03036_),
    .b(_05287_),
    .c(_05288_),
    .o1(_05289_));
 b15aoai13al1n06x5 _30962_ (.a(_03163_),
    .b(_03073_),
    .c(_03157_),
    .d(_03165_),
    .o1(_05290_));
 b15aoai13an1n04x5 _30963_ (.a(net593),
    .b(_03170_),
    .c(_04591_),
    .d(net589),
    .o1(_05291_));
 b15aoi013al1n06x5 _30964_ (.a(_05286_),
    .b(_05289_),
    .c(_05290_),
    .d(_05291_),
    .o1(_05292_));
 b15oai022an1n02x5 _30965_ (.a(_03079_),
    .b(_03053_),
    .c(_03846_),
    .d(net584),
    .o1(_05293_));
 b15aoi112an1n02x5 _30966_ (.a(_03079_),
    .b(_03053_),
    .c(_03836_),
    .d(net591),
    .o1(_05294_));
 b15oai112as1n06x5 _30967_ (.a(_03036_),
    .b(_05293_),
    .c(_05294_),
    .d(_03132_),
    .o1(_05295_));
 b15aoi022aq1n04x5 _30968_ (.a(_03163_),
    .b(_03132_),
    .c(_03150_),
    .d(_03102_),
    .o1(_05297_));
 b15oai112an1n12x5 _30969_ (.a(_03919_),
    .b(_05295_),
    .c(_05297_),
    .d(_04582_),
    .o1(_05298_));
 b15nano23ah1n06x5 _30970_ (.a(_05278_),
    .b(_05282_),
    .c(_05292_),
    .d(_05298_),
    .out0(_05299_));
 b15nandp3as1n24x5 _30971_ (.a(_05236_),
    .b(_05254_),
    .c(_05299_),
    .o1(_05300_));
 b15oai012ar1n02x5 _30972_ (.a(_02742_),
    .b(_02548_),
    .c(_03602_),
    .o1(_05301_));
 b15aoi012ar1n02x5 _30973_ (.a(_04184_),
    .b(_05210_),
    .c(_02569_),
    .o1(_05302_));
 b15nandp2aq1n02x5 _30974_ (.a(_05301_),
    .b(_05302_),
    .o1(_05303_));
 b15aoi012ar1n02x5 _30975_ (.a(_02585_),
    .b(_03602_),
    .c(net836),
    .o1(_05304_));
 b15aoi012ar1n02x5 _30976_ (.a(_02548_),
    .b(_05210_),
    .c(_02573_),
    .o1(_05305_));
 b15oai012ah1n02x5 _30977_ (.a(_05304_),
    .b(_05305_),
    .c(_02541_),
    .o1(_05306_));
 b15aoai13al1n02x5 _30978_ (.a(_02573_),
    .b(_02759_),
    .c(_04411_),
    .d(_03626_),
    .o1(_05308_));
 b15oai112an1n08x5 _30979_ (.a(_02631_),
    .b(_05308_),
    .c(_03362_),
    .d(_02645_),
    .o1(_05309_));
 b15norp02ar1n02x5 _30980_ (.a(_03305_),
    .b(_02602_),
    .o1(_05310_));
 b15aoai13al1n04x5 _30981_ (.a(_02694_),
    .b(_05310_),
    .c(_03305_),
    .d(_02569_),
    .o1(_05311_));
 b15and002ar1n02x5 _30982_ (.a(_03305_),
    .b(_03376_),
    .o(_05312_));
 b15aoi012ar1n04x5 _30983_ (.a(_05312_),
    .b(_03577_),
    .c(net828),
    .o1(_05313_));
 b15oaoi13aq1n08x5 _30984_ (.a(_04174_),
    .b(_05311_),
    .c(_05313_),
    .d(_02670_),
    .o1(_05314_));
 b15oai112ah1n08x5 _30985_ (.a(_05303_),
    .b(_05306_),
    .c(_05309_),
    .d(_05314_),
    .o1(_05315_));
 b15aoi012ar1n02x5 _30986_ (.a(_03602_),
    .b(_02723_),
    .c(_02573_),
    .o1(_05316_));
 b15oai112aq1n04x5 _30987_ (.a(net841),
    .b(_04902_),
    .c(_05316_),
    .d(_02654_),
    .o1(_05317_));
 b15norp02ar1n03x5 _30988_ (.a(_02573_),
    .b(_04440_),
    .o1(_05319_));
 b15aoi022al1n02x5 _30989_ (.a(net834),
    .b(_04411_),
    .c(_05171_),
    .d(_02517_),
    .o1(_05320_));
 b15oaoi13as1n02x5 _30990_ (.a(net832),
    .b(_05320_),
    .c(_03605_),
    .d(_02602_),
    .o1(_05321_));
 b15oai013al1n06x5 _30991_ (.a(_05317_),
    .b(_05319_),
    .c(_05321_),
    .d(net841),
    .o1(_05322_));
 b15aoi022ar1n02x5 _30992_ (.a(_02573_),
    .b(_02548_),
    .c(_03370_),
    .d(_03366_),
    .o1(_05323_));
 b15oaoi13an1n02x5 _30993_ (.a(_02752_),
    .b(_02723_),
    .c(_02664_),
    .d(net836),
    .o1(_05324_));
 b15nand02ar1n02x5 _30994_ (.a(_02554_),
    .b(_02654_),
    .o1(_05325_));
 b15oai022aq1n02x5 _30995_ (.a(net832),
    .b(_05323_),
    .c(_05324_),
    .d(_05325_),
    .o1(_05326_));
 b15nand02ar1n02x5 _30996_ (.a(_03391_),
    .b(_03311_),
    .o1(_05327_));
 b15nandp3ar1n02x5 _30997_ (.a(net832),
    .b(_02637_),
    .c(_03626_),
    .o1(_05328_));
 b15aoi012ar1n02x5 _30998_ (.a(net836),
    .b(_05327_),
    .c(_05328_),
    .o1(_05330_));
 b15and003aq1n04x5 _30999_ (.a(_02566_),
    .b(_02559_),
    .c(_02563_),
    .o(_05331_));
 b15oai022ar1n04x5 _31000_ (.a(_02554_),
    .b(_02593_),
    .c(_05221_),
    .d(_02745_),
    .o1(_05332_));
 b15nor003as1n06x5 _31001_ (.a(_05331_),
    .b(_04410_),
    .c(_05332_),
    .o1(_05333_));
 b15nona23an1n12x5 _31002_ (.a(_05326_),
    .b(_05330_),
    .c(_05333_),
    .d(_03548_),
    .out0(_05334_));
 b15nandp2ar1n05x5 _31003_ (.a(_05225_),
    .b(_02692_),
    .o1(_05335_));
 b15norp02ar1n03x5 _31004_ (.a(_02602_),
    .b(_02748_),
    .o1(_05336_));
 b15aoai13an1n06x5 _31005_ (.a(net840),
    .b(_05336_),
    .c(_02709_),
    .d(_05225_),
    .o1(_05337_));
 b15oai112an1n04x5 _31006_ (.a(net837),
    .b(_02716_),
    .c(_02654_),
    .d(_02748_),
    .o1(_05338_));
 b15norp02as1n02x5 _31007_ (.a(_02507_),
    .b(_02748_),
    .o1(_05339_));
 b15aoi012an1n02x5 _31008_ (.a(net833),
    .b(_02662_),
    .c(_02666_),
    .o1(_05341_));
 b15oai013as1n06x5 _31009_ (.a(_05338_),
    .b(_05339_),
    .c(_05341_),
    .d(net837),
    .o1(_05342_));
 b15oai112as1n16x5 _31010_ (.a(_05335_),
    .b(_05337_),
    .c(_05342_),
    .d(net840),
    .o1(_05343_));
 b15aoi013aq1n02x5 _31011_ (.a(net832),
    .b(_03598_),
    .c(_02649_),
    .d(net835),
    .o1(_05344_));
 b15oai012ar1n02x5 _31012_ (.a(_02593_),
    .b(_03299_),
    .c(net835),
    .o1(_05345_));
 b15aob012ar1n08x5 _31013_ (.a(_05344_),
    .b(_05345_),
    .c(_02665_),
    .out0(_05346_));
 b15oai013ah1n03x5 _31014_ (.a(net832),
    .b(_02515_),
    .c(_03549_),
    .d(net842),
    .o1(_05347_));
 b15norp02an1n04x5 _31015_ (.a(_02635_),
    .b(_03592_),
    .o1(_05348_));
 b15oai022an1n02x5 _31016_ (.a(_02545_),
    .b(_03592_),
    .c(_03341_),
    .d(net835),
    .o1(_05349_));
 b15aoi022an1n06x5 _31017_ (.a(_03395_),
    .b(_05348_),
    .c(_05349_),
    .d(net838),
    .o1(_05350_));
 b15aoai13aq1n04x5 _31018_ (.a(net842),
    .b(_03577_),
    .c(_05348_),
    .d(net835),
    .o1(_05352_));
 b15aoai13al1n08x5 _31019_ (.a(_05346_),
    .b(_05347_),
    .c(_05350_),
    .d(_05352_),
    .o1(_05353_));
 b15aob012ar1n02x5 _31020_ (.a(_02569_),
    .b(_02665_),
    .c(_03351_),
    .out0(_05354_));
 b15norp03as1n04x5 _31021_ (.a(_02631_),
    .b(_02557_),
    .c(_02623_),
    .o1(_05355_));
 b15mdn022ar1n02x5 _31022_ (.a(_03351_),
    .b(_05355_),
    .o1(_05356_),
    .sa(net838));
 b15oab012ah1n03x5 _31023_ (.a(_05354_),
    .b(_05356_),
    .c(_02611_),
    .out0(_05357_));
 b15oai013aq1n02x5 _31024_ (.a(net835),
    .b(_02768_),
    .c(_02611_),
    .d(net838),
    .o1(_05358_));
 b15oaoi13al1n04x5 _31025_ (.a(_05358_),
    .b(net838),
    .c(_04178_),
    .d(_05355_),
    .o1(_05359_));
 b15oai112aq1n16x5 _31026_ (.a(_05343_),
    .b(_05353_),
    .c(_05357_),
    .d(_05359_),
    .o1(_05360_));
 b15nano23aq1n24x5 _31027_ (.a(_05315_),
    .b(_05322_),
    .c(_05334_),
    .d(_05360_),
    .out0(_05361_));
 b15aoi012ar1n02x5 _31028_ (.a(_02325_),
    .b(_02469_),
    .c(_02466_),
    .o1(_05363_));
 b15oai012ar1n02x5 _31029_ (.a(_02367_),
    .b(_02475_),
    .c(_05363_),
    .o1(_05364_));
 b15aoi112as1n08x5 _31030_ (.a(_02279_),
    .b(_04035_),
    .c(_04697_),
    .d(_02300_),
    .o1(_05365_));
 b15aoai13al1n02x5 _31031_ (.a(net715),
    .b(_05365_),
    .c(_02354_),
    .d(_02381_),
    .o1(_05366_));
 b15aoai13ar1n03x5 _31032_ (.a(_05364_),
    .b(_03636_),
    .c(_05052_),
    .d(_05366_),
    .o1(_05367_));
 b15oai012ar1n02x5 _31033_ (.a(_02242_),
    .b(_02311_),
    .c(_04364_),
    .o1(_05368_));
 b15oai012ar1n02x5 _31034_ (.a(_02468_),
    .b(_02367_),
    .c(_02325_),
    .o1(_05369_));
 b15aoi012ar1n02x5 _31035_ (.a(_02298_),
    .b(_02357_),
    .c(_03636_),
    .o1(_05370_));
 b15oai012ar1n02x5 _31036_ (.a(_02425_),
    .b(_05369_),
    .c(_05370_),
    .o1(_05371_));
 b15nand04ar1n02x5 _31037_ (.a(_02393_),
    .b(_05085_),
    .c(_05368_),
    .d(_05371_),
    .o1(_05372_));
 b15aoi022al1n04x5 _31038_ (.a(_04037_),
    .b(_02438_),
    .c(_03680_),
    .d(net711),
    .o1(_05374_));
 b15oai012ah1n02x5 _31039_ (.a(net713),
    .b(_04336_),
    .c(_02438_),
    .o1(_05375_));
 b15aoi022an1n02x5 _31040_ (.a(_02411_),
    .b(_04037_),
    .c(_02438_),
    .d(_02461_),
    .o1(_05376_));
 b15oai112ah1n08x5 _31041_ (.a(_05374_),
    .b(_05375_),
    .c(net703),
    .d(_05376_),
    .o1(_05377_));
 b15oai012an1n02x5 _31042_ (.a(net700),
    .b(net715),
    .c(net708),
    .o1(_05378_));
 b15oai022ar1n02x5 _31043_ (.a(net697),
    .b(_02259_),
    .c(_02366_),
    .d(net715),
    .o1(_05379_));
 b15aoi222as1n04x5 _31044_ (.a(_04044_),
    .b(_03710_),
    .c(_05365_),
    .d(_05378_),
    .e(_05379_),
    .f(_02343_),
    .o1(_05380_));
 b15nona23aq1n08x5 _31045_ (.a(_05367_),
    .b(_05372_),
    .c(_05377_),
    .d(_05380_),
    .out0(_05381_));
 b15nand02ar1n02x5 _31046_ (.a(net707),
    .b(_02376_),
    .o1(_05382_));
 b15oaoi13as1n03x5 _31047_ (.a(_02298_),
    .b(_05382_),
    .c(_04330_),
    .d(net711),
    .o1(_05383_));
 b15nandp2al1n03x5 _31048_ (.a(_02381_),
    .b(_03640_),
    .o1(_05385_));
 b15oai012ah1n08x5 _31049_ (.a(_04019_),
    .b(_05383_),
    .c(_05385_),
    .o1(_05386_));
 b15nand03ar1n02x5 _31050_ (.a(net706),
    .b(_03657_),
    .c(_02462_),
    .o1(_05387_));
 b15oai012an1n04x5 _31051_ (.a(_05387_),
    .b(_04110_),
    .c(net713),
    .o1(_05388_));
 b15aoi012al1n06x5 _31052_ (.a(_03661_),
    .b(_05388_),
    .c(net702),
    .o1(_05389_));
 b15nor002al1n02x5 _31053_ (.a(_03666_),
    .b(_03739_),
    .o1(_05390_));
 b15oai012ah1n02x5 _31054_ (.a(_02259_),
    .b(_02309_),
    .c(net710),
    .o1(_05391_));
 b15aoi013ah1n04x5 _31055_ (.a(_05390_),
    .b(_05391_),
    .c(_04712_),
    .d(_02355_),
    .o1(_05392_));
 b15oai112as1n16x5 _31056_ (.a(_05386_),
    .b(_05389_),
    .c(_05392_),
    .d(net709),
    .o1(_05393_));
 b15nand02ar1n02x5 _31057_ (.a(_04336_),
    .b(_03709_),
    .o1(_05394_));
 b15aoi012ar1n02x5 _31058_ (.a(_02313_),
    .b(_03709_),
    .c(_02242_),
    .o1(_05396_));
 b15oaoi13as1n03x5 _31059_ (.a(net705),
    .b(_05394_),
    .c(_05396_),
    .d(_02300_),
    .o1(_05397_));
 b15norp02ar1n02x5 _31060_ (.a(\us12.a[1] ),
    .b(_02259_),
    .o1(_05398_));
 b15aoi013al1n02x5 _31061_ (.a(_05398_),
    .b(_03657_),
    .c(net695),
    .d(net692),
    .o1(_05399_));
 b15oai022ah1n04x5 _31062_ (.a(_02259_),
    .b(_02427_),
    .c(_05399_),
    .d(_02461_),
    .o1(_05400_));
 b15aoi013an1n08x5 _31063_ (.a(_05397_),
    .b(_05400_),
    .c(_02346_),
    .d(net705),
    .o1(_05401_));
 b15norp02ar1n02x5 _31064_ (.a(_02471_),
    .b(_02457_),
    .o1(_05402_));
 b15oai112as1n04x5 _31065_ (.a(_02461_),
    .b(_02355_),
    .c(_03701_),
    .d(_05402_),
    .o1(_05403_));
 b15aoi012ar1n02x5 _31066_ (.a(net712),
    .b(net706),
    .c(_04706_),
    .o1(_05404_));
 b15oai012aq1n06x5 _31067_ (.a(net705),
    .b(_05404_),
    .c(_02298_),
    .o1(_05405_));
 b15aoi012ar1n02x5 _31068_ (.a(net712),
    .b(_03677_),
    .c(_03651_),
    .o1(_05407_));
 b15oai013an1n02x5 _31069_ (.a(_03677_),
    .b(_03648_),
    .c(_02309_),
    .d(net714),
    .o1(_05408_));
 b15aoi012ar1n04x5 _31070_ (.a(_05407_),
    .b(_05408_),
    .c(_02461_),
    .o1(_05409_));
 b15oai012an1n12x5 _31071_ (.a(_05403_),
    .b(_05405_),
    .c(_05409_),
    .o1(_05410_));
 b15aoi022aq1n02x5 _31072_ (.a(_02411_),
    .b(_02328_),
    .c(_02351_),
    .d(_02461_),
    .o1(_05411_));
 b15oaoi13an1n04x5 _31073_ (.a(net703),
    .b(_04109_),
    .c(_05411_),
    .d(_02242_),
    .o1(_05412_));
 b15oai013as1n04x5 _31074_ (.a(_02251_),
    .b(_02351_),
    .c(_03758_),
    .d(_03755_),
    .o1(_05413_));
 b15aoi022al1n02x5 _31075_ (.a(_02328_),
    .b(_04045_),
    .c(_02475_),
    .d(_02343_),
    .o1(_05414_));
 b15oai112as1n06x5 _31076_ (.a(_05413_),
    .b(_05414_),
    .c(_04037_),
    .d(_02389_),
    .o1(_05415_));
 b15aoi112as1n08x5 _31077_ (.a(_05410_),
    .b(_05412_),
    .c(net713),
    .d(_05415_),
    .o1(_05416_));
 b15nona23as1n32x5 _31078_ (.a(_05381_),
    .b(_05393_),
    .c(_05401_),
    .d(_05416_),
    .out0(_05418_));
 b15xor002an1n16x5 _31079_ (.a(_05361_),
    .b(_05418_),
    .out0(_05419_));
 b15aob012ar1n02x5 _31080_ (.a(net858),
    .b(net860),
    .c(net851),
    .out0(_05420_));
 b15nand04aq1n04x5 _31081_ (.a(_02904_),
    .b(_02899_),
    .c(_03447_),
    .d(_05420_),
    .o1(_05421_));
 b15aoi013ar1n02x5 _31082_ (.a(net855),
    .b(_02899_),
    .c(_02781_),
    .d(_02820_),
    .o1(_05422_));
 b15oai112aq1n02x5 _31083_ (.a(_05421_),
    .b(_05422_),
    .c(_02921_),
    .d(_04539_),
    .o1(_05423_));
 b15nand02ar1n02x5 _31084_ (.a(_02885_),
    .b(_03524_),
    .o1(_05424_));
 b15oaoi13ar1n02x5 _31085_ (.a(_02951_),
    .b(_05424_),
    .c(_02964_),
    .d(_02811_),
    .o1(_05425_));
 b15oai012ar1n02x5 _31086_ (.a(_02811_),
    .b(_02932_),
    .c(_02974_),
    .o1(_05426_));
 b15oaoi13ah1n02x5 _31087_ (.a(net858),
    .b(_05426_),
    .c(_02942_),
    .d(_02820_),
    .o1(_05427_));
 b15oai012an1n02x5 _31088_ (.a(net855),
    .b(_02923_),
    .c(_02942_),
    .o1(_05429_));
 b15oai022al1n04x5 _31089_ (.a(_05423_),
    .b(_05425_),
    .c(_05427_),
    .d(_05429_),
    .o1(_05430_));
 b15nandp2an1n05x5 _31090_ (.a(net850),
    .b(_02885_),
    .o1(_05431_));
 b15obai22an1n04x5 _31091_ (.a(_02985_),
    .b(_05431_),
    .c(_04221_),
    .d(_02867_),
    .out0(_05432_));
 b15aoi012ar1n02x5 _31092_ (.a(net858),
    .b(_02820_),
    .c(_02787_),
    .o1(_05433_));
 b15oai012ar1n02x5 _31093_ (.a(_02864_),
    .b(_03447_),
    .c(_02951_),
    .o1(_05434_));
 b15norp03ah1n03x5 _31094_ (.a(_02929_),
    .b(_05433_),
    .c(_05434_),
    .o1(_05435_));
 b15aoai13ar1n02x5 _31095_ (.a(_03453_),
    .b(net860),
    .c(_02862_),
    .d(_02918_),
    .o1(_05436_));
 b15aoi112aq1n03x5 _31096_ (.a(_05432_),
    .b(_05435_),
    .c(_05436_),
    .d(_02977_),
    .o1(_05437_));
 b15qgbno2an1n10x5 _31097_ (.a(net857),
    .b(_02854_),
    .o1(_05438_));
 b15oaoi13as1n02x5 _31098_ (.a(net850),
    .b(_02954_),
    .c(_02921_),
    .d(_05438_),
    .o1(_05440_));
 b15aoai13aq1n02x5 _31099_ (.a(net857),
    .b(_03002_),
    .c(_02921_),
    .d(_03460_),
    .o1(_05441_));
 b15aoi012al1n04x5 _31100_ (.a(_04285_),
    .b(_05440_),
    .c(_05441_),
    .o1(_05442_));
 b15nand04ah1n06x5 _31101_ (.a(_02833_),
    .b(_02844_),
    .c(_02920_),
    .d(_02882_),
    .o1(_05443_));
 b15nand02al1n06x5 _31102_ (.a(_02915_),
    .b(_03524_),
    .o1(_05444_));
 b15aoi022al1n08x5 _31103_ (.a(net854),
    .b(_02904_),
    .c(_02781_),
    .d(_02989_),
    .o1(_05445_));
 b15oai112al1n16x5 _31104_ (.a(_03516_),
    .b(_05443_),
    .c(_05444_),
    .d(_05445_),
    .o1(_05446_));
 b15oai022an1n02x5 _31105_ (.a(_02873_),
    .b(_02918_),
    .c(_05148_),
    .d(_02940_),
    .o1(_05447_));
 b15aoi012an1n02x5 _31106_ (.a(_05446_),
    .b(_05447_),
    .c(net858),
    .o1(_05448_));
 b15nand04an1n08x5 _31107_ (.a(_05430_),
    .b(_05437_),
    .c(_05442_),
    .d(_05448_),
    .o1(_05449_));
 b15oai022al1n04x5 _31108_ (.a(_02956_),
    .b(_02964_),
    .c(_02921_),
    .d(_02873_),
    .o1(_05451_));
 b15norp02as1n02x5 _31109_ (.a(_04539_),
    .b(_05119_),
    .o1(_05452_));
 b15aoi112al1n02x5 _31110_ (.a(net853),
    .b(_02956_),
    .c(_02918_),
    .d(_02950_),
    .o1(_05453_));
 b15oai013ah1n04x5 _31111_ (.a(net860),
    .b(_05451_),
    .c(_05452_),
    .d(_05453_),
    .o1(_05454_));
 b15aoi022ar1n02x5 _31112_ (.a(_02779_),
    .b(_02781_),
    .c(_02871_),
    .d(_02974_),
    .o1(_05455_));
 b15norp03ah1n03x5 _31113_ (.a(_02873_),
    .b(_02911_),
    .c(_05455_),
    .o1(_05456_));
 b15oai022ar1n02x5 _31114_ (.a(net858),
    .b(_03469_),
    .c(_03460_),
    .d(_02956_),
    .o1(_05457_));
 b15oab012ah1n02x5 _31115_ (.a(_05456_),
    .b(_05457_),
    .c(_02913_),
    .out0(_05458_));
 b15norp02ar1n03x5 _31116_ (.a(_02986_),
    .b(_03020_),
    .o1(_05459_));
 b15oaoi13an1n03x5 _31117_ (.a(_02951_),
    .b(_02862_),
    .c(_02986_),
    .d(net860),
    .o1(_05460_));
 b15norp03al1n08x5 _31118_ (.a(_03470_),
    .b(_05459_),
    .c(_05460_),
    .o1(_05462_));
 b15oai112al1n16x5 _31119_ (.a(_05454_),
    .b(_05458_),
    .c(_05462_),
    .d(_02864_),
    .o1(_05463_));
 b15aoi012ar1n02x5 _31120_ (.a(_03002_),
    .b(_03460_),
    .c(net857),
    .o1(_05464_));
 b15oai112as1n02x5 _31121_ (.a(_02811_),
    .b(_04221_),
    .c(_05464_),
    .d(_02984_),
    .o1(_05465_));
 b15oai022ar1n02x5 _31122_ (.a(net854),
    .b(_02862_),
    .c(_02997_),
    .d(net857),
    .o1(_05466_));
 b15aoi122ah1n02x5 _31123_ (.a(_05465_),
    .b(_03461_),
    .c(_03023_),
    .d(net861),
    .e(_05466_),
    .o1(_05467_));
 b15nandp2ah1n03x5 _31124_ (.a(_02904_),
    .b(_02907_),
    .o1(_05468_));
 b15norp03ar1n02x5 _31125_ (.a(net854),
    .b(net846),
    .c(_03522_),
    .o1(_05469_));
 b15oai012al1n06x5 _31126_ (.a(_02808_),
    .b(_03500_),
    .c(net845),
    .o1(_05470_));
 b15aoi013ar1n02x5 _31127_ (.a(_05469_),
    .b(_05470_),
    .c(_02820_),
    .d(net843),
    .o1(_05471_));
 b15oai012al1n03x5 _31128_ (.a(_05468_),
    .b(_05471_),
    .c(net848),
    .o1(_05473_));
 b15aob012aq1n08x5 _31129_ (.a(_05467_),
    .b(_05473_),
    .c(net857),
    .out0(_05474_));
 b15oaoi13al1n02x5 _31130_ (.a(_04243_),
    .b(_03029_),
    .c(net858),
    .d(_02950_),
    .o1(_05475_));
 b15nand04ar1n02x5 _31131_ (.a(net860),
    .b(net855),
    .c(_02779_),
    .d(_02781_),
    .o1(_05476_));
 b15oaoi13ar1n02x5 _31132_ (.a(_02951_),
    .b(_05476_),
    .c(_03029_),
    .d(net860),
    .o1(_05477_));
 b15nand03an1n12x5 _31133_ (.a(net857),
    .b(_02833_),
    .c(_02920_),
    .o1(_05478_));
 b15aoi122al1n02x5 _31134_ (.a(_03460_),
    .b(_02984_),
    .c(_05478_),
    .d(_03002_),
    .e(net858),
    .o1(_05479_));
 b15nor003an1n03x5 _31135_ (.a(_05475_),
    .b(_05477_),
    .c(_05479_),
    .o1(_05480_));
 b15nand02ar1n02x5 _31136_ (.a(_02954_),
    .b(_04871_),
    .o1(_05481_));
 b15aoai13as1n02x5 _31137_ (.a(_05481_),
    .b(_02882_),
    .c(_02951_),
    .d(_02900_),
    .o1(_05482_));
 b15nand03ah1n06x5 _31138_ (.a(net850),
    .b(_05480_),
    .c(_05482_),
    .o1(_05484_));
 b15aoi112as1n08x5 _31139_ (.a(_05449_),
    .b(_05463_),
    .c(_05474_),
    .d(_05484_),
    .o1(_05485_));
 b15xor002as1n08x5 _31140_ (.a(_05229_),
    .b(_05485_),
    .out0(_05486_));
 b15xor003an1n04x5 _31141_ (.a(_05300_),
    .b(_05419_),
    .c(_05486_),
    .out0(_05487_));
 b15norp02ar1n02x5 _31142_ (.a(net542),
    .b(_05487_),
    .o1(_05488_));
 b15inv040ah1n02x5 _31143_ (.a(\text_in_r[70] ),
    .o1(_05489_));
 b15aoi012ar1n02x5 _31144_ (.a(_05488_),
    .b(_05489_),
    .c(net542),
    .o1(_05490_));
 b15xor002an1n02x5 _31145_ (.a(\u0.w[1][6] ),
    .b(_05490_),
    .out0(_00111_));
 b15aoi112ar1n02x5 _31146_ (.a(net854),
    .b(_03024_),
    .c(_02844_),
    .d(_03523_),
    .o1(_05491_));
 b15aoi022an1n02x5 _31147_ (.a(net850),
    .b(_02799_),
    .c(_02827_),
    .d(_02908_),
    .o1(_05492_));
 b15aoi012as1n02x5 _31148_ (.a(_05491_),
    .b(_05492_),
    .c(net854),
    .o1(_05494_));
 b15nor002as1n02x5 _31149_ (.a(_03522_),
    .b(_03482_),
    .o1(_05495_));
 b15oai012as1n03x5 _31150_ (.a(_05438_),
    .b(_05495_),
    .c(net850),
    .o1(_05496_));
 b15oai012as1n04x5 _31151_ (.a(_02811_),
    .b(_02854_),
    .c(_05495_),
    .o1(_05497_));
 b15oai112ar1n16x5 _31152_ (.a(net861),
    .b(_05496_),
    .c(_05497_),
    .d(_02951_),
    .o1(_05498_));
 b15aoai13ah1n04x5 _31153_ (.a(net861),
    .b(_05494_),
    .c(_05498_),
    .d(_03483_),
    .o1(_05499_));
 b15aoi012ar1n02x5 _31154_ (.a(_03460_),
    .b(_02882_),
    .c(_02951_),
    .o1(_05500_));
 b15oai022ar1n02x5 _31155_ (.a(net857),
    .b(_02834_),
    .c(_02997_),
    .d(_05500_),
    .o1(_05501_));
 b15aoi022ar1n02x5 _31156_ (.a(_03460_),
    .b(_02898_),
    .c(_02974_),
    .d(_03002_),
    .o1(_05502_));
 b15aoai13ar1n02x5 _31157_ (.a(_02951_),
    .b(_02974_),
    .c(_02898_),
    .d(_03002_),
    .o1(_05503_));
 b15nona23al1n04x5 _31158_ (.a(_02811_),
    .b(_05501_),
    .c(_05502_),
    .d(_05503_),
    .out0(_05505_));
 b15aoai13aq1n03x5 _31159_ (.a(_02854_),
    .b(_04480_),
    .c(_02974_),
    .d(_02820_),
    .o1(_05506_));
 b15oab012as1n02x5 _31160_ (.a(_04867_),
    .b(_05119_),
    .c(_02820_),
    .out0(_05507_));
 b15oai012as1n08x5 _31161_ (.a(_05506_),
    .b(_05507_),
    .c(_02951_),
    .o1(_05508_));
 b15aoai13ar1n04x5 _31162_ (.a(_04286_),
    .b(net857),
    .c(_02992_),
    .d(_03427_),
    .o1(_05509_));
 b15oai013aq1n08x5 _31163_ (.a(_05505_),
    .b(_05508_),
    .c(_05509_),
    .d(net850),
    .o1(_05510_));
 b15aob012ar1n02x5 _31164_ (.a(net858),
    .b(_02864_),
    .c(_02858_),
    .out0(_05511_));
 b15nand02ar1n02x5 _31165_ (.a(net860),
    .b(_02864_),
    .o1(_05512_));
 b15aoai13ar1n02x5 _31166_ (.a(_05511_),
    .b(_02900_),
    .c(_02782_),
    .d(_05512_),
    .o1(_05513_));
 b15oaoi13ar1n02x5 _31167_ (.a(net850),
    .b(net855),
    .c(_02782_),
    .d(_02957_),
    .o1(_05514_));
 b15oab012al1n04x5 _31168_ (.a(_04523_),
    .b(_05513_),
    .c(_05514_),
    .out0(_05516_));
 b15aoi012al1n02x5 _31169_ (.a(net858),
    .b(_02864_),
    .c(_04227_),
    .o1(_05517_));
 b15nand04ah1n08x5 _31170_ (.a(net851),
    .b(_02831_),
    .c(_02915_),
    .d(_04265_),
    .o1(_05518_));
 b15oaoi13ar1n08x5 _31171_ (.a(_05517_),
    .b(_05518_),
    .c(_02862_),
    .d(net851),
    .o1(_05519_));
 b15aoi022ar1n02x5 _31172_ (.a(_02908_),
    .b(_03524_),
    .c(_03514_),
    .d(_03024_),
    .o1(_05520_));
 b15nand02an1n02x5 _31173_ (.a(_02951_),
    .b(_05520_),
    .o1(_05521_));
 b15oai022aq1n04x5 _31174_ (.a(_02940_),
    .b(_02954_),
    .c(_02867_),
    .d(_02986_),
    .o1(_05522_));
 b15oaoi13ah1n04x5 _31175_ (.a(_05519_),
    .b(_05521_),
    .c(_05522_),
    .d(_02951_),
    .o1(_05523_));
 b15oaoi13ah1n03x5 _31176_ (.a(net850),
    .b(_04843_),
    .c(_04828_),
    .d(_03029_),
    .o1(_05524_));
 b15oaoi13an1n04x5 _31177_ (.a(_02882_),
    .b(_04542_),
    .c(_02892_),
    .d(_02950_),
    .o1(_05525_));
 b15oai022as1n02x5 _31178_ (.a(_02867_),
    .b(_02876_),
    .c(_02984_),
    .d(_02858_),
    .o1(_05527_));
 b15aoi112as1n04x5 _31179_ (.a(_05524_),
    .b(_05525_),
    .c(_05527_),
    .d(_05438_),
    .o1(_05528_));
 b15norp02ar1n02x5 _31180_ (.a(_02820_),
    .b(_02876_),
    .o1(_05529_));
 b15aoai13al1n02x5 _31181_ (.a(_03469_),
    .b(_05529_),
    .c(_02911_),
    .d(_02782_),
    .o1(_05530_));
 b15aoi112aq1n02x5 _31182_ (.a(_02873_),
    .b(_02877_),
    .c(_02913_),
    .d(_05478_),
    .o1(_05531_));
 b15aoi112as1n02x5 _31183_ (.a(_02811_),
    .b(_02943_),
    .c(_04494_),
    .d(_02918_),
    .o1(_05532_));
 b15nano23al1n06x5 _31184_ (.a(_03471_),
    .b(_05530_),
    .c(_05531_),
    .d(_05532_),
    .out0(_05533_));
 b15nand04as1n16x5 _31185_ (.a(_05516_),
    .b(_05523_),
    .c(_05528_),
    .d(_05533_),
    .o1(_05534_));
 b15aoi012ar1n02x5 _31186_ (.a(_02820_),
    .b(_05468_),
    .c(_05431_),
    .o1(_05535_));
 b15nor003al1n02x5 _31187_ (.a(net861),
    .b(_02940_),
    .c(_02984_),
    .o1(_05536_));
 b15oai022an1n02x5 _31188_ (.a(_02954_),
    .b(_02873_),
    .c(_02948_),
    .d(_02950_),
    .o1(_05538_));
 b15oai013aq1n04x5 _31189_ (.a(net857),
    .b(_05535_),
    .c(_05536_),
    .d(_05538_),
    .o1(_05539_));
 b15orn003an1n02x5 _31190_ (.a(_04302_),
    .b(_03029_),
    .c(_04539_),
    .o(_05540_));
 b15oai012ar1n06x5 _31191_ (.a(_02864_),
    .b(_02787_),
    .c(_02951_),
    .o1(_05541_));
 b15oai122ar1n12x5 _31192_ (.a(_05540_),
    .b(_05541_),
    .c(_02921_),
    .d(_02929_),
    .e(net850),
    .o1(_05542_));
 b15aob012al1n12x5 _31193_ (.a(_05539_),
    .b(_05542_),
    .c(_05498_),
    .out0(_05543_));
 b15nano23as1n24x5 _31194_ (.a(_05499_),
    .b(_05510_),
    .c(_05534_),
    .d(_05543_),
    .out0(_05544_));
 b15nandp2al1n02x5 _31195_ (.a(_02485_),
    .b(_02488_),
    .o1(_05545_));
 b15aoi112aq1n02x5 _31196_ (.a(_02304_),
    .b(_02389_),
    .c(_04035_),
    .d(_04060_),
    .o1(_05546_));
 b15nor004ar1n02x5 _31197_ (.a(net705),
    .b(_02317_),
    .c(_02318_),
    .d(_02300_),
    .o1(_05547_));
 b15oai012ah1n02x5 _31198_ (.a(net712),
    .b(_05546_),
    .c(_05547_),
    .o1(_05549_));
 b15nona23ar1n02x5 _31199_ (.a(\us12.a[4] ),
    .b(net705),
    .c(net709),
    .d(net712),
    .out0(_05550_));
 b15nanb03ar1n02x5 _31200_ (.a(net698),
    .b(net693),
    .c(\us12.a[6] ),
    .out0(_05551_));
 b15oaoi13ar1n03x5 _31201_ (.a(_05550_),
    .b(_05551_),
    .c(_02419_),
    .d(_02259_),
    .o1(_05552_));
 b15nona23ar1n02x5 _31202_ (.a(net698),
    .b(\us12.a[4] ),
    .c(\us12.a[6] ),
    .d(net705),
    .out0(_05553_));
 b15aob012as1n03x5 _31203_ (.a(_05553_),
    .b(_05046_),
    .c(_02437_),
    .out0(_05554_));
 b15aoi013an1n06x5 _31204_ (.a(_05552_),
    .b(_05554_),
    .c(net693),
    .d(_02415_),
    .o1(_05555_));
 b15norp03al1n02x5 _31205_ (.a(net698),
    .b(_02381_),
    .c(_02259_),
    .o1(_05556_));
 b15oai012ar1n02x5 _31206_ (.a(_02418_),
    .b(_04657_),
    .c(net699),
    .o1(_05557_));
 b15oai012ar1n02x5 _31207_ (.a(_03677_),
    .b(_03695_),
    .c(_02317_),
    .o1(_05558_));
 b15aoi022aq1n02x5 _31208_ (.a(_05556_),
    .b(_05557_),
    .c(_05558_),
    .d(_03745_),
    .o1(_05560_));
 b15norp03ar1n02x5 _31209_ (.a(net691),
    .b(_02298_),
    .c(_03695_),
    .o1(_05561_));
 b15aoai13ar1n03x5 _31210_ (.a(_02251_),
    .b(_05561_),
    .c(_02433_),
    .d(_02319_),
    .o1(_05562_));
 b15nand04al1n06x5 _31211_ (.a(_05549_),
    .b(_05555_),
    .c(_05560_),
    .d(_05562_),
    .o1(_05563_));
 b15aoi012ar1n04x5 _31212_ (.a(_03699_),
    .b(_02468_),
    .c(_02324_),
    .o1(_05564_));
 b15aoai13al1n08x5 _31213_ (.a(net715),
    .b(_05564_),
    .c(_03644_),
    .d(_04364_),
    .o1(_05565_));
 b15oaoi13ar1n02x5 _31214_ (.a(\us12.a[2] ),
    .b(_02469_),
    .c(_02471_),
    .d(_03657_),
    .o1(_05566_));
 b15norp03ar1n02x5 _31215_ (.a(_02309_),
    .b(_03657_),
    .c(_03648_),
    .o1(_05567_));
 b15nor003aq1n02x5 _31216_ (.a(_02327_),
    .b(_03695_),
    .c(_04657_),
    .o1(_05568_));
 b15oai013ar1n02x5 _31217_ (.a(_02381_),
    .b(_05566_),
    .c(_05567_),
    .d(_05568_),
    .o1(_05569_));
 b15aoi012ar1n02x5 _31218_ (.a(\us12.a[1] ),
    .b(_02381_),
    .c(_02471_),
    .o1(_05571_));
 b15mdn022an1n02x5 _31219_ (.a(_02492_),
    .b(_02493_),
    .o1(_05572_),
    .sa(_03752_));
 b15aoai13ah1n02x5 _31220_ (.a(_05571_),
    .b(_02381_),
    .c(net692),
    .d(_05572_),
    .o1(_05573_));
 b15oaoi13ar1n02x5 _31221_ (.a(_02390_),
    .b(_04662_),
    .c(_03695_),
    .d(_02327_),
    .o1(_05574_));
 b15oai022ar1n02x5 _31222_ (.a(_02317_),
    .b(_03695_),
    .c(_04662_),
    .d(net715),
    .o1(_05575_));
 b15aoai13ar1n02x5 _31223_ (.a(_02343_),
    .b(_05574_),
    .c(_05575_),
    .d(_02242_),
    .o1(_05576_));
 b15nand04ah1n02x5 _31224_ (.a(_05565_),
    .b(_05569_),
    .c(_05573_),
    .d(_05576_),
    .o1(_05577_));
 b15nor004an1n03x5 _31225_ (.a(_05545_),
    .b(_03747_),
    .c(_05563_),
    .d(_05577_),
    .o1(_05578_));
 b15nand02ar1n02x5 _31226_ (.a(net698),
    .b(\us12.a[6] ),
    .o1(_05579_));
 b15nanb03ar1n02x5 _31227_ (.a(net709),
    .b(net705),
    .c(\us12.a[4] ),
    .out0(_05580_));
 b15oaoi13aq1n03x5 _31228_ (.a(_05579_),
    .b(_05580_),
    .c(\us12.a[4] ),
    .d(_02320_),
    .o1(_05582_));
 b15norp03al1n03x5 _31229_ (.a(\us12.a[6] ),
    .b(_02320_),
    .c(_02318_),
    .o1(_05583_));
 b15oai112as1n08x5 _31230_ (.a(net693),
    .b(_02449_),
    .c(_05582_),
    .d(_05583_),
    .o1(_05584_));
 b15oai022ar1n02x5 _31231_ (.a(_02324_),
    .b(_03657_),
    .c(_02325_),
    .d(_02389_),
    .o1(_05585_));
 b15oai012al1n02x5 _31232_ (.a(_04044_),
    .b(_02392_),
    .c(_05585_),
    .o1(_05586_));
 b15nand02ar1n02x5 _31233_ (.a(_02313_),
    .b(_04016_),
    .o1(_05587_));
 b15aob012al1n06x5 _31234_ (.a(net703),
    .b(_04109_),
    .c(_05587_),
    .out0(_05588_));
 b15oai022ar1n02x5 _31235_ (.a(_02457_),
    .b(_02469_),
    .c(_03673_),
    .d(net705),
    .o1(_05589_));
 b15nand02aq1n02x5 _31236_ (.a(_02412_),
    .b(_05589_),
    .o1(_05590_));
 b15nand04ah1n04x5 _31237_ (.a(_05584_),
    .b(_05586_),
    .c(_05588_),
    .d(_05590_),
    .o1(_05591_));
 b15nandp3ar1n02x5 _31238_ (.a(_02466_),
    .b(_02433_),
    .c(_03699_),
    .o1(_05593_));
 b15oai112ar1n02x5 _31239_ (.a(_02367_),
    .b(_05593_),
    .c(_03697_),
    .d(_02433_),
    .o1(_05594_));
 b15nandp2al1n03x5 _31240_ (.a(_04077_),
    .b(_05594_),
    .o1(_05595_));
 b15oai012aq1n03x5 _31241_ (.a(_03667_),
    .b(_02390_),
    .c(net709),
    .o1(_05596_));
 b15oai022al1n02x5 _31242_ (.a(_02357_),
    .b(_03697_),
    .c(_03764_),
    .d(net703),
    .o1(_05597_));
 b15aoi112an1n04x5 _31243_ (.a(_05596_),
    .b(_05597_),
    .c(_05052_),
    .d(net709),
    .o1(_05598_));
 b15aoi112ar1n02x5 _31244_ (.a(_02320_),
    .b(_02390_),
    .c(_03699_),
    .d(_02469_),
    .o1(_05599_));
 b15aoi022ar1n02x5 _31245_ (.a(_05080_),
    .b(_02415_),
    .c(_04033_),
    .d(_04336_),
    .o1(_05600_));
 b15norp03ar1n02x5 _31246_ (.a(_04060_),
    .b(_04709_),
    .c(_05600_),
    .o1(_05601_));
 b15aoi022as1n06x5 _31247_ (.a(_02426_),
    .b(_04088_),
    .c(_04085_),
    .d(net694),
    .o1(_05602_));
 b15nor004ah1n12x5 _31248_ (.a(net699),
    .b(net691),
    .c(_04359_),
    .d(_05602_),
    .o1(_05604_));
 b15orn003an1n03x5 _31249_ (.a(_05599_),
    .b(_05601_),
    .c(_05604_),
    .o(_05605_));
 b15nor004as1n06x5 _31250_ (.a(_05591_),
    .b(_05595_),
    .c(_05598_),
    .d(_05605_),
    .o1(_05606_));
 b15nand03al1n08x5 _31251_ (.a(_05043_),
    .b(_05578_),
    .c(_05606_),
    .o1(_05607_));
 b15xor002as1n16x5 _31252_ (.a(_03413_),
    .b(net396),
    .out0(_05608_));
 b15aoai13al1n02x5 _31253_ (.a(_03134_),
    .b(_04608_),
    .c(_03075_),
    .d(_03088_),
    .o1(_05609_));
 b15nor002as1n03x5 _31254_ (.a(net576),
    .b(net569),
    .o1(_05610_));
 b15nand03al1n02x5 _31255_ (.a(_05610_),
    .b(_04978_),
    .c(_03984_),
    .o1(_05611_));
 b15oai112ah1n04x5 _31256_ (.a(_03917_),
    .b(_05609_),
    .c(_05611_),
    .d(net580),
    .o1(_05612_));
 b15nor003al1n02x5 _31257_ (.a(net578),
    .b(net572),
    .c(_03253_),
    .o1(_05613_));
 b15and003ar1n02x5 _31258_ (.a(net578),
    .b(net572),
    .c(_03253_),
    .o(_05615_));
 b15oai112al1n06x5 _31259_ (.a(_05610_),
    .b(_03775_),
    .c(_05613_),
    .d(_05615_),
    .o1(_05616_));
 b15oai013ar1n02x5 _31260_ (.a(net581),
    .b(_03281_),
    .c(_03149_),
    .d(net585),
    .o1(_05617_));
 b15aoi012ar1n02x5 _31261_ (.a(net587),
    .b(_03137_),
    .c(_03798_),
    .o1(_05618_));
 b15aoi012ar1n02x5 _31262_ (.a(_03137_),
    .b(_03149_),
    .c(_03067_),
    .o1(_05619_));
 b15oai013aq1n03x5 _31263_ (.a(_05616_),
    .b(_05617_),
    .c(_05618_),
    .d(_05619_),
    .o1(_05620_));
 b15aoai13as1n02x5 _31264_ (.a(net587),
    .b(_04976_),
    .c(_03964_),
    .d(_03807_),
    .o1(_05621_));
 b15oai022an1n04x5 _31265_ (.a(_03123_),
    .b(_03135_),
    .c(_03144_),
    .d(_03086_),
    .o1(_05622_));
 b15nand03ar1n12x5 _31266_ (.a(_03251_),
    .b(_03853_),
    .c(_05622_),
    .o1(_05623_));
 b15norp03al1n02x5 _31267_ (.a(net578),
    .b(net572),
    .c(net586),
    .o1(_05624_));
 b15aoai13aq1n04x5 _31268_ (.a(_05272_),
    .b(_05624_),
    .c(net586),
    .d(_05267_),
    .o1(_05626_));
 b15nandp3ar1n03x5 _31269_ (.a(_05621_),
    .b(_05623_),
    .c(_05626_),
    .o1(_05627_));
 b15oai022as1n02x5 _31270_ (.a(_04582_),
    .b(_04792_),
    .c(_04726_),
    .d(_03100_),
    .o1(_05628_));
 b15nand04an1n08x5 _31271_ (.a(_03223_),
    .b(_03097_),
    .c(_03129_),
    .d(_05628_),
    .o1(_05629_));
 b15norp02ar1n02x5 _31272_ (.a(net581),
    .b(_03187_),
    .o1(_05630_));
 b15aoi012ar1n02x5 _31273_ (.a(_05630_),
    .b(_03962_),
    .c(net581),
    .o1(_05631_));
 b15oai012al1n02x5 _31274_ (.a(_05629_),
    .b(_05631_),
    .c(_03075_),
    .o1(_05632_));
 b15nor004ah1n03x5 _31275_ (.a(_05612_),
    .b(_05620_),
    .c(_05627_),
    .d(_05632_),
    .o1(_05633_));
 b15orn002al1n02x5 _31276_ (.a(net574),
    .b(net584),
    .o(_05634_));
 b15aoi112as1n04x5 _31277_ (.a(_03175_),
    .b(_03782_),
    .c(_03179_),
    .d(_05634_),
    .o1(_05635_));
 b15nor004ah1n03x5 _31278_ (.a(net580),
    .b(_03047_),
    .c(_03192_),
    .d(_05635_),
    .o1(_05637_));
 b15oai012ar1n02x5 _31279_ (.a(net580),
    .b(_03044_),
    .c(_03912_),
    .o1(_05638_));
 b15nanb03ar1n02x5 _31280_ (.a(net577),
    .b(net571),
    .c(net584),
    .out0(_05639_));
 b15nona22ar1n02x5 _31281_ (.a(net571),
    .b(net584),
    .c(net577),
    .out0(_05640_));
 b15aoi112an1n02x5 _31282_ (.a(_03163_),
    .b(_04757_),
    .c(_05639_),
    .d(_05640_),
    .o1(_05641_));
 b15nanb03ar1n02x5 _31283_ (.a(net569),
    .b(net591),
    .c(net576),
    .out0(_05642_));
 b15aoi112ar1n02x5 _31284_ (.a(_03181_),
    .b(_04565_),
    .c(_04792_),
    .d(_05642_),
    .o1(_05643_));
 b15norp03aq1n03x5 _31285_ (.a(_05638_),
    .b(_05641_),
    .c(_05643_),
    .o1(_05644_));
 b15aoai13ah1n02x5 _31286_ (.a(net591),
    .b(_03047_),
    .c(_03171_),
    .d(_03163_),
    .o1(_05645_));
 b15aoi022ar1n02x5 _31287_ (.a(net588),
    .b(_03171_),
    .c(_03199_),
    .d(_03102_),
    .o1(_05646_));
 b15nanb02aq1n02x5 _31288_ (.a(_05646_),
    .b(net584),
    .out0(_05648_));
 b15aoi013an1n04x5 _31289_ (.a(_05637_),
    .b(_05644_),
    .c(_05645_),
    .d(_05648_),
    .o1(_05649_));
 b15oai012as1n04x5 _31290_ (.a(_03036_),
    .b(_03068_),
    .c(_03071_),
    .o1(_05650_));
 b15aoi012aq1n02x5 _31291_ (.a(_03123_),
    .b(_03827_),
    .c(_05650_),
    .o1(_05651_));
 b15aoi013al1n03x5 _31292_ (.a(_03089_),
    .b(_03912_),
    .c(_03827_),
    .d(_04591_),
    .o1(_05652_));
 b15oai012as1n03x5 _31293_ (.a(net580),
    .b(_03079_),
    .c(_03053_),
    .o1(_05653_));
 b15aoai13al1n06x5 _31294_ (.a(_04587_),
    .b(net587),
    .c(_05653_),
    .d(_05650_),
    .o1(_05654_));
 b15aoi112ar1n06x5 _31295_ (.a(_05651_),
    .b(_05652_),
    .c(net591),
    .d(_05654_),
    .o1(_05655_));
 b15oai013ar1n02x5 _31296_ (.a(net580),
    .b(_03079_),
    .c(_03281_),
    .d(_03071_),
    .o1(_05656_));
 b15aoi013aq1n03x5 _31297_ (.a(_05656_),
    .b(_05267_),
    .c(_03984_),
    .d(_05610_),
    .o1(_05657_));
 b15nor004an1n03x5 _31298_ (.a(net574),
    .b(net571),
    .c(_03253_),
    .d(_04006_),
    .o1(_05659_));
 b15aoai13ah1n04x5 _31299_ (.a(_03223_),
    .b(_05659_),
    .c(_04767_),
    .d(_04008_),
    .o1(_05660_));
 b15nano23ar1n02x5 _31300_ (.a(net591),
    .b(_03074_),
    .c(_03087_),
    .d(net569),
    .out0(_05661_));
 b15aoi112ar1n02x5 _31301_ (.a(net580),
    .b(_05661_),
    .c(_03255_),
    .d(_03137_),
    .o1(_05662_));
 b15aoi013as1n02x5 _31302_ (.a(_05657_),
    .b(_05660_),
    .c(_04996_),
    .d(_05662_),
    .o1(_05663_));
 b15nor003ah1n06x5 _31303_ (.a(_05649_),
    .b(_05655_),
    .c(_05663_),
    .o1(_05664_));
 b15nandp3aq1n03x5 _31304_ (.a(_03067_),
    .b(_03057_),
    .c(_03285_),
    .o1(_05665_));
 b15oaoi13aq1n04x5 _31305_ (.a(net581),
    .b(_05665_),
    .c(_03187_),
    .d(_03046_),
    .o1(_05666_));
 b15nor003al1n03x5 _31306_ (.a(net572),
    .b(_03820_),
    .c(_03282_),
    .o1(_05667_));
 b15and002an1n04x5 _31307_ (.a(_03814_),
    .b(_03902_),
    .o(_05668_));
 b15aoai13as1n04x5 _31308_ (.a(net577),
    .b(_05667_),
    .c(_05668_),
    .d(net588),
    .o1(_05670_));
 b15oai012ar1n08x5 _31309_ (.a(_04575_),
    .b(_03217_),
    .c(net569),
    .o1(_05671_));
 b15and003ar1n02x5 _31310_ (.a(_03097_),
    .b(_03204_),
    .c(_05671_),
    .o(_05672_));
 b15aoi112ar1n08x5 _31311_ (.a(_03167_),
    .b(_03964_),
    .c(_03775_),
    .d(net587),
    .o1(_05673_));
 b15nandp2al1n02x5 _31312_ (.a(net591),
    .b(_03219_),
    .o1(_05674_));
 b15aoai13ah1n04x5 _31313_ (.a(_03281_),
    .b(_05672_),
    .c(_05673_),
    .d(_05674_),
    .o1(_05675_));
 b15norp02an1n02x5 _31314_ (.a(_03896_),
    .b(_03827_),
    .o1(_05676_));
 b15aoi022as1n06x5 _31315_ (.a(_03836_),
    .b(_05668_),
    .c(_05676_),
    .d(_03831_),
    .o1(_05677_));
 b15oai112as1n16x5 _31316_ (.a(_05670_),
    .b(_05675_),
    .c(net577),
    .d(_05677_),
    .o1(_05678_));
 b15nano23ar1n12x5 _31317_ (.a(_05633_),
    .b(_05664_),
    .c(_05666_),
    .d(_05678_),
    .out0(_05679_));
 b15xor002an1n02x5 _31318_ (.a(_05361_),
    .b(net395),
    .out0(_05681_));
 b15xor003aq1n03x5 _31319_ (.a(_05544_),
    .b(_05608_),
    .c(_05681_),
    .out0(_05682_));
 b15norp02ar1n02x5 _31320_ (.a(net542),
    .b(_05682_),
    .o1(_05683_));
 b15inv040ah1n02x5 _31321_ (.a(\text_in_r[71] ),
    .o1(_05684_));
 b15aoi012aq1n02x5 _31322_ (.a(_05683_),
    .b(_05684_),
    .c(net542),
    .o1(_05685_));
 b15xor002al1n04x5 _31323_ (.a(\u0.w[1][7] ),
    .b(_05685_),
    .out0(_00112_));
 b15inv020ah1n12x5 _31324_ (.a(\text_in_r[72] ),
    .o1(_05686_));
 b15xnr002as1n16x5 _31325_ (.a(_03034_),
    .b(net395),
    .out0(_05687_));
 b15xor002aq1n03x5 _31326_ (.a(_02772_),
    .b(_05687_),
    .out0(_05688_));
 b15xor002ah1n03x5 _31327_ (.a(_03544_),
    .b(_05688_),
    .out0(_05689_));
 b15mdn022an1n12x5 _31328_ (.a(_05686_),
    .b(_05689_),
    .o1(_05691_),
    .sa(net538));
 b15xor002al1n12x5 _31329_ (.a(\u0.w[1][8] ),
    .b(_05691_),
    .out0(_00073_));
 b15xnr002an1n16x5 _31330_ (.a(net400),
    .b(net395),
    .out0(_05692_));
 b15xor002ar1n02x5 _31331_ (.a(_04319_),
    .b(_05692_),
    .out0(_05693_));
 b15xor002ar1n02x5 _31332_ (.a(_03771_),
    .b(_05693_),
    .out0(_05694_));
 b15cmbn22ar1n02x5 _31333_ (.clk1(\text_in_r[73] ),
    .clk2(_05694_),
    .clkout(_05695_),
    .s(net537));
 b15xor002ar1n02x5 _31334_ (.a(\u0.w[1][9] ),
    .b(_05695_),
    .out0(_00074_));
 b15xor002as1n08x5 _31335_ (.a(net393),
    .b(_04319_),
    .out0(_05696_));
 b15xor002al1n02x5 _31336_ (.a(_04218_),
    .b(_04554_),
    .out0(_05697_));
 b15xor002ar1n02x5 _31337_ (.a(_05696_),
    .b(_05697_),
    .out0(_05698_));
 b15cmbn22aq1n02x5 _31338_ (.clk1(\text_in_r[74] ),
    .clk2(_05698_),
    .clkout(_05700_),
    .s(net536));
 b15qgbxo2an1n05x5 _31339_ (.a(\u0.w[1][10] ),
    .b(_05700_),
    .out0(_00075_));
 b15nand02ar1n02x5 _31340_ (.a(net537),
    .b(\text_in_r[75] ),
    .o1(_05701_));
 b15qgbxo2an1n05x5 _31341_ (.a(_04878_),
    .b(net395),
    .out0(_05702_));
 b15xor002as1n06x5 _31342_ (.a(net392),
    .b(_05702_),
    .out0(_05703_));
 b15xnr002ar1n02x5 _31343_ (.a(_04556_),
    .b(_05703_),
    .out0(_05704_));
 b15oai012ar1n02x5 _31344_ (.a(_05701_),
    .b(_05704_),
    .c(net537),
    .o1(_05705_));
 b15xor002al1n02x5 _31345_ (.a(\u0.w[1][11] ),
    .b(_05705_),
    .out0(_00076_));
 b15xor002al1n02x5 _31346_ (.a(_04956_),
    .b(_05687_),
    .out0(_05706_));
 b15xnr002ar1n02x5 _31347_ (.a(_04721_),
    .b(_05164_),
    .out0(_05707_));
 b15xor002al1n02x5 _31348_ (.a(net397),
    .b(_05707_),
    .out0(_05709_));
 b15xor002ar1n02x5 _31349_ (.a(_05706_),
    .b(_05709_),
    .out0(_05710_));
 b15ztpn00an1n08x5 TAP_412 ();
 b15cmbn22ar1n02x5 _31351_ (.clk1(\text_in_r[76] ),
    .clk2(_05710_),
    .clkout(_05712_),
    .s(ld_r));
 b15xor002al1n02x5 _31352_ (.a(\u0.w[1][12] ),
    .b(_05712_),
    .out0(_00077_));
 b15xor003aq1n06x5 _31353_ (.a(_04800_),
    .b(_05102_),
    .c(_05164_),
    .out0(_05713_));
 b15xor002ar1n02x5 _31354_ (.a(_05486_),
    .b(_05713_),
    .out0(_05714_));
 b15norp02ar1n02x5 _31355_ (.a(net542),
    .b(_05714_),
    .o1(_05715_));
 b15inv040ah1n02x5 _31356_ (.a(\text_in_r[77] ),
    .o1(_05716_));
 b15aoi012ar1n02x5 _31357_ (.a(_05715_),
    .b(_05716_),
    .c(net542),
    .o1(_05717_));
 b15xor002an1n02x5 _31358_ (.a(\u0.w[1][13] ),
    .b(_05717_),
    .out0(_00078_));
 b15xor003an1n02x5 _31359_ (.a(_05030_),
    .b(_05485_),
    .c(_05544_),
    .out0(_05719_));
 b15xor002ar1n02x5 _31360_ (.a(_05419_),
    .b(_05719_),
    .out0(_05720_));
 b15norp02ar1n02x5 _31361_ (.a(net542),
    .b(_05720_),
    .o1(_05721_));
 b15inv040ah1n02x5 _31362_ (.a(\text_in_r[78] ),
    .o1(_05722_));
 b15aoi012ar1n02x5 _31363_ (.a(_05721_),
    .b(_05722_),
    .c(net542),
    .o1(_05723_));
 b15xor002ar1n02x5 _31364_ (.a(\u0.w[1][14] ),
    .b(_05723_),
    .out0(_00079_));
 b15inv000ah1n04x5 _31365_ (.a(\text_in_r[79] ),
    .o1(_05724_));
 b15xor002an1n16x5 _31366_ (.a(_05300_),
    .b(_05544_),
    .out0(_05725_));
 b15xor002an1n06x5 _31367_ (.a(_03034_),
    .b(_05608_),
    .out0(_05726_));
 b15xor002ar1n08x5 _31368_ (.a(_05725_),
    .b(_05726_),
    .out0(_05728_));
 b15mdn022al1n03x5 _31369_ (.a(_05724_),
    .b(_05728_),
    .o1(_05729_),
    .sa(net541));
 b15xor002ar1n03x5 _31370_ (.a(\u0.w[1][15] ),
    .b(_05729_),
    .out0(_00080_));
 b15inv020as1n05x5 _31371_ (.a(\text_in_r[80] ),
    .o1(_05730_));
 b15xor002an1n16x5 _31372_ (.a(net396),
    .b(_05692_),
    .out0(_05731_));
 b15xor002as1n06x5 _31373_ (.a(_02771_),
    .b(_03544_),
    .out0(_05732_));
 b15xor002as1n12x5 _31374_ (.a(_05731_),
    .b(_05732_),
    .out0(_05733_));
 b15mdn022al1n16x5 _31375_ (.a(_05730_),
    .b(_05733_),
    .o1(_05734_),
    .sa(net536));
 b15xor002ah1n16x5 _31376_ (.a(\u0.w[1][16] ),
    .b(_05734_),
    .out0(_00041_));
 b15inv020as1n05x5 _31377_ (.a(\text_in_r[81] ),
    .o1(_05735_));
 b15qgbxo2an1n05x5 _31378_ (.a(net401),
    .b(_03633_),
    .out0(_05737_));
 b15xor003as1n08x5 _31379_ (.a(_05696_),
    .b(_05731_),
    .c(_05737_),
    .out0(_05738_));
 b15mdn022al1n16x5 _31380_ (.a(_05735_),
    .b(_05738_),
    .o1(_05739_),
    .sa(net536));
 b15xor002ah1n16x5 _31381_ (.a(\u0.w[1][17] ),
    .b(_05739_),
    .out0(_00042_));
 b15inv000ah1n04x5 _31382_ (.a(\text_in_r[82] ),
    .o1(_05740_));
 b15xor002al1n16x5 _31383_ (.a(_03769_),
    .b(_04554_),
    .out0(_05741_));
 b15xor002al1n12x5 _31384_ (.a(net392),
    .b(_05741_),
    .out0(_05742_));
 b15xor002as1n06x5 _31385_ (.a(net393),
    .b(_04217_),
    .out0(_05743_));
 b15xor002aq1n16x5 _31386_ (.a(_05742_),
    .b(_05743_),
    .out0(_05744_));
 b15mdn022al1n12x5 _31387_ (.a(_05740_),
    .b(_05744_),
    .o1(_05745_),
    .sa(net536));
 b15xor002as1n12x5 _31388_ (.a(\u0.w[1][18] ),
    .b(_05745_),
    .out0(_00043_));
 b15xor002an1n04x5 _31389_ (.a(_04478_),
    .b(net397),
    .out0(_05747_));
 b15qgbxo2an1n05x5 _31390_ (.a(net399),
    .b(net396),
    .out0(_05748_));
 b15xor002al1n06x5 _31391_ (.a(_05747_),
    .b(_05748_),
    .out0(_05749_));
 b15xor002aq1n08x5 _31392_ (.a(_05703_),
    .b(_05749_),
    .out0(_05750_));
 b15cmbn22al1n08x5 _31393_ (.clk1(\text_in_r[83] ),
    .clk2(_05750_),
    .clkout(_05751_),
    .s(net536));
 b15xor002as1n16x5 _31394_ (.a(\u0.w[1][19] ),
    .b(_05751_),
    .out0(_00044_));
 b15inv000as1n16x5 _31395_ (.a(\text_in_r[84] ),
    .o1(_05752_));
 b15xnr002al1n03x5 _31396_ (.a(_05164_),
    .b(net396),
    .out0(_05753_));
 b15xor002as1n03x5 _31397_ (.a(net398),
    .b(_05753_),
    .out0(_05754_));
 b15xor002ar1n03x5 _31398_ (.a(_04800_),
    .b(_04955_),
    .out0(_05756_));
 b15xor002ar1n02x5 _31399_ (.a(net397),
    .b(net395),
    .out0(_05757_));
 b15xor002an1n02x5 _31400_ (.a(_05756_),
    .b(_05757_),
    .out0(_05758_));
 b15xor002aq1n03x5 _31401_ (.a(_05754_),
    .b(_05758_),
    .out0(_05759_));
 b15mdn022ah1n03x5 _31402_ (.a(_05752_),
    .b(_05759_),
    .o1(_05760_),
    .sa(ld_r));
 b15xor002aq1n06x5 _31403_ (.a(\u0.w[1][20] ),
    .b(_05760_),
    .out0(_00045_));
 b15xor002al1n02x5 _31404_ (.a(_04801_),
    .b(_05030_),
    .out0(_05761_));
 b15xor002ar1n03x5 _31405_ (.a(_05486_),
    .b(_05761_),
    .out0(_05762_));
 b15cmbn22ar1n08x5 _31406_ (.clk1(\text_in_r[85] ),
    .clk2(_05762_),
    .clkout(_05763_),
    .s(net541));
 b15xor002aq1n16x5 _31407_ (.a(\u0.w[1][21] ),
    .b(_05763_),
    .out0(_00046_));
 b15inv020as1n05x5 _31408_ (.a(\text_in_r[86] ),
    .o1(_05765_));
 b15xor002as1n03x5 _31409_ (.a(_05103_),
    .b(_05361_),
    .out0(_05766_));
 b15xor002ah1n06x5 _31410_ (.a(_05725_),
    .b(_05766_),
    .out0(_05767_));
 b15mdn022al1n12x5 _31411_ (.a(_05765_),
    .b(_05767_),
    .o1(_05768_),
    .sa(net541));
 b15xor002aq1n16x5 _31412_ (.a(\u0.w[1][22] ),
    .b(_05768_),
    .out0(_00047_));
 b15xor003as1n08x5 _31413_ (.a(_03413_),
    .b(_05300_),
    .c(_05418_),
    .out0(_05769_));
 b15xor002as1n12x5 _31414_ (.a(_05687_),
    .b(_05769_),
    .out0(_05770_));
 b15nor002an1n06x5 _31415_ (.a(ld_r),
    .b(_05770_),
    .o1(_05771_));
 b15inv020aq1n16x5 _31416_ (.a(\text_in_r[87] ),
    .o1(_05772_));
 b15aoi012as1n16x5 _31417_ (.a(_05771_),
    .b(_05772_),
    .c(ld_r),
    .o1(_05773_));
 b15xor002as1n12x5 _31418_ (.a(\u0.w[1][23] ),
    .b(_05773_),
    .out0(_00048_));
 b15inv020ar1n32x5 _31419_ (.a(\text_in_r[88] ),
    .o1(_05775_));
 b15xor002ah1n04x5 _31420_ (.a(_03544_),
    .b(_05608_),
    .out0(_05776_));
 b15xor002ar1n12x5 _31421_ (.a(net401),
    .b(net400),
    .out0(_05777_));
 b15xor002ar1n12x5 _31422_ (.a(_05776_),
    .b(_05777_),
    .out0(_05778_));
 b15mdn022al1n12x5 _31423_ (.a(_05775_),
    .b(_05778_),
    .o1(_05779_),
    .sa(net537));
 b15xor002ah1n12x5 _31424_ (.a(\u0.w[1][24] ),
    .b(_05779_),
    .out0(_00009_));
 b15xor003an1n04x5 _31425_ (.a(_02772_),
    .b(_03769_),
    .c(_05608_),
    .out0(_05780_));
 b15xor002ar1n04x5 _31426_ (.a(_05696_),
    .b(_05780_),
    .out0(_05781_));
 b15cmbn22ar1n02x5 _31427_ (.clk1(\text_in_r[89] ),
    .clk2(_05781_),
    .clkout(_05782_),
    .s(net536));
 b15xor002ar1n02x5 _31428_ (.a(\u0.w[1][25] ),
    .b(_05782_),
    .out0(_00010_));
 b15xor002al1n03x5 _31429_ (.a(_03633_),
    .b(net399),
    .out0(_05784_));
 b15xor003al1n04x5 _31430_ (.a(net392),
    .b(_05741_),
    .c(_05784_),
    .out0(_05785_));
 b15norp02ar1n02x5 _31431_ (.a(net537),
    .b(_05785_),
    .o1(_05786_));
 b15inv000ar1n24x5 _31432_ (.a(\text_in_r[90] ),
    .o1(_05787_));
 b15aoi012ar1n02x5 _31433_ (.a(_05786_),
    .b(_05787_),
    .c(net537),
    .o1(_05788_));
 b15xor002al1n02x5 _31434_ (.a(\u0.w[1][26] ),
    .b(_05788_),
    .out0(_00011_));
 b15inv040ah1n02x5 _31435_ (.a(\text_in_r[91] ),
    .o1(_05789_));
 b15xor002ah1n03x5 _31436_ (.a(net397),
    .b(_04878_),
    .out0(_05790_));
 b15xor003an1n02x5 _31437_ (.a(net398),
    .b(_05608_),
    .c(_05790_),
    .out0(_05791_));
 b15xor002al1n02x5 _31438_ (.a(_04218_),
    .b(_05791_),
    .out0(_05793_));
 b15ztpn00an1n08x5 TAP_411 ();
 b15mdn022al1n02x5 _31440_ (.a(_05789_),
    .b(_05793_),
    .o1(_05795_),
    .sa(net537));
 b15xor002ar1n02x5 _31441_ (.a(\u0.w[1][27] ),
    .b(_05795_),
    .out0(_00012_));
 b15nand02ar1n02x5 _31442_ (.a(net541),
    .b(\text_in_r[92] ),
    .o1(_05796_));
 b15xor002ar1n02x5 _31443_ (.a(_04803_),
    .b(_05754_),
    .out0(_05797_));
 b15oai012ar1n02x5 _31444_ (.a(_05796_),
    .b(_05797_),
    .c(net541),
    .o1(_05798_));
 b15xor002ar1n02x5 _31445_ (.a(\u0.w[1][28] ),
    .b(_05798_),
    .out0(_00013_));
 b15inv040ah1n02x5 _31446_ (.a(\text_in_r[93] ),
    .o1(_05799_));
 b15xor002ar1n02x5 _31447_ (.a(_04721_),
    .b(_05485_),
    .out0(_05800_));
 b15xor002al1n02x5 _31448_ (.a(_05104_),
    .b(_05800_),
    .out0(_05802_));
 b15mdn022al1n02x5 _31449_ (.a(_05799_),
    .b(_05802_),
    .o1(_05803_),
    .sa(net541));
 b15xor002ar1n02x5 _31450_ (.a(\u0.w[1][29] ),
    .b(_05803_),
    .out0(_00014_));
 b15xor003ar1n03x5 _31451_ (.a(_05102_),
    .b(_05229_),
    .c(_05418_),
    .out0(_05804_));
 b15xor002ar1n02x5 _31452_ (.a(_05725_),
    .b(_05804_),
    .out0(_05805_));
 b15norp02ar1n02x5 _31453_ (.a(net541),
    .b(_05805_),
    .o1(_05806_));
 b15inv040ah1n02x5 _31454_ (.a(\text_in_r[94] ),
    .o1(_05807_));
 b15aoi012ar1n02x5 _31455_ (.a(_05806_),
    .b(_05807_),
    .c(net541),
    .o1(_05808_));
 b15xor002an1n02x5 _31456_ (.a(\u0.w[1][30] ),
    .b(_05808_),
    .out0(_00015_));
 b15xor003ar1n02x5 _31457_ (.a(_05419_),
    .b(net396),
    .c(_05687_),
    .out0(_05809_));
 b15norp02ar1n02x5 _31458_ (.a(ld_r),
    .b(_05809_),
    .o1(_05811_));
 b15inv020ah1n05x5 _31459_ (.a(\text_in_r[95] ),
    .o1(_05812_));
 b15aoi012ar1n02x5 _31460_ (.a(_05811_),
    .b(_05812_),
    .c(ld_r),
    .o1(_05813_));
 b15xor002ar1n02x5 _31461_ (.a(\u0.w[1][31] ),
    .b(_05813_),
    .out0(_00016_));
 b15inv000aq1n06x5 _31462_ (.a(\text_in_r[96] ),
    .o1(_05814_));
 b15ztpn00an1n08x5 TAP_410 ();
 b15ztpn00an1n08x5 TAP_409 ();
 b15ztpn00an1n08x5 TAP_408 ();
 b15ztpn00an1n08x5 TAP_407 ();
 b15ztpn00an1n08x5 TAP_406 ();
 b15inv000as1n48x5 _31468_ (.a(\us00.a[1] ),
    .o1(_05821_));
 b15ztpn00an1n08x5 TAP_405 ();
 b15ztpn00an1n08x5 TAP_404 ();
 b15ztpn00an1n08x5 TAP_403 ();
 b15ztpn00an1n08x5 TAP_402 ();
 b15ztpn00an1n08x5 TAP_401 ();
 b15andc04as1n16x5 _31474_ (.a(net920),
    .b(net923),
    .c(net916),
    .d(net918),
    .o(_05827_));
 b15ztpn00an1n08x5 TAP_400 ();
 b15nonb02as1n16x5 _31476_ (.a(net926),
    .b(net929),
    .out0(_05829_));
 b15ztpn00an1n08x5 TAP_399 ();
 b15nand03al1n02x5 _31478_ (.a(_05821_),
    .b(_05827_),
    .c(_05829_),
    .o1(_05832_));
 b15ztpn00an1n08x5 TAP_398 ();
 b15ztpn00an1n08x5 TAP_397 ();
 b15nanb02as1n24x5 _31481_ (.a(net926),
    .b(net929),
    .out0(_05835_));
 b15ztpn00an1n08x5 TAP_396 ();
 b15ztpn00an1n08x5 TAP_395 ();
 b15ztpn00an1n08x5 TAP_394 ();
 b15nonb02as1n16x5 _31485_ (.a(net915),
    .b(net918),
    .out0(_05839_));
 b15and002al1n32x5 _31486_ (.a(net920),
    .b(net923),
    .o(_05840_));
 b15nandp2aq1n24x5 _31487_ (.a(_05839_),
    .b(_05840_),
    .o1(_05841_));
 b15oai012ar1n06x5 _31488_ (.a(_05832_),
    .b(_05835_),
    .c(_05841_),
    .o1(_05843_));
 b15and002al1n32x5 _31489_ (.a(net916),
    .b(net918),
    .o(_05844_));
 b15ztpn00an1n08x5 TAP_393 ();
 b15nanb02as1n24x5 _31491_ (.a(net927),
    .b(net924),
    .out0(_05846_));
 b15ztpn00an1n08x5 TAP_392 ();
 b15nandp3ar1n02x5 _31493_ (.a(_05835_),
    .b(_05844_),
    .c(_05846_),
    .o1(_05848_));
 b15ztpn00an1n08x5 TAP_391 ();
 b15ztpn00an1n08x5 TAP_390 ();
 b15nand02as1n48x5 _31496_ (.a(net929),
    .b(net926),
    .o1(_05851_));
 b15ztpn00an1n08x5 PHY_389 ();
 b15orn002as1n32x5 _31498_ (.a(net914),
    .b(net917),
    .o(_05854_));
 b15ztpn00an1n08x5 PHY_388 ();
 b15oai012an1n04x5 _31500_ (.a(_05848_),
    .b(_05851_),
    .c(_05854_),
    .o1(_05856_));
 b15ztpn00an1n08x5 PHY_387 ();
 b15ztpn00an1n08x5 PHY_386 ();
 b15ztpn00an1n08x5 PHY_385 ();
 b15nano22ah1n05x5 _31504_ (.a(net920),
    .b(net923),
    .c(net935),
    .out0(_05860_));
 b15aoi022as1n08x5 _31505_ (.a(net935),
    .b(_05843_),
    .c(_05856_),
    .d(_05860_),
    .o1(_05861_));
 b15ztpn00an1n08x5 PHY_384 ();
 b15ztpn00an1n08x5 PHY_383 ();
 b15ztpn00an1n08x5 PHY_382 ();
 b15ztpn00an1n08x5 PHY_381 ();
 b15nonb02as1n16x5 _31510_ (.a(net919),
    .b(net922),
    .out0(_05867_));
 b15ztpn00an1n08x5 PHY_380 ();
 b15ztpn00an1n08x5 PHY_379 ();
 b15nonb02an1n16x5 _31513_ (.a(net916),
    .b(net935),
    .out0(_05870_));
 b15ztpn00an1n08x5 PHY_378 ();
 b15ztpn00an1n08x5 PHY_377 ();
 b15ztpn00an1n08x5 PHY_376 ();
 b15ztpn00an1n08x5 PHY_375 ();
 b15ztpn00an1n08x5 PHY_374 ();
 b15ztpn00an1n08x5 PHY_373 ();
 b15ztpn00an1n08x5 PHY_372 ();
 b15ztpn00an1n08x5 PHY_371 ();
 b15nand03as1n03x5 _31522_ (.a(net917),
    .b(net931),
    .c(net928),
    .o1(_05880_));
 b15nand04ar1n12x5 _31523_ (.a(net925),
    .b(_05867_),
    .c(_05870_),
    .d(_05880_),
    .o1(_05881_));
 b15nandp2ah1n24x5 _31524_ (.a(\us00.a[0] ),
    .b(net932),
    .o1(_05882_));
 b15nanb02as1n24x5 _31525_ (.a(\us00.a[5] ),
    .b(net921),
    .out0(_05883_));
 b15orn002aq1n24x5 _31526_ (.a(net928),
    .b(net925),
    .o(_05884_));
 b15nor003as1n12x5 _31527_ (.a(_05883_),
    .b(_05854_),
    .c(_05884_),
    .o1(_05885_));
 b15nandp2ar1n05x5 _31528_ (.a(_05882_),
    .b(_05885_),
    .o1(_05887_));
 b15ztpn00an1n08x5 PHY_370 ();
 b15ztpn00an1n08x5 PHY_369 ();
 b15ztpn00an1n08x5 PHY_368 ();
 b15nona23ah1n32x5 _31532_ (.a(net914),
    .b(\us00.a[6] ),
    .c(\us00.a[5] ),
    .d(net921),
    .out0(_05891_));
 b15ztpn00an1n08x5 PHY_367 ();
 b15nand02an1n12x5 _31534_ (.a(net931),
    .b(_05829_),
    .o1(_05893_));
 b15orn002al1n32x5 _31535_ (.a(\us00.a[0] ),
    .b(net930),
    .o(_05894_));
 b15and002ah1n16x5 _31536_ (.a(net928),
    .b(net925),
    .o(_05895_));
 b15nandp2as1n05x5 _31537_ (.a(_05894_),
    .b(_05895_),
    .o1(_05896_));
 b15nonb02as1n16x5 _31538_ (.a(net918),
    .b(net916),
    .out0(_05898_));
 b15nandp2as1n32x5 _31539_ (.a(_05898_),
    .b(_05840_),
    .o1(_05899_));
 b15oai022ar1n04x5 _31540_ (.a(_05891_),
    .b(_05893_),
    .c(_05896_),
    .d(_05899_),
    .o1(_05900_));
 b15ztpn00an1n08x5 PHY_366 ();
 b15ztpn00an1n08x5 PHY_365 ();
 b15nanb02aq1n06x5 _31543_ (.a(net922),
    .b(net915),
    .out0(_05903_));
 b15nand02ah1n12x5 _31544_ (.a(net917),
    .b(net932),
    .o1(_05904_));
 b15norp02aq1n08x5 _31545_ (.a(_05903_),
    .b(_05904_),
    .o1(_05905_));
 b15nonb02as1n16x5 _31546_ (.a(net929),
    .b(\us00.a[3] ),
    .out0(_05906_));
 b15ztpn00an1n08x5 PHY_364 ();
 b15aoi012al1n04x5 _31548_ (.a(_05900_),
    .b(_05905_),
    .c(_05906_),
    .o1(_05909_));
 b15nand04aq1n16x5 _31549_ (.a(_05861_),
    .b(_05881_),
    .c(_05887_),
    .d(_05909_),
    .o1(_05910_));
 b15inv020ah1n64x5 _31550_ (.a(net924),
    .o1(_05911_));
 b15ztpn00an1n08x5 PHY_363 ();
 b15ztpn00an1n08x5 PHY_362 ();
 b15ztpn00an1n08x5 PHY_361 ();
 b15nano23as1n24x5 _31554_ (.a(net920),
    .b(net918),
    .c(net916),
    .d(net923),
    .out0(_05915_));
 b15ztpn00an1n08x5 PHY_360 ();
 b15and002al1n16x5 _31556_ (.a(net933),
    .b(net930),
    .o(_05917_));
 b15inv000ah1n48x5 _31557_ (.a(net927),
    .o1(_05918_));
 b15oai012ar1n02x5 _31558_ (.a(_05915_),
    .b(_05917_),
    .c(_05918_),
    .o1(_05920_));
 b15nand04as1n16x5 _31559_ (.a(\us00.a[5] ),
    .b(net921),
    .c(net914),
    .d(net917),
    .o1(_05921_));
 b15ztpn00an1n08x5 PHY_359 ();
 b15oai012ar1n02x5 _31561_ (.a(_05920_),
    .b(_05921_),
    .c(net930),
    .o1(_05923_));
 b15nanb03as1n03x5 _31562_ (.a(net930),
    .b(net927),
    .c(net933),
    .out0(_05924_));
 b15nanb02as1n24x5 _31563_ (.a(\us00.a[0] ),
    .b(net932),
    .out0(_05925_));
 b15ztpn00an1n08x5 PHY_358 ();
 b15oaoi13as1n08x5 _31565_ (.a(net924),
    .b(_05924_),
    .c(_05925_),
    .d(net927),
    .o1(_05927_));
 b15nanb02as1n24x5 _31566_ (.a(net921),
    .b(net919),
    .out0(_05928_));
 b15nandp2an1n48x5 _31567_ (.a(net914),
    .b(net917),
    .o1(_05929_));
 b15ztpn00an1n08x5 PHY_357 ();
 b15norp02ar1n48x5 _31569_ (.a(_05928_),
    .b(_05929_),
    .o1(_05932_));
 b15aoi022an1n04x5 _31570_ (.a(_05911_),
    .b(_05923_),
    .c(_05927_),
    .d(_05932_),
    .o1(_05933_));
 b15nanb02as1n24x5 _31571_ (.a(net914),
    .b(\us00.a[6] ),
    .out0(_05934_));
 b15nandp2ah1n48x5 _31572_ (.a(net919),
    .b(net921),
    .o1(_05935_));
 b15ztpn00an1n08x5 PHY_356 ();
 b15qgbno2an1n10x5 _31574_ (.a(_05934_),
    .b(_05935_),
    .o1(_05937_));
 b15ztpn00an1n08x5 PHY_355 ();
 b15oai022ar1n02x5 _31576_ (.a(net931),
    .b(_05835_),
    .c(_05846_),
    .d(net934),
    .o1(_05939_));
 b15ztpn00an1n08x5 PHY_354 ();
 b15oai012an1n08x5 _31578_ (.a(net924),
    .b(net927),
    .c(net930),
    .o1(_05942_));
 b15ztpn00an1n08x5 PHY_353 ();
 b15ztpn00an1n08x5 PHY_352 ();
 b15aoai13aq1n04x5 _31581_ (.a(_05937_),
    .b(_05939_),
    .c(_05942_),
    .d(net934),
    .o1(_05945_));
 b15inv000as1n08x5 _31582_ (.a(net914),
    .o1(_05946_));
 b15nor002ah1n32x5 _31583_ (.a(net929),
    .b(\us00.a[3] ),
    .o1(_05947_));
 b15ztpn00an1n08x5 PHY_351 ();
 b15nand02al1n04x5 _31585_ (.a(_05946_),
    .b(_05947_),
    .o1(_05949_));
 b15ztpn00an1n08x5 PHY_350 ();
 b15ztpn00an1n08x5 PHY_349 ();
 b15norp03ar1n02x5 _31588_ (.a(\us00.a[6] ),
    .b(_05928_),
    .c(_05917_),
    .o1(_05953_));
 b15nonb02as1n16x5 _31589_ (.a(net933),
    .b(net930),
    .out0(_05954_));
 b15nonb02as1n16x5 _31590_ (.a(net923),
    .b(net920),
    .out0(_05955_));
 b15ztpn00an1n08x5 PHY_348 ();
 b15aoi013an1n03x5 _31592_ (.a(_05953_),
    .b(_05954_),
    .c(_05955_),
    .d(\us00.a[6] ),
    .o1(_05957_));
 b15oai112al1n12x5 _31593_ (.a(_05933_),
    .b(_05945_),
    .c(_05949_),
    .d(_05957_),
    .o1(_05958_));
 b15nona23as1n32x5 _31594_ (.a(net919),
    .b(net914),
    .c(net917),
    .d(net921),
    .out0(_05959_));
 b15ztpn00an1n08x5 PHY_347 ();
 b15ztpn00an1n08x5 PHY_346 ();
 b15oai112al1n02x5 _31597_ (.a(net933),
    .b(_05891_),
    .c(_05959_),
    .d(net930),
    .o1(_05962_));
 b15nor002aq1n08x5 _31598_ (.a(_05821_),
    .b(_05959_),
    .o1(_05964_));
 b15oai112ah1n04x5 _31599_ (.a(_05906_),
    .b(_05962_),
    .c(_05964_),
    .d(net933),
    .o1(_05965_));
 b15orn002aq1n32x5 _31600_ (.a(net919),
    .b(net921),
    .o(_05966_));
 b15nanb02as1n24x5 _31601_ (.a(net917),
    .b(net915),
    .out0(_05967_));
 b15norp02as1n12x5 _31602_ (.a(_05966_),
    .b(_05967_),
    .o1(_05968_));
 b15inv000ah1n48x5 _31603_ (.a(net933),
    .o1(_05969_));
 b15ztpn00an1n08x5 PHY_345 ();
 b15nor002ah1n04x5 _31605_ (.a(_05969_),
    .b(_05835_),
    .o1(_05971_));
 b15nona23as1n32x5 _31606_ (.a(net921),
    .b(\us00.a[6] ),
    .c(net914),
    .d(\us00.a[5] ),
    .out0(_05972_));
 b15ztpn00an1n08x5 PHY_344 ();
 b15norp02as1n48x5 _31608_ (.a(net920),
    .b(net923),
    .o1(_05975_));
 b15ztpn00an1n08x5 PHY_343 ();
 b15nand03as1n08x5 _31610_ (.a(_05918_),
    .b(_05975_),
    .c(_05839_),
    .o1(_05977_));
 b15nandp2ar1n03x5 _31611_ (.a(_05972_),
    .b(_05977_),
    .o1(_05978_));
 b15ztpn00an1n08x5 PHY_342 ();
 b15aoi022al1n02x5 _31613_ (.a(_05968_),
    .b(_05971_),
    .c(_05978_),
    .d(net924),
    .o1(_05980_));
 b15ztpn00an1n08x5 PHY_341 ();
 b15oai012an1n06x5 _31615_ (.a(_05965_),
    .b(_05980_),
    .c(net930),
    .o1(_05982_));
 b15norp02an1n16x5 _31616_ (.a(_05934_),
    .b(_05966_),
    .o1(_05983_));
 b15nand02al1n12x5 _31617_ (.a(net934),
    .b(net928),
    .o1(_05984_));
 b15aoi012an1n02x5 _31618_ (.a(_05821_),
    .b(_05846_),
    .c(_05984_),
    .o1(_05986_));
 b15orn003aq1n08x5 _31619_ (.a(net931),
    .b(net928),
    .c(net925),
    .o(_05987_));
 b15aoi012an1n02x5 _31620_ (.a(_05969_),
    .b(_05851_),
    .c(_05987_),
    .o1(_05988_));
 b15oai012ar1n08x5 _31621_ (.a(_05983_),
    .b(_05986_),
    .c(_05988_),
    .o1(_05989_));
 b15nandp2ah1n05x5 _31622_ (.a(\us00.a[1] ),
    .b(net927),
    .o1(_05990_));
 b15aoi012ar1n02x5 _31623_ (.a(_05969_),
    .b(_05990_),
    .c(_05884_),
    .o1(_05991_));
 b15nanb02ah1n04x5 _31624_ (.a(net926),
    .b(net932),
    .out0(_05992_));
 b15oai012an1n12x5 _31625_ (.a(_05992_),
    .b(_05894_),
    .c(_05911_),
    .o1(_05993_));
 b15ztpn00an1n08x5 PHY_340 ();
 b15aoi012ar1n02x5 _31627_ (.a(_05991_),
    .b(_05993_),
    .c(net927),
    .o1(_05995_));
 b15nona23as1n32x5 _31628_ (.a(net919),
    .b(net917),
    .c(net914),
    .d(net921),
    .out0(_05997_));
 b15oai012an1n02x5 _31629_ (.a(_05989_),
    .b(_05995_),
    .c(_05997_),
    .o1(_05998_));
 b15ztpn00an1n08x5 PHY_339 ();
 b15norp02aq1n16x5 _31631_ (.a(_05883_),
    .b(_05929_),
    .o1(_06000_));
 b15nandp3ar1n02x5 _31632_ (.a(_05969_),
    .b(net930),
    .c(_06000_),
    .o1(_06001_));
 b15oaoi13ar1n02x5 _31633_ (.a(net924),
    .b(_06001_),
    .c(_05841_),
    .d(net930),
    .o1(_06002_));
 b15norp02ah1n32x5 _31634_ (.a(net916),
    .b(net918),
    .o1(_06003_));
 b15ztpn00an1n08x5 PHY_338 ();
 b15nand04aq1n03x5 _31636_ (.a(net930),
    .b(_05867_),
    .c(_06003_),
    .d(_05906_),
    .o1(_06005_));
 b15nonb03as1n06x5 _31637_ (.a(net933),
    .b(net927),
    .c(net924),
    .out0(_06006_));
 b15ztpn00an1n08x5 PHY_337 ();
 b15nonb02as1n03x5 _31639_ (.a(\us00.a[4] ),
    .b(net914),
    .out0(_06009_));
 b15ztpn00an1n08x5 PHY_336 ();
 b15nano22ar1n02x5 _31641_ (.a(\us00.a[6] ),
    .b(net930),
    .c(net919),
    .out0(_06011_));
 b15nonb02aq1n12x5 _31642_ (.a(net920),
    .b(net918),
    .out0(_06012_));
 b15oai112ar1n04x5 _31643_ (.a(_06006_),
    .b(_06009_),
    .c(_06011_),
    .d(_06012_),
    .o1(_06013_));
 b15xnr002an1n08x5 _31644_ (.a(\us00.a[0] ),
    .b(\us00.a[1] ),
    .out0(_06014_));
 b15nand04ah1n02x5 _31645_ (.a(_05975_),
    .b(_05839_),
    .c(_05947_),
    .d(_06014_),
    .o1(_06015_));
 b15and003aq1n04x5 _31646_ (.a(_06005_),
    .b(_06013_),
    .c(_06015_),
    .o(_06016_));
 b15ztpn00an1n08x5 PHY_335 ();
 b15xnr002as1n16x5 _31648_ (.a(net930),
    .b(net928),
    .out0(_06019_));
 b15nonb02ar1n08x5 _31649_ (.a(\us00.a[6] ),
    .b(\us00.a[5] ),
    .out0(_06020_));
 b15nano22ar1n02x5 _31650_ (.a(net921),
    .b(net933),
    .c(net914),
    .out0(_06021_));
 b15nonb02ar1n02x5 _31651_ (.a(net914),
    .b(net921),
    .out0(_06022_));
 b15oai112ar1n02x5 _31652_ (.a(_06019_),
    .b(_06020_),
    .c(_06021_),
    .d(_06022_),
    .o1(_06023_));
 b15nano23ah1n24x5 _31653_ (.a(net914),
    .b(\us00.a[6] ),
    .c(\us00.a[5] ),
    .d(net921),
    .out0(_06024_));
 b15nonb03as1n02x5 _31654_ (.a(net930),
    .b(net927),
    .c(net933),
    .out0(_06025_));
 b15nano23as1n24x5 _31655_ (.a(net921),
    .b(net917),
    .c(net914),
    .d(\us00.a[5] ),
    .out0(_06026_));
 b15aoi022ar1n02x5 _31656_ (.a(_05954_),
    .b(_06024_),
    .c(_06025_),
    .d(_06026_),
    .o1(_06027_));
 b15nandp3aq1n02x5 _31657_ (.a(net924),
    .b(_06023_),
    .c(_06027_),
    .o1(_06028_));
 b15ztpn00an1n08x5 PHY_334 ();
 b15ztpn00an1n08x5 PHY_333 ();
 b15nor004as1n12x5 _31660_ (.a(\us00.a[5] ),
    .b(net921),
    .c(net914),
    .d(\us00.a[6] ),
    .o1(_06032_));
 b15nand02as1n12x5 _31661_ (.a(net927),
    .b(_06032_),
    .o1(_06033_));
 b15nona23aq1n32x5 _31662_ (.a(net919),
    .b(net921),
    .c(net914),
    .d(net917),
    .out0(_06034_));
 b15oaoi13al1n02x5 _31663_ (.a(_05894_),
    .b(_06033_),
    .c(_06034_),
    .d(net927),
    .o1(_06035_));
 b15ztpn00an1n08x5 PHY_332 ();
 b15ornc04as1n24x5 _31665_ (.a(net919),
    .b(net921),
    .c(net915),
    .d(net917),
    .o(_06037_));
 b15nandp3aq1n24x5 _31666_ (.a(net934),
    .b(net931),
    .c(net928),
    .o1(_06038_));
 b15oai012ar1n03x5 _31667_ (.a(_05911_),
    .b(_06037_),
    .c(_06038_),
    .o1(_06039_));
 b15oai012as1n04x5 _31668_ (.a(_06028_),
    .b(_06035_),
    .c(_06039_),
    .o1(_06041_));
 b15nona23aq1n04x5 _31669_ (.a(_05998_),
    .b(_06002_),
    .c(_06016_),
    .d(_06041_),
    .out0(_06042_));
 b15nor004ah1n08x5 _31670_ (.a(_05910_),
    .b(_05958_),
    .c(_05982_),
    .d(_06042_),
    .o1(_06043_));
 b15nanb02as1n24x5 _31671_ (.a(net931),
    .b(net934),
    .out0(_06044_));
 b15norp03ar1n02x5 _31672_ (.a(_05835_),
    .b(_06044_),
    .c(_06034_),
    .o1(_06045_));
 b15nano23as1n24x5 _31673_ (.a(\us00.a[4] ),
    .b(net914),
    .c(\us00.a[6] ),
    .d(\us00.a[5] ),
    .out0(_06046_));
 b15xor002ah1n04x5 _31674_ (.a(net934),
    .b(net931),
    .out0(_06047_));
 b15aoi013an1n03x5 _31675_ (.a(_06045_),
    .b(_05829_),
    .c(_06046_),
    .d(_06047_),
    .o1(_06048_));
 b15nor002ah1n04x5 _31676_ (.a(net931),
    .b(_05884_),
    .o1(_06049_));
 b15nand02aq1n24x5 _31677_ (.a(net931),
    .b(net925),
    .o1(_06050_));
 b15nor003aq1n06x5 _31678_ (.a(_05967_),
    .b(_05935_),
    .c(_06050_),
    .o1(_06052_));
 b15aoi022ah1n06x5 _31679_ (.a(_05932_),
    .b(_06049_),
    .c(_06052_),
    .d(_05984_),
    .o1(_06053_));
 b15nandp2ar1n12x5 _31680_ (.a(_06048_),
    .b(_06053_),
    .o1(_06054_));
 b15ztpn00an1n08x5 PHY_331 ();
 b15norp02an1n48x5 _31682_ (.a(\us00.a[0] ),
    .b(net932),
    .o1(_06056_));
 b15ztpn00an1n08x5 PHY_330 ();
 b15norp02ar1n02x5 _31684_ (.a(net927),
    .b(_05972_),
    .o1(_06058_));
 b15ztpn00an1n08x5 PHY_329 ();
 b15norp02al1n12x5 _31686_ (.a(_05883_),
    .b(_05854_),
    .o1(_06060_));
 b15ztpn00an1n08x5 PHY_328 ();
 b15aoai13ar1n03x5 _31688_ (.a(_06056_),
    .b(_06058_),
    .c(_06060_),
    .d(net927),
    .o1(_06063_));
 b15nand03aq1n02x5 _31689_ (.a(net927),
    .b(_06060_),
    .c(_05917_),
    .o1(_06064_));
 b15aoi012al1n04x5 _31690_ (.a(net924),
    .b(_06063_),
    .c(_06064_),
    .o1(_06065_));
 b15norp02aq1n04x5 _31691_ (.a(_06054_),
    .b(_06065_),
    .o1(_06066_));
 b15nandp2as1n08x5 _31692_ (.a(_05955_),
    .b(_05844_),
    .o1(_06067_));
 b15norp02ar1n02x5 _31693_ (.a(net930),
    .b(_06067_),
    .o1(_06068_));
 b15ztpn00an1n08x5 PHY_327 ();
 b15oai112al1n02x5 _31695_ (.a(net927),
    .b(_05882_),
    .c(_06068_),
    .d(_06032_),
    .o1(_06070_));
 b15ztpn00an1n08x5 PHY_326 ();
 b15and002al1n32x5 _31697_ (.a(net932),
    .b(net929),
    .o(_06072_));
 b15oaoi13ar1n02x5 _31698_ (.a(_05854_),
    .b(_05883_),
    .c(_05928_),
    .d(_06072_),
    .o1(_06074_));
 b15nor003ar1n06x5 _31699_ (.a(net930),
    .b(_05883_),
    .c(_05854_),
    .o1(_06075_));
 b15nonb02al1n16x5 _31700_ (.a(net930),
    .b(net927),
    .out0(_06076_));
 b15oai013ar1n02x5 _31701_ (.a(_06074_),
    .b(_06075_),
    .c(_06076_),
    .d(net933),
    .o1(_06077_));
 b15nona23as1n32x5 _31702_ (.a(net921),
    .b(net915),
    .c(net917),
    .d(net919),
    .out0(_06078_));
 b15oai112an1n04x5 _31703_ (.a(_06070_),
    .b(_06077_),
    .c(_05990_),
    .d(_06078_),
    .o1(_06079_));
 b15ztpn00an1n08x5 PHY_325 ();
 b15norp02ah1n12x5 _31705_ (.a(net932),
    .b(net929),
    .o1(_06081_));
 b15nandp2al1n03x5 _31706_ (.a(_06081_),
    .b(_05915_),
    .o1(_06082_));
 b15ztpn00an1n08x5 PHY_324 ();
 b15oai012ar1n02x5 _31708_ (.a(net930),
    .b(_06000_),
    .c(_05932_),
    .o1(_06085_));
 b15aoi012ar1n02x5 _31709_ (.a(_05969_),
    .b(_06082_),
    .c(_06085_),
    .o1(_06086_));
 b15norp02as1n04x5 _31710_ (.a(_06079_),
    .b(_06086_),
    .o1(_06087_));
 b15oai112as1n16x5 _31711_ (.a(_06043_),
    .b(_06066_),
    .c(_06087_),
    .d(_05911_),
    .o1(_06088_));
 b15inv000as1n48x5 _31712_ (.a(net558),
    .o1(_06089_));
 b15ztpn00an1n08x5 PHY_323 ();
 b15orn002aq1n32x5 _31714_ (.a(\us33.a[5] ),
    .b(\us33.a[4] ),
    .o(_06091_));
 b15ztpn00an1n08x5 PHY_322 ();
 b15ztpn00an1n08x5 PHY_321 ();
 b15ztpn00an1n08x5 PHY_320 ();
 b15nanb02as1n24x5 _31718_ (.a(\us33.a[7] ),
    .b(net546),
    .out0(_06096_));
 b15ztpn00an1n08x5 PHY_319 ();
 b15ztpn00an1n08x5 PHY_318 ();
 b15ztpn00an1n08x5 PHY_317 ();
 b15nandp2as1n24x5 _31722_ (.a(net566),
    .b(net556),
    .o1(_06100_));
 b15nor004aq1n02x5 _31723_ (.a(_06089_),
    .b(_06091_),
    .c(_06096_),
    .d(_06100_),
    .o1(_06101_));
 b15ztpn00an1n08x5 PHY_316 ();
 b15orn002al1n08x5 _31725_ (.a(net553),
    .b(\us33.a[6] ),
    .o(_06103_));
 b15ztpn00an1n08x5 PHY_315 ();
 b15nandp2aq1n32x5 _31727_ (.a(net553),
    .b(net558),
    .o1(_06105_));
 b15ztpn00an1n08x5 PHY_314 ();
 b15inv040as1n12x5 _31729_ (.a(\us33.a[6] ),
    .o1(_06108_));
 b15oai012an1n04x5 _31730_ (.a(_06103_),
    .b(_06105_),
    .c(_06108_),
    .o1(_06109_));
 b15ztpn00an1n08x5 PHY_313 ();
 b15inv000as1n48x5 _31732_ (.a(net567),
    .o1(_06111_));
 b15ztpn00an1n08x5 PHY_312 ();
 b15ztpn00an1n08x5 PHY_311 ();
 b15nor002ah1n04x5 _31735_ (.a(_06111_),
    .b(\us33.a[7] ),
    .o1(_06114_));
 b15ztpn00an1n08x5 PHY_310 ();
 b15ztpn00an1n08x5 PHY_309 ();
 b15and002ah1n32x5 _31738_ (.a(\us33.a[5] ),
    .b(net551),
    .o(_06118_));
 b15aoi013ar1n04x5 _31739_ (.a(_06101_),
    .b(_06109_),
    .c(_06114_),
    .d(_06118_),
    .o1(_06119_));
 b15ztpn00an1n08x5 PHY_308 ();
 b15nanb02aq1n24x5 _31741_ (.a(net564),
    .b(net555),
    .out0(_06121_));
 b15ztpn00an1n08x5 PHY_307 ();
 b15ztpn00an1n08x5 PHY_306 ();
 b15ztpn00an1n08x5 PHY_305 ();
 b15nona23ah1n32x5 _31745_ (.a(net552),
    .b(net546),
    .c(net543),
    .d(\us33.a[5] ),
    .out0(_06125_));
 b15ztpn00an1n08x5 PHY_304 ();
 b15orn002ah1n24x5 _31747_ (.a(net556),
    .b(net559),
    .o(_06127_));
 b15ztpn00an1n08x5 PHY_303 ();
 b15ztpn00an1n08x5 PHY_302 ();
 b15ztpn00an1n08x5 PHY_301 ();
 b15ztpn00an1n08x5 PHY_300 ();
 b15nona23as1n32x5 _31752_ (.a(net552),
    .b(net543),
    .c(net546),
    .d(net548),
    .out0(_06133_));
 b15oai022as1n04x5 _31753_ (.a(_06121_),
    .b(_06125_),
    .c(_06127_),
    .d(_06133_),
    .o1(_06134_));
 b15nanb02as1n24x5 _31754_ (.a(net549),
    .b(net552),
    .out0(_06135_));
 b15ztpn00an1n08x5 PHY_299 ();
 b15ztpn00an1n08x5 PHY_298 ();
 b15ztpn00an1n08x5 PHY_297 ();
 b15norp02as1n02x5 _31758_ (.a(net553),
    .b(net545),
    .o1(_06140_));
 b15ztpn00an1n08x5 PHY_296 ();
 b15ztpn00an1n08x5 PHY_295 ();
 b15and002al1n12x5 _31761_ (.a(net563),
    .b(net558),
    .o(_06143_));
 b15nor004as1n02x5 _31762_ (.a(net544),
    .b(_06135_),
    .c(_06140_),
    .d(_06143_),
    .o1(_06144_));
 b15nanb02as1n24x5 _31763_ (.a(net553),
    .b(net565),
    .out0(_06145_));
 b15qgbna2an1n05x5 _31764_ (.o1(_06146_),
    .a(\us33.a[6] ),
    .b(_06145_));
 b15aoi012al1n04x5 _31765_ (.a(_06134_),
    .b(_06144_),
    .c(_06146_),
    .o1(_06147_));
 b15ztpn00an1n08x5 PHY_294 ();
 b15ztpn00an1n08x5 PHY_293 ();
 b15ztpn00an1n08x5 PHY_292 ();
 b15ztpn00an1n08x5 PHY_291 ();
 b15ztpn00an1n08x5 PHY_290 ();
 b15ztpn00an1n08x5 PHY_289 ();
 b15nanb02as1n24x5 _31772_ (.a(net559),
    .b(\us33.a[3] ),
    .out0(_06155_));
 b15norp03an1n04x5 _31773_ (.a(_06111_),
    .b(_06133_),
    .c(_06155_),
    .o1(_06156_));
 b15ztpn00an1n08x5 PHY_288 ();
 b15andc04as1n16x5 _31775_ (.a(net548),
    .b(net552),
    .c(net543),
    .d(net546),
    .o(_06158_));
 b15ztpn00an1n08x5 PHY_287 ();
 b15ztpn00an1n08x5 PHY_286 ();
 b15ztpn00an1n08x5 PHY_285 ();
 b15nonb02as1n12x5 _31779_ (.a(net559),
    .b(net556),
    .out0(_06163_));
 b15aoi012as1n08x5 _31780_ (.a(_06156_),
    .b(_06158_),
    .c(_06163_),
    .o1(_06164_));
 b15oai112ar1n16x5 _31781_ (.a(_06119_),
    .b(_06147_),
    .c(net563),
    .d(_06164_),
    .o1(_06165_));
 b15nanb02ah1n12x5 _31782_ (.a(net554),
    .b(\us33.a[5] ),
    .out0(_06166_));
 b15nor002an1n03x5 _31783_ (.a(_06108_),
    .b(_06166_),
    .o1(_06167_));
 b15ztpn00an1n08x5 PHY_284 ();
 b15nor002ah1n06x5 _31785_ (.a(\us33.a[5] ),
    .b(\us33.a[6] ),
    .o1(_06169_));
 b15ztpn00an1n08x5 PHY_283 ();
 b15and002ah1n04x5 _31787_ (.a(net558),
    .b(\us33.a[4] ),
    .o(_06171_));
 b15aoai13ar1n02x5 _31788_ (.a(_06114_),
    .b(_06167_),
    .c(_06169_),
    .d(_06171_),
    .o1(_06173_));
 b15nanb02as1n24x5 _31789_ (.a(net551),
    .b(net547),
    .out0(_06174_));
 b15ztpn00an1n08x5 PHY_282 ();
 b15oai012ah1n06x5 _31791_ (.a(_06174_),
    .b(_06135_),
    .c(_06111_),
    .o1(_06176_));
 b15norp02ar1n02x5 _31792_ (.a(_06105_),
    .b(_06096_),
    .o1(_06177_));
 b15aob012an1n02x5 _31793_ (.a(_06173_),
    .b(_06176_),
    .c(_06177_),
    .out0(_06178_));
 b15inv000ah1n64x5 _31794_ (.a(net563),
    .o1(_06179_));
 b15ztpn00an1n08x5 PHY_281 ();
 b15ztpn00an1n08x5 PHY_280 ();
 b15ztpn00an1n08x5 PHY_279 ();
 b15ztpn00an1n08x5 PHY_278 ();
 b15ztpn00an1n08x5 PHY_277 ();
 b15ztpn00an1n08x5 PHY_276 ();
 b15nanb02as1n03x5 _31801_ (.a(net558),
    .b(\us33.a[5] ),
    .out0(_06187_));
 b15oai013ah1n03x5 _31802_ (.a(_06179_),
    .b(_06145_),
    .c(_06096_),
    .d(_06187_),
    .o1(_06188_));
 b15aoi012ar1n06x5 _31803_ (.a(_06165_),
    .b(_06178_),
    .c(_06188_),
    .o1(_06189_));
 b15ztpn00an1n08x5 PHY_275 ();
 b15ztpn00an1n08x5 PHY_274 ();
 b15ztpn00an1n08x5 PHY_273 ();
 b15nonb02as1n16x5 _31807_ (.a(\us33.a[6] ),
    .b(net544),
    .out0(_06193_));
 b15nand02ah1n48x5 _31808_ (.a(_06193_),
    .b(_06118_),
    .o1(_06195_));
 b15ztpn00an1n08x5 PHY_272 ();
 b15nona23as1n32x5 _31810_ (.a(net549),
    .b(net543),
    .c(net546),
    .d(net550),
    .out0(_06197_));
 b15ztpn00an1n08x5 PHY_271 ();
 b15nand02ah1n06x5 _31812_ (.a(net562),
    .b(_06163_),
    .o1(_06199_));
 b15oai022ar1n02x5 _31813_ (.a(_06155_),
    .b(_06195_),
    .c(_06197_),
    .d(_06199_),
    .o1(_06200_));
 b15inv020as1n56x5 _31814_ (.a(net554),
    .o1(_06201_));
 b15ztpn00an1n08x5 PHY_270 ();
 b15qgbna2an1n05x5 _31816_ (.o1(_06203_),
    .a(_06201_),
    .b(net544));
 b15ztpn00an1n08x5 PHY_269 ();
 b15nor002ah1n06x5 _31818_ (.a(net551),
    .b(net545),
    .o1(_06206_));
 b15nor002as1n24x5 _31819_ (.a(net560),
    .b(net557),
    .o1(_06207_));
 b15nandp3aq1n02x5 _31820_ (.a(net549),
    .b(_06206_),
    .c(_06207_),
    .o1(_06208_));
 b15ztpn00an1n08x5 PHY_268 ();
 b15nandp2al1n08x5 _31822_ (.a(net551),
    .b(net545),
    .o1(_06210_));
 b15inv000al1n20x5 _31823_ (.a(net547),
    .o1(_06211_));
 b15nand02ah1n03x5 _31824_ (.a(net560),
    .b(_06211_),
    .o1(_06212_));
 b15oaoi13aq1n08x5 _31825_ (.a(_06203_),
    .b(_06208_),
    .c(_06210_),
    .d(_06212_),
    .o1(_06213_));
 b15oab012al1n03x5 _31826_ (.a(net566),
    .b(_06200_),
    .c(_06213_),
    .out0(_06214_));
 b15nonb02ah1n16x5 _31827_ (.a(net549),
    .b(net550),
    .out0(_06215_));
 b15nor002an1n24x5 _31828_ (.a(net544),
    .b(net545),
    .o1(_06217_));
 b15nandp2aq1n32x5 _31829_ (.a(net544),
    .b(\us33.a[6] ),
    .o1(_06218_));
 b15nor002ah1n04x5 _31830_ (.a(net555),
    .b(_06218_),
    .o1(_06219_));
 b15and002aq1n24x5 _31831_ (.a(net554),
    .b(net558),
    .o(_06220_));
 b15norp02ah1n48x5 _31832_ (.a(net554),
    .b(\us33.a[2] ),
    .o1(_06221_));
 b15ztpn00an1n08x5 PHY_267 ();
 b15aoi012al1n06x5 _31834_ (.a(_06220_),
    .b(_06221_),
    .c(net566),
    .o1(_06223_));
 b15oai122ar1n12x5 _31835_ (.a(_06215_),
    .b(_06217_),
    .c(_06219_),
    .d(_06223_),
    .e(_06179_),
    .o1(_06224_));
 b15ztpn00an1n08x5 PHY_266 ();
 b15ztpn00an1n08x5 PHY_265 ();
 b15and002as1n24x5 _31838_ (.a(net544),
    .b(net545),
    .o(_06228_));
 b15ztpn00an1n08x5 PHY_264 ();
 b15nand02as1n24x5 _31840_ (.a(_06228_),
    .b(_06215_),
    .o1(_06230_));
 b15aoi022ar1n02x5 _31841_ (.a(_06111_),
    .b(_06127_),
    .c(_06230_),
    .d(_06163_),
    .o1(_06231_));
 b15norp02an1n02x5 _31842_ (.a(net561),
    .b(_06231_),
    .o1(_06232_));
 b15oab012al1n08x5 _31843_ (.c(_06232_),
    .a(_06214_),
    .b(_06224_),
    .out0(_06233_));
 b15ztpn00an1n08x5 PHY_263 ();
 b15orn002aq1n12x5 _31845_ (.a(net558),
    .b(\us33.a[5] ),
    .o(_06235_));
 b15nanb02as1n24x5 _31846_ (.a(net546),
    .b(net543),
    .out0(_06236_));
 b15ztpn00an1n08x5 PHY_262 ();
 b15nor004an1n03x5 _31848_ (.a(net550),
    .b(_06145_),
    .c(_06235_),
    .d(_06236_),
    .o1(_06239_));
 b15nano23as1n24x5 _31849_ (.a(net543),
    .b(net546),
    .c(net549),
    .d(net552),
    .out0(_06240_));
 b15aoi112an1n04x5 _31850_ (.a(_06179_),
    .b(_06239_),
    .c(_06220_),
    .d(_06240_),
    .o1(_06241_));
 b15nonb02as1n16x5 _31851_ (.a(\us33.a[0] ),
    .b(net559),
    .out0(_06242_));
 b15nano23as1n24x5 _31852_ (.a(net552),
    .b(net543),
    .c(net546),
    .d(net549),
    .out0(_06243_));
 b15nand02as1n48x5 _31853_ (.a(\us33.a[5] ),
    .b(net552),
    .o1(_06244_));
 b15nor002ah1n32x5 _31854_ (.a(_06236_),
    .b(_06244_),
    .o1(_06245_));
 b15ztpn00an1n08x5 PHY_261 ();
 b15ztpn00an1n08x5 PHY_260 ();
 b15aoi022an1n06x5 _31857_ (.a(_06242_),
    .b(_06243_),
    .c(_06245_),
    .d(_06201_),
    .o1(_06248_));
 b15ztpn00an1n08x5 PHY_259 ();
 b15ztpn00an1n08x5 PHY_258 ();
 b15ztpn00an1n08x5 PHY_257 ();
 b15nanb02as1n24x5 _31861_ (.a(net567),
    .b(\us33.a[2] ),
    .out0(_06253_));
 b15aoi013ar1n02x5 _31862_ (.a(net561),
    .b(net553),
    .c(_06240_),
    .d(_06253_),
    .o1(_06254_));
 b15nand02as1n08x5 _31863_ (.a(net553),
    .b(net550),
    .o1(_06255_));
 b15ztpn00an1n08x5 PHY_256 ();
 b15norp02an1n12x5 _31865_ (.a(net567),
    .b(\us33.a[5] ),
    .o1(_06257_));
 b15norp03ar1n02x5 _31866_ (.a(net558),
    .b(_06257_),
    .c(_06096_),
    .o1(_06258_));
 b15nonb02ar1n12x5 _31867_ (.a(\us33.a[7] ),
    .b(\us33.a[6] ),
    .out0(_06259_));
 b15ztpn00an1n08x5 PHY_255 ();
 b15aoi013as1n02x5 _31869_ (.a(_06258_),
    .b(_06257_),
    .c(_06259_),
    .d(net558),
    .o1(_06262_));
 b15oai112al1n02x5 _31870_ (.a(_06248_),
    .b(_06254_),
    .c(_06255_),
    .d(_06262_),
    .o1(_06263_));
 b15nor002as1n24x5 _31871_ (.a(net567),
    .b(net554),
    .o1(_06264_));
 b15nonb03an1n12x5 _31872_ (.a(net543),
    .b(net546),
    .c(net550),
    .out0(_06265_));
 b15norp02aq1n24x5 _31873_ (.a(net558),
    .b(net547),
    .o1(_06266_));
 b15aoi013aq1n03x5 _31874_ (.a(_06263_),
    .b(_06264_),
    .c(_06265_),
    .d(_06266_),
    .o1(_06267_));
 b15oai112an1n12x5 _31875_ (.a(_06189_),
    .b(_06233_),
    .c(_06241_),
    .d(_06267_),
    .o1(_06268_));
 b15nand02ar1n48x5 _31876_ (.a(net551),
    .b(\us33.a[7] ),
    .o1(_06269_));
 b15qgbno2an1n10x5 _31877_ (.a(\us33.a[6] ),
    .b(_06269_),
    .o1(_06270_));
 b15nandp2as1n16x5 _31878_ (.a(_06259_),
    .b(_06118_),
    .o1(_06272_));
 b15aoai13an1n06x5 _31879_ (.a(_06111_),
    .b(_06221_),
    .c(_06272_),
    .d(_06220_),
    .o1(_06273_));
 b15nand02aq1n16x5 _31880_ (.a(net558),
    .b(\us33.a[5] ),
    .o1(_06274_));
 b15ztpn00an1n08x5 PHY_254 ();
 b15oai012ar1n02x5 _31882_ (.a(_06274_),
    .b(_06235_),
    .c(_06201_),
    .o1(_06276_));
 b15nand02an1n04x5 _31883_ (.a(net567),
    .b(_06276_),
    .o1(_06277_));
 b15nand04ar1n16x5 _31884_ (.a(_06166_),
    .b(_06270_),
    .c(_06273_),
    .d(_06277_),
    .o1(_06278_));
 b15inv020ah1n12x5 _31885_ (.a(net550),
    .o1(_06279_));
 b15ztpn00an1n08x5 PHY_253 ();
 b15ztpn00an1n08x5 PHY_252 ();
 b15ztpn00an1n08x5 PHY_251 ();
 b15qgbno2an1n05x5 _31889_ (.o1(_06284_),
    .a(net558),
    .b(_06096_));
 b15ztpn00an1n08x5 PHY_250 ();
 b15aoai13aq1n02x5 _31891_ (.a(net567),
    .b(_06284_),
    .c(_06259_),
    .d(net558),
    .o1(_06286_));
 b15orn002al1n32x5 _31892_ (.a(\us33.a[7] ),
    .b(\us33.a[6] ),
    .o(_06287_));
 b15ztpn00an1n08x5 PHY_249 ();
 b15oai112ar1n02x5 _31894_ (.a(_06279_),
    .b(_06286_),
    .c(_06287_),
    .d(_06253_),
    .o1(_06289_));
 b15ztpn00an1n08x5 PHY_248 ();
 b15oai012ar1n02x5 _31896_ (.a(net550),
    .b(_06287_),
    .c(\us33.a[2] ),
    .o1(_06291_));
 b15nand04as1n04x5 _31897_ (.a(_06201_),
    .b(_06211_),
    .c(_06289_),
    .d(_06291_),
    .o1(_06292_));
 b15norp02an1n16x5 _31898_ (.a(_06201_),
    .b(\us33.a[2] ),
    .o1(_06294_));
 b15nor002ah1n24x5 _31899_ (.a(_06236_),
    .b(_06091_),
    .o1(_06295_));
 b15aoi012ar1n04x5 _31900_ (.a(net561),
    .b(_06294_),
    .c(_06295_),
    .o1(_06296_));
 b15aoi022ah1n08x5 _31901_ (.a(net561),
    .b(_06278_),
    .c(_06292_),
    .d(_06296_),
    .o1(_06297_));
 b15nona23as1n32x5 _31902_ (.a(net544),
    .b(net545),
    .c(\us33.a[5] ),
    .d(net551),
    .out0(_06298_));
 b15ztpn00an1n08x5 PHY_247 ();
 b15nand02aq1n04x5 _31904_ (.a(net563),
    .b(net555),
    .o1(_06300_));
 b15norp02ar1n02x5 _31905_ (.a(_06298_),
    .b(_06300_),
    .o1(_06301_));
 b15nor002ah1n04x5 _31906_ (.a(_06135_),
    .b(_06287_),
    .o1(_06302_));
 b15aoi112as1n02x5 _31907_ (.a(\us33.a[2] ),
    .b(_06301_),
    .c(_06302_),
    .d(_06264_),
    .o1(_06303_));
 b15ztpn00an1n08x5 PHY_246 ();
 b15nona22al1n24x5 _31909_ (.a(\us33.a[4] ),
    .b(\us33.a[7] ),
    .c(\us33.a[6] ),
    .out0(_06306_));
 b15orn003an1n04x5 _31910_ (.a(_06179_),
    .b(net547),
    .c(_06306_),
    .o(_06307_));
 b15aoi012ar1n02x5 _31911_ (.a(_06145_),
    .b(_06272_),
    .c(_06307_),
    .o1(_06308_));
 b15ztpn00an1n08x5 PHY_245 ();
 b15nand04ah1n02x5 _31913_ (.a(net549),
    .b(net550),
    .c(net544),
    .d(net545),
    .o1(_06310_));
 b15aoi012ar1n02x5 _31914_ (.a(_06121_),
    .b(_06298_),
    .c(_06310_),
    .o1(_06311_));
 b15and002ah1n16x5 _31915_ (.a(net562),
    .b(\us33.a[0] ),
    .o(_06312_));
 b15nor004as1n12x5 _31916_ (.a(net548),
    .b(net552),
    .c(net543),
    .d(net546),
    .o1(_06313_));
 b15ztpn00an1n08x5 PHY_244 ();
 b15aoi013aq1n04x5 _31918_ (.a(_06311_),
    .b(_06312_),
    .c(_06313_),
    .d(_06201_),
    .o1(_06316_));
 b15aoi012ah1n02x5 _31919_ (.a(_06167_),
    .b(_06257_),
    .c(_06108_),
    .o1(_06317_));
 b15nanb02an1n24x5 _31920_ (.a(net544),
    .b(net551),
    .out0(_06318_));
 b15oai013ar1n02x5 _31921_ (.a(_06316_),
    .b(_06317_),
    .c(_06318_),
    .d(net560),
    .o1(_06319_));
 b15norp02aq1n02x5 _31922_ (.a(_06308_),
    .b(_06319_),
    .o1(_06320_));
 b15aoi012aq1n06x5 _31923_ (.a(_06303_),
    .b(_06320_),
    .c(\us33.a[2] ),
    .o1(_06321_));
 b15ztpn00an1n08x5 PHY_243 ();
 b15ztpn00an1n08x5 PHY_242 ();
 b15nor002al1n16x5 _31926_ (.a(net547),
    .b(net551),
    .o1(_06324_));
 b15nandp2al1n24x5 _31927_ (.a(_06324_),
    .b(_06228_),
    .o1(_06325_));
 b15nor002aq1n12x5 _31928_ (.a(net561),
    .b(net566),
    .o1(_06327_));
 b15oai012aq1n06x5 _31929_ (.a(net557),
    .b(_06325_),
    .c(_06327_),
    .o1(_06328_));
 b15ztpn00an1n08x5 PHY_241 ();
 b15aoai13ar1n02x5 _31931_ (.a(_06179_),
    .b(_06118_),
    .c(_06324_),
    .d(_06111_),
    .o1(_06330_));
 b15oaoi13an1n02x5 _31932_ (.a(_06218_),
    .b(_06330_),
    .c(_06244_),
    .d(net564),
    .o1(_06331_));
 b15oaoi13as1n03x5 _31933_ (.a(net555),
    .b(_06328_),
    .c(_06331_),
    .d(net557),
    .o1(_06332_));
 b15nonb02as1n12x5 _31934_ (.a(net563),
    .b(net558),
    .out0(_06333_));
 b15nand02ar1n02x5 _31935_ (.a(net564),
    .b(net551),
    .o1(_06334_));
 b15nand04al1n03x5 _31936_ (.a(_06211_),
    .b(_06193_),
    .c(_06333_),
    .d(_06334_),
    .o1(_06335_));
 b15nand02ah1n03x5 _31937_ (.a(net560),
    .b(net557),
    .o1(_06336_));
 b15oai112an1n04x5 _31938_ (.a(net555),
    .b(_06335_),
    .c(_06195_),
    .d(_06336_),
    .o1(_06338_));
 b15nand02al1n16x5 _31939_ (.a(net557),
    .b(_06313_),
    .o1(_06339_));
 b15oab012aq1n03x5 _31940_ (.a(_06338_),
    .b(_06339_),
    .c(_06312_),
    .out0(_06340_));
 b15nor002al1n16x5 _31941_ (.a(_06218_),
    .b(_06174_),
    .o1(_06341_));
 b15aoi012an1n02x5 _31942_ (.a(_06218_),
    .b(_06135_),
    .c(_06174_),
    .o1(_06342_));
 b15aoi022ar1n02x5 _31943_ (.a(_06089_),
    .b(_06341_),
    .c(_06342_),
    .d(net564),
    .o1(_06343_));
 b15nanb02ar1n06x5 _31944_ (.a(_06343_),
    .b(net560),
    .out0(_06344_));
 b15nanb02an1n16x5 _31945_ (.a(net547),
    .b(net558),
    .out0(_06345_));
 b15nanb03ar1n12x5 _31946_ (.a(net558),
    .b(net547),
    .c(net565),
    .out0(_06346_));
 b15aoi012ah1n02x5 _31947_ (.a(_06210_),
    .b(_06345_),
    .c(_06346_),
    .o1(_06347_));
 b15ztpn00an1n08x5 PHY_240 ();
 b15aoi012aq1n02x5 _31949_ (.a(_06174_),
    .b(\us33.a[6] ),
    .c(net564),
    .o1(_06350_));
 b15oai112an1n12x5 _31950_ (.a(_06179_),
    .b(net544),
    .c(_06347_),
    .d(_06350_),
    .o1(_06351_));
 b15aoi013as1n08x5 _31951_ (.a(_06332_),
    .b(_06340_),
    .c(_06344_),
    .d(_06351_),
    .o1(_06352_));
 b15nor004as1n12x5 _31952_ (.a(_06268_),
    .b(_06297_),
    .c(_06321_),
    .d(_06352_),
    .o1(_06353_));
 b15xor002ah1n16x5 _31953_ (.a(_06088_),
    .b(_06353_),
    .out0(_06354_));
 b15ztpn00an1n08x5 PHY_239 ();
 b15oai022ar1n02x5 _31955_ (.a(net931),
    .b(_05972_),
    .c(_06050_),
    .d(_06037_),
    .o1(_06356_));
 b15aoi012al1n02x5 _31956_ (.a(net934),
    .b(net928),
    .c(_06356_),
    .o1(_06357_));
 b15nanb02an1n08x5 _31957_ (.a(net917),
    .b(net920),
    .out0(_06358_));
 b15ztpn00an1n08x5 PHY_238 ();
 b15nanb02ah1n02x5 _31959_ (.a(net915),
    .b(net922),
    .out0(_06361_));
 b15aoi112al1n06x5 _31960_ (.a(_05851_),
    .b(_06358_),
    .c(_06361_),
    .d(_05903_),
    .o1(_06362_));
 b15oai013as1n12x5 _31961_ (.a(net935),
    .b(_05966_),
    .c(_05967_),
    .d(_05835_),
    .o1(_06363_));
 b15nanb02aq1n16x5 _31962_ (.a(net932),
    .b(\us00.a[3] ),
    .out0(_06364_));
 b15orn002as1n04x5 _31963_ (.a(net922),
    .b(net918),
    .o(_06365_));
 b15norp02as1n03x5 _31964_ (.a(_06364_),
    .b(_06365_),
    .o1(_06366_));
 b15nand02an1n03x5 _31965_ (.a(net920),
    .b(net916),
    .o1(_06367_));
 b15nor002as1n08x5 _31966_ (.a(net920),
    .b(net916),
    .o1(_06368_));
 b15aob012al1n06x5 _31967_ (.a(_06367_),
    .b(_06368_),
    .c(net929),
    .out0(_06369_));
 b15aoi112as1n08x5 _31968_ (.a(_06362_),
    .b(_06363_),
    .c(_06366_),
    .d(_06369_),
    .o1(_06371_));
 b15norp02ar1n02x5 _31969_ (.a(_05911_),
    .b(_06034_),
    .o1(_06372_));
 b15aoi012aq1n02x5 _31970_ (.a(_06372_),
    .b(_05964_),
    .c(_05911_),
    .o1(_06373_));
 b15ztpn00an1n08x5 PHY_237 ();
 b15oaoi13aq1n04x5 _31972_ (.a(_06357_),
    .b(_06371_),
    .c(_06373_),
    .d(net928),
    .o1(_06375_));
 b15ztpn00an1n08x5 PHY_236 ();
 b15oaoi13ar1n02x5 _31974_ (.a(_05954_),
    .b(net928),
    .c(_05928_),
    .d(_05854_),
    .o1(_06377_));
 b15nonb02ar1n16x5 _31975_ (.a(net930),
    .b(\us00.a[0] ),
    .out0(_06378_));
 b15nor003al1n03x5 _31976_ (.a(_05883_),
    .b(_05854_),
    .c(_06378_),
    .o1(_06379_));
 b15oai112aq1n02x5 _31977_ (.a(net924),
    .b(_06377_),
    .c(_06379_),
    .d(net928),
    .o1(_06380_));
 b15nanb02as1n24x5 _31978_ (.a(net927),
    .b(\us00.a[0] ),
    .out0(_06382_));
 b15aoi012ar1n02x5 _31979_ (.a(_06382_),
    .b(_05891_),
    .c(_05921_),
    .o1(_06383_));
 b15aoi013ar1n02x5 _31980_ (.a(_06383_),
    .b(_05932_),
    .c(_06382_),
    .d(_05821_),
    .o1(_06384_));
 b15oai012aq1n04x5 _31981_ (.a(_06380_),
    .b(_06384_),
    .c(net924),
    .o1(_06385_));
 b15nanb02an1n24x5 _31982_ (.a(net916),
    .b(net920),
    .out0(_06386_));
 b15ztpn00an1n08x5 PHY_235 ();
 b15nonb02aq1n16x5 _31984_ (.a(net918),
    .b(\us00.a[3] ),
    .out0(_06388_));
 b15nand03ar1n08x5 _31985_ (.a(net923),
    .b(_06388_),
    .c(_05925_),
    .o1(_06389_));
 b15nonb02ar1n08x5 _31986_ (.a(\us00.a[3] ),
    .b(net918),
    .out0(_06390_));
 b15nanb03as1n04x5 _31987_ (.a(net923),
    .b(_05894_),
    .c(_06390_),
    .out0(_06391_));
 b15aoi112as1n08x5 _31988_ (.a(net929),
    .b(_06386_),
    .c(_06389_),
    .d(_06391_),
    .o1(_06393_));
 b15ztpn00an1n08x5 PHY_234 ();
 b15aoi022ar1n02x5 _31990_ (.a(_05918_),
    .b(_06032_),
    .c(_05827_),
    .d(_05969_),
    .o1(_06395_));
 b15nor003ah1n03x5 _31991_ (.a(_05911_),
    .b(_06056_),
    .c(_06395_),
    .o1(_06396_));
 b15nand02an1n24x5 _31992_ (.a(net931),
    .b(_05947_),
    .o1(_06397_));
 b15oai022an1n06x5 _31993_ (.a(_06034_),
    .b(_05851_),
    .c(_05997_),
    .d(_06397_),
    .o1(_06398_));
 b15aoi112aq1n08x5 _31994_ (.a(_06393_),
    .b(_06396_),
    .c(_06398_),
    .d(_05969_),
    .o1(_06399_));
 b15ztpn00an1n08x5 PHY_233 ();
 b15nano23aq1n03x5 _31996_ (.a(net920),
    .b(\us00.a[3] ),
    .c(\us00.a[0] ),
    .d(net923),
    .out0(_06401_));
 b15nonb03an1n03x5 _31997_ (.a(net923),
    .b(\us00.a[3] ),
    .c(net920),
    .out0(_06402_));
 b15oai112an1n12x5 _31998_ (.a(\us00.a[1] ),
    .b(_05898_),
    .c(_06401_),
    .d(_06402_),
    .o1(_06404_));
 b15nand02ah1n24x5 _31999_ (.a(_05975_),
    .b(_05839_),
    .o1(_06405_));
 b15oaoi13as1n08x5 _32000_ (.a(_05918_),
    .b(_06404_),
    .c(_06405_),
    .d(_05993_),
    .o1(_06406_));
 b15ztpn00an1n08x5 PHY_232 ();
 b15nand03al1n02x5 _32002_ (.a(_05894_),
    .b(_05906_),
    .c(_06032_),
    .o1(_06408_));
 b15aoi112aq1n03x5 _32003_ (.a(net919),
    .b(_05854_),
    .c(_06397_),
    .d(_06408_),
    .o1(_06409_));
 b15oaoi13as1n02x5 _32004_ (.a(_05846_),
    .b(_05921_),
    .c(_06378_),
    .d(_06078_),
    .o1(_06410_));
 b15nand03al1n02x5 _32005_ (.a(_06056_),
    .b(_05947_),
    .c(_06032_),
    .o1(_06411_));
 b15nand04ah1n02x5 _32006_ (.a(_05955_),
    .b(_06003_),
    .c(_05906_),
    .d(_06047_),
    .o1(_06412_));
 b15oai112an1n06x5 _32007_ (.a(_06411_),
    .b(_06412_),
    .c(_05841_),
    .d(_06397_),
    .o1(_06413_));
 b15nor004as1n06x5 _32008_ (.a(_06406_),
    .b(_06409_),
    .c(_06410_),
    .d(_06413_),
    .o1(_06415_));
 b15nona23aq1n24x5 _32009_ (.a(_06375_),
    .b(_06385_),
    .c(_06399_),
    .d(_06415_),
    .out0(_06416_));
 b15nand02ar1n02x5 _32010_ (.a(_05898_),
    .b(_05971_),
    .o1(_06417_));
 b15ztpn00an1n08x5 PHY_231 ();
 b15norp03ar1n02x5 _32012_ (.a(net914),
    .b(_05911_),
    .c(_05894_),
    .o1(_06419_));
 b15norp02ar1n02x5 _32013_ (.a(net914),
    .b(_05925_),
    .o1(_06420_));
 b15norp03al1n02x5 _32014_ (.a(_05946_),
    .b(_05918_),
    .c(_06378_),
    .o1(_06421_));
 b15oaoi13aq1n02x5 _32015_ (.a(_06419_),
    .b(_05911_),
    .c(_06420_),
    .d(_06421_),
    .o1(_06422_));
 b15oaoi13an1n03x5 _32016_ (.a(_05935_),
    .b(_06417_),
    .c(_06422_),
    .d(\us00.a[6] ),
    .o1(_06423_));
 b15nonb02as1n12x5 _32017_ (.a(net934),
    .b(net928),
    .out0(_06424_));
 b15aoi022ah1n06x5 _32018_ (.a(_06072_),
    .b(_06046_),
    .c(_06424_),
    .d(_05968_),
    .o1(_06426_));
 b15norp03ar1n02x5 _32019_ (.a(_05928_),
    .b(_05854_),
    .c(_05925_),
    .o1(_06427_));
 b15oai022ar1n02x5 _32020_ (.a(_05928_),
    .b(_05854_),
    .c(_05929_),
    .d(_05883_),
    .o1(_06428_));
 b15aoai13ar1n02x5 _32021_ (.a(net927),
    .b(_06427_),
    .c(_06428_),
    .d(_05954_),
    .o1(_06429_));
 b15aoi012ar1n02x5 _32022_ (.a(net924),
    .b(_06000_),
    .c(_06025_),
    .o1(_06430_));
 b15aoi022an1n04x5 _32023_ (.a(net924),
    .b(_06426_),
    .c(_06429_),
    .d(_06430_),
    .o1(_06431_));
 b15nonb03al1n08x5 _32024_ (.a(net929),
    .b(net932),
    .c(\us00.a[0] ),
    .out0(_06432_));
 b15nand03ar1n02x5 _32025_ (.a(_05911_),
    .b(_06432_),
    .c(_05827_),
    .o1(_06433_));
 b15orn002al1n12x5 _32026_ (.a(\us00.a[0] ),
    .b(\us00.a[2] ),
    .o(_06434_));
 b15nand04as1n16x5 _32027_ (.a(_05898_),
    .b(_05975_),
    .c(_06434_),
    .d(_06038_),
    .o1(_06435_));
 b15nandp3ar1n03x5 _32028_ (.a(_05839_),
    .b(_05840_),
    .c(_06432_),
    .o1(_06437_));
 b15aoai13ah1n03x5 _32029_ (.a(_06433_),
    .b(_05911_),
    .c(_06435_),
    .d(_06437_),
    .o1(_06438_));
 b15aoi013ar1n03x5 _32030_ (.a(\us00.a[3] ),
    .b(_06081_),
    .c(_06368_),
    .d(net918),
    .o1(_06439_));
 b15nand03as1n08x5 _32031_ (.a(_05918_),
    .b(_05839_),
    .c(_05840_),
    .o1(_06440_));
 b15nandp3as1n04x5 _32032_ (.a(_05821_),
    .b(_05898_),
    .c(_05975_),
    .o1(_06441_));
 b15aoai13ar1n08x5 _32033_ (.a(_06439_),
    .b(net935),
    .c(_06440_),
    .d(_06441_),
    .o1(_06442_));
 b15norp02an1n03x5 _32034_ (.a(net933),
    .b(_06072_),
    .o1(_06443_));
 b15aoi112ah1n06x5 _32035_ (.a(_05899_),
    .b(_06443_),
    .c(_06019_),
    .d(net933),
    .o1(_06444_));
 b15oai013ah1n04x5 _32036_ (.a(\us00.a[3] ),
    .b(_05959_),
    .c(_05969_),
    .d(net927),
    .o1(_06445_));
 b15oaoi13as1n08x5 _32037_ (.a(_06438_),
    .b(_06442_),
    .c(_06444_),
    .d(_06445_),
    .o1(_06446_));
 b15aoi122an1n06x5 _32038_ (.a(net930),
    .b(_06024_),
    .c(_05895_),
    .d(_06046_),
    .e(_06006_),
    .o1(_06448_));
 b15orn002as1n03x5 _32039_ (.a(net921),
    .b(net933),
    .o(_06449_));
 b15nand04ah1n04x5 _32040_ (.a(net919),
    .b(_05947_),
    .c(_05844_),
    .d(_06449_),
    .o1(_06450_));
 b15nand03an1n04x5 _32041_ (.a(net934),
    .b(net925),
    .c(_06026_),
    .o1(_06451_));
 b15aoi013an1n06x5 _32042_ (.a(_06448_),
    .b(_06450_),
    .c(_06451_),
    .d(net931),
    .o1(_06452_));
 b15nor002ar1n24x5 _32043_ (.a(\us00.a[0] ),
    .b(\us00.a[2] ),
    .o1(_06453_));
 b15ztpn00an1n08x5 PHY_230 ();
 b15norp02ar1n02x5 _32045_ (.a(net923),
    .b(\us00.a[3] ),
    .o1(_06455_));
 b15nona23al1n05x5 _32046_ (.a(_06453_),
    .b(_06386_),
    .c(_06455_),
    .d(net918),
    .out0(_06456_));
 b15nano23ar1n12x5 _32047_ (.a(net916),
    .b(net932),
    .c(net935),
    .d(net920),
    .out0(_06457_));
 b15norp02aq1n03x5 _32048_ (.a(net920),
    .b(net918),
    .o1(_06459_));
 b15aoi012aq1n06x5 _32049_ (.a(net916),
    .b(net935),
    .c(net932),
    .o1(_06460_));
 b15aoi122aq1n08x5 _32050_ (.a(_06457_),
    .b(_05870_),
    .c(_06459_),
    .d(_06460_),
    .e(_06012_),
    .o1(_06461_));
 b15oai013ah1n12x5 _32051_ (.a(_06456_),
    .b(_06461_),
    .c(net923),
    .d(_05884_),
    .o1(_06462_));
 b15orn002ah1n04x5 _32052_ (.a(net931),
    .b(net928),
    .o(_06463_));
 b15aoi012an1n02x5 _32053_ (.a(_06463_),
    .b(_05844_),
    .c(_05955_),
    .o1(_06464_));
 b15nand02an1n24x5 _32054_ (.a(_05867_),
    .b(_05844_),
    .o1(_06465_));
 b15aoai13as1n04x5 _32055_ (.a(net934),
    .b(_06464_),
    .c(_06465_),
    .d(_06072_),
    .o1(_06466_));
 b15oai112aq1n02x5 _32056_ (.a(net925),
    .b(_05844_),
    .c(_05867_),
    .d(_05955_),
    .o1(_06467_));
 b15nonb02al1n16x5 _32057_ (.a(net928),
    .b(net934),
    .out0(_06468_));
 b15ztpn00an1n08x5 PHY_229 ();
 b15oaoi13an1n04x5 _32059_ (.a(_06467_),
    .b(_06468_),
    .c(_05821_),
    .d(_06067_),
    .o1(_06471_));
 b15aoi112as1n08x5 _32060_ (.a(_06452_),
    .b(_06462_),
    .c(_06466_),
    .d(_06471_),
    .o1(_06472_));
 b15nona23aq1n16x5 _32061_ (.a(_06423_),
    .b(_06431_),
    .c(_06446_),
    .d(_06472_),
    .out0(_06473_));
 b15norp02ar1n48x5 _32062_ (.a(_06416_),
    .b(_06473_),
    .o1(_06474_));
 b15ztpn00an1n08x5 PHY_228 ();
 b15inv020aq1n80x5 _32064_ (.a(net821),
    .o1(_06476_));
 b15ztpn00an1n08x5 PHY_227 ();
 b15ztpn00an1n08x5 PHY_226 ();
 b15ztpn00an1n08x5 PHY_225 ();
 b15ztpn00an1n08x5 PHY_224 ();
 b15ztpn00an1n08x5 PHY_223 ();
 b15ztpn00an1n08x5 PHY_222 ();
 b15ztpn00an1n08x5 PHY_221 ();
 b15ztpn00an1n08x5 PHY_220 ();
 b15ztpn00an1n08x5 PHY_219 ();
 b15ztpn00an1n08x5 PHY_218 ();
 b15nandp2ah1n48x5 _32075_ (.a(\us11.a[5] ),
    .b(net806),
    .o1(_06488_));
 b15ztpn00an1n08x5 PHY_217 ();
 b15ztpn00an1n08x5 PHY_216 ();
 b15ztpn00an1n08x5 PHY_215 ();
 b15ztpn00an1n08x5 PHY_214 ();
 b15ztpn00an1n08x5 PHY_213 ();
 b15xor002an1n04x5 _32081_ (.a(net800),
    .b(net812),
    .out0(_06495_));
 b15nor004al1n02x5 _32082_ (.a(net798),
    .b(net808),
    .c(_06488_),
    .d(_06495_),
    .o1(_06496_));
 b15ztpn00an1n08x5 PHY_212 ();
 b15ztpn00an1n08x5 PHY_211 ();
 b15nonb02as1n16x5 _32085_ (.a(net808),
    .b(net812),
    .out0(_06499_));
 b15ztpn00an1n08x5 PHY_210 ();
 b15norp02an1n32x5 _32087_ (.a(net802),
    .b(net804),
    .o1(_06501_));
 b15aoi013ar1n02x5 _32088_ (.a(_06496_),
    .b(_06499_),
    .c(_06501_),
    .d(net798),
    .o1(_06503_));
 b15ztpn00an1n08x5 PHY_209 ();
 b15ztpn00an1n08x5 PHY_208 ();
 b15ztpn00an1n08x5 PHY_207 ();
 b15ztpn00an1n08x5 PHY_206 ();
 b15ztpn00an1n08x5 PHY_205 ();
 b15nor004as1n12x5 _32094_ (.a(net803),
    .b(net807),
    .c(\us11.a[7] ),
    .d(net800),
    .o1(_06509_));
 b15ztpn00an1n08x5 PHY_204 ();
 b15ztpn00an1n08x5 PHY_203 ();
 b15ztpn00an1n08x5 PHY_202 ();
 b15nonb02as1n16x5 _32098_ (.a(net812),
    .b(net815),
    .out0(_06514_));
 b15ztpn00an1n08x5 PHY_201 ();
 b15nandp3ar1n02x5 _32100_ (.a(net808),
    .b(_06509_),
    .c(_06514_),
    .o1(_06516_));
 b15aoi012an1n02x5 _32101_ (.a(_06476_),
    .b(_06503_),
    .c(_06516_),
    .o1(_06517_));
 b15and002ar1n24x5 _32102_ (.a(net817),
    .b(net813),
    .o(_06518_));
 b15nandp2aq1n08x5 _32103_ (.a(net819),
    .b(net810),
    .o1(_06519_));
 b15and003ar1n04x5 _32104_ (.a(_06509_),
    .b(_06518_),
    .c(_06519_),
    .o(_06520_));
 b15ztpn00an1n08x5 PHY_200 ();
 b15nanb02aq1n12x5 _32106_ (.a(net804),
    .b(net799),
    .out0(_06522_));
 b15ztpn00an1n08x5 PHY_199 ();
 b15nanb02an1n16x5 _32108_ (.a(net799),
    .b(net805),
    .out0(_06525_));
 b15ztpn00an1n08x5 PHY_198 ();
 b15nanb02as1n24x5 _32110_ (.a(\us11.a[0] ),
    .b(net818),
    .out0(_06527_));
 b15ztpn00an1n08x5 PHY_197 ();
 b15oai012ah1n03x5 _32112_ (.a(_06522_),
    .b(_06525_),
    .c(_06527_),
    .o1(_06529_));
 b15nonb02as1n16x5 _32113_ (.a(net812),
    .b(net808),
    .out0(_06530_));
 b15ztpn00an1n08x5 PHY_196 ();
 b15ztpn00an1n08x5 PHY_195 ();
 b15nonb02ah1n12x5 _32116_ (.a(net803),
    .b(net797),
    .out0(_06533_));
 b15aoi013as1n06x5 _32117_ (.a(_06520_),
    .b(_06529_),
    .c(_06530_),
    .d(_06533_),
    .o1(_06534_));
 b15inv040an1n60x5 _32118_ (.a(net808),
    .o1(_06536_));
 b15ztpn00an1n08x5 PHY_194 ();
 b15and002al1n24x5 _32120_ (.a(net798),
    .b(net800),
    .o(_06538_));
 b15nonb02as1n16x5 _32121_ (.a(net803),
    .b(net805),
    .out0(_06539_));
 b15ztpn00an1n08x5 PHY_193 ();
 b15nandp3as1n03x5 _32123_ (.a(_06536_),
    .b(_06538_),
    .c(_06539_),
    .o1(_06541_));
 b15nanb02as1n24x5 _32124_ (.a(net815),
    .b(net812),
    .out0(_06542_));
 b15ztpn00an1n08x5 PHY_192 ();
 b15ztpn00an1n08x5 PHY_191 ();
 b15nonb02as1n16x5 _32127_ (.a(net805),
    .b(net803),
    .out0(_06545_));
 b15ztpn00an1n08x5 PHY_190 ();
 b15norp02an1n32x5 _32129_ (.a(net815),
    .b(net808),
    .o1(_06548_));
 b15nand04al1n02x5 _32130_ (.a(net798),
    .b(net821),
    .c(_06545_),
    .d(_06548_),
    .o1(_06549_));
 b15oai122ah1n04x5 _32131_ (.a(_06534_),
    .b(_06541_),
    .c(_06542_),
    .d(_06495_),
    .e(_06549_),
    .o1(_06550_));
 b15ztpn00an1n08x5 PHY_189 ();
 b15inv000ah1n16x5 _32133_ (.a(net797),
    .o1(_06552_));
 b15nonb03as1n12x5 _32134_ (.a(net799),
    .b(net804),
    .c(net802),
    .out0(_06553_));
 b15nandp2as1n12x5 _32135_ (.a(_06552_),
    .b(_06553_),
    .o1(_06554_));
 b15and002as1n32x5 _32136_ (.a(net802),
    .b(net804),
    .o(_06555_));
 b15nonb02as1n16x5 _32137_ (.a(net798),
    .b(net801),
    .out0(_06556_));
 b15nand02ah1n32x5 _32138_ (.a(_06555_),
    .b(_06556_),
    .o1(_06558_));
 b15ztpn00an1n08x5 PHY_188 ();
 b15aoi012ar1n02x5 _32140_ (.a(net809),
    .b(_06554_),
    .c(_06558_),
    .o1(_06560_));
 b15ztpn00an1n08x5 PHY_187 ();
 b15ztpn00an1n08x5 PHY_186 ();
 b15ztpn00an1n08x5 PHY_185 ();
 b15ztpn00an1n08x5 PHY_184 ();
 b15nonb02aq1n16x5 _32145_ (.a(net812),
    .b(net821),
    .out0(_06565_));
 b15oai012ar1n04x5 _32146_ (.a(net815),
    .b(_06558_),
    .c(_06565_),
    .o1(_06566_));
 b15norp02ah1n48x5 _32147_ (.a(net818),
    .b(net814),
    .o1(_06567_));
 b15ztpn00an1n08x5 PHY_183 ();
 b15ztpn00an1n08x5 PHY_182 ();
 b15ztpn00an1n08x5 PHY_181 ();
 b15aoi022al1n02x5 _32151_ (.a(_06567_),
    .b(_06554_),
    .c(_06558_),
    .d(net812),
    .o1(_06572_));
 b15oai112ah1n06x5 _32152_ (.a(_06560_),
    .b(_06566_),
    .c(_06476_),
    .d(_06572_),
    .o1(_06573_));
 b15inv040ah1n40x5 _32153_ (.a(net812),
    .o1(_06574_));
 b15ztpn00an1n08x5 PHY_180 ();
 b15ztpn00an1n08x5 PHY_179 ();
 b15nonb02as1n16x5 _32156_ (.a(net815),
    .b(net821),
    .out0(_06577_));
 b15ztpn00an1n08x5 PHY_178 ();
 b15nano23as1n24x5 _32158_ (.a(net798),
    .b(net801),
    .c(\us11.a[5] ),
    .d(net806),
    .out0(_06580_));
 b15nand02al1n02x5 _32159_ (.a(_06577_),
    .b(_06580_),
    .o1(_06581_));
 b15ztpn00an1n08x5 PHY_177 ();
 b15ztpn00an1n08x5 PHY_176 ();
 b15aoi013an1n02x5 _32162_ (.a(net809),
    .b(_06501_),
    .c(_06556_),
    .d(_06476_),
    .o1(_06584_));
 b15ztpn00an1n08x5 PHY_175 ();
 b15nonb02al1n08x5 _32164_ (.a(net801),
    .b(net798),
    .out0(_06586_));
 b15nandp2ah1n16x5 _32165_ (.a(_06586_),
    .b(_06555_),
    .o1(_06587_));
 b15oai112ar1n08x5 _32166_ (.a(_06581_),
    .b(_06584_),
    .c(_06587_),
    .d(_06577_),
    .o1(_06588_));
 b15nandp2ar1n32x5 _32167_ (.a(_06538_),
    .b(_06545_),
    .o1(_06589_));
 b15ztpn00an1n08x5 PHY_174 ();
 b15ztpn00an1n08x5 PHY_173 ();
 b15nona23as1n32x5 _32170_ (.a(net807),
    .b(\us11.a[7] ),
    .c(net801),
    .d(\us11.a[5] ),
    .out0(_06593_));
 b15oai012al1n03x5 _32171_ (.a(_06589_),
    .b(_06593_),
    .c(_06577_),
    .o1(_06594_));
 b15ztpn00an1n08x5 PHY_172 ();
 b15oai112aq1n08x5 _32173_ (.a(_06574_),
    .b(_06588_),
    .c(_06594_),
    .d(_06536_),
    .o1(_06596_));
 b15nona23aq1n12x5 _32174_ (.a(_06517_),
    .b(_06550_),
    .c(_06573_),
    .d(_06596_),
    .out0(_06597_));
 b15ztpn00an1n08x5 PHY_171 ();
 b15ztpn00an1n08x5 PHY_170 ();
 b15nona23as1n32x5 _32177_ (.a(\us11.a[5] ),
    .b(net798),
    .c(net801),
    .d(net806),
    .out0(_06600_));
 b15nonb02as1n16x5 _32178_ (.a(net815),
    .b(net812),
    .out0(_06602_));
 b15ztpn00an1n08x5 PHY_169 ();
 b15nor004aq1n08x5 _32180_ (.a(net809),
    .b(_06514_),
    .c(_06600_),
    .d(_06602_),
    .o1(_06604_));
 b15nanb02as1n24x5 _32181_ (.a(net814),
    .b(net815),
    .out0(_06605_));
 b15nano23ah1n24x5 _32182_ (.a(\us11.a[5] ),
    .b(net798),
    .c(net801),
    .d(net806),
    .out0(_06606_));
 b15ztpn00an1n08x5 PHY_168 ();
 b15oai112an1n06x5 _32184_ (.a(_06605_),
    .b(_06606_),
    .c(net820),
    .d(_06514_),
    .o1(_06608_));
 b15nor002aq1n12x5 _32185_ (.a(net820),
    .b(net818),
    .o1(_06609_));
 b15nandp2ah1n24x5 _32186_ (.a(_06501_),
    .b(_06556_),
    .o1(_06610_));
 b15ztpn00an1n08x5 PHY_167 ();
 b15oai013ah1n08x5 _32188_ (.a(_06608_),
    .b(_06609_),
    .c(_06610_),
    .d(_06574_),
    .o1(_06613_));
 b15aoi012al1n16x5 _32189_ (.a(_06604_),
    .b(_06613_),
    .c(net809),
    .o1(_06614_));
 b15orn002ah1n08x5 _32190_ (.a(\us11.a[5] ),
    .b(net806),
    .o(_06615_));
 b15nor002al1n24x5 _32191_ (.a(\us11.a[0] ),
    .b(net813),
    .o1(_06616_));
 b15ztpn00an1n08x5 PHY_166 ();
 b15ztpn00an1n08x5 PHY_165 ();
 b15nandp3as1n03x5 _32194_ (.a(\us11.a[0] ),
    .b(net818),
    .c(net813),
    .o1(_06619_));
 b15nano22ah1n12x5 _32195_ (.a(net801),
    .b(\us11.a[3] ),
    .c(net798),
    .out0(_06620_));
 b15nona23al1n05x5 _32196_ (.a(_06615_),
    .b(_06616_),
    .c(_06619_),
    .d(_06620_),
    .out0(_06621_));
 b15ztpn00an1n08x5 PHY_164 ();
 b15nor004an1n03x5 _32198_ (.a(net806),
    .b(net801),
    .c(\us11.a[0] ),
    .d(net818),
    .o1(_06623_));
 b15and002ar1n32x5 _32199_ (.a(\us11.a[0] ),
    .b(net818),
    .o(_06624_));
 b15ztpn00an1n08x5 PHY_163 ();
 b15aoi013aq1n06x5 _32201_ (.a(_06623_),
    .b(_06624_),
    .c(net801),
    .d(net806),
    .o1(_06626_));
 b15orn002aq1n12x5 _32202_ (.a(net802),
    .b(net797),
    .o(_06627_));
 b15orn002al1n32x5 _32203_ (.a(net814),
    .b(net809),
    .o(_06628_));
 b15ztpn00an1n08x5 PHY_162 ();
 b15oai013ah1n12x5 _32205_ (.a(_06621_),
    .b(_06626_),
    .c(_06627_),
    .d(_06628_),
    .o1(_06630_));
 b15orn002ar1n24x5 _32206_ (.a(net817),
    .b(net813),
    .o(_06631_));
 b15inv000al1n56x5 _32207_ (.a(net818),
    .o1(_06632_));
 b15ztpn00an1n08x5 PHY_161 ();
 b15oai012ar1n02x5 _32209_ (.a(_06476_),
    .b(_06632_),
    .c(_06499_),
    .o1(_06635_));
 b15and003ar1n02x5 _32210_ (.a(_06631_),
    .b(_06619_),
    .c(_06635_),
    .o(_06636_));
 b15nanb03al1n08x5 _32211_ (.a(net798),
    .b(net801),
    .c(\us11.a[3] ),
    .out0(_06637_));
 b15norp02al1n32x5 _32212_ (.a(net798),
    .b(net801),
    .o1(_06638_));
 b15nand02an1n32x5 _32213_ (.a(_06545_),
    .b(_06638_),
    .o1(_06639_));
 b15oai022al1n02x5 _32214_ (.a(_06488_),
    .b(_06637_),
    .c(_06639_),
    .d(net809),
    .o1(_06640_));
 b15aoi012an1n04x5 _32215_ (.a(_06630_),
    .b(_06636_),
    .c(_06640_),
    .o1(_06641_));
 b15nanb02as1n24x5 _32216_ (.a(net815),
    .b(net821),
    .out0(_06642_));
 b15nand02aq1n32x5 _32217_ (.a(\us11.a[7] ),
    .b(net800),
    .o1(_06643_));
 b15nanb02as1n24x5 _32218_ (.a(net803),
    .b(net805),
    .out0(_06645_));
 b15ztpn00an1n08x5 PHY_160 ();
 b15norp02ar1n08x5 _32220_ (.a(_06643_),
    .b(_06645_),
    .o1(_06647_));
 b15aoi022as1n04x5 _32221_ (.a(net809),
    .b(_06647_),
    .c(_06509_),
    .d(_06530_),
    .o1(_06648_));
 b15oai112as1n16x5 _32222_ (.a(_06614_),
    .b(_06641_),
    .c(_06642_),
    .d(_06648_),
    .o1(_06649_));
 b15and002an1n32x5 _32223_ (.a(net814),
    .b(net808),
    .o(_06650_));
 b15ztpn00an1n08x5 PHY_159 ();
 b15nano23as1n24x5 _32225_ (.a(\us11.a[5] ),
    .b(net806),
    .c(net798),
    .d(net801),
    .out0(_06652_));
 b15nand02as1n08x5 _32226_ (.a(_06650_),
    .b(_06652_),
    .o1(_06653_));
 b15inv000an1n16x5 _32227_ (.a(net805),
    .o1(_06654_));
 b15ztpn00an1n08x5 PHY_158 ();
 b15nand02ar1n02x5 _32229_ (.a(net802),
    .b(net820),
    .o1(_06657_));
 b15nand04ar1n02x5 _32230_ (.a(_06654_),
    .b(_06556_),
    .c(_06530_),
    .d(_06657_),
    .o1(_06658_));
 b15nanb02as1n24x5 _32231_ (.a(net812),
    .b(net808),
    .out0(_06659_));
 b15ztpn00an1n08x5 PHY_157 ();
 b15ornc04as1n24x5 _32233_ (.a(\us11.a[5] ),
    .b(net806),
    .c(net798),
    .d(net801),
    .o(_06661_));
 b15ztpn00an1n08x5 PHY_156 ();
 b15oai112aq1n02x5 _32235_ (.a(_06653_),
    .b(_06658_),
    .c(_06659_),
    .d(_06661_),
    .o1(_06663_));
 b15ztpn00an1n08x5 PHY_155 ();
 b15ztpn00an1n08x5 PHY_154 ();
 b15oai013aq1n03x5 _32238_ (.a(_06663_),
    .b(_06602_),
    .c(_06514_),
    .d(net820),
    .o1(_06667_));
 b15nanb02aq1n06x5 _32239_ (.a(net809),
    .b(net816),
    .out0(_06668_));
 b15nor002ah1n08x5 _32240_ (.a(_06661_),
    .b(_06668_),
    .o1(_06669_));
 b15ztpn00an1n08x5 PHY_153 ();
 b15nanb02aq1n02x5 _32242_ (.a(net816),
    .b(net809),
    .out0(_06671_));
 b15norp03ar1n03x5 _32243_ (.a(net820),
    .b(_06671_),
    .c(_06639_),
    .o1(_06672_));
 b15nonb02aq1n16x5 _32244_ (.a(net815),
    .b(net808),
    .out0(_06673_));
 b15xor002ar1n02x5 _32245_ (.a(_06476_),
    .b(_06673_),
    .out0(_06674_));
 b15nanb02as1n24x5 _32246_ (.a(net805),
    .b(net803),
    .out0(_06675_));
 b15nor002al1n32x5 _32247_ (.a(_06643_),
    .b(_06675_),
    .o1(_06676_));
 b15aoi112aq1n03x5 _32248_ (.a(_06669_),
    .b(_06672_),
    .c(_06674_),
    .d(_06676_),
    .o1(_06678_));
 b15ztpn00an1n08x5 PHY_152 ();
 b15ztpn00an1n08x5 PHY_151 ();
 b15oai012ah1n06x5 _32251_ (.a(_06667_),
    .b(_06678_),
    .c(net814),
    .o1(_06681_));
 b15norp02al1n12x5 _32252_ (.a(net799),
    .b(net815),
    .o1(_06682_));
 b15ztpn00an1n08x5 PHY_150 ();
 b15aoi012ar1n02x5 _32254_ (.a(_06553_),
    .b(_06682_),
    .c(_06555_),
    .o1(_06684_));
 b15nor004aq1n02x5 _32255_ (.a(_06552_),
    .b(net820),
    .c(_06574_),
    .d(_06684_),
    .o1(_06685_));
 b15nandp2aq1n24x5 _32256_ (.a(_06538_),
    .b(_06539_),
    .o1(_06686_));
 b15oaoi13ar1n02x5 _32257_ (.a(_06567_),
    .b(_06686_),
    .c(_06639_),
    .d(net814),
    .o1(_06687_));
 b15ztpn00an1n08x5 PHY_149 ();
 b15aoi112ah1n02x5 _32259_ (.a(_06536_),
    .b(_06685_),
    .c(_06687_),
    .d(net820),
    .o1(_06690_));
 b15and002al1n08x5 _32260_ (.a(net805),
    .b(net797),
    .o(_06691_));
 b15nandp2aq1n02x5 _32261_ (.a(_06476_),
    .b(_06691_),
    .o1(_06692_));
 b15and002al1n08x5 _32262_ (.a(net803),
    .b(net799),
    .o(_06693_));
 b15nand02an1n02x5 _32263_ (.a(_06514_),
    .b(_06693_),
    .o1(_06694_));
 b15ztpn00an1n08x5 PHY_148 ();
 b15ztpn00an1n08x5 PHY_147 ();
 b15oaoi13aq1n08x5 _32266_ (.a(_06692_),
    .b(_06694_),
    .c(_06605_),
    .d(net803),
    .o1(_06697_));
 b15nonb02as1n16x5 _32267_ (.a(net821),
    .b(net812),
    .out0(_06698_));
 b15andc04aq1n16x5 _32268_ (.a(net802),
    .b(net804),
    .c(net797),
    .d(net799),
    .o(_06700_));
 b15aoi112al1n06x5 _32269_ (.a(net808),
    .b(_06697_),
    .c(_06698_),
    .d(_06700_),
    .o1(_06701_));
 b15oai112an1n04x5 _32270_ (.a(_06555_),
    .b(_06602_),
    .c(_06638_),
    .d(_06538_),
    .o1(_06702_));
 b15nandp2ar1n32x5 _32271_ (.a(net821),
    .b(net815),
    .o1(_06703_));
 b15nandp3as1n04x5 _32272_ (.a(_06539_),
    .b(_06638_),
    .c(_06703_),
    .o1(_06704_));
 b15orn002as1n24x5 _32273_ (.a(net819),
    .b(net817),
    .o(_06705_));
 b15norp02al1n12x5 _32274_ (.a(_06574_),
    .b(_06705_),
    .o1(_06706_));
 b15oai122al1n08x5 _32275_ (.a(_06702_),
    .b(_06704_),
    .c(_06706_),
    .d(_06593_),
    .e(_06476_),
    .o1(_06707_));
 b15norp02as1n03x5 _32276_ (.a(net808),
    .b(_06707_),
    .o1(_06708_));
 b15nona23ah1n32x5 _32277_ (.a(\us11.a[5] ),
    .b(net801),
    .c(\us11.a[7] ),
    .d(net806),
    .out0(_06709_));
 b15oai012ar1n02x5 _32278_ (.a(_06709_),
    .b(_06593_),
    .c(net819),
    .o1(_06711_));
 b15ztpn00an1n08x5 PHY_146 ();
 b15nonb02aq1n06x5 _32280_ (.a(net817),
    .b(\us11.a[7] ),
    .out0(_06713_));
 b15nor002ah1n12x5 _32281_ (.a(net800),
    .b(net813),
    .o1(_06714_));
 b15and002an1n02x5 _32282_ (.a(net800),
    .b(net819),
    .o(_06715_));
 b15ao0022ar1n02x5 _32283_ (.a(_06539_),
    .b(_06714_),
    .c(_06715_),
    .d(_06545_),
    .o(_06716_));
 b15aoi022al1n02x5 _32284_ (.a(_06518_),
    .b(_06711_),
    .c(_06713_),
    .d(_06716_),
    .o1(_06717_));
 b15nanb02an1n04x5 _32285_ (.a(net811),
    .b(net802),
    .out0(_06718_));
 b15ztpn00an1n08x5 PHY_145 ();
 b15nandp3al1n04x5 _32287_ (.a(net805),
    .b(net797),
    .c(net800),
    .o1(_06720_));
 b15orn002al1n32x5 _32288_ (.a(\us11.a[7] ),
    .b(net800),
    .o(_06722_));
 b15ztpn00an1n08x5 PHY_144 ();
 b15nanb02ah1n24x5 _32290_ (.a(net805),
    .b(net819),
    .out0(_06724_));
 b15oaoi13an1n02x5 _32291_ (.a(_06718_),
    .b(_06720_),
    .c(_06722_),
    .d(_06724_),
    .o1(_06725_));
 b15nor002an1n08x5 _32292_ (.a(_06675_),
    .b(_06722_),
    .o1(_06726_));
 b15aoi012ar1n02x5 _32293_ (.a(_06725_),
    .b(_06726_),
    .c(_06518_),
    .o1(_06727_));
 b15nona23as1n32x5 _32294_ (.a(\us11.a[5] ),
    .b(net806),
    .c(net798),
    .d(net801),
    .out0(_06728_));
 b15nanb02aq1n12x5 _32295_ (.a(net814),
    .b(net821),
    .out0(_06729_));
 b15oai022al1n16x5 _32296_ (.a(_06728_),
    .b(_06542_),
    .c(_06600_),
    .d(_06729_),
    .o1(_06730_));
 b15oai012ar1n02x5 _32297_ (.a(net810),
    .b(_06527_),
    .c(_06720_),
    .o1(_06731_));
 b15nanb02ah1n03x5 _32298_ (.a(net805),
    .b(net811),
    .out0(_06733_));
 b15oai012an1n08x5 _32299_ (.a(_06733_),
    .b(_06631_),
    .c(_06654_),
    .o1(_06734_));
 b15ztpn00an1n08x5 PHY_143 ();
 b15nanb02as1n03x5 _32301_ (.a(net798),
    .b(\us11.a[5] ),
    .out0(_06736_));
 b15norp03ar1n08x5 _32302_ (.a(net801),
    .b(\us11.a[0] ),
    .c(_06736_),
    .o1(_06737_));
 b15aoi112ar1n02x5 _32303_ (.a(_06730_),
    .b(_06731_),
    .c(_06734_),
    .d(_06737_),
    .o1(_06738_));
 b15and003aq1n08x5 _32304_ (.a(_06717_),
    .b(_06727_),
    .c(_06738_),
    .o(_06739_));
 b15oai022al1n08x5 _32305_ (.a(_06690_),
    .b(_06701_),
    .c(_06708_),
    .d(_06739_),
    .o1(_06740_));
 b15nor004as1n12x5 _32306_ (.a(_06597_),
    .b(_06649_),
    .c(_06681_),
    .d(_06740_),
    .o1(_06741_));
 b15ztpn00an1n08x5 PHY_142 ();
 b15ztpn00an1n08x5 PHY_141 ();
 b15ztpn00an1n08x5 PHY_140 ();
 b15ztpn00an1n08x5 PHY_139 ();
 b15ztpn00an1n08x5 PHY_138 ();
 b15nandp2ah1n48x5 _32312_ (.a(net688),
    .b(net686),
    .o1(_06748_));
 b15ztpn00an1n08x5 PHY_137 ();
 b15ztpn00an1n08x5 PHY_136 ();
 b15ztpn00an1n08x5 PHY_135 ();
 b15ztpn00an1n08x5 PHY_134 ();
 b15ztpn00an1n08x5 PHY_133 ();
 b15ztpn00an1n08x5 PHY_132 ();
 b15nano23aq1n24x5 _32319_ (.a(net674),
    .b(net676),
    .c(\us22.a[7] ),
    .d(net671),
    .out0(_06756_));
 b15ztpn00an1n08x5 PHY_131 ();
 b15inv040al1n40x5 _32321_ (.a(net681),
    .o1(_06758_));
 b15ztpn00an1n08x5 PHY_130 ();
 b15aoi012ar1n02x5 _32323_ (.a(_06748_),
    .b(_06756_),
    .c(_06758_),
    .o1(_06760_));
 b15norp02aq1n48x5 _32324_ (.a(\us22.a[0] ),
    .b(net687),
    .o1(_06761_));
 b15ztpn00an1n08x5 PHY_129 ();
 b15ztpn00an1n08x5 PHY_128 ();
 b15ztpn00an1n08x5 PHY_127 ();
 b15ztpn00an1n08x5 PHY_126 ();
 b15norp02as1n48x5 _32329_ (.a(net669),
    .b(net672),
    .o1(_06767_));
 b15nonb02as1n16x5 _32330_ (.a(\us22.a[5] ),
    .b(\us22.a[4] ),
    .out0(_06768_));
 b15nandp2as1n32x5 _32331_ (.a(_06767_),
    .b(_06768_),
    .o1(_06769_));
 b15ztpn00an1n08x5 PHY_125 ();
 b15oaoi13ar1n02x5 _32333_ (.a(_06760_),
    .b(_06761_),
    .c(net680),
    .d(_06769_),
    .o1(_06771_));
 b15ztpn00an1n08x5 PHY_124 ();
 b15ztpn00an1n08x5 PHY_123 ();
 b15ztpn00an1n08x5 PHY_122 ();
 b15nonb02as1n16x5 _32337_ (.a(net680),
    .b(net685),
    .out0(_06775_));
 b15and002as1n32x5 _32338_ (.a(\us22.a[5] ),
    .b(\us22.a[4] ),
    .o(_06777_));
 b15nand02as1n16x5 _32339_ (.a(_06777_),
    .b(_06767_),
    .o1(_06778_));
 b15norp02ar1n02x5 _32340_ (.a(_06775_),
    .b(_06778_),
    .o1(_06779_));
 b15ztpn00an1n08x5 PHY_121 ();
 b15orn002al1n16x5 _32342_ (.a(net670),
    .b(net671),
    .o(_06781_));
 b15ztpn00an1n08x5 PHY_120 ();
 b15nanb02aq1n24x5 _32344_ (.a(net676),
    .b(net674),
    .out0(_06783_));
 b15norp02as1n08x5 _32345_ (.a(_06781_),
    .b(_06783_),
    .o1(_06784_));
 b15oai022ah1n02x5 _32346_ (.a(net677),
    .b(_06771_),
    .c(_06779_),
    .d(_06784_),
    .o1(_06785_));
 b15inv040as1n60x5 _32347_ (.a(net688),
    .o1(_06786_));
 b15ztpn00an1n08x5 PHY_119 ();
 b15ztpn00an1n08x5 PHY_118 ();
 b15orn002aq1n24x5 _32350_ (.a(\us22.a[1] ),
    .b(net680),
    .o(_06790_));
 b15ztpn00an1n08x5 PHY_117 ();
 b15inv000al1n80x5 _32352_ (.a(net685),
    .o1(_06792_));
 b15ztpn00an1n08x5 PHY_116 ();
 b15ztpn00an1n08x5 PHY_115 ();
 b15oai122al1n08x5 _32355_ (.a(_06786_),
    .b(_06756_),
    .c(_06790_),
    .d(_06784_),
    .e(_06792_),
    .o1(_06795_));
 b15ztpn00an1n08x5 PHY_114 ();
 b15ztpn00an1n08x5 PHY_113 ();
 b15ztpn00an1n08x5 PHY_112 ();
 b15nanb02as1n24x5 _32359_ (.a(net686),
    .b(net682),
    .out0(_06800_));
 b15ztpn00an1n08x5 PHY_111 ();
 b15ztpn00an1n08x5 PHY_110 ();
 b15ztpn00an1n08x5 PHY_109 ();
 b15oai112ah1n04x5 _32363_ (.a(net689),
    .b(_06800_),
    .c(_06784_),
    .d(net680),
    .o1(_06804_));
 b15aoi013ah1n04x5 _32364_ (.a(_06785_),
    .b(_06795_),
    .c(_06804_),
    .d(net677),
    .o1(_06805_));
 b15ztpn00an1n08x5 PHY_108 ();
 b15nano23as1n24x5 _32366_ (.a(net674),
    .b(net671),
    .c(\us22.a[7] ),
    .d(net676),
    .out0(_06807_));
 b15ztpn00an1n08x5 PHY_107 ();
 b15ztpn00an1n08x5 PHY_106 ();
 b15ztpn00an1n08x5 PHY_105 ();
 b15ztpn00an1n08x5 PHY_104 ();
 b15nonb02aq1n06x5 _32371_ (.a(net677),
    .b(net684),
    .out0(_06813_));
 b15ztpn00an1n08x5 PHY_103 ();
 b15ztpn00an1n08x5 PHY_102 ();
 b15ztpn00an1n08x5 PHY_101 ();
 b15oai112an1n06x5 _32375_ (.a(_06758_),
    .b(_06807_),
    .c(_06813_),
    .d(net689),
    .o1(_06817_));
 b15ztpn00an1n08x5 PHY_100 ();
 b15ztpn00an1n08x5 PHY_99 ();
 b15nand02as1n06x5 _32378_ (.a(_06786_),
    .b(_06807_),
    .o1(_06821_));
 b15nonb02as1n16x5 _32379_ (.a(net670),
    .b(net672),
    .out0(_06822_));
 b15nonb02as1n16x5 _32380_ (.a(\us22.a[4] ),
    .b(\us22.a[5] ),
    .out0(_06823_));
 b15nand02ar1n32x5 _32381_ (.a(_06822_),
    .b(_06823_),
    .o1(_06824_));
 b15ztpn00an1n08x5 PHY_98 ();
 b15inv000ah1n64x5 _32383_ (.a(net677),
    .o1(_06826_));
 b15ztpn00an1n08x5 PHY_97 ();
 b15oaoi13as1n02x5 _32385_ (.a(_06792_),
    .b(_06821_),
    .c(_06824_),
    .d(_06826_),
    .o1(_06828_));
 b15ztpn00an1n08x5 PHY_96 ();
 b15ztpn00an1n08x5 PHY_95 ();
 b15aoai13an1n06x5 _32388_ (.a(net680),
    .b(_06828_),
    .c(_06807_),
    .d(_06826_),
    .o1(_06832_));
 b15ztpn00an1n08x5 PHY_94 ();
 b15ztpn00an1n08x5 PHY_93 ();
 b15ztpn00an1n08x5 PHY_92 ();
 b15and003as1n02x5 _32392_ (.a(net675),
    .b(net669),
    .c(\us22.a[6] ),
    .o(_06836_));
 b15nanb02aq1n24x5 _32393_ (.a(\us22.a[0] ),
    .b(net678),
    .out0(_06837_));
 b15nanb02ar1n16x5 _32394_ (.a(net679),
    .b(net688),
    .out0(_06838_));
 b15norp02as1n48x5 _32395_ (.a(\us22.a[5] ),
    .b(\us22.a[4] ),
    .o1(_06839_));
 b15ztpn00an1n08x5 PHY_91 ();
 b15nand03ah1n24x5 _32397_ (.a(net682),
    .b(_06822_),
    .c(_06839_),
    .o1(_06841_));
 b15obai22ar1n16x5 _32398_ (.a(_06836_),
    .b(_06837_),
    .c(_06838_),
    .d(_06841_),
    .out0(_06843_));
 b15nano23as1n24x5 _32399_ (.a(net676),
    .b(net671),
    .c(net670),
    .d(net674),
    .out0(_06844_));
 b15ztpn00an1n08x5 PHY_90 ();
 b15aoi012ar1n04x5 _32401_ (.a(_06843_),
    .b(_06844_),
    .c(net689),
    .o1(_06846_));
 b15oai112al1n12x5 _32402_ (.a(_06817_),
    .b(_06832_),
    .c(_06846_),
    .d(_06792_),
    .o1(_06847_));
 b15ztpn00an1n08x5 PHY_89 ();
 b15nor002ar1n32x5 _32404_ (.a(net682),
    .b(net679),
    .o1(_06849_));
 b15nanb02as1n24x5 _32405_ (.a(\us22.a[1] ),
    .b(net690),
    .out0(_06850_));
 b15nand04al1n08x5 _32406_ (.a(_06777_),
    .b(_06822_),
    .c(_06849_),
    .d(_06850_),
    .o1(_06851_));
 b15nonb02as1n16x5 _32407_ (.a(net671),
    .b(net670),
    .out0(_06852_));
 b15nand02ah1n24x5 _32408_ (.a(_06852_),
    .b(_06839_),
    .o1(_06854_));
 b15ztpn00an1n08x5 PHY_88 ();
 b15ztpn00an1n08x5 PHY_87 ();
 b15ztpn00an1n08x5 PHY_86 ();
 b15orn002al1n08x5 _32412_ (.a(net689),
    .b(net681),
    .o(_06858_));
 b15nandp2aq1n24x5 _32413_ (.a(net684),
    .b(net681),
    .o1(_06859_));
 b15oai112aq1n12x5 _32414_ (.a(net678),
    .b(_06858_),
    .c(_06859_),
    .d(_06786_),
    .o1(_06860_));
 b15oai012aq1n12x5 _32415_ (.a(_06851_),
    .b(_06854_),
    .c(_06860_),
    .o1(_06861_));
 b15nandp2ah1n12x5 _32416_ (.a(net677),
    .b(_06756_),
    .o1(_06862_));
 b15nanb02as1n24x5 _32417_ (.a(net682),
    .b(net686),
    .out0(_06863_));
 b15ztpn00an1n08x5 PHY_85 ();
 b15nor004as1n12x5 _32419_ (.a(net673),
    .b(net675),
    .c(net669),
    .d(net672),
    .o1(_06866_));
 b15nandp2an1n08x5 _32420_ (.a(_06826_),
    .b(_06866_),
    .o1(_06867_));
 b15oai022ah1n06x5 _32421_ (.a(_06800_),
    .b(_06862_),
    .c(_06863_),
    .d(_06867_),
    .o1(_06868_));
 b15nanb02as1n24x5 _32422_ (.a(net679),
    .b(net682),
    .out0(_06869_));
 b15ztpn00an1n08x5 PHY_84 ();
 b15ztpn00an1n08x5 PHY_83 ();
 b15and002al1n08x5 _32425_ (.a(net671),
    .b(net690),
    .o(_06872_));
 b15ztpn00an1n08x5 PHY_82 ();
 b15ztpn00an1n08x5 PHY_81 ();
 b15nano22an1n12x5 _32428_ (.a(net673),
    .b(net675),
    .c(net669),
    .out0(_06876_));
 b15nand02ar1n02x5 _32429_ (.a(_06872_),
    .b(_06876_),
    .o1(_06877_));
 b15nand02an1n48x5 _32430_ (.a(_06822_),
    .b(_06839_),
    .o1(_06878_));
 b15ztpn00an1n08x5 PHY_80 ();
 b15ztpn00an1n08x5 PHY_79 ();
 b15oaoi13al1n02x5 _32433_ (.a(_06869_),
    .b(_06877_),
    .c(_06878_),
    .d(net684),
    .o1(_06881_));
 b15inv040ah1n20x5 _32434_ (.a(net669),
    .o1(_06882_));
 b15ztpn00an1n08x5 PHY_78 ();
 b15ztpn00an1n08x5 PHY_77 ();
 b15ztpn00an1n08x5 PHY_76 ();
 b15ztpn00an1n08x5 PHY_75 ();
 b15and003ar1n08x5 _32439_ (.a(\us22.a[5] ),
    .b(\us22.a[4] ),
    .c(net672),
    .o(_06888_));
 b15and002ah1n12x5 _32440_ (.a(net682),
    .b(net679),
    .o(_06889_));
 b15ztpn00an1n08x5 PHY_74 ();
 b15norp03ar1n02x5 _32442_ (.a(net673),
    .b(net675),
    .c(\us22.a[6] ),
    .o1(_06891_));
 b15aoi022aq1n02x5 _32443_ (.a(_06849_),
    .b(_06888_),
    .c(_06889_),
    .d(_06891_),
    .o1(_06892_));
 b15nor003an1n06x5 _32444_ (.a(_06882_),
    .b(_06892_),
    .c(_06761_),
    .o1(_06893_));
 b15nor004ah1n03x5 _32445_ (.a(_06861_),
    .b(_06868_),
    .c(_06881_),
    .d(_06893_),
    .o1(_06894_));
 b15ztpn00an1n08x5 PHY_73 ();
 b15and002as1n32x5 _32447_ (.a(net670),
    .b(net672),
    .o(_06896_));
 b15ztpn00an1n08x5 PHY_72 ();
 b15nandp3ar1n02x5 _32449_ (.a(_06823_),
    .b(_06896_),
    .c(_06813_),
    .o1(_06899_));
 b15ztpn00an1n08x5 PHY_71 ();
 b15nona23aq1n24x5 _32451_ (.a(net674),
    .b(\us22.a[7] ),
    .c(net671),
    .d(net675),
    .out0(_06901_));
 b15ztpn00an1n08x5 PHY_70 ();
 b15oai112aq1n02x5 _32453_ (.a(net689),
    .b(_06899_),
    .c(_06901_),
    .d(net683),
    .o1(_06903_));
 b15nonb02as1n16x5 _32454_ (.a(net685),
    .b(net680),
    .out0(_06904_));
 b15nand04ar1n02x5 _32455_ (.a(_06826_),
    .b(_06904_),
    .c(_06823_),
    .d(_06896_),
    .o1(_06905_));
 b15nand02as1n48x5 _32456_ (.a(_06777_),
    .b(_06822_),
    .o1(_06906_));
 b15ztpn00an1n08x5 PHY_69 ();
 b15oai013ar1n03x5 _32458_ (.a(_06905_),
    .b(_06800_),
    .c(_06906_),
    .d(_06826_),
    .o1(_06909_));
 b15oai012ah1n04x5 _32459_ (.a(_06903_),
    .b(_06909_),
    .c(net689),
    .o1(_06910_));
 b15nonb02as1n16x5 _32460_ (.a(net688),
    .b(net687),
    .out0(_06911_));
 b15nonb02as1n16x5 _32461_ (.a(net679),
    .b(net682),
    .out0(_06912_));
 b15nand03as1n12x5 _32462_ (.a(_06896_),
    .b(_06768_),
    .c(_06912_),
    .o1(_06913_));
 b15nonb02ar1n16x5 _32463_ (.a(net683),
    .b(net679),
    .out0(_06914_));
 b15nanb02as1n24x5 _32464_ (.a(net688),
    .b(net686),
    .out0(_06915_));
 b15ztpn00an1n08x5 PHY_68 ();
 b15nand02al1n04x5 _32466_ (.a(_06914_),
    .b(_06915_),
    .o1(_06917_));
 b15oai022aq1n12x5 _32467_ (.a(_06911_),
    .b(_06913_),
    .c(_06917_),
    .d(_06906_),
    .o1(_06918_));
 b15ztpn00an1n08x5 PHY_67 ();
 b15orn002al1n16x5 _32469_ (.a(\us22.a[5] ),
    .b(\us22.a[4] ),
    .o(_06921_));
 b15nanb02aq1n16x5 _32470_ (.a(net672),
    .b(net687),
    .out0(_06922_));
 b15nor003al1n06x5 _32471_ (.a(net669),
    .b(_06921_),
    .c(_06922_),
    .o1(_06923_));
 b15andc04as1n16x5 _32472_ (.a(net674),
    .b(net676),
    .c(net670),
    .d(net671),
    .o(_06924_));
 b15aoai13al1n08x5 _32473_ (.a(_06914_),
    .b(_06923_),
    .c(_06924_),
    .d(_06761_),
    .o1(_06925_));
 b15nonb02aq1n06x5 _32474_ (.a(net670),
    .b(net680),
    .out0(_06926_));
 b15and002ah1n16x5 _32475_ (.a(net672),
    .b(net679),
    .o(_06927_));
 b15ztpn00an1n08x5 PHY_66 ();
 b15aoi112ar1n02x5 _32477_ (.a(net671),
    .b(net677),
    .c(_06850_),
    .d(_06915_),
    .o1(_06929_));
 b15oai112ah1n02x5 _32478_ (.a(_06823_),
    .b(_06926_),
    .c(_06927_),
    .d(_06929_),
    .o1(_06931_));
 b15nanb03aq1n06x5 _32479_ (.a(_06918_),
    .b(_06925_),
    .c(_06931_),
    .out0(_06932_));
 b15nandp2ar1n32x5 _32480_ (.a(net674),
    .b(net676),
    .o1(_06933_));
 b15nanb03as1n16x5 _32481_ (.a(net670),
    .b(net671),
    .c(\us22.a[3] ),
    .out0(_06934_));
 b15nor004aq1n02x5 _32482_ (.a(_06792_),
    .b(_06758_),
    .c(_06933_),
    .d(_06934_),
    .o1(_06935_));
 b15nandp2an1n24x5 _32483_ (.a(net670),
    .b(net671),
    .o1(_06936_));
 b15nor003ar1n12x5 _32484_ (.a(net677),
    .b(_06936_),
    .c(_06783_),
    .o1(_06937_));
 b15aoi112an1n03x5 _32485_ (.a(net690),
    .b(_06935_),
    .c(_06937_),
    .d(_06792_),
    .o1(_06938_));
 b15nor004ar1n02x5 _32486_ (.a(\us22.a[1] ),
    .b(_06758_),
    .c(_06933_),
    .d(_06934_),
    .o1(_06939_));
 b15qbfno2bn1n16x5 _32487_ (.a(_06933_),
    .b(_06934_),
    .o1(_06940_));
 b15oaoi13as1n02x5 _32488_ (.a(_06939_),
    .b(_06904_),
    .c(_06937_),
    .d(_06940_),
    .o1(_06942_));
 b15aoi012as1n06x5 _32489_ (.a(_06938_),
    .b(_06942_),
    .c(net690),
    .o1(_06943_));
 b15nano23aq1n08x5 _32490_ (.a(_06894_),
    .b(_06910_),
    .c(_06932_),
    .d(_06943_),
    .out0(_06944_));
 b15nandp2aq1n16x5 _32491_ (.a(\us22.a[3] ),
    .b(_06924_),
    .o1(_06945_));
 b15ztpn00an1n08x5 PHY_65 ();
 b15ztpn00an1n08x5 PHY_64 ();
 b15nand04as1n03x5 _32494_ (.a(_06826_),
    .b(_06777_),
    .c(_06852_),
    .d(_06915_),
    .o1(_06948_));
 b15aoi012al1n06x5 _32495_ (.a(net680),
    .b(_06945_),
    .c(_06948_),
    .o1(_06949_));
 b15nonb02ah1n06x5 _32496_ (.a(net679),
    .b(net672),
    .out0(_06950_));
 b15ztpn00an1n08x5 PHY_63 ();
 b15aoai13al1n06x5 _32498_ (.a(_06950_),
    .b(net688),
    .c(_06882_),
    .d(net687),
    .o1(_06953_));
 b15nanb02ah1n16x5 _32499_ (.a(net687),
    .b(net672),
    .out0(_06954_));
 b15norp02ah1n12x5 _32500_ (.a(net690),
    .b(\us22.a[3] ),
    .o1(_06955_));
 b15nandp3al1n04x5 _32501_ (.a(net669),
    .b(_06954_),
    .c(_06955_),
    .o1(_06956_));
 b15aoi112ah1n06x5 _32502_ (.a(net683),
    .b(_06921_),
    .c(_06953_),
    .d(_06956_),
    .o1(_06957_));
 b15ztpn00an1n08x5 PHY_62 ();
 b15nor003as1n12x5 _32504_ (.a(net669),
    .b(net678),
    .c(_06921_),
    .o1(_06959_));
 b15nor002an1n08x5 _32505_ (.a(\us22.a[6] ),
    .b(net680),
    .o1(_06960_));
 b15nandp3as1n03x5 _32506_ (.a(_06761_),
    .b(_06959_),
    .c(_06960_),
    .o1(_06961_));
 b15nor002ar1n12x5 _32507_ (.a(_06901_),
    .b(_06790_),
    .o1(_06962_));
 b15ztpn00an1n08x5 PHY_61 ();
 b15orn002ah1n04x5 _32509_ (.a(net676),
    .b(\us22.a[3] ),
    .o(_06965_));
 b15and002as1n16x5 _32510_ (.a(net690),
    .b(net680),
    .o(_06966_));
 b15norp03as1n04x5 _32511_ (.a(\us22.a[1] ),
    .b(_06965_),
    .c(_06966_),
    .o1(_06967_));
 b15ztpn00an1n08x5 PHY_60 ();
 b15nanb02ah1n12x5 _32513_ (.a(\us22.a[7] ),
    .b(net671),
    .out0(_06969_));
 b15norp02ar1n02x5 _32514_ (.a(net673),
    .b(_06969_),
    .o1(_06970_));
 b15aoi022as1n04x5 _32515_ (.a(_06826_),
    .b(_06962_),
    .c(_06967_),
    .d(_06970_),
    .o1(_06971_));
 b15nona23ah1n12x5 _32516_ (.a(_06949_),
    .b(_06957_),
    .c(_06961_),
    .d(_06971_),
    .out0(_06972_));
 b15nand02ar1n24x5 _32517_ (.a(_06839_),
    .b(_06896_),
    .o1(_06973_));
 b15nand02aq1n16x5 _32518_ (.a(net681),
    .b(_06866_),
    .o1(_06975_));
 b15oaoi13ah1n04x5 _32519_ (.a(_06860_),
    .b(_06973_),
    .c(_06975_),
    .d(_06761_),
    .o1(_06976_));
 b15nano23aq1n06x5 _32520_ (.a(net673),
    .b(net669),
    .c(net672),
    .d(net675),
    .out0(_06977_));
 b15ztpn00an1n08x5 PHY_59 ();
 b15aoai13as1n02x5 _32522_ (.a(_06977_),
    .b(_06775_),
    .c(net688),
    .d(_06863_),
    .o1(_06979_));
 b15nandp2ar1n32x5 _32523_ (.a(net688),
    .b(net682),
    .o1(_06980_));
 b15nandp2ah1n48x5 _32524_ (.a(_06896_),
    .b(_06768_),
    .o1(_06981_));
 b15ztpn00an1n08x5 PHY_58 ();
 b15oaoi13as1n08x5 _32526_ (.a(_06826_),
    .b(_06979_),
    .c(_06980_),
    .d(_06981_),
    .o1(_06983_));
 b15nanb02aq1n24x5 _32527_ (.a(net674),
    .b(net676),
    .out0(_06984_));
 b15nor002an1n08x5 _32528_ (.a(_06781_),
    .b(_06984_),
    .o1(_06986_));
 b15ztpn00an1n08x5 PHY_57 ();
 b15oai112ar1n04x5 _32530_ (.a(net690),
    .b(_06863_),
    .c(_06869_),
    .d(net685),
    .o1(_06988_));
 b15ztpn00an1n08x5 PHY_56 ();
 b15nanb02as1n24x5 _32532_ (.a(\us22.a[3] ),
    .b(\us22.a[1] ),
    .out0(_06990_));
 b15oai112al1n02x5 _32533_ (.a(_06786_),
    .b(_06990_),
    .c(_06790_),
    .d(_06826_),
    .o1(_06991_));
 b15nand03as1n04x5 _32534_ (.a(_06986_),
    .b(_06988_),
    .c(_06991_),
    .o1(_06992_));
 b15nor002ah1n04x5 _32535_ (.a(_06901_),
    .b(_06990_),
    .o1(_06993_));
 b15norp03ah1n02x5 _32536_ (.a(_06850_),
    .b(_06984_),
    .c(_06936_),
    .o1(_06994_));
 b15nanb03ah1n04x5 _32537_ (.a(\us22.a[6] ),
    .b(net670),
    .c(net674),
    .out0(_06995_));
 b15nor004as1n06x5 _32538_ (.a(\us22.a[1] ),
    .b(_06965_),
    .c(_06966_),
    .d(_06995_),
    .o1(_06997_));
 b15oai013ah1n04x5 _32539_ (.a(net683),
    .b(_06993_),
    .c(_06994_),
    .d(_06997_),
    .o1(_06998_));
 b15inv020aq1n40x5 _32540_ (.a(net672),
    .o1(_06999_));
 b15ztpn00an1n08x5 PHY_55 ();
 b15aoi013ah1n03x5 _32542_ (.a(_06937_),
    .b(_06959_),
    .c(_06999_),
    .d(net690),
    .o1(_07001_));
 b15oai112aq1n16x5 _32543_ (.a(_06992_),
    .b(_06998_),
    .c(_06800_),
    .d(_07001_),
    .o1(_07002_));
 b15nor004as1n12x5 _32544_ (.a(_06972_),
    .b(_06976_),
    .c(_06983_),
    .d(_07002_),
    .o1(_07003_));
 b15nona23as1n32x5 _32545_ (.a(_06805_),
    .b(_06847_),
    .c(_06944_),
    .d(_07003_),
    .out0(_07004_));
 b15xor002an1n16x5 _32546_ (.a(_06741_),
    .b(_07004_),
    .out0(_07005_));
 b15qgbxo2an1n05x5 _32547_ (.a(_06474_),
    .b(_07005_),
    .out0(_07006_));
 b15xor002aq1n08x5 _32548_ (.a(_06354_),
    .b(_07006_),
    .out0(_07008_));
 b15mdn022ar1n16x5 _32549_ (.a(_05814_),
    .b(_07008_),
    .o1(_07009_),
    .sa(net536));
 b15xor002an1n16x5 _32550_ (.a(\u0.w[0][0] ),
    .b(_07009_),
    .out0(_00097_));
 b15nand02as1n32x5 _32551_ (.a(\us33.a[0] ),
    .b(net559),
    .o1(_07010_));
 b15nanb02an1n08x5 _32552_ (.a(net548),
    .b(net554),
    .out0(_07011_));
 b15norp02ah1n32x5 _32553_ (.a(net566),
    .b(net557),
    .o1(_07012_));
 b15ztpn00an1n08x5 PHY_54 ();
 b15nor003as1n06x5 _32555_ (.a(_06306_),
    .b(_07011_),
    .c(_07012_),
    .o1(_07014_));
 b15oai022an1n06x5 _32556_ (.a(net549),
    .b(_06096_),
    .c(_06274_),
    .d(_06236_),
    .o1(_07015_));
 b15orn002aq1n12x5 _32557_ (.a(net561),
    .b(net553),
    .o(_07016_));
 b15nor002as1n03x5 _32558_ (.a(net550),
    .b(_07016_),
    .o1(_07018_));
 b15aoai13an1n06x5 _32559_ (.a(_07010_),
    .b(_07014_),
    .c(_07015_),
    .d(_07018_),
    .o1(_07019_));
 b15nandp2ar1n04x5 _32560_ (.a(net555),
    .b(net549),
    .o1(_07020_));
 b15aoi112ar1n02x5 _32561_ (.a(_07012_),
    .b(_07020_),
    .c(net561),
    .d(_07010_),
    .o1(_07021_));
 b15aoai13al1n02x5 _32562_ (.a(_06265_),
    .b(_07021_),
    .c(_06264_),
    .d(_06266_),
    .o1(_07022_));
 b15ztpn00an1n08x5 PHY_53 ();
 b15norp02an1n03x5 _32564_ (.a(\us33.a[3] ),
    .b(_06133_),
    .o1(_07024_));
 b15nano23aq1n24x5 _32565_ (.a(net552),
    .b(net546),
    .c(net543),
    .d(net548),
    .out0(_07025_));
 b15nanb02ah1n16x5 _32566_ (.a(net562),
    .b(net559),
    .out0(_07026_));
 b15and003ar1n02x5 _32567_ (.a(\us33.a[3] ),
    .b(_07025_),
    .c(_07026_),
    .o(_07027_));
 b15oai012ar1n08x5 _32568_ (.a(\us33.a[0] ),
    .b(_07024_),
    .c(_07027_),
    .o1(_07029_));
 b15nand02aq1n12x5 _32569_ (.a(_06179_),
    .b(_06111_),
    .o1(_07030_));
 b15ztpn00an1n08x5 PHY_52 ();
 b15ornc04as1n24x5 _32571_ (.a(net548),
    .b(net552),
    .c(net543),
    .d(net546),
    .o(_07032_));
 b15and002aq1n24x5 _32572_ (.a(net566),
    .b(net557),
    .o(_07033_));
 b15oaoi13ar1n02x5 _32573_ (.a(net555),
    .b(_07032_),
    .c(_07033_),
    .d(_06298_),
    .o1(_07034_));
 b15orn002as1n04x5 _32574_ (.a(net560),
    .b(net557),
    .o(_07035_));
 b15nano23ah1n08x5 _32575_ (.a(net548),
    .b(net552),
    .c(net543),
    .d(net546),
    .out0(_07036_));
 b15oai112as1n02x5 _32576_ (.a(_07030_),
    .b(_07034_),
    .c(_07035_),
    .d(_07036_),
    .o1(_07037_));
 b15nand04aq1n06x5 _32577_ (.a(_07019_),
    .b(_07022_),
    .c(_07029_),
    .d(_07037_),
    .o1(_07038_));
 b15nand02as1n16x5 _32578_ (.a(_06324_),
    .b(_06193_),
    .o1(_07040_));
 b15oa0022al1n02x5 _32579_ (.a(_06127_),
    .b(_06195_),
    .c(_07040_),
    .d(_06100_),
    .o(_07041_));
 b15and002al1n08x5 _32580_ (.a(net549),
    .b(net544),
    .o(_07042_));
 b15nor004al1n02x5 _32581_ (.a(net550),
    .b(net545),
    .c(_06155_),
    .d(_07042_),
    .o1(_07043_));
 b15oab012al1n03x5 _32582_ (.a(_07043_),
    .b(_06195_),
    .c(net556),
    .out0(_07044_));
 b15nanb03al1n06x5 _32583_ (.a(net559),
    .b(\us33.a[3] ),
    .c(net562),
    .out0(_07045_));
 b15oab012ah1n03x5 _32584_ (.a(\us33.a[0] ),
    .b(_07032_),
    .c(_07045_),
    .out0(_07046_));
 b15oai022ah1n04x5 _32585_ (.a(net561),
    .b(_07041_),
    .c(_07044_),
    .d(_07046_),
    .o1(_07047_));
 b15nonb02as1n16x5 _32586_ (.a(net551),
    .b(net544),
    .out0(_07048_));
 b15xor002aq1n03x5 _32587_ (.a(net562),
    .b(_07033_),
    .out0(_07049_));
 b15norp03ar1n02x5 _32588_ (.a(net553),
    .b(net549),
    .c(net546),
    .o1(_07051_));
 b15nandp2an1n08x5 _32589_ (.a(net549),
    .b(net546),
    .o1(_07052_));
 b15norp03ar1n02x5 _32590_ (.a(_06201_),
    .b(_07052_),
    .c(_07012_),
    .o1(_07053_));
 b15oai112an1n04x5 _32591_ (.a(_07048_),
    .b(_07049_),
    .c(_07051_),
    .d(_07053_),
    .o1(_07054_));
 b15oai022ar1n02x5 _32592_ (.a(_06211_),
    .b(_06096_),
    .c(_07011_),
    .d(_06236_),
    .o1(_07055_));
 b15nand03ar1n04x5 _32593_ (.a(\us33.a[2] ),
    .b(_06279_),
    .c(_07055_),
    .o1(_07056_));
 b15nanb02ah1n24x5 _32594_ (.a(net567),
    .b(net563),
    .out0(_07057_));
 b15nandp2al1n03x5 _32595_ (.a(net554),
    .b(_07057_),
    .o1(_07058_));
 b15aoi012al1n02x5 _32596_ (.a(_07058_),
    .b(_06295_),
    .c(net565),
    .o1(_07059_));
 b15oa0012ar1n08x5 _32597_ (.a(_07054_),
    .b(_07056_),
    .c(_07059_),
    .o(_07060_));
 b15nonb03as1n12x5 _32598_ (.a(net557),
    .b(net564),
    .c(net560),
    .out0(_07062_));
 b15orn003al1n16x5 _32599_ (.a(net551),
    .b(_06166_),
    .c(_06287_),
    .o(_07063_));
 b15nonb02as1n04x5 _32600_ (.a(net555),
    .b(net549),
    .out0(_07064_));
 b15nand03ah1n03x5 _32601_ (.a(net550),
    .b(_06228_),
    .c(_07064_),
    .o1(_07065_));
 b15aoi122ar1n06x5 _32602_ (.a(_07062_),
    .b(_07063_),
    .c(_07065_),
    .d(_06155_),
    .e(_06312_),
    .o1(_07066_));
 b15norp02an1n12x5 _32603_ (.a(net563),
    .b(_06111_),
    .o1(_07067_));
 b15ztpn00an1n08x5 PHY_51 ();
 b15nano22aq1n06x5 _32605_ (.a(net543),
    .b(net546),
    .c(net559),
    .out0(_07069_));
 b15oai112as1n02x5 _32606_ (.a(net555),
    .b(_06215_),
    .c(_06217_),
    .d(_07069_),
    .o1(_07070_));
 b15aoi112al1n03x5 _32607_ (.a(_07067_),
    .b(_07070_),
    .c(_06230_),
    .d(_06207_),
    .o1(_07071_));
 b15ztpn00an1n08x5 PHY_50 ();
 b15nandp3al1n08x5 _32609_ (.a(_06108_),
    .b(_06266_),
    .c(_07048_),
    .o1(_07074_));
 b15xnr002ah1n12x5 _32610_ (.a(net562),
    .b(\us33.a[0] ),
    .out0(_07075_));
 b15mdn022ar1n06x5 _32611_ (.a(_07074_),
    .b(_06339_),
    .o1(_07076_),
    .sa(_07075_));
 b15aoi112ah1n04x5 _32612_ (.a(_07066_),
    .b(_07071_),
    .c(net555),
    .d(_07076_),
    .o1(_07077_));
 b15nona23as1n12x5 _32613_ (.a(_07038_),
    .b(_07047_),
    .c(_07060_),
    .d(_07077_),
    .out0(_07078_));
 b15nandp3al1n08x5 _32614_ (.a(net551),
    .b(net544),
    .c(net545),
    .o1(_07079_));
 b15norp03al1n08x5 _32615_ (.a(_06145_),
    .b(_06345_),
    .c(_07079_),
    .o1(_07080_));
 b15oai013ar1n02x5 _32616_ (.a(_06179_),
    .b(net559),
    .c(_06121_),
    .d(_06298_),
    .o1(_07081_));
 b15norp02as1n02x5 _32617_ (.a(_07080_),
    .b(_07081_),
    .o1(_07082_));
 b15nor003aq1n06x5 _32618_ (.a(net554),
    .b(net558),
    .c(\us33.a[5] ),
    .o1(_07084_));
 b15oab012ar1n02x5 _32619_ (.a(_07084_),
    .b(_07052_),
    .c(_06201_),
    .out0(_07085_));
 b15orn003ah1n04x5 _32620_ (.a(net565),
    .b(_06269_),
    .c(_07085_),
    .o(_07086_));
 b15aoai13ar1n02x5 _32621_ (.a(_06220_),
    .b(_06243_),
    .c(_07036_),
    .d(net566),
    .o1(_07087_));
 b15aoi013al1n02x5 _32622_ (.a(_07082_),
    .b(_07086_),
    .c(_07087_),
    .d(net561),
    .o1(_07088_));
 b15oaoi13an1n03x5 _32623_ (.a(_06179_),
    .b(net565),
    .c(_06089_),
    .d(_06295_),
    .o1(_07089_));
 b15nanb02an1n24x5 _32624_ (.a(net551),
    .b(net544),
    .out0(_07090_));
 b15aob012as1n02x5 _32625_ (.a(_07052_),
    .b(_06169_),
    .c(net557),
    .out0(_07091_));
 b15nanb02an1n06x5 _32626_ (.a(_07090_),
    .b(_07091_),
    .out0(_07092_));
 b15nanb02as1n24x5 _32627_ (.a(net561),
    .b(net566),
    .out0(_07093_));
 b15norp02as1n03x5 _32628_ (.a(net557),
    .b(_07093_),
    .o1(_07095_));
 b15nor004as1n06x5 _32629_ (.a(net554),
    .b(_07089_),
    .c(_07092_),
    .d(_07095_),
    .o1(_07096_));
 b15nonb02as1n16x5 _32630_ (.a(\us33.a[1] ),
    .b(net567),
    .out0(_07097_));
 b15norp03ar1n02x5 _32631_ (.a(_06133_),
    .b(_06155_),
    .c(_07097_),
    .o1(_07098_));
 b15aoi013an1n03x5 _32632_ (.a(_07098_),
    .b(_06327_),
    .c(_06313_),
    .d(_06221_),
    .o1(_07099_));
 b15nand02ar1n24x5 _32633_ (.a(_06179_),
    .b(net556),
    .o1(_07100_));
 b15oai122ah1n02x5 _32634_ (.a(net559),
    .b(_06100_),
    .c(_06230_),
    .d(_06298_),
    .e(_07100_),
    .o1(_07101_));
 b15ztpn00an1n08x5 PHY_49 ();
 b15nor002aq1n04x5 _32636_ (.a(net556),
    .b(_07093_),
    .o1(_07103_));
 b15aoi022ar1n02x5 _32637_ (.a(net556),
    .b(_06158_),
    .c(_07103_),
    .d(_06243_),
    .o1(_07104_));
 b15aob012ar1n04x5 _32638_ (.a(_07101_),
    .b(_07104_),
    .c(_06089_),
    .out0(_07106_));
 b15nona23ah1n08x5 _32639_ (.a(_07088_),
    .b(_07096_),
    .c(_07099_),
    .d(_07106_),
    .out0(_07107_));
 b15nanb02ah1n12x5 _32640_ (.a(net559),
    .b(net566),
    .out0(_07108_));
 b15aoi022ar1n04x5 _32641_ (.a(_06143_),
    .b(_07025_),
    .c(_06333_),
    .d(_06158_),
    .o1(_07109_));
 b15nonb02ar1n12x5 _32642_ (.a(net557),
    .b(net564),
    .out0(_07110_));
 b15ztpn00an1n08x5 PHY_48 ();
 b15aoi022al1n02x5 _32644_ (.a(_07110_),
    .b(_06158_),
    .c(_07025_),
    .d(_06089_),
    .o1(_07112_));
 b15oai112as1n06x5 _32645_ (.a(_07108_),
    .b(_07109_),
    .c(_07112_),
    .d(net561),
    .o1(_07113_));
 b15norp03aq1n03x5 _32646_ (.a(net555),
    .b(_06279_),
    .c(_06108_),
    .o1(_07114_));
 b15nor002an1n08x5 _32647_ (.a(net549),
    .b(net544),
    .o1(_07115_));
 b15oai112aq1n12x5 _32648_ (.a(_07113_),
    .b(_07114_),
    .c(_07115_),
    .d(_07042_),
    .o1(_07117_));
 b15nandp2an1n05x5 _32649_ (.a(net562),
    .b(_06253_),
    .o1(_07118_));
 b15oai013as1n03x5 _32650_ (.a(_07118_),
    .b(_06272_),
    .c(_06242_),
    .d(net562),
    .o1(_07119_));
 b15oaoi13as1n03x5 _32651_ (.a(net555),
    .b(_07119_),
    .c(_06245_),
    .d(_06111_),
    .o1(_07120_));
 b15oai112an1n04x5 _32652_ (.a(net561),
    .b(net555),
    .c(_06325_),
    .d(_07033_),
    .o1(_07121_));
 b15aoai13an1n02x5 _32653_ (.a(net555),
    .b(_07012_),
    .c(_06325_),
    .d(net566),
    .o1(_07122_));
 b15oai112ar1n08x5 _32654_ (.a(_07121_),
    .b(_07122_),
    .c(_06240_),
    .d(_06245_),
    .o1(_07123_));
 b15oai012as1n08x5 _32655_ (.a(_07117_),
    .b(_07120_),
    .c(_07123_),
    .o1(_07124_));
 b15norp03as1n24x5 _32656_ (.a(_07078_),
    .b(_07107_),
    .c(_07124_),
    .o1(_07125_));
 b15xnr002aq1n12x5 _32657_ (.a(_06474_),
    .b(_07125_),
    .out0(_07126_));
 b15nand03an1n06x5 _32658_ (.a(\us11.a[3] ),
    .b(_06545_),
    .c(_06713_),
    .o1(_07128_));
 b15ztpn00an1n08x5 PHY_47 ();
 b15nandp2ah1n16x5 _32660_ (.a(net819),
    .b(net813),
    .o1(_07130_));
 b15nanb02al1n02x5 _32661_ (.a(_07128_),
    .b(_07130_),
    .out0(_07131_));
 b15nanb02as1n12x5 _32662_ (.a(net797),
    .b(net811),
    .out0(_07132_));
 b15orn003ah1n03x5 _32663_ (.a(\us11.a[3] ),
    .b(_06488_),
    .c(_07132_),
    .o(_07133_));
 b15oaoi13ah1n04x5 _32664_ (.a(net800),
    .b(_07131_),
    .c(_07133_),
    .d(_06476_),
    .o1(_07134_));
 b15nor003ah1n06x5 _32665_ (.a(_06675_),
    .b(_06722_),
    .c(_06605_),
    .o1(_07135_));
 b15oab012an1n06x5 _32666_ (.a(_07135_),
    .b(_06619_),
    .c(_06600_),
    .out0(_07136_));
 b15nor002ah1n08x5 _32667_ (.a(_06645_),
    .b(_06722_),
    .o1(_07137_));
 b15norp02ar1n02x5 _32668_ (.a(_06574_),
    .b(_06624_),
    .o1(_07139_));
 b15aoi022aq1n02x5 _32669_ (.a(_06567_),
    .b(_07137_),
    .c(_07139_),
    .d(_06509_),
    .o1(_07140_));
 b15nanb02aq1n16x5 _32670_ (.a(\us11.a[7] ),
    .b(net800),
    .out0(_07141_));
 b15nor002ah1n06x5 _32671_ (.a(_07141_),
    .b(_06645_),
    .o1(_07142_));
 b15aoi022al1n06x5 _32672_ (.a(_06567_),
    .b(_07142_),
    .c(_07137_),
    .d(net813),
    .o1(_07143_));
 b15oai112aq1n12x5 _32673_ (.a(_07136_),
    .b(_07140_),
    .c(_07143_),
    .d(net819),
    .o1(_07144_));
 b15oai022as1n06x5 _32674_ (.a(_06705_),
    .b(_07133_),
    .c(_07128_),
    .d(_07130_),
    .o1(_07145_));
 b15aoi122as1n08x5 _32675_ (.a(_07134_),
    .b(_07144_),
    .c(_06536_),
    .d(net800),
    .e(_07145_),
    .o1(_07146_));
 b15nonb02aq1n12x5 _32676_ (.a(net808),
    .b(net815),
    .out0(_07147_));
 b15nanb02as1n24x5 _32677_ (.a(\us11.a[6] ),
    .b(\us11.a[7] ),
    .out0(_07148_));
 b15nor004ah1n06x5 _32678_ (.a(_06476_),
    .b(net811),
    .c(_06615_),
    .d(_07148_),
    .o1(_07150_));
 b15aoai13ar1n02x5 _32679_ (.a(_07147_),
    .b(_07150_),
    .c(_06565_),
    .d(_06647_),
    .o1(_07151_));
 b15xor002as1n16x5 _32680_ (.a(net821),
    .b(net815),
    .out0(_07152_));
 b15nand04ar1n02x5 _32681_ (.a(_06555_),
    .b(_06556_),
    .c(_06650_),
    .d(_07152_),
    .o1(_07153_));
 b15oai013ar1n02x5 _32682_ (.a(_07153_),
    .b(_07152_),
    .c(_06628_),
    .d(_06728_),
    .o1(_07154_));
 b15nandp2ar1n24x5 _32683_ (.a(net817),
    .b(net810),
    .o1(_07155_));
 b15nanb02as1n08x5 _32684_ (.a(net821),
    .b(net814),
    .out0(_07156_));
 b15nand02an1n24x5 _32685_ (.a(_07156_),
    .b(_06729_),
    .o1(_07157_));
 b15aoi112al1n02x5 _32686_ (.a(_07155_),
    .b(_07157_),
    .c(_06610_),
    .d(_06589_),
    .o1(_07158_));
 b15ztpn00an1n08x5 PHY_46 ();
 b15nand02ar1n48x5 _32688_ (.a(net813),
    .b(\us11.a[3] ),
    .o1(_07161_));
 b15nor004ar1n02x5 _32689_ (.a(\us11.a[0] ),
    .b(net816),
    .c(_06600_),
    .d(_07161_),
    .o1(_07162_));
 b15nor003al1n02x5 _32690_ (.a(_07154_),
    .b(_07158_),
    .c(_07162_),
    .o1(_07163_));
 b15ztpn00an1n08x5 PHY_45 ();
 b15nor004ar1n02x5 _32692_ (.a(_06536_),
    .b(_06643_),
    .c(_06675_),
    .d(_06605_),
    .o1(_07165_));
 b15aoi012an1n02x5 _32693_ (.a(_07165_),
    .b(_06726_),
    .c(_06536_),
    .o1(_07166_));
 b15nona22an1n24x5 _32694_ (.a(\us11.a[5] ),
    .b(net806),
    .c(net801),
    .out0(_07167_));
 b15nor004al1n03x5 _32695_ (.a(net798),
    .b(_06632_),
    .c(_06536_),
    .d(_07167_),
    .o1(_07168_));
 b15nor003al1n08x5 _32696_ (.a(_06632_),
    .b(_06488_),
    .c(_07148_),
    .o1(_07169_));
 b15aoi012al1n04x5 _32697_ (.a(_07168_),
    .b(_07169_),
    .c(_06536_),
    .o1(_07170_));
 b15aoi012ar1n06x5 _32698_ (.a(net819),
    .b(_07166_),
    .c(_07170_),
    .o1(_07172_));
 b15nor002ah1n32x5 _32699_ (.a(net812),
    .b(net808),
    .o1(_07173_));
 b15ztpn00an1n08x5 PHY_44 ();
 b15nand03an1n02x5 _32701_ (.a(_06509_),
    .b(_06609_),
    .c(_07173_),
    .o1(_07175_));
 b15nand04ar1n06x5 _32702_ (.a(_06586_),
    .b(_06555_),
    .c(_06705_),
    .d(_06650_),
    .o1(_07176_));
 b15nand02aq1n06x5 _32703_ (.a(net809),
    .b(_06567_),
    .o1(_07177_));
 b15oai112aq1n08x5 _32704_ (.a(_07175_),
    .b(_07176_),
    .c(_07177_),
    .d(_06709_),
    .o1(_07178_));
 b15norp03ar1n02x5 _32705_ (.a(_06645_),
    .b(_06637_),
    .c(_06624_),
    .o1(_07179_));
 b15oab012ar1n02x5 _32706_ (.a(net811),
    .b(_06669_),
    .c(_07179_),
    .out0(_07180_));
 b15nor002aq1n02x5 _32707_ (.a(net799),
    .b(_06567_),
    .o1(_07181_));
 b15nanb02ah1n12x5 _32708_ (.a(net797),
    .b(net810),
    .out0(_07183_));
 b15nor003as1n03x5 _32709_ (.a(net817),
    .b(_06488_),
    .c(_07183_),
    .o1(_07184_));
 b15orn002ar1n08x5 _32710_ (.a(net817),
    .b(net810),
    .o(_07185_));
 b15nand02al1n24x5 _32711_ (.a(net805),
    .b(net797),
    .o1(_07186_));
 b15oai022aq1n06x5 _32712_ (.a(_07185_),
    .b(_07186_),
    .c(_07183_),
    .d(net805),
    .o1(_07187_));
 b15inv000aq1n08x5 _32713_ (.a(net803),
    .o1(_07188_));
 b15aoai13as1n08x5 _32714_ (.a(_07181_),
    .b(_07184_),
    .c(_07187_),
    .d(_07188_),
    .o1(_07189_));
 b15ztpn00an1n08x5 PHY_43 ();
 b15nano23aq1n24x5 _32716_ (.a(\us11.a[5] ),
    .b(net801),
    .c(net798),
    .d(net806),
    .out0(_07191_));
 b15nandp3ar1n02x5 _32717_ (.a(_06476_),
    .b(net809),
    .c(_07191_),
    .o1(_07192_));
 b15nand04al1n02x5 _32718_ (.a(net814),
    .b(_06536_),
    .c(_06538_),
    .d(_06545_),
    .o1(_07194_));
 b15aob012ah1n04x5 _32719_ (.a(net818),
    .b(_07192_),
    .c(_07194_),
    .out0(_07195_));
 b15nona23al1n04x5 _32720_ (.a(_07178_),
    .b(_07180_),
    .c(_07189_),
    .d(_07195_),
    .out0(_07196_));
 b15nano23an1n05x5 _32721_ (.a(_07151_),
    .b(_07163_),
    .c(_07172_),
    .d(_07196_),
    .out0(_07197_));
 b15nand04as1n16x5 _32722_ (.a(net803),
    .b(net805),
    .c(\us11.a[7] ),
    .d(net800),
    .o1(_07198_));
 b15oai122ar1n08x5 _32723_ (.a(\us11.a[0] ),
    .b(_06593_),
    .c(_06628_),
    .d(_07198_),
    .e(_07155_),
    .o1(_07199_));
 b15qgbna2an1n05x5 _32724_ (.o1(_07200_),
    .a(net816),
    .b(_07173_));
 b15and003al1n02x5 _32725_ (.a(_06536_),
    .b(_06555_),
    .c(_06714_),
    .o(_07201_));
 b15and002ar1n08x5 _32726_ (.a(net799),
    .b(net811),
    .o(_07202_));
 b15aoi013ah1n04x5 _32727_ (.a(_07201_),
    .b(_07202_),
    .c(_06501_),
    .d(net809),
    .o1(_07203_));
 b15oai122an1n08x5 _32728_ (.a(_06653_),
    .b(_06709_),
    .c(_07200_),
    .d(_07203_),
    .e(_06552_),
    .o1(_07205_));
 b15norp02ar1n48x5 _32729_ (.a(_07141_),
    .b(_06488_),
    .o1(_07206_));
 b15ztpn00an1n08x5 PHY_42 ();
 b15nandp3aq1n02x5 _32731_ (.a(net810),
    .b(_07206_),
    .c(_06602_),
    .o1(_07208_));
 b15norp02al1n16x5 _32732_ (.a(net805),
    .b(net797),
    .o1(_07209_));
 b15nand02as1n06x5 _32733_ (.a(\us11.a[7] ),
    .b(net816),
    .o1(_07210_));
 b15oab012al1n04x5 _32734_ (.a(_07209_),
    .b(_07210_),
    .c(_06488_),
    .out0(_07211_));
 b15nand02an1n04x5 _32735_ (.a(net800),
    .b(net813),
    .o1(_07212_));
 b15oai013ar1n08x5 _32736_ (.a(_07208_),
    .b(_07211_),
    .c(_07212_),
    .d(net810),
    .o1(_07213_));
 b15oai013as1n06x5 _32737_ (.a(_07199_),
    .b(_07205_),
    .c(_07213_),
    .d(\us11.a[0] ),
    .o1(_07214_));
 b15nandp2aq1n04x5 _32738_ (.a(_06671_),
    .b(_06668_),
    .o1(_07216_));
 b15nand04an1n06x5 _32739_ (.a(_06476_),
    .b(net814),
    .c(_06676_),
    .d(_07216_),
    .o1(_07217_));
 b15nonb02aq1n16x5 _32740_ (.a(net799),
    .b(net810),
    .out0(_07218_));
 b15nand04al1n03x5 _32741_ (.a(net799),
    .b(net816),
    .c(net811),
    .d(net810),
    .o1(_07219_));
 b15oai012as1n03x5 _32742_ (.a(_07219_),
    .b(_06659_),
    .c(net799),
    .o1(_07220_));
 b15aoi022as1n08x5 _32743_ (.a(_06545_),
    .b(_07218_),
    .c(_07220_),
    .d(_06539_),
    .o1(_07221_));
 b15oai013al1n12x5 _32744_ (.a(_07217_),
    .b(_07221_),
    .c(_06476_),
    .d(_06552_),
    .o1(_07222_));
 b15nor002as1n03x5 _32745_ (.a(net798),
    .b(_07167_),
    .o1(_07223_));
 b15aoi022ar1n12x5 _32746_ (.a(net811),
    .b(_06580_),
    .c(_07223_),
    .d(_06632_),
    .o1(_07224_));
 b15nanb02aq1n12x5 _32747_ (.a(net809),
    .b(net820),
    .out0(_07225_));
 b15aoi022ar1n02x5 _32748_ (.a(_07206_),
    .b(_06698_),
    .c(_06700_),
    .d(_06514_),
    .o1(_07227_));
 b15oai022as1n04x5 _32749_ (.a(_07224_),
    .b(_07225_),
    .c(_07227_),
    .d(net809),
    .o1(_07228_));
 b15norp03al1n12x5 _32750_ (.a(\us11.a[7] ),
    .b(net810),
    .c(_07167_),
    .o1(_07229_));
 b15nonb02an1n16x5 _32751_ (.a(net810),
    .b(net799),
    .out0(_07230_));
 b15aoai13aq1n06x5 _32752_ (.a(_06698_),
    .b(_07229_),
    .c(_07230_),
    .d(_06555_),
    .o1(_07231_));
 b15nonb03an1n04x5 _32753_ (.a(net802),
    .b(net804),
    .c(net797),
    .out0(_07232_));
 b15and002aq1n03x5 _32754_ (.a(net797),
    .b(net810),
    .o(_07233_));
 b15aoi022ar1n02x5 _32755_ (.a(_06548_),
    .b(_07232_),
    .c(_07233_),
    .d(_06545_),
    .o1(_07234_));
 b15orn003aq1n02x5 _32756_ (.a(net799),
    .b(_06574_),
    .c(_07234_),
    .o(_07235_));
 b15nanb03ar1n03x5 _32757_ (.a(net816),
    .b(net797),
    .c(net802),
    .out0(_07236_));
 b15aoi112ah1n02x5 _32758_ (.a(_06659_),
    .b(_06522_),
    .c(_06627_),
    .d(_07236_),
    .o1(_07238_));
 b15xor002an1n02x5 _32759_ (.a(net814),
    .b(_06577_),
    .out0(_07239_));
 b15norp02ar1n32x5 _32760_ (.a(_06615_),
    .b(_07148_),
    .o1(_07240_));
 b15aoi013as1n04x5 _32761_ (.a(_07238_),
    .b(_07239_),
    .c(_06536_),
    .d(_07240_),
    .o1(_07241_));
 b15nonb02ah1n04x5 _32762_ (.a(net803),
    .b(net799),
    .out0(_07242_));
 b15xor002al1n04x5 _32763_ (.a(net804),
    .b(net797),
    .out0(_07243_));
 b15and003ar1n03x5 _32764_ (.a(_06705_),
    .b(_07173_),
    .c(_06652_),
    .o(_07244_));
 b15nonb03aq1n12x5 _32765_ (.a(net810),
    .b(net814),
    .c(net816),
    .out0(_07245_));
 b15oai112al1n12x5 _32766_ (.a(_07242_),
    .b(_07243_),
    .c(_07244_),
    .d(_07245_),
    .o1(_07246_));
 b15nand04as1n12x5 _32767_ (.a(_07231_),
    .b(_07235_),
    .c(_07241_),
    .d(_07246_),
    .o1(_07247_));
 b15and002al1n12x5 _32768_ (.a(net799),
    .b(net808),
    .o(_07249_));
 b15norp02an1n24x5 _32769_ (.a(net803),
    .b(net797),
    .o1(_07250_));
 b15and002aq1n08x5 _32770_ (.a(net803),
    .b(net797),
    .o(_07251_));
 b15nor002al1n16x5 _32771_ (.a(net799),
    .b(net810),
    .o1(_07252_));
 b15aoi022an1n02x5 _32772_ (.a(_07249_),
    .b(_07250_),
    .c(_07251_),
    .d(_07252_),
    .o1(_07253_));
 b15nanb02al1n03x5 _32773_ (.a(_06724_),
    .b(_06632_),
    .out0(_07254_));
 b15aoi022an1n02x5 _32774_ (.a(_06650_),
    .b(_06691_),
    .c(_07209_),
    .d(_07173_),
    .o1(_07255_));
 b15nand02aq1n03x5 _32775_ (.a(net816),
    .b(_06693_),
    .o1(_07256_));
 b15oai022an1n08x5 _32776_ (.a(_07253_),
    .b(_07254_),
    .c(_07255_),
    .d(_07256_),
    .o1(_07257_));
 b15nona23as1n24x5 _32777_ (.a(net806),
    .b(net801),
    .c(net798),
    .d(\us11.a[5] ),
    .out0(_07258_));
 b15norp02aq1n02x5 _32778_ (.a(_07258_),
    .b(_07200_),
    .o1(_07260_));
 b15nandp3ar1n03x5 _32779_ (.a(net809),
    .b(_07191_),
    .c(_06602_),
    .o1(_07261_));
 b15norp03ar1n02x5 _32780_ (.a(_07167_),
    .b(_06519_),
    .c(_07210_),
    .o1(_07262_));
 b15nonb02ah1n12x5 _32781_ (.a(\us11.a[0] ),
    .b(\us11.a[1] ),
    .out0(_07263_));
 b15aoi013al1n03x5 _32782_ (.a(_07262_),
    .b(_07263_),
    .c(_06499_),
    .d(_07206_),
    .o1(_07264_));
 b15nona23ar1n08x5 _32783_ (.a(_07257_),
    .b(_07260_),
    .c(_07261_),
    .d(_07264_),
    .out0(_07265_));
 b15nor004an1n12x5 _32784_ (.a(_07222_),
    .b(_07228_),
    .c(_07247_),
    .d(_07265_),
    .o1(_07266_));
 b15nand04as1n16x5 _32785_ (.a(_07146_),
    .b(_07197_),
    .c(_07214_),
    .d(_07266_),
    .o1(_07267_));
 b15ztpn00an1n08x5 PHY_41 ();
 b15nand02ar1n48x5 _32787_ (.a(_06767_),
    .b(_06823_),
    .o1(_07269_));
 b15ztpn00an1n08x5 PHY_40 ();
 b15oaoi13aq1n03x5 _32789_ (.a(net684),
    .b(_06841_),
    .c(_07269_),
    .d(net681),
    .o1(_07272_));
 b15nandp3as1n08x5 _32790_ (.a(net681),
    .b(_06767_),
    .c(_06823_),
    .o1(_07273_));
 b15oaoi13ah1n03x5 _32791_ (.a(net689),
    .b(_07273_),
    .c(_06878_),
    .d(_06863_),
    .o1(_07274_));
 b15nor002ah1n02x5 _32792_ (.a(_06786_),
    .b(_06841_),
    .o1(_07275_));
 b15nor004ar1n08x5 _32793_ (.a(net678),
    .b(_07272_),
    .c(_07274_),
    .d(_07275_),
    .o1(_07276_));
 b15nonb02aq1n08x5 _32794_ (.a(net680),
    .b(net690),
    .out0(_07277_));
 b15nand03as1n03x5 _32795_ (.a(_07277_),
    .b(_06823_),
    .c(_06896_),
    .o1(_07278_));
 b15nanb02ah1n24x5 _32796_ (.a(net681),
    .b(net689),
    .out0(_07279_));
 b15oai112ah1n02x5 _32797_ (.a(_06792_),
    .b(_07278_),
    .c(_07279_),
    .d(_06878_),
    .o1(_07280_));
 b15nand02as1n32x5 _32798_ (.a(_06823_),
    .b(_06896_),
    .o1(_07282_));
 b15ztpn00an1n08x5 PHY_39 ();
 b15aoi022ar1n08x5 _32800_ (.a(_06878_),
    .b(_07282_),
    .c(_06980_),
    .d(_06858_),
    .o1(_07284_));
 b15oai012ah1n06x5 _32801_ (.a(_07280_),
    .b(_07284_),
    .c(_06792_),
    .o1(_07285_));
 b15aoi012al1n12x5 _32802_ (.a(_07276_),
    .b(_07285_),
    .c(net678),
    .o1(_07286_));
 b15nanb02ah1n12x5 _32803_ (.a(net677),
    .b(net671),
    .out0(_07287_));
 b15nonb02aq1n12x5 _32804_ (.a(net669),
    .b(net675),
    .out0(_07288_));
 b15nand02ar1n02x5 _32805_ (.a(_06790_),
    .b(_07288_),
    .o1(_07289_));
 b15ztpn00an1n08x5 PHY_38 ();
 b15and002al1n24x5 _32807_ (.a(net686),
    .b(net682),
    .o(_07291_));
 b15aoai13ar1n02x5 _32808_ (.a(net676),
    .b(_06926_),
    .c(_07291_),
    .d(_06882_),
    .o1(_07293_));
 b15aoi112an1n02x5 _32809_ (.a(net674),
    .b(_07287_),
    .c(_07289_),
    .d(_07293_),
    .o1(_07294_));
 b15aoai13ar1n04x5 _32810_ (.a(net689),
    .b(_07294_),
    .c(_06912_),
    .d(_06756_),
    .o1(_07295_));
 b15ztpn00an1n08x5 PHY_37 ();
 b15xor002ar1n03x5 _32812_ (.a(_06786_),
    .b(_07291_),
    .out0(_07297_));
 b15oai122ar1n08x5 _32813_ (.a(net677),
    .b(_06904_),
    .c(_06824_),
    .d(_07297_),
    .e(_06906_),
    .o1(_07298_));
 b15nandp3ar1n02x5 _32814_ (.a(net680),
    .b(_06924_),
    .c(_06748_),
    .o1(_07299_));
 b15oai013ah1n02x5 _32815_ (.a(_07299_),
    .b(_06775_),
    .c(_06906_),
    .d(net689),
    .o1(_07300_));
 b15oai012al1n06x5 _32816_ (.a(_07298_),
    .b(_07300_),
    .c(net677),
    .o1(_07301_));
 b15nanb02an1n24x5 _32817_ (.a(net672),
    .b(net669),
    .out0(_07302_));
 b15aoi022ar1n04x5 _32818_ (.a(_06914_),
    .b(_06823_),
    .c(_06768_),
    .d(_06912_),
    .o1(_07304_));
 b15norp03ar1n08x5 _32819_ (.a(net686),
    .b(_07302_),
    .c(_07304_),
    .o1(_07305_));
 b15and002al1n24x5 _32820_ (.a(net688),
    .b(net686),
    .o(_07306_));
 b15ztpn00an1n08x5 PHY_36 ();
 b15nand03an1n04x5 _32822_ (.a(net675),
    .b(\us22.a[6] ),
    .c(_06914_),
    .o1(_07308_));
 b15nonb02ar1n16x5 _32823_ (.a(net669),
    .b(\us22.a[5] ),
    .out0(_07309_));
 b15nonb02as1n06x5 _32824_ (.a(net673),
    .b(net669),
    .out0(_07310_));
 b15aoi022ar1n08x5 _32825_ (.a(net687),
    .b(_07309_),
    .c(_07310_),
    .d(_06761_),
    .o1(_07311_));
 b15oai022ah1n08x5 _32826_ (.a(_06913_),
    .b(_07306_),
    .c(_07308_),
    .d(_07311_),
    .o1(_07312_));
 b15norp03ar1n08x5 _32827_ (.a(_06868_),
    .b(_07305_),
    .c(_07312_),
    .o1(_07313_));
 b15ztpn00an1n08x5 PHY_35 ();
 b15nor004ah1n02x5 _32829_ (.a(net676),
    .b(net671),
    .c(net680),
    .d(\us22.a[3] ),
    .o1(_07316_));
 b15nonb02al1n04x5 _32830_ (.a(net680),
    .b(net670),
    .out0(_07317_));
 b15aoi013ar1n06x5 _32831_ (.a(_07316_),
    .b(_07317_),
    .c(_06927_),
    .d(net676),
    .o1(_07318_));
 b15inv040as1n12x5 _32832_ (.a(net674),
    .o1(_07319_));
 b15oai122an1n16x5 _32833_ (.a(\us22.a[1] ),
    .b(_06945_),
    .c(_06786_),
    .d(_07318_),
    .e(_07319_),
    .o1(_07320_));
 b15nand02ar1n02x5 _32834_ (.a(_06844_),
    .b(_06955_),
    .o1(_07321_));
 b15aoi012al1n02x5 _32835_ (.a(net680),
    .b(_06862_),
    .c(_07321_),
    .o1(_07322_));
 b15ztpn00an1n08x5 PHY_34 ();
 b15nor003ar1n02x5 _32837_ (.a(_06758_),
    .b(\us22.a[3] ),
    .c(_06769_),
    .o1(_07324_));
 b15oai013an1n04x5 _32838_ (.a(_07320_),
    .b(_07322_),
    .c(_07324_),
    .d(net685),
    .o1(_07326_));
 b15nand04as1n08x5 _32839_ (.a(_07295_),
    .b(_07301_),
    .c(_07313_),
    .d(_07326_),
    .o1(_07327_));
 b15norp03ar1n02x5 _32840_ (.a(net685),
    .b(_06826_),
    .c(_06844_),
    .o1(_07328_));
 b15nor002ar1n24x5 _32841_ (.a(net676),
    .b(net670),
    .o1(_07329_));
 b15oai112an1n08x5 _32842_ (.a(net671),
    .b(_07329_),
    .c(\us22.a[3] ),
    .d(_07319_),
    .o1(_07330_));
 b15aoi112ar1n02x5 _32843_ (.a(net689),
    .b(_07328_),
    .c(_07330_),
    .d(net685),
    .o1(_07331_));
 b15nandp3al1n04x5 _32844_ (.a(_06792_),
    .b(_06852_),
    .c(_06839_),
    .o1(_07332_));
 b15nand03al1n03x5 _32845_ (.a(net685),
    .b(net677),
    .c(_06844_),
    .o1(_07333_));
 b15aoi012ar1n04x5 _32846_ (.a(_06786_),
    .b(_07332_),
    .c(_07333_),
    .o1(_07334_));
 b15norp03aq1n02x5 _32847_ (.a(_06758_),
    .b(_07331_),
    .c(_07334_),
    .o1(_07335_));
 b15ztpn00an1n08x5 PHY_33 ();
 b15nandp2al1n24x5 _32849_ (.a(\us22.a[1] ),
    .b(\us22.a[3] ),
    .o1(_07338_));
 b15nonb02aq1n03x5 _32850_ (.a(net676),
    .b(\us22.a[3] ),
    .out0(_07339_));
 b15oai022ar1n04x5 _32851_ (.a(net676),
    .b(_07338_),
    .c(_07339_),
    .d(net674),
    .o1(_07340_));
 b15aoi012ar1n02x5 _32852_ (.a(_06955_),
    .b(_07306_),
    .c(_07330_),
    .o1(_07341_));
 b15oai112ar1n08x5 _32853_ (.a(_06852_),
    .b(_07340_),
    .c(_07341_),
    .d(net680),
    .o1(_07342_));
 b15nor002aq1n04x5 _32854_ (.a(_07335_),
    .b(_07342_),
    .o1(_07343_));
 b15nona23al1n32x5 _32855_ (.a(net675),
    .b(net669),
    .c(net672),
    .d(net673),
    .out0(_07344_));
 b15aoi012as1n02x5 _32856_ (.a(net678),
    .b(_06904_),
    .c(_07344_),
    .o1(_07345_));
 b15aoai13al1n04x5 _32857_ (.a(net688),
    .b(_07291_),
    .c(_07344_),
    .d(_06758_),
    .o1(_07346_));
 b15oab012ar1n12x5 _32858_ (.c(net688),
    .a(net682),
    .b(net686),
    .out0(_07348_));
 b15oai112ah1n12x5 _32859_ (.a(_07345_),
    .b(_07346_),
    .c(_06866_),
    .d(_07348_),
    .o1(_07349_));
 b15nand03ah1n04x5 _32860_ (.a(\us22.a[5] ),
    .b(\us22.a[2] ),
    .c(\us22.a[3] ),
    .o1(_07350_));
 b15nona23ar1n08x5 _32861_ (.a(\us22.a[4] ),
    .b(\us22.a[1] ),
    .c(\us22.a[6] ),
    .d(net670),
    .out0(_07351_));
 b15nona23ar1n08x5 _32862_ (.a(net670),
    .b(\us22.a[6] ),
    .c(\us22.a[1] ),
    .d(\us22.a[4] ),
    .out0(_07352_));
 b15aoi112as1n08x5 _32863_ (.a(net690),
    .b(_07350_),
    .c(_07351_),
    .d(_07352_),
    .o1(_07353_));
 b15nand03as1n16x5 _32864_ (.a(\us22.a[1] ),
    .b(net680),
    .c(\us22.a[3] ),
    .o1(_07354_));
 b15norp03as1n04x5 _32865_ (.a(_06936_),
    .b(_06783_),
    .c(_07354_),
    .o1(_07355_));
 b15orn002ah1n12x5 _32866_ (.a(net683),
    .b(net679),
    .o(_07356_));
 b15nor003ar1n06x5 _32867_ (.a(_06933_),
    .b(_07356_),
    .c(_06969_),
    .o1(_07357_));
 b15oaoi13as1n08x5 _32868_ (.a(_07353_),
    .b(net690),
    .c(_07355_),
    .d(_07357_),
    .o1(_07359_));
 b15nand02ar1n02x5 _32869_ (.a(net683),
    .b(_06940_),
    .o1(_07360_));
 b15norp02ah1n24x5 _32870_ (.a(net687),
    .b(\us22.a[3] ),
    .o1(_07361_));
 b15oaoi13an1n03x5 _32871_ (.a(_06786_),
    .b(_06977_),
    .c(_07361_),
    .d(_06912_),
    .o1(_07362_));
 b15nonb03as1n12x5 _32872_ (.a(net686),
    .b(net682),
    .c(net679),
    .out0(_07363_));
 b15nano23aq1n24x5 _32873_ (.a(net675),
    .b(net669),
    .c(net672),
    .d(net673),
    .out0(_07364_));
 b15nonb02an1n08x5 _32874_ (.a(\us22.a[7] ),
    .b(\us22.a[1] ),
    .out0(_07365_));
 b15nor002aq1n08x5 _32875_ (.a(_06783_),
    .b(_07365_),
    .o1(_07366_));
 b15nano22an1n08x5 _32876_ (.a(net672),
    .b(net683),
    .c(net679),
    .out0(_07367_));
 b15aoi022ar1n02x5 _32877_ (.a(_07363_),
    .b(_07364_),
    .c(_07366_),
    .d(_07367_),
    .o1(_07368_));
 b15nanb02al1n02x5 _32878_ (.a(net673),
    .b(net669),
    .out0(_07370_));
 b15nor004ar1n03x5 _32879_ (.a(net675),
    .b(_07356_),
    .c(_06954_),
    .d(_07370_),
    .o1(_07371_));
 b15nano23as1n24x5 _32880_ (.a(net669),
    .b(net672),
    .c(net673),
    .d(net675),
    .out0(_07372_));
 b15aoi112al1n02x5 _32881_ (.a(net688),
    .b(_07371_),
    .c(_07372_),
    .d(_06889_),
    .o1(_07373_));
 b15ao0022an1n04x5 _32882_ (.a(_07360_),
    .b(_07362_),
    .c(_07368_),
    .d(_07373_),
    .o(_07374_));
 b15orn003an1n02x5 _32883_ (.a(_06954_),
    .b(_06838_),
    .c(_07370_),
    .o(_07375_));
 b15nand02an1n04x5 _32884_ (.a(net672),
    .b(_07310_),
    .o1(_07376_));
 b15nanb02aq1n24x5 _32885_ (.a(net682),
    .b(net679),
    .out0(_07377_));
 b15nonb02aq1n12x5 _32886_ (.a(net686),
    .b(net688),
    .out0(_07378_));
 b15nor002ah1n04x5 _32887_ (.a(_06911_),
    .b(_07378_),
    .o1(_07379_));
 b15oai013as1n08x5 _32888_ (.a(_07375_),
    .b(_07376_),
    .c(_07377_),
    .d(_07379_),
    .o1(_07381_));
 b15oai012aq1n03x5 _32889_ (.a(_06756_),
    .b(_06904_),
    .c(net689),
    .o1(_07382_));
 b15oai112al1n12x5 _32890_ (.a(_06826_),
    .b(_07382_),
    .c(_06769_),
    .d(net689),
    .o1(_07383_));
 b15nandp2aq1n16x5 _32891_ (.a(_06777_),
    .b(_06896_),
    .o1(_07384_));
 b15oai122al1n16x5 _32892_ (.a(net678),
    .b(_06859_),
    .c(_07384_),
    .d(_06973_),
    .e(_06748_),
    .o1(_07385_));
 b15aoi012al1n02x5 _32893_ (.a(net686),
    .b(net682),
    .c(_06866_),
    .o1(_07386_));
 b15nand02as1n12x5 _32894_ (.a(_06839_),
    .b(_06767_),
    .o1(_07387_));
 b15oaoi13an1n04x5 _32895_ (.a(_07386_),
    .b(_07387_),
    .c(_06966_),
    .d(_07269_),
    .o1(_07388_));
 b15aoi222an1n12x5 _32896_ (.a(net675),
    .b(_07381_),
    .c(_07383_),
    .d(_07385_),
    .e(_07388_),
    .f(net678),
    .o1(_07389_));
 b15nand04aq1n16x5 _32897_ (.a(_07349_),
    .b(_07359_),
    .c(_07374_),
    .d(_07389_),
    .o1(_07390_));
 b15nor004as1n12x5 _32898_ (.a(_07286_),
    .b(_07327_),
    .c(_07343_),
    .d(_07390_),
    .o1(_07392_));
 b15xor002an1n12x5 _32899_ (.a(_07267_),
    .b(_07392_),
    .out0(_07393_));
 b15nor004ah1n04x5 _32900_ (.a(net930),
    .b(net927),
    .c(_05934_),
    .d(_05935_),
    .o1(_07394_));
 b15aoai13ar1n04x5 _32901_ (.a(net933),
    .b(_07394_),
    .c(_06000_),
    .d(_06072_),
    .o1(_07395_));
 b15oai013as1n03x5 _32902_ (.a(_07395_),
    .b(_06067_),
    .c(_06019_),
    .d(net933),
    .o1(_07396_));
 b15nandp2ah1n05x5 _32903_ (.a(net918),
    .b(_05975_),
    .o1(_07397_));
 b15aoi012al1n02x5 _32904_ (.a(_05946_),
    .b(_06434_),
    .c(_06044_),
    .o1(_07398_));
 b15nonb02ar1n08x5 _32905_ (.a(\us00.a[2] ),
    .b(\us00.a[7] ),
    .out0(_07399_));
 b15aoi112aq1n03x5 _32906_ (.a(_07397_),
    .b(_07398_),
    .c(_06014_),
    .d(_07399_),
    .o1(_07400_));
 b15norp03ar1n02x5 _32907_ (.a(\us00.a[5] ),
    .b(\us00.a[4] ),
    .c(net918),
    .o1(_07401_));
 b15aoi013an1n02x5 _32908_ (.a(_07401_),
    .b(_06453_),
    .c(_05840_),
    .d(net918),
    .o1(_07403_));
 b15oai013ar1n02x5 _32909_ (.a(_06033_),
    .b(_07403_),
    .c(\us00.a[7] ),
    .d(_05821_),
    .o1(_07404_));
 b15nand03al1n04x5 _32910_ (.a(\us00.a[5] ),
    .b(net923),
    .c(\us00.a[7] ),
    .o1(_07405_));
 b15nandp3ar1n02x5 _32911_ (.a(net918),
    .b(\us00.a[1] ),
    .c(_06434_),
    .o1(_07406_));
 b15oaoi13ar1n02x5 _32912_ (.a(_07405_),
    .b(_07406_),
    .c(_06382_),
    .d(net918),
    .o1(_07407_));
 b15orn003ar1n02x5 _32913_ (.a(_07400_),
    .b(_07404_),
    .c(_07407_),
    .o(_07408_));
 b15oai012ar1n04x5 _32914_ (.a(\us00.a[3] ),
    .b(_07396_),
    .c(_07408_),
    .o1(_07409_));
 b15norp02aq1n08x5 _32915_ (.a(\us00.a[2] ),
    .b(_05959_),
    .o1(_07410_));
 b15nor003ar1n08x5 _32916_ (.a(_05918_),
    .b(_05934_),
    .c(_05935_),
    .o1(_07411_));
 b15oai012ar1n03x5 _32917_ (.a(_06056_),
    .b(_07410_),
    .c(_07411_),
    .o1(_07412_));
 b15nanb02ar1n02x5 _32918_ (.a(net927),
    .b(\us00.a[5] ),
    .out0(_07414_));
 b15oai012ar1n02x5 _32919_ (.a(_07414_),
    .b(_05990_),
    .c(\us00.a[5] ),
    .o1(_07415_));
 b15nand04aq1n03x5 _32920_ (.a(\us00.a[6] ),
    .b(\us00.a[0] ),
    .c(_06009_),
    .d(_07415_),
    .o1(_07416_));
 b15aboi22ah1n04x5 _32921_ (.a(_07400_),
    .b(net924),
    .c(_07412_),
    .d(_07416_),
    .out0(_07417_));
 b15aoai13ah1n03x5 _32922_ (.a(net935),
    .b(_06072_),
    .c(_05829_),
    .d(_05821_),
    .o1(_07418_));
 b15nonb03al1n08x5 _32923_ (.a(net929),
    .b(net926),
    .c(net932),
    .out0(_07419_));
 b15nor002ah1n02x5 _32924_ (.a(_05925_),
    .b(_05846_),
    .o1(_07420_));
 b15nor002as1n03x5 _32925_ (.a(_07419_),
    .b(_07420_),
    .o1(_07421_));
 b15aoi012aq1n06x5 _32926_ (.a(_06405_),
    .b(_07418_),
    .c(_07421_),
    .o1(_07422_));
 b15aoai13ar1n02x5 _32927_ (.a(\us00.a[3] ),
    .b(_05882_),
    .c(_05932_),
    .d(net927),
    .o1(_07423_));
 b15oai012ar1n02x5 _32928_ (.a(_05932_),
    .b(_06014_),
    .c(_05918_),
    .o1(_07425_));
 b15oaoi13ar1n03x5 _32929_ (.a(_07423_),
    .b(_07425_),
    .c(_05891_),
    .d(_05918_),
    .o1(_07426_));
 b15orn002al1n08x5 _32930_ (.a(_06034_),
    .b(_05987_),
    .o(_07427_));
 b15nano22ar1n02x5 _32931_ (.a(net931),
    .b(net925),
    .c(net915),
    .out0(_07428_));
 b15nonb03as1n03x5 _32932_ (.a(net922),
    .b(net917),
    .c(net919),
    .out0(_07429_));
 b15aoai13al1n02x5 _32933_ (.a(_07428_),
    .b(_07429_),
    .c(_05867_),
    .d(net917),
    .o1(_07430_));
 b15aoi012ar1n02x5 _32934_ (.a(net934),
    .b(_07427_),
    .c(_07430_),
    .o1(_07431_));
 b15nonb03al1n08x5 _32935_ (.a(net919),
    .b(net915),
    .c(net917),
    .out0(_07432_));
 b15nand02ar1n02x5 _32936_ (.a(_05821_),
    .b(_07432_),
    .o1(_07433_));
 b15nand02ar1n02x5 _32937_ (.a(net922),
    .b(_05829_),
    .o1(_07434_));
 b15oaoi13ar1n03x5 _32938_ (.a(_07433_),
    .b(_07434_),
    .c(_05835_),
    .d(net922),
    .o1(_07436_));
 b15nonb02aq1n03x5 _32939_ (.a(net935),
    .b(net926),
    .out0(_07437_));
 b15oai012ar1n04x5 _32940_ (.a(_07437_),
    .b(net929),
    .c(net922),
    .o1(_07438_));
 b15nor004ah1n04x5 _32941_ (.a(net920),
    .b(_06072_),
    .c(_05929_),
    .d(_07438_),
    .o1(_07439_));
 b15orn003al1n08x5 _32942_ (.a(_07431_),
    .b(_07436_),
    .c(_07439_),
    .o(_07440_));
 b15nor004ah1n03x5 _32943_ (.a(_07417_),
    .b(_07422_),
    .c(_07426_),
    .d(_07440_),
    .o1(_07441_));
 b15mdn022an1n04x5 _32944_ (.a(_05959_),
    .b(_06078_),
    .o1(_07442_),
    .sa(net925));
 b15nand02ar1n02x5 _32945_ (.a(net928),
    .b(_06050_),
    .o1(_07443_));
 b15aob012ar1n03x5 _32946_ (.a(net934),
    .b(_05893_),
    .c(_07443_),
    .out0(_07444_));
 b15aoi012aq1n02x5 _32947_ (.a(_06049_),
    .b(_05895_),
    .c(net931),
    .o1(_07445_));
 b15oai112al1n08x5 _32948_ (.a(_07442_),
    .b(_07444_),
    .c(_07445_),
    .d(net934),
    .o1(_07447_));
 b15nand02ah1n24x5 _32949_ (.a(_05867_),
    .b(_06003_),
    .o1(_07448_));
 b15oai022al1n12x5 _32950_ (.a(_06397_),
    .b(_07448_),
    .c(_05896_),
    .d(_05899_),
    .o1(_07449_));
 b15nonb02aq1n12x5 _32951_ (.a(net929),
    .b(net932),
    .out0(_07450_));
 b15nor002aq1n12x5 _32952_ (.a(net935),
    .b(net926),
    .o1(_07451_));
 b15nona23ar1n04x5 _32953_ (.a(_07450_),
    .b(_06367_),
    .c(_07451_),
    .d(_06365_),
    .out0(_07452_));
 b15oaoi13an1n04x5 _32954_ (.a(_07452_),
    .b(net918),
    .c(net923),
    .d(_05918_),
    .o1(_07453_));
 b15norp03ar1n04x5 _32955_ (.a(net923),
    .b(net918),
    .c(net929),
    .o1(_07454_));
 b15nor004aq1n04x5 _32956_ (.a(net920),
    .b(net916),
    .c(net935),
    .d(\us00.a[3] ),
    .o1(_07455_));
 b15and003an1n02x5 _32957_ (.a(net920),
    .b(net916),
    .c(\us00.a[3] ),
    .o(_07456_));
 b15oai112an1n12x5 _32958_ (.a(_05925_),
    .b(_07454_),
    .c(_07455_),
    .d(_07456_),
    .o1(_07458_));
 b15aoi012al1n02x5 _32959_ (.a(_05860_),
    .b(_05975_),
    .c(net935),
    .o1(_07459_));
 b15nand03aq1n02x5 _32960_ (.a(net932),
    .b(_05906_),
    .c(_05844_),
    .o1(_07460_));
 b15oai012an1n06x5 _32961_ (.a(_07458_),
    .b(_07459_),
    .c(_07460_),
    .o1(_07461_));
 b15oai012ar1n06x5 _32962_ (.a(_07419_),
    .b(_06046_),
    .c(_05827_),
    .o1(_07462_));
 b15nano23ah1n06x5 _32963_ (.a(net920),
    .b(net923),
    .c(net916),
    .d(net918),
    .out0(_07463_));
 b15oai112as1n08x5 _32964_ (.a(net935),
    .b(_07463_),
    .c(_05829_),
    .d(_05906_),
    .o1(_07464_));
 b15nanb02as1n24x5 _32965_ (.a(net928),
    .b(net931),
    .out0(_07465_));
 b15aoi022an1n06x5 _32966_ (.a(_06072_),
    .b(_06388_),
    .c(_06390_),
    .d(_07465_),
    .o1(_07466_));
 b15nandp2al1n03x5 _32967_ (.a(net916),
    .b(_05955_),
    .o1(_07467_));
 b15oai112al1n12x5 _32968_ (.a(_07462_),
    .b(_07464_),
    .c(_07466_),
    .d(_07467_),
    .o1(_07469_));
 b15nor004al1n12x5 _32969_ (.a(_07449_),
    .b(_07453_),
    .c(_07461_),
    .d(_07469_),
    .o1(_07470_));
 b15nona23ar1n02x5 _32970_ (.a(net915),
    .b(net917),
    .c(net925),
    .d(net922),
    .out0(_07471_));
 b15nanb03an1n06x5 _32971_ (.a(net922),
    .b(net915),
    .c(net917),
    .out0(_07472_));
 b15nanb02as1n06x5 _32972_ (.a(net925),
    .b(net934),
    .out0(_07473_));
 b15oaoi13as1n02x5 _32973_ (.a(net919),
    .b(_07471_),
    .c(_07472_),
    .d(_07473_),
    .o1(_07474_));
 b15norp02as1n03x5 _32974_ (.a(_05911_),
    .b(_06078_),
    .o1(_07475_));
 b15oai012ar1n08x5 _32975_ (.a(_06076_),
    .b(_07474_),
    .c(_07475_),
    .o1(_07476_));
 b15nor003aq1n02x5 _32976_ (.a(net934),
    .b(_05928_),
    .c(_05854_),
    .o1(_07477_));
 b15aoi012al1n02x5 _32977_ (.a(_05972_),
    .b(_06044_),
    .c(_07465_),
    .o1(_07478_));
 b15oai012al1n06x5 _32978_ (.a(_05911_),
    .b(_07477_),
    .c(_07478_),
    .o1(_07480_));
 b15nor002aq1n02x5 _32979_ (.a(net918),
    .b(_05884_),
    .o1(_07481_));
 b15nor002aq1n03x5 _32980_ (.a(_06056_),
    .b(_06386_),
    .o1(_07482_));
 b15aoai13as1n08x5 _32981_ (.a(_07481_),
    .b(_06457_),
    .c(net923),
    .d(_07482_),
    .o1(_07483_));
 b15norp02aq1n02x5 _32982_ (.a(net925),
    .b(_06037_),
    .o1(_07484_));
 b15nor004as1n02x5 _32983_ (.a(_05967_),
    .b(_06056_),
    .c(_05935_),
    .d(_05851_),
    .o1(_07485_));
 b15oai112as1n06x5 _32984_ (.a(_06463_),
    .b(_06038_),
    .c(_07484_),
    .d(_07485_),
    .o1(_07486_));
 b15nand04ah1n12x5 _32985_ (.a(_07476_),
    .b(_07480_),
    .c(_07483_),
    .d(_07486_),
    .o1(_07487_));
 b15oai012al1n06x5 _32986_ (.a(_06060_),
    .b(_06468_),
    .c(_06081_),
    .o1(_07488_));
 b15aoi012al1n08x5 _32987_ (.a(net925),
    .b(_06435_),
    .c(_07488_),
    .o1(_07489_));
 b15nano23ar1n12x5 _32988_ (.a(_07447_),
    .b(_07470_),
    .c(_07487_),
    .d(_07489_),
    .out0(_07491_));
 b15and003as1n12x5 _32989_ (.a(_07409_),
    .b(_07441_),
    .c(_07491_),
    .o(_07492_));
 b15xor002as1n02x5 _32990_ (.a(_07393_),
    .b(_07492_),
    .out0(_07493_));
 b15xor003aq1n02x5 _32991_ (.a(_06354_),
    .b(_07126_),
    .c(_07493_),
    .out0(_07494_));
 b15cmbn22as1n04x5 _32992_ (.clk1(\text_in_r[97] ),
    .clk2(_07494_),
    .clkout(_07495_),
    .s(net536));
 b15xor002an1n12x5 _32993_ (.a(net532),
    .b(_07495_),
    .out0(_00098_));
 b15ztpn00an1n08x5 PHY_32 ();
 b15aoi012ar1n02x5 _32995_ (.a(_06839_),
    .b(_06777_),
    .c(_06792_),
    .o1(_07497_));
 b15oai013an1n03x5 _32996_ (.a(net680),
    .b(\us22.a[3] ),
    .c(_06936_),
    .d(_07497_),
    .o1(_07498_));
 b15ztpn00an1n08x5 PHY_31 ();
 b15oai112ar1n04x5 _32998_ (.a(net670),
    .b(_06768_),
    .c(_06792_),
    .d(net671),
    .o1(_07501_));
 b15oai022al1n02x5 _32999_ (.a(\us22.a[1] ),
    .b(_06981_),
    .c(_07501_),
    .d(_06786_),
    .o1(_07502_));
 b15aoi012aq1n04x5 _33000_ (.a(_07498_),
    .b(_07502_),
    .c(\us22.a[3] ),
    .o1(_07503_));
 b15nonb02as1n03x5 _33001_ (.a(net690),
    .b(\us22.a[3] ),
    .out0(_07504_));
 b15nandp3ar1n02x5 _33002_ (.a(\us22.a[1] ),
    .b(_06844_),
    .c(_07504_),
    .o1(_07505_));
 b15aob012al1n02x5 _33003_ (.a(_07505_),
    .b(_06940_),
    .c(_06792_),
    .out0(_07506_));
 b15oab012ar1n12x5 _33004_ (.c(net680),
    .a(_07503_),
    .b(_07506_),
    .out0(_07507_));
 b15nona22aq1n12x5 _33005_ (.a(net688),
    .b(net686),
    .c(net682),
    .out0(_07508_));
 b15nand04ah1n04x5 _33006_ (.a(net673),
    .b(_06999_),
    .c(_06826_),
    .d(_07508_),
    .o1(_07509_));
 b15oai012an1n04x5 _33007_ (.a(net682),
    .b(_06977_),
    .c(_06786_),
    .o1(_07510_));
 b15nanb02ar1n24x5 _33008_ (.a(net669),
    .b(net675),
    .out0(_07512_));
 b15nand02aq1n02x5 _33009_ (.a(net683),
    .b(_07288_),
    .o1(_07513_));
 b15aoi122as1n04x5 _33010_ (.a(_07509_),
    .b(_07510_),
    .c(net686),
    .d(_07512_),
    .e(_07513_),
    .o1(_07514_));
 b15nor003ar1n08x5 _33011_ (.a(_06786_),
    .b(_06954_),
    .c(_07512_),
    .o1(_07515_));
 b15nand02al1n02x5 _33012_ (.a(net673),
    .b(net679),
    .o1(_07516_));
 b15oai012an1n06x5 _33013_ (.a(_07516_),
    .b(_06869_),
    .c(net673),
    .o1(_07517_));
 b15nandp2al1n08x5 _33014_ (.a(net683),
    .b(net677),
    .o1(_07518_));
 b15oai022ah1n08x5 _33015_ (.a(_06906_),
    .b(_07518_),
    .c(_06990_),
    .d(_07387_),
    .o1(_07519_));
 b15aoi122ah1n08x5 _33016_ (.a(_07514_),
    .b(_07515_),
    .c(_07517_),
    .d(_07519_),
    .e(_06786_),
    .o1(_07520_));
 b15nanb02al1n06x5 _33017_ (.a(\us22.a[5] ),
    .b(net687),
    .out0(_07521_));
 b15and002al1n12x5 _33018_ (.a(\us22.a[4] ),
    .b(net670),
    .o(_07523_));
 b15nandp2aq1n02x5 _33019_ (.a(_07523_),
    .b(_07367_),
    .o1(_07524_));
 b15aoi022ah1n08x5 _33020_ (.a(_06767_),
    .b(_06914_),
    .c(_06896_),
    .d(_06912_),
    .o1(_07525_));
 b15oaoi13as1n08x5 _33021_ (.a(_07521_),
    .b(_07524_),
    .c(_07525_),
    .d(net675),
    .o1(_07526_));
 b15oai012as1n03x5 _33022_ (.a(net683),
    .b(net678),
    .c(_06906_),
    .o1(_07527_));
 b15oai012ah1n04x5 _33023_ (.a(_06906_),
    .b(_06761_),
    .c(_06981_),
    .o1(_07528_));
 b15nor002an1n03x5 _33024_ (.a(_06849_),
    .b(_07306_),
    .o1(_07529_));
 b15aoi013ah1n06x5 _33025_ (.a(_07526_),
    .b(_07527_),
    .c(_07528_),
    .d(_07529_),
    .o1(_07530_));
 b15nanb02al1n06x5 _33026_ (.a(\us22.a[6] ),
    .b(net673),
    .out0(_07531_));
 b15oai022ar1n02x5 _33027_ (.a(_07531_),
    .b(_06837_),
    .c(_07287_),
    .d(net673),
    .o1(_07532_));
 b15nandp3al1n04x5 _33028_ (.a(net686),
    .b(_07288_),
    .c(_07532_),
    .o1(_07534_));
 b15nor003an1n12x5 _33029_ (.a(net689),
    .b(net684),
    .c(net681),
    .o1(_07535_));
 b15oai112ar1n02x5 _33030_ (.a(net678),
    .b(_06756_),
    .c(_06966_),
    .d(_07535_),
    .o1(_07536_));
 b15oai013an1n02x5 _33031_ (.a(_06851_),
    .b(_07377_),
    .c(_06769_),
    .d(_07306_),
    .o1(_07537_));
 b15nandp2an1n03x5 _33032_ (.a(_07363_),
    .b(_07364_),
    .o1(_07538_));
 b15nandp3ah1n03x5 _33033_ (.a(_06866_),
    .b(_07378_),
    .c(_06912_),
    .o1(_07539_));
 b15nand02aq1n04x5 _33034_ (.a(net678),
    .b(_06915_),
    .o1(_07540_));
 b15oai112al1n16x5 _33035_ (.a(_07538_),
    .b(_07539_),
    .c(_06975_),
    .d(_07540_),
    .o1(_07541_));
 b15nano23aq1n05x5 _33036_ (.a(_07534_),
    .b(_07536_),
    .c(_07537_),
    .d(_07541_),
    .out0(_07542_));
 b15aoi013an1n02x5 _33037_ (.a(_06826_),
    .b(_06822_),
    .c(_06859_),
    .d(_06839_),
    .o1(_07543_));
 b15nandp2ah1n16x5 _33038_ (.a(_06777_),
    .b(_06852_),
    .o1(_07545_));
 b15norp02as1n24x5 _33039_ (.a(net687),
    .b(net683),
    .o1(_07546_));
 b15oaoi13an1n04x5 _33040_ (.a(_07543_),
    .b(_06878_),
    .c(_07545_),
    .d(_07546_),
    .o1(_07547_));
 b15oai012ah1n04x5 _33041_ (.a(_06786_),
    .b(_07363_),
    .c(_06878_),
    .o1(_07548_));
 b15oai112as1n04x5 _33042_ (.a(net684),
    .b(_07279_),
    .c(_06869_),
    .d(net689),
    .o1(_07549_));
 b15aoi012as1n02x5 _33043_ (.a(_07269_),
    .b(_07377_),
    .c(_06792_),
    .o1(_07550_));
 b15aoi022ah1n08x5 _33044_ (.a(_07547_),
    .b(_07548_),
    .c(_07549_),
    .d(_07550_),
    .o1(_07551_));
 b15nand04ah1n16x5 _33045_ (.a(_07520_),
    .b(_07530_),
    .c(_07542_),
    .d(_07551_),
    .o1(_07552_));
 b15nand03an1n16x5 _33046_ (.a(net689),
    .b(net679),
    .c(_07372_),
    .o1(_07553_));
 b15aoi013ar1n02x5 _33047_ (.a(net684),
    .b(_06849_),
    .c(_06924_),
    .d(_06786_),
    .o1(_07554_));
 b15nand02aq1n04x5 _33048_ (.a(_07553_),
    .b(_07554_),
    .o1(_07556_));
 b15nand03ar1n06x5 _33049_ (.a(_06786_),
    .b(_06912_),
    .c(_06844_),
    .o1(_07557_));
 b15oai112ar1n12x5 _33050_ (.a(net684),
    .b(_07557_),
    .c(_06981_),
    .d(_06869_),
    .o1(_07558_));
 b15aoi012ar1n02x5 _33051_ (.a(_06786_),
    .b(_06800_),
    .c(_06863_),
    .o1(_07559_));
 b15oai013an1n04x5 _33052_ (.a(net679),
    .b(_07282_),
    .c(_07559_),
    .d(_07535_),
    .o1(_07560_));
 b15aoi112ar1n02x5 _33053_ (.a(net689),
    .b(_06863_),
    .c(_06823_),
    .d(_06896_),
    .o1(_07561_));
 b15nand03ar1n03x5 _33054_ (.a(_06869_),
    .b(_06823_),
    .c(_06896_),
    .o1(_07562_));
 b15oaoi13aq1n03x5 _33055_ (.a(_07561_),
    .b(_06769_),
    .c(_07562_),
    .d(_07535_),
    .o1(_07563_));
 b15aoi022aq1n12x5 _33056_ (.a(_07556_),
    .b(_07558_),
    .c(_07560_),
    .d(_07563_),
    .o1(_07564_));
 b15oai022an1n02x5 _33057_ (.a(_06867_),
    .b(_06790_),
    .c(_06769_),
    .d(_07354_),
    .o1(_07565_));
 b15nandp3ar1n02x5 _33058_ (.a(_06826_),
    .b(_06863_),
    .c(_06768_),
    .o1(_07567_));
 b15oaoi13as1n02x5 _33059_ (.a(_06969_),
    .b(_07567_),
    .c(_06984_),
    .d(_07518_),
    .o1(_07568_));
 b15oai012an1n06x5 _33060_ (.a(net689),
    .b(_07565_),
    .c(_07568_),
    .o1(_07569_));
 b15aoi012an1n02x5 _33061_ (.a(_06786_),
    .b(_06863_),
    .c(_07518_),
    .o1(_07570_));
 b15aoai13aq1n06x5 _33062_ (.a(_06924_),
    .b(_07570_),
    .c(_06912_),
    .d(net684),
    .o1(_07571_));
 b15aoi112al1n02x5 _33063_ (.a(_06826_),
    .b(_06824_),
    .c(_07279_),
    .d(net684),
    .o1(_07572_));
 b15aoi013aq1n04x5 _33064_ (.a(_07572_),
    .b(_06986_),
    .c(_06813_),
    .d(net683),
    .o1(_07573_));
 b15nand04al1n16x5 _33065_ (.a(_07564_),
    .b(_07569_),
    .c(_07571_),
    .d(_07573_),
    .o1(_07574_));
 b15aoi012ar1n02x5 _33066_ (.a(_07354_),
    .b(_06821_),
    .c(_06854_),
    .o1(_07575_));
 b15nandp2an1n12x5 _33067_ (.a(net677),
    .b(_06807_),
    .o1(_07576_));
 b15oai012ar1n03x5 _33068_ (.a(_07576_),
    .b(_06854_),
    .c(net677),
    .o1(_07578_));
 b15aoi013al1n03x5 _33069_ (.a(_07575_),
    .b(_07578_),
    .c(_06911_),
    .d(net680),
    .o1(_07579_));
 b15nandp2aq1n16x5 _33070_ (.a(_06786_),
    .b(_06792_),
    .o1(_07580_));
 b15norp03al1n08x5 _33071_ (.a(_07580_),
    .b(_06783_),
    .c(_06934_),
    .o1(_07581_));
 b15nor002ar1n06x5 _33072_ (.a(_06854_),
    .b(_06915_),
    .o1(_07582_));
 b15norp02ar1n02x5 _33073_ (.a(_06748_),
    .b(_07576_),
    .o1(_07583_));
 b15nor003an1n03x5 _33074_ (.a(_07581_),
    .b(_07582_),
    .c(_07583_),
    .o1(_07584_));
 b15oai012ar1n08x5 _33075_ (.a(_07579_),
    .b(_07584_),
    .c(net680),
    .o1(_07585_));
 b15nor004as1n12x5 _33076_ (.a(_07507_),
    .b(_07552_),
    .c(_07574_),
    .d(_07585_),
    .o1(_07586_));
 b15nandp2aq1n04x5 _33077_ (.a(net934),
    .b(_07442_),
    .o1(_07587_));
 b15nand02an1n03x5 _33078_ (.a(net925),
    .b(_05915_),
    .o1(_07589_));
 b15oai112aq1n06x5 _33079_ (.a(net928),
    .b(_07587_),
    .c(_07589_),
    .d(_05925_),
    .o1(_07590_));
 b15nanb03al1n04x5 _33080_ (.a(net920),
    .b(net916),
    .c(net926),
    .out0(_07591_));
 b15orn003ar1n02x5 _33081_ (.a(_05969_),
    .b(net926),
    .c(_06386_),
    .o(_07592_));
 b15aoi012ar1n02x5 _33082_ (.a(_06365_),
    .b(_07591_),
    .c(_07592_),
    .o1(_07593_));
 b15nand03ah1n06x5 _33083_ (.a(net925),
    .b(_05955_),
    .c(_05844_),
    .o1(_07594_));
 b15oaoi13an1n08x5 _33084_ (.a(_06044_),
    .b(_07594_),
    .c(net925),
    .d(_06037_),
    .o1(_07595_));
 b15norp03aq1n03x5 _33085_ (.a(net929),
    .b(_07593_),
    .c(_07595_),
    .o1(_07596_));
 b15nandp2ar1n05x5 _33086_ (.a(net918),
    .b(\us00.a[0] ),
    .o1(_07597_));
 b15and002ar1n02x5 _33087_ (.a(net916),
    .b(\us00.a[3] ),
    .o(_07598_));
 b15aoi022as1n06x5 _33088_ (.a(_05840_),
    .b(_07399_),
    .c(_07598_),
    .d(_05975_),
    .o1(_07600_));
 b15mdn022aq1n06x5 _33089_ (.a(_06032_),
    .b(_05827_),
    .o1(_07601_),
    .sa(\us00.a[3] ));
 b15oai222as1n16x5 _33090_ (.a(_05899_),
    .b(_05846_),
    .c(_07597_),
    .d(_07600_),
    .e(_07601_),
    .f(_05918_),
    .o1(_07602_));
 b15oai012aq1n02x5 _33091_ (.a(_06024_),
    .b(_07602_),
    .c(net932),
    .o1(_07603_));
 b15aob012ah1n03x5 _33092_ (.a(_07590_),
    .b(_07596_),
    .c(_07603_),
    .out0(_07604_));
 b15inv040ah1n10x5 _33093_ (.a(net919),
    .o1(_07605_));
 b15nand04ar1n02x5 _33094_ (.a(net922),
    .b(net915),
    .c(net918),
    .d(_05954_),
    .o1(_07606_));
 b15oai013ar1n02x5 _33095_ (.a(_07606_),
    .b(_05925_),
    .c(_05854_),
    .d(net922),
    .o1(_07607_));
 b15and003ar1n03x5 _33096_ (.a(_07605_),
    .b(_05947_),
    .c(_07607_),
    .o(_07608_));
 b15oaoi13aq1n04x5 _33097_ (.a(_06365_),
    .b(_07591_),
    .c(net926),
    .d(_06386_),
    .o1(_07609_));
 b15nano23ar1n02x5 _33098_ (.a(net923),
    .b(_06368_),
    .c(_05925_),
    .d(net918),
    .out0(_07611_));
 b15oai012al1n02x5 _33099_ (.a(_05906_),
    .b(_07609_),
    .c(_07611_),
    .o1(_07612_));
 b15aob012al1n04x5 _33100_ (.a(_07612_),
    .b(_07602_),
    .c(_05821_),
    .out0(_07613_));
 b15nor004an1n06x5 _33101_ (.a(_05821_),
    .b(_05934_),
    .c(_05966_),
    .d(_06424_),
    .o1(_07614_));
 b15aoai13ah1n08x5 _33102_ (.a(net925),
    .b(_07614_),
    .c(_06060_),
    .d(_06081_),
    .o1(_07615_));
 b15nanb02al1n06x5 _33103_ (.a(net920),
    .b(net915),
    .out0(_07616_));
 b15orn002al1n02x5 _33104_ (.a(net917),
    .b(net932),
    .o(_07617_));
 b15oai022an1n02x5 _33105_ (.a(_05904_),
    .b(_07616_),
    .c(_07617_),
    .d(_06386_),
    .o1(_07618_));
 b15nand04as1n06x5 _33106_ (.a(net922),
    .b(_05969_),
    .c(_05829_),
    .d(_07618_),
    .o1(_07619_));
 b15oai012ar1n02x5 _33107_ (.a(_05929_),
    .b(_05854_),
    .c(_05821_),
    .o1(_07620_));
 b15nandp3al1n02x5 _33108_ (.a(_05975_),
    .b(_05906_),
    .c(_07620_),
    .o1(_07622_));
 b15norp02ar1n08x5 _33109_ (.a(net926),
    .b(_05882_),
    .o1(_07623_));
 b15aoi222an1n06x5 _33110_ (.a(_05821_),
    .b(_07609_),
    .c(_07623_),
    .d(_05937_),
    .e(_06032_),
    .f(_07420_),
    .o1(_07624_));
 b15nand04aq1n06x5 _33111_ (.a(_07615_),
    .b(_07619_),
    .c(_07622_),
    .d(_07624_),
    .o1(_07625_));
 b15and003al1n02x5 _33112_ (.a(net921),
    .b(_06003_),
    .c(_06047_),
    .o(_07626_));
 b15oai112as1n06x5 _33113_ (.a(net919),
    .b(_05906_),
    .c(_05905_),
    .d(_07626_),
    .o1(_07627_));
 b15aoi012ah1n02x5 _33114_ (.a(net928),
    .b(_05925_),
    .c(_05915_),
    .o1(_07628_));
 b15oai112an1n06x5 _33115_ (.a(net925),
    .b(_06044_),
    .c(_06000_),
    .d(_05918_),
    .o1(_07629_));
 b15oai012as1n08x5 _33116_ (.a(_07627_),
    .b(_07628_),
    .c(_07629_),
    .o1(_07630_));
 b15nor004ar1n08x5 _33117_ (.a(_07608_),
    .b(_07613_),
    .c(_07625_),
    .d(_07630_),
    .o1(_07631_));
 b15nand03an1n06x5 _33118_ (.a(net931),
    .b(net926),
    .c(_07410_),
    .o1(_07633_));
 b15norp02ar1n08x5 _33119_ (.a(\us00.a[1] ),
    .b(\us00.a[3] ),
    .o1(_07634_));
 b15aoi012ar1n04x5 _33120_ (.a(\us00.a[0] ),
    .b(_05827_),
    .c(_07634_),
    .o1(_07635_));
 b15norp02ar1n32x5 _33121_ (.a(_05967_),
    .b(_05935_),
    .o1(_07636_));
 b15nano23ah1n12x5 _33122_ (.a(net920),
    .b(net915),
    .c(net918),
    .d(net923),
    .out0(_07637_));
 b15aoi022ar1n02x5 _33123_ (.a(_07636_),
    .b(_05851_),
    .c(_07637_),
    .d(_05894_),
    .o1(_07638_));
 b15oai112aq1n06x5 _33124_ (.a(_07633_),
    .b(_07635_),
    .c(_07638_),
    .d(_05947_),
    .o1(_07639_));
 b15nanb02ar1n02x5 _33125_ (.a(_05992_),
    .b(_07637_),
    .out0(_07640_));
 b15aoi022ar1n02x5 _33126_ (.a(_05911_),
    .b(_07636_),
    .c(_07637_),
    .d(net934),
    .o1(_07641_));
 b15oaoi13an1n03x5 _33127_ (.a(_05918_),
    .b(_07640_),
    .c(_07641_),
    .d(net932),
    .o1(_07642_));
 b15nandp3ar1n02x5 _33128_ (.a(_05975_),
    .b(_06003_),
    .c(_05895_),
    .o1(_07643_));
 b15oai013aq1n02x5 _33129_ (.a(_07643_),
    .b(_05846_),
    .c(_05841_),
    .d(net931),
    .o1(_07644_));
 b15ztpn00an1n08x5 PHY_30 ();
 b15nand02ar1n24x5 _33131_ (.a(_05955_),
    .b(_06003_),
    .o1(_07646_));
 b15oai012al1n02x5 _33132_ (.a(net934),
    .b(_06397_),
    .c(_07646_),
    .o1(_07647_));
 b15oai013as1n04x5 _33133_ (.a(_07639_),
    .b(_07642_),
    .c(_07644_),
    .d(_07647_),
    .o1(_07648_));
 b15oai012ah1n12x5 _33134_ (.a(_05911_),
    .b(_06044_),
    .c(_06078_),
    .o1(_07649_));
 b15nor003aq1n03x5 _33135_ (.a(net929),
    .b(_06386_),
    .c(_07617_),
    .o1(_07650_));
 b15xor002ar1n02x5 _33136_ (.a(net917),
    .b(net929),
    .out0(_07651_));
 b15norp03as1n03x5 _33137_ (.a(_05821_),
    .b(_07616_),
    .c(_07651_),
    .o1(_07652_));
 b15oaoi13al1n04x5 _33138_ (.a(_07649_),
    .b(net922),
    .c(_07650_),
    .d(_07652_),
    .o1(_07654_));
 b15oai012ar1n03x5 _33139_ (.a(net931),
    .b(_06468_),
    .c(_06424_),
    .o1(_07655_));
 b15nor003aq1n06x5 _33140_ (.a(net934),
    .b(net931),
    .c(net928),
    .o1(_07656_));
 b15oai022ah1n02x5 _33141_ (.a(_07450_),
    .b(_05854_),
    .c(_05929_),
    .d(_07656_),
    .o1(_07657_));
 b15nandp3as1n03x5 _33142_ (.a(_05867_),
    .b(_07655_),
    .c(_07657_),
    .o1(_07658_));
 b15oai122aq1n12x5 _33143_ (.a(_07429_),
    .b(_06424_),
    .c(_05821_),
    .d(net915),
    .e(_06463_),
    .o1(_07659_));
 b15norp02ar1n02x5 _33144_ (.a(net917),
    .b(_05935_),
    .o1(_07660_));
 b15xor002al1n02x5 _33145_ (.a(net915),
    .b(net934),
    .out0(_07661_));
 b15aoi013an1n03x5 _33146_ (.a(_05911_),
    .b(_07660_),
    .c(_07661_),
    .d(net929),
    .o1(_07662_));
 b15aoi013an1n06x5 _33147_ (.a(_07654_),
    .b(_07658_),
    .c(_07659_),
    .d(_07662_),
    .o1(_07663_));
 b15nor003ar1n02x5 _33148_ (.a(\us00.a[3] ),
    .b(_07465_),
    .c(_05921_),
    .o1(_07665_));
 b15nor002an1n03x5 _33149_ (.a(net932),
    .b(_05851_),
    .o1(_07666_));
 b15aoai13aq1n04x5 _33150_ (.a(net935),
    .b(_07665_),
    .c(_07666_),
    .d(_05915_),
    .o1(_07667_));
 b15nand02aq1n12x5 _33151_ (.a(net921),
    .b(net914),
    .o1(_07668_));
 b15norp02as1n04x5 _33152_ (.a(_05884_),
    .b(_07668_),
    .o1(_07669_));
 b15oai022ah1n12x5 _33153_ (.a(_05954_),
    .b(_06358_),
    .c(_05904_),
    .d(net920),
    .o1(_07670_));
 b15norp02as1n03x5 _33154_ (.a(_06019_),
    .b(_07473_),
    .o1(_07671_));
 b15aoi222as1n12x5 _33155_ (.a(_05983_),
    .b(_05927_),
    .c(_07669_),
    .d(_07670_),
    .e(_07671_),
    .f(_06026_),
    .o1(_07672_));
 b15norp02ar1n03x5 _33156_ (.a(_05921_),
    .b(_05942_),
    .o1(_07673_));
 b15aoi012ah1n04x5 _33157_ (.a(_07673_),
    .b(_05968_),
    .c(_05911_),
    .o1(_07674_));
 b15aoi012ar1n02x5 _33158_ (.a(net934),
    .b(_06397_),
    .c(_05851_),
    .o1(_07676_));
 b15oai112an1n02x5 _33159_ (.a(_07667_),
    .b(_07672_),
    .c(_07674_),
    .d(_07676_),
    .o1(_07677_));
 b15norp02ah1n04x5 _33160_ (.a(_07663_),
    .b(_07677_),
    .o1(_07678_));
 b15andc04as1n16x5 _33161_ (.a(_07604_),
    .b(_07631_),
    .c(_07648_),
    .d(_07678_),
    .o(_07679_));
 b15nand02aq1n16x5 _33162_ (.a(_06545_),
    .b(_06620_),
    .o1(_07680_));
 b15nonb02as1n03x5 _33163_ (.a(net799),
    .b(net803),
    .out0(_07681_));
 b15aoi022al1n08x5 _33164_ (.a(net803),
    .b(_07252_),
    .c(_07681_),
    .d(_06650_),
    .o1(_07682_));
 b15oai122an1n16x5 _33165_ (.a(_06476_),
    .b(_06605_),
    .c(_07680_),
    .d(_07682_),
    .e(_07186_),
    .o1(_07683_));
 b15oai012an1n06x5 _33166_ (.a(_06553_),
    .b(_06530_),
    .c(_07233_),
    .o1(_07684_));
 b15oaoi13an1n02x5 _33167_ (.a(net816),
    .b(_07684_),
    .c(_07161_),
    .d(_07258_),
    .o1(_07685_));
 b15nanb02al1n08x5 _33168_ (.a(net813),
    .b(net797),
    .out0(_07687_));
 b15nand03an1n08x5 _33169_ (.a(_06539_),
    .b(_07252_),
    .c(_07687_),
    .o1(_07688_));
 b15oai112aq1n02x5 _33170_ (.a(net819),
    .b(_07688_),
    .c(_06628_),
    .d(_06589_),
    .o1(_07689_));
 b15norp03an1n04x5 _33171_ (.a(net809),
    .b(_06645_),
    .c(_06722_),
    .o1(_07690_));
 b15and002ar1n02x5 _33172_ (.a(_06602_),
    .b(_07690_),
    .o(_07691_));
 b15oai013aq1n04x5 _33173_ (.a(_07683_),
    .b(_07685_),
    .c(_07689_),
    .d(_07691_),
    .o1(_07692_));
 b15norp03ar1n02x5 _33174_ (.a(_06661_),
    .b(_06628_),
    .c(_06642_),
    .o1(_07693_));
 b15xor002ar1n02x5 _33175_ (.a(net811),
    .b(_06673_),
    .out0(_07694_));
 b15aoi013an1n02x5 _33176_ (.a(_07693_),
    .b(_07694_),
    .c(_07142_),
    .d(net819),
    .o1(_07695_));
 b15nand04aq1n02x5 _33177_ (.a(net803),
    .b(net805),
    .c(net797),
    .d(net816),
    .o1(_07696_));
 b15nor004ah1n03x5 _33178_ (.a(net811),
    .b(_07230_),
    .c(_07696_),
    .d(_07218_),
    .o1(_07698_));
 b15nanb02ah1n04x5 _33179_ (.a(net810),
    .b(net797),
    .out0(_07699_));
 b15oai022ah1n06x5 _33180_ (.a(_06724_),
    .b(_07183_),
    .c(_07699_),
    .d(_06654_),
    .o1(_07700_));
 b15aoi013an1n08x5 _33181_ (.a(_07698_),
    .b(_07700_),
    .c(_06514_),
    .d(_06693_),
    .o1(_07701_));
 b15nand02al1n03x5 _33182_ (.a(net806),
    .b(net809),
    .o1(_07702_));
 b15aob012as1n03x5 _33183_ (.a(\us11.a[5] ),
    .b(net806),
    .c(\us11.a[0] ),
    .out0(_07703_));
 b15nand04as1n08x5 _33184_ (.a(_06538_),
    .b(_06602_),
    .c(_07702_),
    .d(_07703_),
    .o1(_07704_));
 b15nandp3as1n02x5 _33185_ (.a(_06533_),
    .b(_07161_),
    .c(_06682_),
    .o1(_07705_));
 b15ztpn00an1n08x5 PHY_29 ();
 b15aoai13as1n02x5 _33187_ (.a(_07704_),
    .b(_07705_),
    .c(net805),
    .d(_06628_),
    .o1(_07707_));
 b15oaoi13al1n02x5 _33188_ (.a(_06659_),
    .b(_06610_),
    .c(_06527_),
    .d(_06686_),
    .o1(_07709_));
 b15nano23ah1n03x5 _33189_ (.a(_07695_),
    .b(_07701_),
    .c(_07707_),
    .d(_07709_),
    .out0(_07710_));
 b15ztpn00an1n08x5 PHY_28 ();
 b15nand02ar1n02x5 _33191_ (.a(_06577_),
    .b(_07209_),
    .o1(_07712_));
 b15nand02ar1n02x5 _33192_ (.a(net803),
    .b(_07230_),
    .o1(_07713_));
 b15nand02al1n12x5 _33193_ (.a(net801),
    .b(_06536_),
    .o1(_07714_));
 b15oaoi13ah1n03x5 _33194_ (.a(_07712_),
    .b(_07713_),
    .c(net803),
    .d(_07714_),
    .o1(_07715_));
 b15nandp3ar1n08x5 _33195_ (.a(net819),
    .b(_06533_),
    .c(_07218_),
    .o1(_07716_));
 b15oai012ah1n03x5 _33196_ (.a(_07716_),
    .b(_07198_),
    .c(_06519_),
    .o1(_07717_));
 b15oai012an1n06x5 _33197_ (.a(net811),
    .b(_06558_),
    .c(_07185_),
    .o1(_07718_));
 b15oai022ah1n08x5 _33198_ (.a(net811),
    .b(_07715_),
    .c(_07717_),
    .d(_07718_),
    .o1(_07720_));
 b15nano23as1n24x5 _33199_ (.a(net804),
    .b(net797),
    .c(net799),
    .d(net802),
    .out0(_07721_));
 b15nor002al1n06x5 _33200_ (.a(_06659_),
    .b(_06703_),
    .o1(_07722_));
 b15aoi022ah1n06x5 _33201_ (.a(_06580_),
    .b(_06530_),
    .c(_07721_),
    .d(_07722_),
    .o1(_07723_));
 b15nand04aq1n16x5 _33202_ (.a(_07692_),
    .b(_07710_),
    .c(_07720_),
    .d(_07723_),
    .o1(_07724_));
 b15norp02as1n04x5 _33203_ (.a(_06488_),
    .b(_07148_),
    .o1(_07725_));
 b15aoi022ar1n02x5 _33204_ (.a(net811),
    .b(_07725_),
    .c(_06652_),
    .d(_06567_),
    .o1(_07726_));
 b15oai012ar1n02x5 _33205_ (.a(net818),
    .b(net813),
    .c(_06661_),
    .o1(_07727_));
 b15oaoi13aq1n02x5 _33206_ (.a(net819),
    .b(_07727_),
    .c(_06676_),
    .d(_06509_),
    .o1(_07728_));
 b15nandp2ah1n04x5 _33207_ (.a(_06574_),
    .b(_06527_),
    .o1(_07729_));
 b15oai013al1n02x5 _33208_ (.a(_07729_),
    .b(_06652_),
    .c(_06676_),
    .d(_06509_),
    .o1(_07731_));
 b15oai022ah1n04x5 _33209_ (.a(net819),
    .b(_07726_),
    .c(_07728_),
    .d(_07731_),
    .o1(_07732_));
 b15orn002al1n02x5 _33210_ (.a(net800),
    .b(net817),
    .o(_07733_));
 b15aoi112an1n06x5 _33211_ (.a(_06645_),
    .b(_07733_),
    .c(_07132_),
    .d(_07687_),
    .o1(_07734_));
 b15aoi013ar1n02x5 _33212_ (.a(_07734_),
    .b(_07157_),
    .c(_07191_),
    .d(net816),
    .o1(_07735_));
 b15aoi112al1n02x5 _33213_ (.a(net803),
    .b(_07148_),
    .c(_06574_),
    .d(net805),
    .o1(_07736_));
 b15nanb02aq1n16x5 _33214_ (.a(net797),
    .b(net805),
    .out0(_07737_));
 b15oai012aq1n03x5 _33215_ (.a(_07737_),
    .b(_07687_),
    .c(net805),
    .o1(_07738_));
 b15aoi013aq1n04x5 _33216_ (.a(_07736_),
    .b(_07738_),
    .c(_06715_),
    .d(net803),
    .o1(_07739_));
 b15oai012ar1n04x5 _33217_ (.a(_07735_),
    .b(_07739_),
    .c(net816),
    .o1(_07740_));
 b15oab012ar1n08x5 _33218_ (.c(_07740_),
    .a(_06536_),
    .b(_07732_),
    .out0(_07742_));
 b15nor002ah1n02x5 _33219_ (.a(_06632_),
    .b(_07716_),
    .o1(_07743_));
 b15nand03al1n02x5 _33220_ (.a(net799),
    .b(_06533_),
    .c(_07147_),
    .o1(_07744_));
 b15nand03al1n03x5 _33221_ (.a(_07188_),
    .b(_06556_),
    .c(_06673_),
    .o1(_07745_));
 b15aoi012ar1n04x5 _33222_ (.a(net811),
    .b(_07744_),
    .c(_07745_),
    .o1(_07746_));
 b15nonb02ah1n12x5 _33223_ (.a(net797),
    .b(net803),
    .out0(_07747_));
 b15nand03al1n03x5 _33224_ (.a(net799),
    .b(_06499_),
    .c(_07747_),
    .o1(_07748_));
 b15inv000aq1n06x5 _33225_ (.a(net800),
    .o1(_07749_));
 b15nand03as1n03x5 _33226_ (.a(_07749_),
    .b(_06533_),
    .c(_06530_),
    .o1(_07750_));
 b15aoi022an1n04x5 _33227_ (.a(_06527_),
    .b(_06642_),
    .c(_07748_),
    .d(_07750_),
    .o1(_07751_));
 b15oai013ar1n08x5 _33228_ (.a(net804),
    .b(_07743_),
    .c(_07746_),
    .d(_07751_),
    .o1(_07753_));
 b15orn002an1n16x5 _33229_ (.a(net819),
    .b(\us11.a[3] ),
    .o(_07754_));
 b15oaoi13aq1n03x5 _33230_ (.a(net803),
    .b(_06720_),
    .c(_07754_),
    .d(_06722_),
    .o1(_07755_));
 b15oai022ar1n02x5 _33231_ (.a(net810),
    .b(_06643_),
    .c(_06722_),
    .d(_06519_),
    .o1(_07756_));
 b15ao0022ar1n03x5 _33232_ (.a(_07250_),
    .b(_07252_),
    .c(_07756_),
    .d(net803),
    .o(_07757_));
 b15aoai13an1n08x5 _33233_ (.a(_06518_),
    .b(_07755_),
    .c(_07757_),
    .d(_06654_),
    .o1(_07758_));
 b15nandp2ah1n02x5 _33234_ (.a(net798),
    .b(_06632_),
    .o1(_07759_));
 b15norp03al1n02x5 _33235_ (.a(\us11.a[5] ),
    .b(net806),
    .c(net801),
    .o1(_07760_));
 b15aoi013al1n03x5 _33236_ (.a(_07760_),
    .b(_06555_),
    .c(_06476_),
    .d(net801),
    .o1(_07761_));
 b15oai122aq1n12x5 _33237_ (.a(_06536_),
    .b(_06610_),
    .c(_06616_),
    .d(_07759_),
    .e(_07761_),
    .o1(_07762_));
 b15nandp3aq1n12x5 _33238_ (.o1(_07764_),
    .a(_06552_),
    .b(net815),
    .c(_06553_));
 b15oaoi13ar1n08x5 _33239_ (.a(_06698_),
    .b(_07764_),
    .c(net811),
    .d(_06558_),
    .o1(_07765_));
 b15oai022ar1n06x5 _33240_ (.a(_06527_),
    .b(_07258_),
    .c(_06639_),
    .d(_07729_),
    .o1(_07766_));
 b15oai013as1n06x5 _33241_ (.a(_07762_),
    .b(_07765_),
    .c(_07766_),
    .d(_06536_),
    .o1(_07767_));
 b15nandp3ar1n02x5 _33242_ (.a(_06476_),
    .b(_06509_),
    .c(_07173_),
    .o1(_07768_));
 b15oai112aq1n04x5 _33243_ (.a(net816),
    .b(_07768_),
    .c(_07688_),
    .d(_06574_),
    .o1(_07769_));
 b15oaoi13as1n02x5 _33244_ (.a(_06593_),
    .b(_07716_),
    .c(_06659_),
    .d(net819),
    .o1(_07770_));
 b15nor002ar1n02x5 _33245_ (.a(_06659_),
    .b(_06558_),
    .o1(_07771_));
 b15oai013an1n06x5 _33246_ (.a(_07769_),
    .b(_07770_),
    .c(_07771_),
    .d(net816),
    .o1(_07772_));
 b15nand04aq1n16x5 _33247_ (.a(_07753_),
    .b(_07758_),
    .c(_07767_),
    .d(_07772_),
    .o1(_07773_));
 b15norp03as1n24x5 _33248_ (.a(_07724_),
    .b(_07742_),
    .c(_07773_),
    .o1(_07775_));
 b15xnr002an1n16x5 _33249_ (.a(_07679_),
    .b(_07775_),
    .out0(_07776_));
 b15oai013ar1n02x5 _33250_ (.a(_06111_),
    .b(_06105_),
    .c(_06197_),
    .d(net561),
    .o1(_07777_));
 b15aoi012aq1n02x5 _33251_ (.a(_07777_),
    .b(_06221_),
    .c(_06245_),
    .o1(_07778_));
 b15nona22an1n16x5 _33252_ (.a(net555),
    .b(net547),
    .c(\us33.a[6] ),
    .out0(_07779_));
 b15xor002aq1n02x5 _33253_ (.a(net557),
    .b(net544),
    .out0(_07780_));
 b15nor003al1n02x5 _33254_ (.a(net551),
    .b(_07779_),
    .c(_07780_),
    .o1(_07781_));
 b15oai012ar1n02x5 _33255_ (.a(net564),
    .b(_06195_),
    .c(_07035_),
    .o1(_07782_));
 b15nor002aq1n02x5 _33256_ (.a(_07781_),
    .b(_07782_),
    .o1(_07783_));
 b15nandp2an1n08x5 _33257_ (.a(net557),
    .b(net545),
    .o1(_07784_));
 b15oai022ar1n02x5 _33258_ (.a(net557),
    .b(_06236_),
    .c(_07784_),
    .d(net544),
    .o1(_07786_));
 b15nand03ah1n03x5 _33259_ (.a(net555),
    .b(_06118_),
    .c(_07786_),
    .o1(_07787_));
 b15nand04aq1n04x5 _33260_ (.a(net560),
    .b(net555),
    .c(net557),
    .d(_06342_),
    .o1(_07788_));
 b15aoi013ah1n04x5 _33261_ (.a(_07778_),
    .b(_07783_),
    .c(_07787_),
    .d(_07788_),
    .o1(_07789_));
 b15oai022ar1n02x5 _33262_ (.a(_06127_),
    .b(_06298_),
    .c(_07040_),
    .d(_06253_),
    .o1(_07790_));
 b15nonb02aq1n16x5 _33263_ (.a(net550),
    .b(net549),
    .out0(_07791_));
 b15nand03al1n03x5 _33264_ (.a(_06089_),
    .b(_06108_),
    .c(_07791_),
    .o1(_07792_));
 b15oaoi13an1n04x5 _33265_ (.a(_06203_),
    .b(_07792_),
    .c(_06174_),
    .d(_07784_),
    .o1(_07793_));
 b15aoai13an1n02x5 _33266_ (.a(net561),
    .b(_07790_),
    .c(_07793_),
    .d(_06111_),
    .o1(_07794_));
 b15oai112ar1n02x5 _33267_ (.a(_06228_),
    .b(_07062_),
    .c(_06215_),
    .d(_07791_),
    .o1(_07795_));
 b15nand02an1n24x5 _33268_ (.a(net563),
    .b(net564),
    .o1(_07797_));
 b15nand03an1n06x5 _33269_ (.a(net545),
    .b(_07797_),
    .c(_07042_),
    .o1(_07798_));
 b15oai013ar1n02x5 _33270_ (.a(_07795_),
    .b(_07798_),
    .c(net557),
    .d(net551),
    .o1(_07799_));
 b15nor004an1n02x5 _33271_ (.a(_06179_),
    .b(_06211_),
    .c(_07012_),
    .d(_07079_),
    .o1(_07800_));
 b15nandp3ar1n08x5 _33272_ (.a(_06089_),
    .b(_07036_),
    .c(_07057_),
    .o1(_07801_));
 b15oai012ah1n02x5 _33273_ (.a(_07801_),
    .b(_06195_),
    .c(_06336_),
    .o1(_07802_));
 b15oai013aq1n03x5 _33274_ (.a(net556),
    .b(_07799_),
    .c(_07800_),
    .d(_07802_),
    .o1(_07803_));
 b15nanb02as1n24x5 _33275_ (.a(net554),
    .b(net559),
    .out0(_07804_));
 b15aoi022ar1n02x5 _33276_ (.a(net557),
    .b(_07115_),
    .c(_07042_),
    .d(net561),
    .o1(_07805_));
 b15nand02ar1n02x5 _33277_ (.a(_06108_),
    .b(_06264_),
    .o1(_07806_));
 b15oai022ar1n02x5 _33278_ (.a(_07804_),
    .b(_07798_),
    .c(_07805_),
    .d(_07806_),
    .o1(_07808_));
 b15nandp2al1n02x5 _33279_ (.a(net551),
    .b(_07808_),
    .o1(_07809_));
 b15oai112al1n02x5 _33280_ (.a(_06217_),
    .b(_07064_),
    .c(_07010_),
    .d(_06279_),
    .o1(_07810_));
 b15aoi012as1n02x5 _33281_ (.a(_07810_),
    .b(_06339_),
    .c(_06179_),
    .o1(_07811_));
 b15nano23aq1n24x5 _33282_ (.a(net548),
    .b(net546),
    .c(net543),
    .d(net552),
    .out0(_07812_));
 b15oab012al1n08x5 _33283_ (.c(net561),
    .a(net559),
    .b(net566),
    .out0(_07813_));
 b15oai022as1n02x5 _33284_ (.a(_07108_),
    .b(_07812_),
    .c(_06313_),
    .d(_07813_),
    .o1(_07814_));
 b15oaoi13ah1n03x5 _33285_ (.a(_06179_),
    .b(_07010_),
    .c(_07812_),
    .d(net559),
    .o1(_07815_));
 b15norp03al1n12x5 _33286_ (.a(net556),
    .b(_07814_),
    .c(_07815_),
    .o1(_07816_));
 b15nandp2aq1n12x5 _33287_ (.a(_06215_),
    .b(_06217_),
    .o1(_07817_));
 b15oai022ah1n02x5 _33288_ (.a(_06325_),
    .b(_06100_),
    .c(_06127_),
    .d(_07817_),
    .o1(_07819_));
 b15aoi112as1n04x5 _33289_ (.a(_07811_),
    .b(_07816_),
    .c(net561),
    .d(_07819_),
    .o1(_07820_));
 b15nand04ah1n06x5 _33290_ (.a(_07794_),
    .b(_07803_),
    .c(_07809_),
    .d(_07820_),
    .o1(_07821_));
 b15nanb02an1n03x5 _33291_ (.a(\us33.a[6] ),
    .b(net558),
    .out0(_07822_));
 b15nona22ah1n02x5 _33292_ (.a(net551),
    .b(net544),
    .c(net547),
    .out0(_07823_));
 b15oaoi13ar1n03x5 _33293_ (.a(_07822_),
    .b(_07823_),
    .c(_06269_),
    .d(net547),
    .o1(_07824_));
 b15norp02ah1n02x5 _33294_ (.a(net564),
    .b(net551),
    .o1(_07825_));
 b15and003ar1n02x5 _33295_ (.a(_06266_),
    .b(_06228_),
    .c(_07825_),
    .o(_07826_));
 b15oai012al1n06x5 _33296_ (.a(_06179_),
    .b(_07824_),
    .c(_07826_),
    .o1(_07827_));
 b15nanb02an1n08x5 _33297_ (.a(\us33.a[6] ),
    .b(net564),
    .out0(_07828_));
 b15nanb03ar1n02x5 _33298_ (.a(net544),
    .b(net551),
    .c(net547),
    .out0(_07830_));
 b15oaoi13an1n03x5 _33299_ (.a(_07828_),
    .b(_07830_),
    .c(_07090_),
    .d(_06345_),
    .o1(_07831_));
 b15oai013al1n06x5 _33300_ (.a(_07032_),
    .b(_06091_),
    .c(_06236_),
    .d(net564),
    .o1(_07832_));
 b15aoi112an1n04x5 _33301_ (.a(net555),
    .b(_07831_),
    .c(_07832_),
    .d(_06333_),
    .o1(_07833_));
 b15nor002as1n04x5 _33302_ (.a(_06298_),
    .b(_07026_),
    .o1(_07834_));
 b15norp02aq1n08x5 _33303_ (.a(_06218_),
    .b(_06135_),
    .o1(_07835_));
 b15aoi013an1n08x5 _33304_ (.a(_07834_),
    .b(_07835_),
    .c(_07097_),
    .d(_06089_),
    .o1(_07836_));
 b15aoi022ah1n08x5 _33305_ (.a(_07827_),
    .b(_07833_),
    .c(_07836_),
    .d(net555),
    .o1(_07837_));
 b15nand02ar1n32x5 _33306_ (.a(_06228_),
    .b(_07791_),
    .o1(_07838_));
 b15nona23as1n32x5 _33307_ (.a(net548),
    .b(net546),
    .c(net543),
    .d(net552),
    .out0(_07839_));
 b15oai022as1n06x5 _33308_ (.a(_06145_),
    .b(_07838_),
    .c(_07100_),
    .d(_07839_),
    .o1(_07841_));
 b15nor003ah1n04x5 _33309_ (.a(_06279_),
    .b(_06096_),
    .c(_07057_),
    .o1(_07842_));
 b15and002ar1n03x5 _33310_ (.a(_06179_),
    .b(_06265_),
    .o(_07843_));
 b15oai112ah1n12x5 _33311_ (.a(net547),
    .b(_06294_),
    .c(_07842_),
    .d(_07843_),
    .o1(_07844_));
 b15nonb02an1n04x5 _33312_ (.a(\us33.a[6] ),
    .b(net558),
    .out0(_07845_));
 b15nanb02al1n02x5 _33313_ (.a(net544),
    .b(net547),
    .out0(_07846_));
 b15norp03aq1n02x5 _33314_ (.a(net555),
    .b(_07845_),
    .c(_07846_),
    .o1(_07847_));
 b15norp03al1n02x5 _33315_ (.a(net547),
    .b(_06105_),
    .c(_06218_),
    .o1(_07848_));
 b15oai012an1n04x5 _33316_ (.a(_07825_),
    .b(_07847_),
    .c(_07848_),
    .o1(_07849_));
 b15nanb03an1n08x5 _33317_ (.a(_07841_),
    .b(_07844_),
    .c(_07849_),
    .out0(_07850_));
 b15oai012ar1n02x5 _33318_ (.a(_06201_),
    .b(_06125_),
    .c(_07093_),
    .o1(_07852_));
 b15nanb02an1n06x5 _33319_ (.a(net545),
    .b(net547),
    .out0(_07853_));
 b15nanb02ar1n12x5 _33320_ (.a(net547),
    .b(net545),
    .out0(_07854_));
 b15oai012as1n02x5 _33321_ (.a(_07853_),
    .b(_07854_),
    .c(_06111_),
    .o1(_07855_));
 b15nanb02an1n06x5 _33322_ (.a(net557),
    .b(net561),
    .out0(_07856_));
 b15norp02ar1n03x5 _33323_ (.a(_07090_),
    .b(_07856_),
    .o1(_07857_));
 b15aoi012aq1n02x5 _33324_ (.a(_07852_),
    .b(_07855_),
    .c(_07857_),
    .o1(_07858_));
 b15aoi013an1n03x5 _33325_ (.a(_06201_),
    .b(_07812_),
    .c(_07010_),
    .d(net561),
    .o1(_07859_));
 b15norp03ah1n03x5 _33326_ (.a(_06179_),
    .b(_06242_),
    .c(_07110_),
    .o1(_07860_));
 b15oai012aq1n04x5 _33327_ (.a(_06295_),
    .b(_07095_),
    .c(_07860_),
    .o1(_07861_));
 b15aoi012as1n06x5 _33328_ (.a(_07858_),
    .b(_07859_),
    .c(_07861_),
    .o1(_07863_));
 b15nona23ar1n02x5 _33329_ (.a(net553),
    .b(net544),
    .c(\us33.a[6] ),
    .d(net551),
    .out0(_07864_));
 b15nanb02ar1n16x5 _33330_ (.a(\us33.a[6] ),
    .b(net553),
    .out0(_07865_));
 b15oaoi13al1n03x5 _33331_ (.a(_06346_),
    .b(_07864_),
    .c(_07090_),
    .d(_07865_),
    .o1(_07866_));
 b15nonb02al1n16x5 _33332_ (.a(net553),
    .b(net565),
    .out0(_07867_));
 b15oai112al1n02x5 _33333_ (.a(_06266_),
    .b(_07048_),
    .c(_07867_),
    .d(_06179_),
    .o1(_07868_));
 b15oab012ah1n03x5 _33334_ (.a(_07866_),
    .b(_07868_),
    .c(_06146_),
    .out0(_07869_));
 b15aoi012an1n02x5 _33335_ (.a(_06105_),
    .b(_07093_),
    .c(\us33.a[5] ),
    .o1(_07870_));
 b15oai012aq1n02x5 _33336_ (.a(net558),
    .b(_07867_),
    .c(net563),
    .o1(_07871_));
 b15nor003al1n03x5 _33337_ (.a(_06091_),
    .b(_06096_),
    .c(_06221_),
    .o1(_07872_));
 b15aoi022as1n06x5 _33338_ (.a(_06270_),
    .b(_07870_),
    .c(_07871_),
    .d(_07872_),
    .o1(_07874_));
 b15oai022ar1n06x5 _33339_ (.a(_06100_),
    .b(_06197_),
    .c(_07779_),
    .d(_06269_),
    .o1(_07875_));
 b15oai022an1n08x5 _33340_ (.a(_06145_),
    .b(_07854_),
    .c(_07853_),
    .d(_06121_),
    .o1(_07876_));
 b15aoai13al1n08x5 _33341_ (.a(_06143_),
    .b(_07875_),
    .c(_07876_),
    .d(_07048_),
    .o1(_07877_));
 b15norp02as1n02x5 _33342_ (.a(_06244_),
    .b(_06253_),
    .o1(_07878_));
 b15oai022as1n02x5 _33343_ (.a(_06236_),
    .b(_06300_),
    .c(_07016_),
    .d(_06096_),
    .o1(_07879_));
 b15nor003ah1n02x5 _33344_ (.a(\us33.a[5] ),
    .b(net545),
    .c(_07016_),
    .o1(_07880_));
 b15mdn022al1n04x5 _33345_ (.a(_07090_),
    .b(_06318_),
    .o1(_07881_),
    .sa(net558));
 b15aoi022an1n08x5 _33346_ (.a(_07878_),
    .b(_07879_),
    .c(_07880_),
    .d(_07881_),
    .o1(_07882_));
 b15nand04al1n16x5 _33347_ (.a(_07869_),
    .b(_07874_),
    .c(_07877_),
    .d(_07882_),
    .o1(_07883_));
 b15nor004as1n12x5 _33348_ (.a(_07837_),
    .b(_07850_),
    .c(_07863_),
    .d(_07883_),
    .o1(_07885_));
 b15nona22aq1n32x5 _33349_ (.a(_07789_),
    .b(_07821_),
    .c(_07885_),
    .out0(_07886_));
 b15xnr002an1n16x5 _33350_ (.a(_07492_),
    .b(_07886_),
    .out0(_07887_));
 b15xor003al1n02x5 _33351_ (.a(_07586_),
    .b(_07776_),
    .c(_07887_),
    .out0(_07888_));
 b15nor002ar1n03x5 _33352_ (.a(net535),
    .b(_07888_),
    .o1(_07889_));
 b15inv000aq1n06x5 _33353_ (.a(\text_in_r[98] ),
    .o1(_07890_));
 b15aoi012al1n08x5 _33354_ (.a(_07889_),
    .b(_07890_),
    .c(net535),
    .o1(_07891_));
 b15xor002ar1n02x5 _33355_ (.a(\u0.w[0][2] ),
    .b(_07891_),
    .out0(_00099_));
 b15inv040as1n04x5 _33356_ (.a(\text_in_r[99] ),
    .o1(_07892_));
 b15oai012an1n02x5 _33357_ (.a(\us22.a[3] ),
    .b(_06854_),
    .c(net680),
    .o1(_07893_));
 b15nand02an1n02x5 _33358_ (.a(_06981_),
    .b(_06769_),
    .o1(_07895_));
 b15oai112al1n08x5 _33359_ (.a(_06911_),
    .b(_07893_),
    .c(_07895_),
    .d(\us22.a[3] ),
    .o1(_07896_));
 b15norp03aq1n02x5 _33360_ (.a(_06869_),
    .b(_07580_),
    .c(_07384_),
    .o1(_07897_));
 b15oai022al1n04x5 _33361_ (.a(net677),
    .b(_06936_),
    .c(_07338_),
    .d(_06781_),
    .o1(_07898_));
 b15nonb02aq1n03x5 _33362_ (.a(net690),
    .b(net680),
    .out0(_07899_));
 b15aoi013ar1n04x5 _33363_ (.a(_07897_),
    .b(_07898_),
    .c(_07899_),
    .d(_06839_),
    .o1(_07900_));
 b15nonb02ah1n16x5 _33364_ (.a(net684),
    .b(net679),
    .out0(_07901_));
 b15nand04aq1n04x5 _33365_ (.a(_06758_),
    .b(_06872_),
    .c(_06876_),
    .d(_07901_),
    .o1(_07902_));
 b15nandp3ar1n08x5 _33366_ (.a(_07896_),
    .b(_07900_),
    .c(_07902_),
    .o1(_07903_));
 b15nanb02aq1n06x5 _33367_ (.a(\us22.a[0] ),
    .b(net669),
    .out0(_07904_));
 b15and002ar1n16x5 _33368_ (.a(\us22.a[1] ),
    .b(\us22.a[3] ),
    .o(_07906_));
 b15nor003ah1n04x5 _33369_ (.a(net672),
    .b(net687),
    .c(\us22.a[3] ),
    .o1(_07907_));
 b15aoi022ar1n04x5 _33370_ (.a(_06888_),
    .b(_07906_),
    .c(_07907_),
    .d(_06839_),
    .o1(_07908_));
 b15nor002ar1n06x5 _33371_ (.a(_07904_),
    .b(_07908_),
    .o1(_07909_));
 b15nand02as1n24x5 _33372_ (.a(_06822_),
    .b(_06768_),
    .o1(_07910_));
 b15oai013al1n06x5 _33373_ (.a(_06901_),
    .b(_07910_),
    .c(net689),
    .d(_06863_),
    .o1(_07911_));
 b15aoi012as1n02x5 _33374_ (.a(_07909_),
    .b(_07911_),
    .c(net677),
    .o1(_07912_));
 b15aoi012aq1n02x5 _33375_ (.a(net683),
    .b(_06786_),
    .c(_06999_),
    .o1(_07913_));
 b15oai112an1n12x5 _33376_ (.a(_06959_),
    .b(_07913_),
    .c(_06999_),
    .d(_06850_),
    .o1(_07914_));
 b15aoi022ar1n08x5 _33377_ (.a(_06866_),
    .b(_06889_),
    .c(_07372_),
    .d(_07361_),
    .o1(_07915_));
 b15aoi022ar1n08x5 _33378_ (.a(net688),
    .b(_06844_),
    .c(_06807_),
    .d(_06849_),
    .o1(_07917_));
 b15oai022ah1n06x5 _33379_ (.a(net688),
    .b(_07915_),
    .c(_07917_),
    .d(_06792_),
    .o1(_07918_));
 b15nand03ah1n02x5 _33380_ (.a(net688),
    .b(_06800_),
    .c(_06863_),
    .o1(_07919_));
 b15aoi112as1n04x5 _33381_ (.a(net679),
    .b(_07282_),
    .c(_07919_),
    .d(_07508_),
    .o1(_07920_));
 b15oai012aq1n02x5 _33382_ (.a(_06786_),
    .b(net682),
    .c(_07901_),
    .o1(_07921_));
 b15nand03an1n02x5 _33383_ (.a(net679),
    .b(_06800_),
    .c(_06863_),
    .o1(_07922_));
 b15aoi012al1n04x5 _33384_ (.a(_06981_),
    .b(_07921_),
    .c(_07922_),
    .o1(_07923_));
 b15norp03ar1n16x5 _33385_ (.a(_07918_),
    .b(_07920_),
    .c(_07923_),
    .o1(_07924_));
 b15and003ar1n02x5 _33386_ (.a(net675),
    .b(net669),
    .c(net687),
    .o(_07925_));
 b15aoi013al1n02x5 _33387_ (.a(_07925_),
    .b(_06768_),
    .c(_06911_),
    .d(_06882_),
    .o1(_07926_));
 b15nonb02an1n04x5 _33388_ (.a(net672),
    .b(net688),
    .out0(_07928_));
 b15aoi022ar1n02x5 _33389_ (.a(net675),
    .b(_06822_),
    .c(_07329_),
    .d(_07928_),
    .o1(_07929_));
 b15oai022ah1n04x5 _33390_ (.a(net672),
    .b(_07926_),
    .c(_07929_),
    .d(net673),
    .o1(_07930_));
 b15nonb03aq1n03x5 _33391_ (.a(net673),
    .b(net669),
    .c(net672),
    .out0(_07931_));
 b15aoi022ar1n02x5 _33392_ (.a(_06927_),
    .b(_07309_),
    .c(_07931_),
    .d(_06914_),
    .o1(_07932_));
 b15aoi022ar1n02x5 _33393_ (.a(_06950_),
    .b(_07309_),
    .c(_07310_),
    .d(_07367_),
    .o1(_07933_));
 b15oai022aq1n04x5 _33394_ (.a(_06748_),
    .b(_07932_),
    .c(_07933_),
    .d(_07379_),
    .o1(_07934_));
 b15aoi022ah1n08x5 _33395_ (.a(_06889_),
    .b(_07930_),
    .c(_07934_),
    .d(net675),
    .o1(_07935_));
 b15nand04aq1n16x5 _33396_ (.a(_07912_),
    .b(_07914_),
    .c(_07924_),
    .d(_07935_),
    .o1(_07936_));
 b15nor002ar1n06x5 _33397_ (.a(_06915_),
    .b(_07377_),
    .o1(_07937_));
 b15nand02ar1n02x5 _33398_ (.a(net677),
    .b(_07372_),
    .o1(_07939_));
 b15oaoi13an1n02x5 _33399_ (.a(_07937_),
    .b(_07939_),
    .c(_07269_),
    .d(_07291_),
    .o1(_07940_));
 b15aoai13aq1n02x5 _33400_ (.a(_06911_),
    .b(_06849_),
    .c(net677),
    .d(_06973_),
    .o1(_07941_));
 b15norp02ar1n08x5 _33401_ (.a(net671),
    .b(net678),
    .o1(_07942_));
 b15and002ah1n08x5 _33402_ (.a(net674),
    .b(\us22.a[7] ),
    .o(_07943_));
 b15nandp3al1n08x5 _33403_ (.a(_06850_),
    .b(_07942_),
    .c(_07943_),
    .o1(_07944_));
 b15oai012ah1n02x5 _33404_ (.a(_06913_),
    .b(_07944_),
    .c(net675),
    .o1(_07945_));
 b15aoi022an1n06x5 _33405_ (.a(_07940_),
    .b(_07941_),
    .c(_07945_),
    .d(net689),
    .o1(_07946_));
 b15nand04ar1n02x5 _33406_ (.a(\us22.a[7] ),
    .b(_06777_),
    .c(_06872_),
    .d(_07901_),
    .o1(_07947_));
 b15inv040an1n12x5 _33407_ (.a(\us22.a[4] ),
    .o1(_07948_));
 b15oai012aq1n02x5 _33408_ (.a(_07947_),
    .b(_07944_),
    .c(_07948_),
    .o1(_07950_));
 b15oaoi13an1n03x5 _33409_ (.a(_06761_),
    .b(_07576_),
    .c(_07306_),
    .d(_06867_),
    .o1(_07951_));
 b15oai012ah1n02x5 _33410_ (.a(net680),
    .b(_07950_),
    .c(_07951_),
    .o1(_07952_));
 b15norp02ar1n02x5 _33411_ (.a(_07910_),
    .b(_07338_),
    .o1(_07953_));
 b15aoi022aq1n02x5 _33412_ (.a(_06756_),
    .b(_06761_),
    .c(_07953_),
    .d(net689),
    .o1(_07954_));
 b15oai112as1n08x5 _33413_ (.a(_07946_),
    .b(_07952_),
    .c(_06758_),
    .d(_07954_),
    .o1(_07955_));
 b15oai022ar1n02x5 _33414_ (.a(net690),
    .b(_06921_),
    .c(_07279_),
    .d(_06933_),
    .o1(_07956_));
 b15and003ar1n02x5 _33415_ (.a(net685),
    .b(_06822_),
    .c(_07956_),
    .o(_07957_));
 b15nanb02ar1n02x5 _33416_ (.a(net669),
    .b(\us22.a[0] ),
    .out0(_07958_));
 b15nand03ah1n02x5 _33417_ (.a(_06888_),
    .b(_07904_),
    .c(_07958_),
    .o1(_07959_));
 b15nand02al1n06x5 _33418_ (.a(net669),
    .b(_06839_),
    .o1(_07961_));
 b15oaoi13aq1n04x5 _33419_ (.a(net683),
    .b(_07959_),
    .c(_06922_),
    .d(_07961_),
    .o1(_07962_));
 b15aoi112an1n04x5 _33420_ (.a(_06758_),
    .b(_06850_),
    .c(_06878_),
    .d(_07545_),
    .o1(_07963_));
 b15oai013ah1n04x5 _33421_ (.a(net678),
    .b(_07957_),
    .c(_07962_),
    .d(_07963_),
    .o1(_07964_));
 b15oai022aq1n12x5 _33422_ (.a(_06859_),
    .b(_07282_),
    .c(_07344_),
    .d(_07279_),
    .o1(_07965_));
 b15aoi022ar1n04x5 _33423_ (.a(_06904_),
    .b(_06924_),
    .c(_06966_),
    .d(_07364_),
    .o1(_07966_));
 b15nandp3al1n04x5 _33424_ (.a(\us22.a[6] ),
    .b(_06775_),
    .c(_07329_),
    .o1(_07967_));
 b15nandp3al1n04x5 _33425_ (.a(_06999_),
    .b(_07523_),
    .c(_06904_),
    .o1(_07968_));
 b15aoai13ar1n08x5 _33426_ (.a(_07966_),
    .b(net673),
    .c(_07967_),
    .d(_07968_),
    .o1(_07969_));
 b15nandp2aq1n03x5 _33427_ (.a(net671),
    .b(_06786_),
    .o1(_07970_));
 b15aoi022ar1n02x5 _33428_ (.a(_06777_),
    .b(_06926_),
    .c(_07317_),
    .d(_06839_),
    .o1(_07972_));
 b15oai012an1n04x5 _33429_ (.a(_06826_),
    .b(_07970_),
    .c(_07972_),
    .o1(_07973_));
 b15oai022an1n06x5 _33430_ (.a(_06826_),
    .b(_07965_),
    .c(_07969_),
    .d(_07973_),
    .o1(_07974_));
 b15aoai13as1n02x5 _33431_ (.a(net676),
    .b(_07504_),
    .c(_06761_),
    .d(\us22.a[3] ),
    .o1(_07975_));
 b15oaoi13al1n04x5 _33432_ (.a(net680),
    .b(_07975_),
    .c(_06990_),
    .d(net676),
    .o1(_07976_));
 b15norp03an1n04x5 _33433_ (.a(net676),
    .b(_06869_),
    .c(_07580_),
    .o1(_07977_));
 b15oai112al1n12x5 _33434_ (.a(_06999_),
    .b(_07943_),
    .c(_07976_),
    .d(_07977_),
    .o1(_07978_));
 b15and002ah1n02x5 _33435_ (.a(\us22.a[5] ),
    .b(net680),
    .o(_07979_));
 b15norp03al1n02x5 _33436_ (.a(net676),
    .b(net670),
    .c(\us22.a[3] ),
    .o1(_07980_));
 b15aoai13al1n03x5 _33437_ (.a(_07979_),
    .b(_07980_),
    .c(\us22.a[3] ),
    .d(_07523_),
    .o1(_07981_));
 b15oaoi13as1n02x5 _33438_ (.a(\us22.a[6] ),
    .b(_07981_),
    .c(_07961_),
    .d(_07356_),
    .o1(_07983_));
 b15nandp2aq1n08x5 _33439_ (.a(net681),
    .b(_06844_),
    .o1(_07984_));
 b15aob012an1n12x5 _33440_ (.a(_07984_),
    .b(_07361_),
    .c(_06807_),
    .out0(_07985_));
 b15oai012aq1n08x5 _33441_ (.a(net690),
    .b(_07983_),
    .c(_07985_),
    .o1(_07986_));
 b15nand04an1n16x5 _33442_ (.a(_07964_),
    .b(_07974_),
    .c(_07978_),
    .d(_07986_),
    .o1(_07987_));
 b15nor004as1n12x5 _33443_ (.a(_07903_),
    .b(_07936_),
    .c(_07955_),
    .d(_07987_),
    .o1(_07988_));
 b15nand03an1n08x5 _33444_ (.a(net809),
    .b(_06555_),
    .c(_06556_),
    .o1(_07989_));
 b15nor003aq1n06x5 _33445_ (.a(\us11.a[0] ),
    .b(net818),
    .c(_07989_),
    .o1(_07990_));
 b15nor002aq1n04x5 _33446_ (.a(\us11.a[3] ),
    .b(_06661_),
    .o1(_07991_));
 b15aoi112al1n03x5 _33447_ (.a(net813),
    .b(_07990_),
    .c(_07991_),
    .d(\us11.a[0] ),
    .o1(_07992_));
 b15nand02aq1n04x5 _33448_ (.a(_06476_),
    .b(_06669_),
    .o1(_07994_));
 b15nor002aq1n04x5 _33449_ (.a(_06736_),
    .b(_07714_),
    .o1(_07995_));
 b15nor002as1n03x5 _33450_ (.a(_06536_),
    .b(_06610_),
    .o1(_07996_));
 b15oai013ar1n08x5 _33451_ (.a(_07263_),
    .b(_07991_),
    .c(_07995_),
    .d(_07996_),
    .o1(_07997_));
 b15aoi013al1n06x5 _33452_ (.a(_07992_),
    .b(_07994_),
    .c(_07997_),
    .d(net813),
    .o1(_07998_));
 b15ztpn00an1n08x5 PHY_27 ();
 b15norp03ar1n02x5 _33454_ (.a(net813),
    .b(\us11.a[3] ),
    .c(_06587_),
    .o1(_08000_));
 b15aoai13ar1n03x5 _33455_ (.a(\us11.a[0] ),
    .b(_08000_),
    .c(_06650_),
    .d(_06606_),
    .o1(_08001_));
 b15oaoi13ar1n02x5 _33456_ (.a(\us11.a[0] ),
    .b(_06610_),
    .c(_07258_),
    .d(net813),
    .o1(_08002_));
 b15aoai13as1n02x5 _33457_ (.a(\us11.a[3] ),
    .b(_08002_),
    .c(_07240_),
    .d(_06574_),
    .o1(_08003_));
 b15nandp3ah1n02x5 _33458_ (.a(_06536_),
    .b(_07206_),
    .c(_06565_),
    .o1(_08005_));
 b15aoi013an1n04x5 _33459_ (.a(_06632_),
    .b(_08001_),
    .c(_08003_),
    .d(_08005_),
    .o1(_08006_));
 b15norp03aq1n04x5 _33460_ (.a(_06567_),
    .b(_06600_),
    .c(_07225_),
    .o1(_08007_));
 b15nanb02as1n24x5 _33461_ (.a(net808),
    .b(net812),
    .out0(_08008_));
 b15norp03ah1n03x5 _33462_ (.a(_08008_),
    .b(_07258_),
    .c(_07152_),
    .o1(_08009_));
 b15aoi112ah1n06x5 _33463_ (.a(_08007_),
    .b(_08009_),
    .c(_06676_),
    .d(_07722_),
    .o1(_08010_));
 b15oai112ar1n02x5 _33464_ (.a(net821),
    .b(_07191_),
    .c(net809),
    .d(_06574_),
    .o1(_08011_));
 b15nand04ar1n02x5 _33465_ (.a(_06538_),
    .b(_06539_),
    .c(_07173_),
    .d(_07152_),
    .o1(_08012_));
 b15orn003ar1n02x5 _33466_ (.a(_08008_),
    .b(_07198_),
    .c(_07152_),
    .o(_08013_));
 b15and003an1n03x5 _33467_ (.a(_08011_),
    .b(_08012_),
    .c(_08013_),
    .o(_08014_));
 b15nand04ar1n02x5 _33468_ (.a(net820),
    .b(_06539_),
    .c(_06638_),
    .d(_06605_),
    .o1(_08016_));
 b15oaoi13ar1n02x5 _33469_ (.a(net809),
    .b(_08016_),
    .c(_07258_),
    .d(_06605_),
    .o1(_08017_));
 b15aoai13ar1n02x5 _33470_ (.a(_06476_),
    .b(_07173_),
    .c(_06650_),
    .d(net815),
    .o1(_08018_));
 b15aoi012ar1n02x5 _33471_ (.a(_07198_),
    .b(_07200_),
    .c(_08018_),
    .o1(_08019_));
 b15nano23aq1n03x5 _33472_ (.a(_08010_),
    .b(_08014_),
    .c(_08017_),
    .d(_08019_),
    .out0(_08020_));
 b15nor004an1n06x5 _33473_ (.a(net802),
    .b(_06632_),
    .c(_06659_),
    .d(_06724_),
    .o1(_08021_));
 b15aoai13ar1n02x5 _33474_ (.a(_06555_),
    .b(_06609_),
    .c(_06673_),
    .d(net820),
    .o1(_08022_));
 b15norp02ah1n04x5 _33475_ (.a(net821),
    .b(_06536_),
    .o1(_08023_));
 b15aob012ar1n04x5 _33476_ (.a(_08022_),
    .b(_08023_),
    .c(_06501_),
    .out0(_08024_));
 b15aoai13ar1n06x5 _33477_ (.a(_06638_),
    .b(_08021_),
    .c(_08024_),
    .d(net814),
    .o1(_08025_));
 b15norp02as1n04x5 _33478_ (.a(net797),
    .b(net808),
    .o1(_08027_));
 b15oai022aq1n12x5 _33479_ (.a(_06724_),
    .b(_07183_),
    .c(_07754_),
    .d(_07186_),
    .o1(_08028_));
 b15aoi022an1n08x5 _33480_ (.a(_06545_),
    .b(_08027_),
    .c(_08028_),
    .d(net802),
    .o1(_08029_));
 b15norp03ar1n16x5 _33481_ (.a(net799),
    .b(_06542_),
    .c(_08029_),
    .o1(_08030_));
 b15nandp2aq1n02x5 _33482_ (.a(net815),
    .b(_07690_),
    .o1(_08031_));
 b15nand03ar1n04x5 _33483_ (.a(_06632_),
    .b(net809),
    .c(_06676_),
    .o1(_08032_));
 b15aoi012an1n06x5 _33484_ (.a(net814),
    .b(_08031_),
    .c(_08032_),
    .o1(_08033_));
 b15nano23an1n16x5 _33485_ (.a(_08020_),
    .b(_08025_),
    .c(_08030_),
    .d(_08033_),
    .out0(_08034_));
 b15norp03ar1n08x5 _33486_ (.a(net810),
    .b(_06643_),
    .c(_06645_),
    .o1(_08035_));
 b15aoi122ar1n04x5 _33487_ (.a(\us11.a[0] ),
    .b(_07206_),
    .c(_06499_),
    .d(_06514_),
    .e(_08035_),
    .o1(_08036_));
 b15norp03an1n02x5 _33488_ (.a(_06643_),
    .b(_06645_),
    .c(_06628_),
    .o1(_08038_));
 b15aoai13aq1n04x5 _33489_ (.a(_06632_),
    .b(_08038_),
    .c(_06650_),
    .d(_07206_),
    .o1(_08039_));
 b15nand02an1n04x5 _33490_ (.a(_06518_),
    .b(_08035_),
    .o1(_08040_));
 b15aoi013aq1n08x5 _33491_ (.a(_08036_),
    .b(_08039_),
    .c(\us11.a[0] ),
    .d(_08040_),
    .o1(_08041_));
 b15oai013as1n04x5 _33492_ (.a(_06718_),
    .b(_06616_),
    .c(_06632_),
    .d(net802),
    .o1(_08042_));
 b15nand04as1n06x5 _33493_ (.a(net799),
    .b(_06705_),
    .c(_06691_),
    .d(_08042_),
    .o1(_08043_));
 b15oai022ar1n02x5 _33494_ (.a(_06522_),
    .b(_06642_),
    .c(_07152_),
    .d(_06525_),
    .o1(_08044_));
 b15nandp3ah1n02x5 _33495_ (.a(_06574_),
    .b(_07250_),
    .c(_08044_),
    .o1(_08045_));
 b15aoi012al1n06x5 _33496_ (.a(_06536_),
    .b(_08043_),
    .c(_08045_),
    .o1(_08046_));
 b15nand03as1n08x5 _33497_ (.a(net809),
    .b(_07191_),
    .c(_06518_),
    .o1(_08047_));
 b15nanb02an1n06x5 _33498_ (.a(net800),
    .b(net808),
    .out0(_08049_));
 b15nand03ah1n03x5 _33499_ (.a(\us11.a[7] ),
    .b(_06501_),
    .c(_08049_),
    .o1(_08050_));
 b15aoi012ah1n02x5 _33500_ (.a(_06609_),
    .b(_06698_),
    .c(_07749_),
    .o1(_08051_));
 b15aobi12ah1n02x5 _33501_ (.a(_06522_),
    .b(_06682_),
    .c(net804),
    .out0(_08052_));
 b15nand03an1n04x5 _33502_ (.a(net809),
    .b(_06565_),
    .c(_07250_),
    .o1(_08053_));
 b15oai122ar1n12x5 _33503_ (.a(_08047_),
    .b(_08050_),
    .c(_08051_),
    .d(_08052_),
    .e(_08053_),
    .o1(_08054_));
 b15aoi012ar1n02x5 _33504_ (.a(_06553_),
    .b(_07252_),
    .c(_06555_),
    .o1(_08055_));
 b15nand02ar1n02x5 _33505_ (.a(net797),
    .b(_06698_),
    .o1(_08056_));
 b15aoi012ar1n02x5 _33506_ (.a(net816),
    .b(_06476_),
    .c(_07188_),
    .o1(_08057_));
 b15nand03ar1n03x5 _33507_ (.a(net799),
    .b(_07173_),
    .c(_07209_),
    .o1(_08058_));
 b15oai022as1n02x5 _33508_ (.a(_08055_),
    .b(_08056_),
    .c(_08057_),
    .d(_08058_),
    .o1(_08060_));
 b15norp03ar1n02x5 _33509_ (.a(_06567_),
    .b(_06558_),
    .c(_06519_),
    .o1(_08061_));
 b15oai013ar1n02x5 _33510_ (.a(_07680_),
    .b(_06624_),
    .c(_08008_),
    .d(_06554_),
    .o1(_08062_));
 b15ornc04an1n06x5 _33511_ (.a(_08054_),
    .b(_08060_),
    .c(_08061_),
    .d(_08062_),
    .o(_08063_));
 b15and003ar1n02x5 _33512_ (.a(net802),
    .b(net797),
    .c(net814),
    .o(_08064_));
 b15aob012ar1n02x5 _33513_ (.a(_08064_),
    .b(_06525_),
    .c(_06522_),
    .out0(_08065_));
 b15norp02ar1n02x5 _33514_ (.a(_06476_),
    .b(_06548_),
    .o1(_08066_));
 b15oaoi13ar1n02x5 _33515_ (.a(_08065_),
    .b(_07155_),
    .c(_06686_),
    .d(_08066_),
    .o1(_08067_));
 b15nand02al1n02x5 _33516_ (.a(_06602_),
    .b(_07721_),
    .o1(_08068_));
 b15oaoi13al1n04x5 _33517_ (.a(net819),
    .b(_08068_),
    .c(_06639_),
    .d(_07185_),
    .o1(_08069_));
 b15oai122ar1n12x5 _33518_ (.a(_07721_),
    .b(_07216_),
    .c(net814),
    .d(_06650_),
    .e(net820),
    .o1(_08071_));
 b15norp02ar1n02x5 _33519_ (.a(_06552_),
    .b(_06574_),
    .o1(_08072_));
 b15norp03al1n02x5 _33520_ (.a(net799),
    .b(_06488_),
    .c(_06668_),
    .o1(_08073_));
 b15aoai13ar1n04x5 _33521_ (.a(_08072_),
    .b(_08073_),
    .c(_06501_),
    .d(_07249_),
    .o1(_08074_));
 b15nona23an1n08x5 _33522_ (.a(_08067_),
    .b(_08069_),
    .c(_08071_),
    .d(_08074_),
    .out0(_08075_));
 b15nor004as1n12x5 _33523_ (.a(_08041_),
    .b(_08046_),
    .c(_08063_),
    .d(_08075_),
    .o1(_08076_));
 b15nona23as1n32x5 _33524_ (.a(_07998_),
    .b(_08006_),
    .c(_08034_),
    .d(_08076_),
    .out0(_08077_));
 b15xnr002an1n16x5 _33525_ (.a(_07988_),
    .b(_08077_),
    .out0(_08078_));
 b15nand02ah1n02x5 _33526_ (.a(net918),
    .b(net926),
    .o1(_08079_));
 b15nor002aq1n04x5 _33527_ (.a(_07616_),
    .b(_08079_),
    .o1(_08080_));
 b15norp03ar1n02x5 _33528_ (.a(_07605_),
    .b(_05854_),
    .c(_05835_),
    .o1(_08082_));
 b15oab012al1n03x5 _33529_ (.a(net922),
    .b(_08080_),
    .c(_08082_),
    .out0(_08083_));
 b15nand04aq1n03x5 _33530_ (.a(_05911_),
    .b(_05955_),
    .c(_06019_),
    .d(_05844_),
    .o1(_08084_));
 b15oai112aq1n06x5 _33531_ (.a(net934),
    .b(_08084_),
    .c(_05893_),
    .d(_05841_),
    .o1(_08085_));
 b15oai022ar1n02x5 _33532_ (.a(_05841_),
    .b(_05835_),
    .c(_06050_),
    .d(_06405_),
    .o1(_08086_));
 b15oai022as1n04x5 _33533_ (.a(_08083_),
    .b(_08085_),
    .c(_08086_),
    .d(net935),
    .o1(_08087_));
 b15oaoi13aq1n03x5 _33534_ (.a(_05972_),
    .b(_06434_),
    .c(_05969_),
    .d(_05829_),
    .o1(_08088_));
 b15norp03aq1n02x5 _33535_ (.a(net928),
    .b(net925),
    .c(_05921_),
    .o1(_08089_));
 b15nor002ar1n02x5 _33536_ (.a(_05918_),
    .b(_07589_),
    .o1(_08090_));
 b15oai013ah1n04x5 _33537_ (.a(net931),
    .b(_08088_),
    .c(_08089_),
    .d(_08090_),
    .o1(_08091_));
 b15norp02ar1n02x5 _33538_ (.a(_05997_),
    .b(_07451_),
    .o1(_08093_));
 b15oai012ar1n02x5 _33539_ (.a(net928),
    .b(_06052_),
    .c(_08093_),
    .o1(_08094_));
 b15orn002aq1n04x5 _33540_ (.a(net930),
    .b(net925),
    .o(_08095_));
 b15nor003ar1n08x5 _33541_ (.a(net917),
    .b(_05966_),
    .c(_08095_),
    .o1(_08096_));
 b15norp02ar1n02x5 _33542_ (.a(_05935_),
    .b(_05904_),
    .o1(_08097_));
 b15aoai13ar1n02x5 _33543_ (.a(_05870_),
    .b(_08096_),
    .c(_08097_),
    .d(net925),
    .o1(_08098_));
 b15norp02ar1n02x5 _33544_ (.a(net922),
    .b(net932),
    .o1(_08099_));
 b15aoai13ar1n06x5 _33545_ (.a(_08099_),
    .b(_08080_),
    .c(_07432_),
    .d(_07437_),
    .o1(_08100_));
 b15oai022ar1n08x5 _33546_ (.a(_07465_),
    .b(_05997_),
    .c(_05984_),
    .d(_05959_),
    .o1(_08101_));
 b15aoi022ah1n12x5 _33547_ (.a(_06044_),
    .b(_05885_),
    .c(_08101_),
    .d(_05911_),
    .o1(_08102_));
 b15andc04aq1n03x5 _33548_ (.a(_08094_),
    .b(_08098_),
    .c(_08100_),
    .d(_08102_),
    .o(_08104_));
 b15nandp3ar1n02x5 _33549_ (.a(_05955_),
    .b(_07450_),
    .c(_06003_),
    .o1(_08105_));
 b15oaoi13as1n03x5 _33550_ (.a(net925),
    .b(_08105_),
    .c(_06382_),
    .d(_05841_),
    .o1(_08106_));
 b15oai013ah1n06x5 _33551_ (.a(_07427_),
    .b(_06078_),
    .c(_05846_),
    .d(_05969_),
    .o1(_08107_));
 b15aoi012ar1n06x5 _33552_ (.a(net934),
    .b(_06050_),
    .c(_05987_),
    .o1(_08108_));
 b15nor004ar1n06x5 _33553_ (.a(_05895_),
    .b(_06465_),
    .c(_07623_),
    .d(_08108_),
    .o1(_08109_));
 b15aoi022ar1n02x5 _33554_ (.a(_07605_),
    .b(_05844_),
    .c(_05954_),
    .d(_07432_),
    .o1(_08110_));
 b15nor003ah1n03x5 _33555_ (.a(net922),
    .b(_05851_),
    .c(_08110_),
    .o1(_08111_));
 b15nor004ar1n08x5 _33556_ (.a(_08106_),
    .b(_08107_),
    .c(_08109_),
    .d(_08111_),
    .o1(_08112_));
 b15nand04as1n12x5 _33557_ (.a(_08087_),
    .b(_08091_),
    .c(_08104_),
    .d(_08112_),
    .o1(_08113_));
 b15nanb02al1n06x5 _33558_ (.a(net930),
    .b(net921),
    .out0(_08115_));
 b15oa0022as1n03x5 _33559_ (.a(_05911_),
    .b(_05966_),
    .c(_08115_),
    .d(_07605_),
    .o(_08116_));
 b15nand02an1n03x5 _33560_ (.a(net928),
    .b(_06003_),
    .o1(_08117_));
 b15oai122ar1n12x5 _33561_ (.a(_05969_),
    .b(_05997_),
    .c(_05893_),
    .d(_08116_),
    .e(_08117_),
    .o1(_08118_));
 b15aoi022ar1n02x5 _33562_ (.a(_05975_),
    .b(_05947_),
    .c(_05895_),
    .d(_05840_),
    .o1(_08119_));
 b15oai022ar1n04x5 _33563_ (.a(_07465_),
    .b(_05959_),
    .c(_08119_),
    .d(_05967_),
    .o1(_08120_));
 b15oai012ar1n06x5 _33564_ (.a(_08118_),
    .b(_08120_),
    .c(_05969_),
    .o1(_08121_));
 b15aoi022ar1n02x5 _33565_ (.a(net928),
    .b(_05867_),
    .c(_06434_),
    .d(_05955_),
    .o1(_08122_));
 b15aoi012ar1n02x5 _33566_ (.a(net931),
    .b(_06468_),
    .c(_05932_),
    .o1(_08123_));
 b15nona23al1n05x5 _33567_ (.a(_08122_),
    .b(_08123_),
    .c(net925),
    .d(_05844_),
    .out0(_08124_));
 b15qgbno2an1n10x5 _33568_ (.a(_05821_),
    .b(_05846_),
    .o1(_08126_));
 b15aoi012aq1n02x5 _33569_ (.a(_05870_),
    .b(_07465_),
    .c(net934),
    .o1(_08127_));
 b15aoi022ah1n04x5 _33570_ (.a(_05839_),
    .b(_08126_),
    .c(_08127_),
    .d(_06388_),
    .o1(_08128_));
 b15oai112ah1n12x5 _33571_ (.a(_08121_),
    .b(_08124_),
    .c(_05966_),
    .d(_08128_),
    .o1(_08129_));
 b15norp03ar1n04x5 _33572_ (.a(net932),
    .b(_05835_),
    .c(_06365_),
    .o1(_08130_));
 b15nor003ah1n03x5 _33573_ (.a(net920),
    .b(net915),
    .c(_05969_),
    .o1(_08131_));
 b15aoai13as1n08x5 _33574_ (.a(_08130_),
    .b(_08131_),
    .c(_05870_),
    .d(net920),
    .o1(_08132_));
 b15nandp3aq1n04x5 _33575_ (.a(net931),
    .b(_05947_),
    .c(_05915_),
    .o1(_08133_));
 b15aoi022ar1n02x5 _33576_ (.a(_05829_),
    .b(_06012_),
    .c(_06020_),
    .d(_05906_),
    .o1(_08134_));
 b15orn003aq1n04x5 _33577_ (.a(_05894_),
    .b(_07668_),
    .c(_08134_),
    .o(_08135_));
 b15oai022al1n02x5 _33578_ (.a(_05935_),
    .b(_05835_),
    .c(_05846_),
    .d(_05966_),
    .o1(_08137_));
 b15nand03an1n06x5 _33579_ (.a(_06003_),
    .b(_05917_),
    .c(_08137_),
    .o1(_08138_));
 b15nand04an1n12x5 _33580_ (.a(_08132_),
    .b(_08133_),
    .c(_08135_),
    .d(_08138_),
    .o1(_08139_));
 b15nandp2ah1n02x5 _33581_ (.a(_06056_),
    .b(_05906_),
    .o1(_08140_));
 b15aoi012aq1n06x5 _33582_ (.a(_05829_),
    .b(_05906_),
    .c(net932),
    .o1(_08141_));
 b15oaoi13al1n08x5 _33583_ (.a(_05921_),
    .b(_08140_),
    .c(_08141_),
    .d(_05969_),
    .o1(_08142_));
 b15norp03ar1n03x5 _33584_ (.a(net934),
    .b(net928),
    .c(_05921_),
    .o1(_08143_));
 b15aoi112ar1n04x5 _33585_ (.a(net926),
    .b(_08143_),
    .c(_06072_),
    .d(_07636_),
    .o1(_08144_));
 b15oai013al1n04x5 _33586_ (.a(_05959_),
    .b(_06044_),
    .c(_05997_),
    .d(net927),
    .o1(_08145_));
 b15norp02ah1n02x5 _33587_ (.a(_05911_),
    .b(_08145_),
    .o1(_08146_));
 b15norp03as1n04x5 _33588_ (.a(_05969_),
    .b(_05911_),
    .c(_06078_),
    .o1(_08148_));
 b15oab012ar1n02x5 _33589_ (.a(_08148_),
    .b(_06441_),
    .c(net926),
    .out0(_08149_));
 b15oai022aq1n06x5 _33590_ (.a(_08144_),
    .b(_08146_),
    .c(_08149_),
    .d(_05918_),
    .o1(_08150_));
 b15nor003ah1n08x5 _33591_ (.a(_08139_),
    .b(_08142_),
    .c(_08150_),
    .o1(_08151_));
 b15norp02aq1n02x5 _33592_ (.a(net933),
    .b(_06075_),
    .o1(_08152_));
 b15norp03ah1n03x5 _33593_ (.a(net928),
    .b(_05883_),
    .c(_05854_),
    .o1(_08153_));
 b15aoi022aq1n02x5 _33594_ (.a(_05968_),
    .b(_07450_),
    .c(_08153_),
    .d(net931),
    .o1(_08154_));
 b15aoi012ar1n06x5 _33595_ (.a(_08152_),
    .b(_08154_),
    .c(net933),
    .o1(_08155_));
 b15aoai13as1n03x5 _33596_ (.a(_05954_),
    .b(_07411_),
    .c(_05918_),
    .d(_05983_),
    .o1(_08156_));
 b15nor003ar1n08x5 _33597_ (.a(net927),
    .b(_05934_),
    .c(_05935_),
    .o1(_08157_));
 b15aoi012an1n04x5 _33598_ (.a(_08157_),
    .b(_05983_),
    .c(net927),
    .o1(_08159_));
 b15oai112al1n16x5 _33599_ (.a(net924),
    .b(_08156_),
    .c(_08159_),
    .d(net933),
    .o1(_08160_));
 b15norp02ar1n02x5 _33600_ (.a(net930),
    .b(_06034_),
    .o1(_08161_));
 b15aoai13aq1n03x5 _33601_ (.a(_06468_),
    .b(_08161_),
    .c(net930),
    .d(_06032_),
    .o1(_08162_));
 b15nandp2ar1n02x5 _33602_ (.a(_06032_),
    .b(_06424_),
    .o1(_08163_));
 b15nona23al1n05x5 _33603_ (.a(_06444_),
    .b(_07649_),
    .c(_08162_),
    .d(_08163_),
    .out0(_08164_));
 b15aoi022ah1n12x5 _33604_ (.a(\us00.a[3] ),
    .b(_08155_),
    .c(_08160_),
    .d(_08164_),
    .o1(_08165_));
 b15nona23an1n32x5 _33605_ (.a(_08113_),
    .b(_08129_),
    .c(_08151_),
    .d(_08165_),
    .out0(_08166_));
 b15oai012ar1n02x5 _33606_ (.a(_07033_),
    .b(_06217_),
    .c(_06228_),
    .o1(_08167_));
 b15aoi022ar1n02x5 _33607_ (.a(net561),
    .b(_06228_),
    .c(_06217_),
    .d(_06327_),
    .o1(_08168_));
 b15oai012ar1n02x5 _33608_ (.a(_08167_),
    .b(_08168_),
    .c(net557),
    .o1(_08170_));
 b15nand03aq1n02x5 _33609_ (.a(net556),
    .b(_06118_),
    .c(_08170_),
    .o1(_08171_));
 b15oai022as1n02x5 _33610_ (.a(_06089_),
    .b(_06236_),
    .c(_06096_),
    .d(net555),
    .o1(_08172_));
 b15aoi022as1n06x5 _33611_ (.a(_06228_),
    .b(_07064_),
    .c(_08172_),
    .d(net549),
    .o1(_08173_));
 b15oai013an1n08x5 _33612_ (.a(_08171_),
    .b(_08173_),
    .c(_07093_),
    .d(net550),
    .o1(_08174_));
 b15aoi022ar1n02x5 _33613_ (.a(net557),
    .b(_07791_),
    .c(_06215_),
    .d(_07012_),
    .o1(_08175_));
 b15nand02ar1n02x5 _33614_ (.a(net556),
    .b(_06228_),
    .o1(_08176_));
 b15oai022al1n02x5 _33615_ (.a(_06145_),
    .b(_06195_),
    .c(_08175_),
    .d(_08176_),
    .o1(_08177_));
 b15aoi012aq1n02x5 _33616_ (.a(_07110_),
    .b(_06266_),
    .c(net564),
    .o1(_08178_));
 b15oai013an1n08x5 _33617_ (.a(net560),
    .b(_06103_),
    .c(_06318_),
    .d(_08178_),
    .o1(_08179_));
 b15nor003ah1n02x5 _33618_ (.a(_07793_),
    .b(_08177_),
    .c(_08179_),
    .o1(_08181_));
 b15nand02ah1n06x5 _33619_ (.a(_07854_),
    .b(_07853_),
    .o1(_08182_));
 b15oai013aq1n08x5 _33620_ (.a(_06179_),
    .b(_06155_),
    .c(_06318_),
    .d(_08182_),
    .o1(_08183_));
 b15oaoi13ar1n02x5 _33621_ (.a(_07010_),
    .b(_06195_),
    .c(net556),
    .d(_06298_),
    .o1(_08184_));
 b15oab012an1n04x5 _33622_ (.a(_08181_),
    .b(_08183_),
    .c(_08184_),
    .out0(_08185_));
 b15ztpn00an1n08x5 PHY_26 ();
 b15oai022ar1n02x5 _33624_ (.a(_06133_),
    .b(_07804_),
    .c(_07035_),
    .d(_07838_),
    .o1(_08187_));
 b15nand02al1n04x5 _33625_ (.a(net564),
    .b(_08187_),
    .o1(_08188_));
 b15norp02ah1n16x5 _33626_ (.a(_06269_),
    .b(_07779_),
    .o1(_08189_));
 b15aoi012ar1n02x5 _33627_ (.a(_06125_),
    .b(_06121_),
    .c(_07804_),
    .o1(_08190_));
 b15norp02ar1n02x5 _33628_ (.a(net557),
    .b(_06325_),
    .o1(_08192_));
 b15oai013aq1n04x5 _33629_ (.a(net561),
    .b(_08189_),
    .c(_08190_),
    .d(_08192_),
    .o1(_08193_));
 b15aoai13an1n06x5 _33630_ (.a(net563),
    .b(_06220_),
    .c(_06091_),
    .d(net567),
    .o1(_08194_));
 b15oaoi13ah1n04x5 _33631_ (.a(_06201_),
    .b(_06091_),
    .c(_06244_),
    .d(\us33.a[2] ),
    .o1(_08195_));
 b15aoi012al1n04x5 _33632_ (.a(_06091_),
    .b(_07097_),
    .c(_06089_),
    .o1(_08196_));
 b15oai112as1n16x5 _33633_ (.a(_06259_),
    .b(_08194_),
    .c(_08195_),
    .d(_08196_),
    .o1(_08197_));
 b15norp03ar1n03x5 _33634_ (.a(net547),
    .b(net544),
    .c(_06145_),
    .o1(_08198_));
 b15norp02aq1n03x5 _33635_ (.a(_06089_),
    .b(_06210_),
    .o1(_08199_));
 b15nand02ar1n02x5 _33636_ (.a(_06179_),
    .b(_08199_),
    .o1(_08200_));
 b15and002al1n04x5 _33637_ (.a(net551),
    .b(\us33.a[6] ),
    .o(_08201_));
 b15aoi022ar1n02x5 _33638_ (.a(_06206_),
    .b(_06207_),
    .c(_08201_),
    .d(_06333_),
    .o1(_08203_));
 b15aob012ar1n08x5 _33639_ (.a(_08198_),
    .b(_08200_),
    .c(_08203_),
    .out0(_08204_));
 b15nand04ah1n12x5 _33640_ (.a(_08188_),
    .b(_08193_),
    .c(_08197_),
    .d(_08204_),
    .o1(_08205_));
 b15xnr002ar1n02x5 _33641_ (.a(net556),
    .b(net550),
    .out0(_08206_));
 b15oai022ar1n02x5 _33642_ (.a(net550),
    .b(_06121_),
    .c(_08206_),
    .d(net561),
    .o1(_08207_));
 b15aoi013aq1n02x5 _33643_ (.a(net557),
    .b(net549),
    .c(_06217_),
    .d(_08207_),
    .o1(_08208_));
 b15nanb02ar1n03x5 _33644_ (.a(_07040_),
    .b(_07103_),
    .out0(_08209_));
 b15nand02al1n02x5 _33645_ (.a(_06245_),
    .b(_07867_),
    .o1(_08210_));
 b15aoi013ah1n03x5 _33646_ (.a(_08208_),
    .b(_08209_),
    .c(_08210_),
    .d(net557),
    .o1(_08211_));
 b15oai012ah1n03x5 _33647_ (.a(net561),
    .b(_06220_),
    .c(_07012_),
    .o1(_08212_));
 b15nand04as1n02x5 _33648_ (.a(net550),
    .b(_06217_),
    .c(_07035_),
    .d(_07064_),
    .o1(_08214_));
 b15aob012al1n12x5 _33649_ (.a(_08212_),
    .b(_08214_),
    .c(_07063_),
    .out0(_08215_));
 b15nor004ar1n06x5 _33650_ (.a(_06105_),
    .b(_06174_),
    .c(_06287_),
    .d(_07797_),
    .o1(_08216_));
 b15nor004ah1n03x5 _33651_ (.a(_06235_),
    .b(_06218_),
    .c(_06255_),
    .d(_07057_),
    .o1(_08217_));
 b15oai012aq1n03x5 _33652_ (.a(_06135_),
    .b(_06174_),
    .c(net563),
    .o1(_08218_));
 b15nor003an1n03x5 _33653_ (.a(_06089_),
    .b(_06096_),
    .c(_06100_),
    .o1(_08219_));
 b15aoi112ah1n04x5 _33654_ (.a(_08216_),
    .b(_08217_),
    .c(_08218_),
    .d(_08219_),
    .o1(_08220_));
 b15mdn022an1n04x5 _33655_ (.a(_06135_),
    .b(_06174_),
    .o1(_08221_),
    .sa(_06089_));
 b15norp03aq1n04x5 _33656_ (.a(_06201_),
    .b(_06096_),
    .c(_07057_),
    .o1(_08222_));
 b15nandp3al1n08x5 _33657_ (.a(net565),
    .b(_07856_),
    .c(_07026_),
    .o1(_08223_));
 b15aoi112ar1n06x5 _33658_ (.a(_06166_),
    .b(_06269_),
    .c(_07097_),
    .d(\us33.a[6] ),
    .o1(_08225_));
 b15aoi022ah1n08x5 _33659_ (.a(_08221_),
    .b(_08222_),
    .c(_08223_),
    .d(_08225_),
    .o1(_08226_));
 b15norp02an1n04x5 _33660_ (.a(\us33.a[7] ),
    .b(_06091_),
    .o1(_08227_));
 b15nand04an1n08x5 _33661_ (.a(\us33.a[6] ),
    .b(_08227_),
    .c(_06221_),
    .d(_07097_),
    .o1(_08228_));
 b15nand04an1n16x5 _33662_ (.a(_08215_),
    .b(_08220_),
    .c(_08226_),
    .d(_08228_),
    .o1(_08229_));
 b15oaoi13aq1n02x5 _33663_ (.a(_06242_),
    .b(_06307_),
    .c(_07838_),
    .d(_06253_),
    .o1(_08230_));
 b15aoi012aq1n08x5 _33664_ (.a(_07012_),
    .b(_07010_),
    .c(net561),
    .o1(_08231_));
 b15aoai13as1n04x5 _33665_ (.a(net555),
    .b(_08230_),
    .c(_08231_),
    .d(_06341_),
    .o1(_08232_));
 b15aoi022ar1n02x5 _33666_ (.a(net559),
    .b(_06240_),
    .c(_06313_),
    .d(net562),
    .o1(_08233_));
 b15oai012aq1n04x5 _33667_ (.a(_06201_),
    .b(_06242_),
    .c(_08233_),
    .o1(_08234_));
 b15nor002aq1n03x5 _33668_ (.a(_07839_),
    .b(_07026_),
    .o1(_08236_));
 b15aoai13al1n04x5 _33669_ (.a(_06313_),
    .b(_07033_),
    .c(_07097_),
    .d(_06089_),
    .o1(_08237_));
 b15mdn022ar1n08x5 _33670_ (.a(_06243_),
    .b(_06313_),
    .o1(_08238_),
    .sa(_06089_));
 b15oai112ah1n12x5 _33671_ (.a(net556),
    .b(_08237_),
    .c(_08238_),
    .d(net562),
    .o1(_08239_));
 b15oai012al1n02x5 _33672_ (.a(_06312_),
    .b(_07812_),
    .c(_06243_),
    .o1(_08240_));
 b15oaoi13aq1n04x5 _33673_ (.a(net559),
    .b(_08240_),
    .c(_07030_),
    .d(_06133_),
    .o1(_08241_));
 b15oai013ar1n12x5 _33674_ (.a(_08234_),
    .b(_08236_),
    .c(_08239_),
    .d(_08241_),
    .o1(_08242_));
 b15nona23an1n08x5 _33675_ (.a(_08211_),
    .b(_08229_),
    .c(_08232_),
    .d(_08242_),
    .out0(_08243_));
 b15nor004as1n12x5 _33676_ (.a(_08174_),
    .b(_08185_),
    .c(_08205_),
    .d(_08243_),
    .o1(_08244_));
 b15xor002an1n02x5 _33677_ (.a(_08166_),
    .b(_08244_),
    .out0(_08245_));
 b15xor002al1n03x5 _33678_ (.a(_07679_),
    .b(_08245_),
    .out0(_08247_));
 b15xor003as1n04x5 _33679_ (.a(_06354_),
    .b(_08078_),
    .c(_08247_),
    .out0(_08248_));
 b15mdn022al1n12x5 _33680_ (.a(_07892_),
    .b(_08248_),
    .o1(_08249_),
    .sa(net535));
 b15xor002an1n16x5 _33681_ (.a(\u0.w[0][3] ),
    .b(_08249_),
    .out0(_00100_));
 b15ztpn00an1n08x5 PHY_25 ();
 b15nand03al1n02x5 _33683_ (.a(_06574_),
    .b(_06661_),
    .c(_07764_),
    .o1(_08251_));
 b15oai012ar1n02x5 _33684_ (.a(net811),
    .b(_06558_),
    .c(net817),
    .o1(_08252_));
 b15nand03aq1n02x5 _33685_ (.a(net819),
    .b(_08251_),
    .c(_08252_),
    .o1(_08253_));
 b15nor003ar1n08x5 _33686_ (.a(net798),
    .b(_06574_),
    .c(_07167_),
    .o1(_08254_));
 b15nor002ah1n06x5 _33687_ (.a(net818),
    .b(_06587_),
    .o1(_08255_));
 b15and002ar1n03x5 _33688_ (.a(_06574_),
    .b(_07169_),
    .o(_08257_));
 b15oai013ar1n12x5 _33689_ (.a(_06476_),
    .b(_08254_),
    .c(_08255_),
    .d(_08257_),
    .o1(_08258_));
 b15aoi022ar1n04x5 _33690_ (.a(net811),
    .b(_07206_),
    .c(_06509_),
    .d(_06602_),
    .o1(_08259_));
 b15aoi013an1n04x5 _33691_ (.a(net810),
    .b(_08253_),
    .c(_08258_),
    .d(_08259_),
    .o1(_08260_));
 b15nanb02ar1n02x5 _33692_ (.a(net811),
    .b(net799),
    .out0(_08261_));
 b15oai022ar1n02x5 _33693_ (.a(_06675_),
    .b(_08261_),
    .c(_06525_),
    .d(net803),
    .o1(_08262_));
 b15nand03ar1n04x5 _33694_ (.a(_06536_),
    .b(_06713_),
    .c(_08262_),
    .o1(_08263_));
 b15oai013ar1n02x5 _33695_ (.a(net819),
    .b(_06643_),
    .c(_06675_),
    .d(_07161_),
    .o1(_08264_));
 b15aoi013ar1n02x5 _33696_ (.a(_08264_),
    .b(_07230_),
    .c(_06734_),
    .d(_07250_),
    .o1(_08265_));
 b15nor004an1n03x5 _33697_ (.a(net810),
    .b(_06593_),
    .c(_06514_),
    .d(_06602_),
    .o1(_08266_));
 b15aoi112ah1n04x5 _33698_ (.a(net819),
    .b(_08266_),
    .c(_07137_),
    .d(_06650_),
    .o1(_08268_));
 b15nandp3ar1n02x5 _33699_ (.a(_06632_),
    .b(_06499_),
    .c(_06509_),
    .o1(_08269_));
 b15aoi022ar1n02x5 _33700_ (.a(_08263_),
    .b(_08265_),
    .c(_08268_),
    .d(_08269_),
    .o1(_08270_));
 b15nandp3ar1n02x5 _33701_ (.a(net817),
    .b(_07230_),
    .c(_07747_),
    .o1(_08271_));
 b15nand02ar1n02x5 _33702_ (.a(net819),
    .b(_06539_),
    .o1(_08272_));
 b15aoi012ar1n06x5 _33703_ (.a(_06620_),
    .b(_06548_),
    .c(_06556_),
    .o1(_08273_));
 b15oaoi13al1n02x5 _33704_ (.a(net811),
    .b(_08271_),
    .c(_08272_),
    .d(_08273_),
    .o1(_08274_));
 b15nand04al1n02x5 _33705_ (.a(net811),
    .b(net810),
    .c(_06527_),
    .d(_07721_),
    .o1(_08275_));
 b15norp03an1n02x5 _33706_ (.a(net805),
    .b(net799),
    .c(net810),
    .o1(_08276_));
 b15aoai13aq1n04x5 _33707_ (.a(_06533_),
    .b(_08276_),
    .c(_07249_),
    .d(net805),
    .o1(_08277_));
 b15nand03al1n02x5 _33708_ (.a(net799),
    .b(_07173_),
    .c(_07747_),
    .o1(_08279_));
 b15nand03al1n03x5 _33709_ (.a(net811),
    .b(_06509_),
    .c(_07225_),
    .o1(_08280_));
 b15aoi013al1n03x5 _33710_ (.a(net816),
    .b(_08277_),
    .c(_08279_),
    .d(_08280_),
    .o1(_08281_));
 b15aoi022ar1n02x5 _33711_ (.a(_06577_),
    .b(_06545_),
    .c(_06539_),
    .d(net819),
    .o1(_08282_));
 b15oai022aq1n02x5 _33712_ (.a(_06488_),
    .b(_07183_),
    .c(_07699_),
    .d(_08282_),
    .o1(_08283_));
 b15aoi012ar1n02x5 _33713_ (.a(_08281_),
    .b(_08283_),
    .c(_07202_),
    .o1(_08284_));
 b15nona23al1n04x5 _33714_ (.a(_08270_),
    .b(_08274_),
    .c(_08275_),
    .d(_08284_),
    .out0(_08285_));
 b15oai012ar1n02x5 _33715_ (.a(_06714_),
    .b(net810),
    .c(_06654_),
    .o1(_08286_));
 b15oai012al1n02x5 _33716_ (.a(_07251_),
    .b(_06536_),
    .c(net805),
    .o1(_08287_));
 b15oaoi13ar1n02x5 _33717_ (.a(net819),
    .b(_07680_),
    .c(_08286_),
    .d(_08287_),
    .o1(_08288_));
 b15oa0022ar1n02x5 _33718_ (.a(_06654_),
    .b(_07183_),
    .c(_07699_),
    .d(_06724_),
    .o(_08290_));
 b15nand02al1n02x5 _33719_ (.a(net811),
    .b(_07242_),
    .o1(_08291_));
 b15oai022ar1n02x5 _33720_ (.a(net811),
    .b(_07680_),
    .c(_08290_),
    .d(_08291_),
    .o1(_08292_));
 b15oai012as1n03x5 _33721_ (.a(net816),
    .b(_08288_),
    .c(_08292_),
    .o1(_08293_));
 b15norp02ar1n03x5 _33722_ (.a(_06536_),
    .b(_07198_),
    .o1(_08294_));
 b15oai022ar1n02x5 _33723_ (.a(net810),
    .b(_06639_),
    .c(_07198_),
    .d(net819),
    .o1(_08295_));
 b15aoi112ar1n02x5 _33724_ (.a(_06574_),
    .b(_08294_),
    .c(_08295_),
    .d(_06632_),
    .o1(_08296_));
 b15nor002al1n04x5 _33725_ (.a(net809),
    .b(_06686_),
    .o1(_08297_));
 b15oai012ar1n08x5 _33726_ (.a(_06541_),
    .b(_06589_),
    .c(_06536_),
    .o1(_08298_));
 b15aoi022an1n16x5 _33727_ (.a(net815),
    .b(_08297_),
    .c(_08298_),
    .d(net821),
    .o1(_08299_));
 b15aoai13an1n04x5 _33728_ (.a(_08293_),
    .b(_08296_),
    .c(_08299_),
    .d(_06574_),
    .o1(_08301_));
 b15oai022ar1n02x5 _33729_ (.a(_06476_),
    .b(_07186_),
    .c(_07132_),
    .d(net805),
    .o1(_08302_));
 b15nand03ar1n03x5 _33730_ (.a(_06703_),
    .b(_06693_),
    .c(_08302_),
    .o1(_08303_));
 b15nand04al1n02x5 _33731_ (.a(net799),
    .b(net817),
    .c(_06733_),
    .d(_07747_),
    .o1(_08304_));
 b15aob012ar1n08x5 _33732_ (.a(net810),
    .b(_08303_),
    .c(_08304_),
    .out0(_08305_));
 b15oai012al1n02x5 _33733_ (.a(_08277_),
    .b(_08008_),
    .c(_06728_),
    .o1(_08306_));
 b15oai012ar1n02x5 _33734_ (.a(net820),
    .b(_06530_),
    .c(_07245_),
    .o1(_08307_));
 b15oai012ar1n02x5 _33735_ (.a(_08307_),
    .b(_08008_),
    .c(net816),
    .o1(_08308_));
 b15aoi022aq1n02x5 _33736_ (.a(_06476_),
    .b(_08306_),
    .c(_08308_),
    .d(_06652_),
    .o1(_08309_));
 b15and002ar1n02x5 _33737_ (.a(_07263_),
    .b(_07681_),
    .o(_08310_));
 b15obai22ar1n02x5 _33738_ (.a(_07233_),
    .b(net804),
    .c(_08008_),
    .d(_07737_),
    .out0(_08312_));
 b15aoi112ah1n03x5 _33739_ (.a(_06675_),
    .b(_06722_),
    .c(_07152_),
    .d(_06574_),
    .o1(_08313_));
 b15aoi022al1n02x5 _33740_ (.a(_08310_),
    .b(_08312_),
    .c(_08313_),
    .d(net810),
    .o1(_08314_));
 b15nandp3ar1n02x5 _33741_ (.a(net820),
    .b(_07147_),
    .c(_07242_),
    .o1(_08315_));
 b15nand02ar1n02x5 _33742_ (.a(_07173_),
    .b(_07681_),
    .o1(_08316_));
 b15oaoi13aq1n03x5 _33743_ (.a(_07186_),
    .b(_08315_),
    .c(_08316_),
    .d(net820),
    .o1(_08317_));
 b15and003al1n02x5 _33744_ (.a(_06673_),
    .b(_07721_),
    .c(_07157_),
    .o(_08318_));
 b15nano23al1n06x5 _33745_ (.a(_07241_),
    .b(_08314_),
    .c(_08317_),
    .d(_08318_),
    .out0(_08319_));
 b15nand04aq1n12x5 _33746_ (.a(_06614_),
    .b(_08305_),
    .c(_08309_),
    .d(_08319_),
    .o1(_08320_));
 b15nor004an1n08x5 _33747_ (.a(_08260_),
    .b(_08285_),
    .c(_08301_),
    .d(_08320_),
    .o1(_08321_));
 b15ao0022al1n03x5 _33748_ (.a(_05917_),
    .b(_05885_),
    .c(_08126_),
    .d(_05968_),
    .o(_08323_));
 b15oaoi13al1n03x5 _33749_ (.a(net924),
    .b(_05918_),
    .c(_06037_),
    .d(_06056_),
    .o1(_08324_));
 b15norp03aq1n02x5 _33750_ (.a(net930),
    .b(_05928_),
    .c(_05854_),
    .o1(_08325_));
 b15nanb02aq1n04x5 _33751_ (.a(_08325_),
    .b(net927),
    .out0(_08326_));
 b15oaoi13al1n04x5 _33752_ (.a(net933),
    .b(_07448_),
    .c(_06037_),
    .d(net930),
    .o1(_08327_));
 b15oaoi13as1n08x5 _33753_ (.a(_08323_),
    .b(_08324_),
    .c(_08326_),
    .d(_08327_),
    .o1(_08328_));
 b15oab012ar1n02x5 _33754_ (.a(_06364_),
    .b(_07636_),
    .c(_08153_),
    .out0(_08329_));
 b15nonb03aq1n04x5 _33755_ (.a(_08133_),
    .b(_08329_),
    .c(_06363_),
    .out0(_08330_));
 b15oai122al1n16x5 _33756_ (.a(\us00.a[3] ),
    .b(_06440_),
    .c(_05821_),
    .d(_07646_),
    .e(_05918_),
    .o1(_08331_));
 b15nand02ar1n02x5 _33757_ (.a(net927),
    .b(_05915_),
    .o1(_08332_));
 b15aoai13an1n02x5 _33758_ (.a(_06082_),
    .b(_05821_),
    .c(_05977_),
    .d(_08332_),
    .o1(_08334_));
 b15oaoi13as1n03x5 _33759_ (.a(net933),
    .b(_08331_),
    .c(_08334_),
    .d(net925),
    .o1(_08335_));
 b15oai012an1n08x5 _33760_ (.a(_08328_),
    .b(_08330_),
    .c(_08335_),
    .o1(_08336_));
 b15oab012aq1n06x5 _33761_ (.a(net919),
    .b(_05893_),
    .c(_07472_),
    .out0(_08337_));
 b15nandp3ar1n02x5 _33762_ (.a(net923),
    .b(net916),
    .c(net929),
    .o1(_08338_));
 b15xnr002ar1n02x5 _33763_ (.a(net916),
    .b(net929),
    .out0(_08339_));
 b15oai013ar1n03x5 _33764_ (.a(_08338_),
    .b(_08339_),
    .c(net923),
    .d(net932),
    .o1(_08340_));
 b15nanb02aq1n04x5 _33765_ (.a(_08079_),
    .b(_08340_),
    .out0(_08341_));
 b15and003as1n03x5 _33766_ (.a(net923),
    .b(net918),
    .c(net926),
    .o(_08342_));
 b15norp03al1n08x5 _33767_ (.a(net923),
    .b(net918),
    .c(net926),
    .o1(_08343_));
 b15oai112an1n12x5 _33768_ (.a(_05918_),
    .b(_06460_),
    .c(_08342_),
    .d(_08343_),
    .o1(_08345_));
 b15aoi013ah1n08x5 _33769_ (.a(_08337_),
    .b(_08341_),
    .c(_08345_),
    .d(net920),
    .o1(_08346_));
 b15aoi022as1n08x5 _33770_ (.a(_05840_),
    .b(_06388_),
    .c(_06390_),
    .d(_05975_),
    .o1(_08347_));
 b15nandp2al1n02x5 _33771_ (.a(_05946_),
    .b(_06056_),
    .o1(_08348_));
 b15aoi022ar1n04x5 _33772_ (.a(_05969_),
    .b(_05906_),
    .c(_05829_),
    .d(_05946_),
    .o1(_08349_));
 b15oai022al1n06x5 _33773_ (.a(_08347_),
    .b(_08348_),
    .c(_08349_),
    .d(_07397_),
    .o1(_08350_));
 b15oai012al1n02x5 _33774_ (.a(_07473_),
    .b(_05947_),
    .c(net931),
    .o1(_08351_));
 b15oai022an1n04x5 _33775_ (.a(_05918_),
    .b(_05899_),
    .c(_06067_),
    .d(_08351_),
    .o1(_08352_));
 b15aoi112ar1n06x5 _33776_ (.a(_08350_),
    .b(_08352_),
    .c(_07636_),
    .d(_05927_),
    .o1(_08353_));
 b15oab012ar1n04x5 _33777_ (.a(net933),
    .b(_05964_),
    .c(_08325_),
    .out0(_08354_));
 b15oai022ah1n04x5 _33778_ (.a(_07465_),
    .b(_05959_),
    .c(_07448_),
    .d(_05918_),
    .o1(_08356_));
 b15oai012ar1n12x5 _33779_ (.a(net924),
    .b(_08354_),
    .c(_08356_),
    .o1(_08357_));
 b15nona23ar1n12x5 _33780_ (.a(_06406_),
    .b(_08346_),
    .c(_08353_),
    .d(_08357_),
    .out0(_08358_));
 b15oai012ar1n02x5 _33781_ (.a(_05851_),
    .b(_06382_),
    .c(_05972_),
    .o1(_08359_));
 b15oaoi13ah1n03x5 _33782_ (.a(net931),
    .b(_08359_),
    .c(_07637_),
    .d(_06046_),
    .o1(_08360_));
 b15oai022ar1n04x5 _33783_ (.a(_05911_),
    .b(_05921_),
    .c(_06067_),
    .d(net927),
    .o1(_08361_));
 b15aoi022ah1n06x5 _33784_ (.a(_05827_),
    .b(_06468_),
    .c(_08361_),
    .d(net933),
    .o1(_08362_));
 b15nor003aq1n02x5 _33785_ (.a(_07605_),
    .b(net922),
    .c(net928),
    .o1(_08363_));
 b15and003ar1n02x5 _33786_ (.a(_07605_),
    .b(net922),
    .c(net928),
    .o(_08364_));
 b15oai112aq1n08x5 _33787_ (.a(_05839_),
    .b(_07451_),
    .c(_08363_),
    .d(_08364_),
    .o1(_08365_));
 b15aoi112al1n02x5 _33788_ (.a(_05906_),
    .b(_05997_),
    .c(_05846_),
    .d(_05969_),
    .o1(_08367_));
 b15and002as1n04x5 _33789_ (.a(net933),
    .b(net927),
    .o(_08368_));
 b15aoi112aq1n03x5 _33790_ (.a(_05821_),
    .b(_08367_),
    .c(_08368_),
    .d(_07637_),
    .o1(_08369_));
 b15aoi022ar1n12x5 _33791_ (.a(_08360_),
    .b(_08362_),
    .c(_08365_),
    .d(_08369_),
    .o1(_08370_));
 b15nand02an1n04x5 _33792_ (.a(_05906_),
    .b(_06379_),
    .o1(_08371_));
 b15oai112ah1n06x5 _33793_ (.a(_05846_),
    .b(_05932_),
    .c(net934),
    .d(_06076_),
    .o1(_08372_));
 b15oai112an1n16x5 _33794_ (.a(_08371_),
    .b(_08372_),
    .c(_05959_),
    .d(_05987_),
    .o1(_08373_));
 b15nandp3ar1n02x5 _33795_ (.a(net929),
    .b(_06364_),
    .c(_05992_),
    .o1(_08374_));
 b15aob012an1n08x5 _33796_ (.a(_07463_),
    .b(_07418_),
    .c(_08374_),
    .out0(_08375_));
 b15nand02ar1n02x5 _33797_ (.a(_06026_),
    .b(_07419_),
    .o1(_08376_));
 b15oai012al1n02x5 _33798_ (.a(_08376_),
    .b(_07448_),
    .c(_06050_),
    .o1(_08378_));
 b15oa0022ar1n02x5 _33799_ (.a(net917),
    .b(_05851_),
    .c(_05904_),
    .d(_05884_),
    .o(_08379_));
 b15oai022aq1n04x5 _33800_ (.a(_06364_),
    .b(_05929_),
    .c(_08379_),
    .d(net915),
    .o1(_08380_));
 b15aoai13ah1n03x5 _33801_ (.a(net935),
    .b(_08378_),
    .c(_08380_),
    .d(_05975_),
    .o1(_08381_));
 b15nona23an1n12x5 _33802_ (.a(_08107_),
    .b(_08373_),
    .c(_08375_),
    .d(_08381_),
    .out0(_08382_));
 b15nor004as1n12x5 _33803_ (.a(_08336_),
    .b(_08358_),
    .c(_08370_),
    .d(_08382_),
    .o1(_08383_));
 b15xor002as1n06x5 _33804_ (.a(net394),
    .b(_08383_),
    .out0(_08384_));
 b15norp02ar1n02x5 _33805_ (.a(_06145_),
    .b(_07052_),
    .o1(_08385_));
 b15aoai13ar1n02x5 _33806_ (.a(\us33.a[2] ),
    .b(_08385_),
    .c(_08182_),
    .d(net553),
    .o1(_08386_));
 b15aob012an1n02x5 _33807_ (.a(_08386_),
    .b(_06221_),
    .c(_06169_),
    .out0(_08387_));
 b15nand04as1n06x5 _33808_ (.a(net561),
    .b(net550),
    .c(net543),
    .d(_08387_),
    .o1(_08389_));
 b15aoai13an1n08x5 _33809_ (.a(_07115_),
    .b(_08199_),
    .c(_06221_),
    .d(_06206_),
    .o1(_08390_));
 b15oai112al1n16x5 _33810_ (.a(net564),
    .b(_08390_),
    .c(_07804_),
    .d(_07839_),
    .o1(_08391_));
 b15nor002ar1n02x5 _33811_ (.a(_06179_),
    .b(_06255_),
    .o1(_08392_));
 b15oai112al1n06x5 _33812_ (.a(net543),
    .b(_06169_),
    .c(_07018_),
    .d(_08392_),
    .o1(_08393_));
 b15oai122ar1n08x5 _33813_ (.a(_08393_),
    .b(_06195_),
    .c(_06155_),
    .d(_06272_),
    .e(_07804_),
    .o1(_08394_));
 b15oai012as1n04x5 _33814_ (.a(_08391_),
    .b(_08394_),
    .c(net565),
    .o1(_08395_));
 b15nandp3ah1n12x5 _33815_ (.o1(_08396_),
    .a(net564),
    .b(_06193_),
    .c(_06118_));
 b15nandp2as1n03x5 _33816_ (.a(net560),
    .b(_06201_),
    .o1(_08397_));
 b15oai022ar1n02x5 _33817_ (.a(_07100_),
    .b(_08396_),
    .c(_08397_),
    .d(_06272_),
    .o1(_08398_));
 b15and002al1n02x5 _33818_ (.a(net557),
    .b(_08398_),
    .o(_08400_));
 b15aoi012ar1n02x5 _33819_ (.a(net560),
    .b(net564),
    .c(_07804_),
    .o1(_08401_));
 b15aoai13ar1n02x5 _33820_ (.a(_06302_),
    .b(_08401_),
    .c(_06333_),
    .d(_06121_),
    .o1(_08402_));
 b15oai022al1n02x5 _33821_ (.a(_06253_),
    .b(_07040_),
    .c(_07093_),
    .d(_07839_),
    .o1(_08403_));
 b15aob012al1n04x5 _33822_ (.a(_08402_),
    .b(_08403_),
    .c(net555),
    .out0(_08404_));
 b15nor004ar1n02x5 _33823_ (.a(_06089_),
    .b(_06091_),
    .c(_06096_),
    .d(_06312_),
    .o1(_08405_));
 b15aoai13ar1n02x5 _33824_ (.a(_06201_),
    .b(_08405_),
    .c(_06245_),
    .d(_06242_),
    .o1(_08406_));
 b15aoi012ar1n02x5 _33825_ (.a(net557),
    .b(_06240_),
    .c(_07057_),
    .o1(_08407_));
 b15oai112aq1n02x5 _33826_ (.a(net555),
    .b(_06228_),
    .c(_07093_),
    .d(_06211_),
    .o1(_08408_));
 b15oai013aq1n02x5 _33827_ (.a(_08406_),
    .b(_08407_),
    .c(_08408_),
    .d(net550),
    .o1(_08409_));
 b15nor004al1n04x5 _33828_ (.a(net554),
    .b(_06096_),
    .c(_06244_),
    .d(_07012_),
    .o1(_08411_));
 b15aoai13an1n06x5 _33829_ (.a(_07049_),
    .b(_08411_),
    .c(net553),
    .d(_06295_),
    .o1(_08412_));
 b15oai022ar1n02x5 _33830_ (.a(_06236_),
    .b(_06274_),
    .c(_07854_),
    .d(_06179_),
    .o1(_08413_));
 b15aoi022ar1n02x5 _33831_ (.a(_06211_),
    .b(_06193_),
    .c(_08413_),
    .d(net565),
    .o1(_08414_));
 b15oai012aq1n03x5 _33832_ (.a(_08412_),
    .b(_08414_),
    .c(_06255_),
    .o1(_08415_));
 b15nor004ah1n04x5 _33833_ (.a(_08400_),
    .b(_08404_),
    .c(_08409_),
    .d(_08415_),
    .o1(_08416_));
 b15nano23ah1n24x5 _33834_ (.a(net548),
    .b(net543),
    .c(net546),
    .d(net552),
    .out0(_08417_));
 b15nor002as1n04x5 _33835_ (.a(net557),
    .b(_07097_),
    .o1(_08418_));
 b15aoi122an1n02x5 _33836_ (.a(_06201_),
    .b(_08417_),
    .c(_07860_),
    .d(_08418_),
    .e(_06341_),
    .o1(_08419_));
 b15mdn022aq1n04x5 _33837_ (.a(_06125_),
    .b(_07032_),
    .o1(_08420_),
    .sa(_06253_));
 b15aoai13as1n08x5 _33838_ (.a(net563),
    .b(_08420_),
    .c(_06176_),
    .d(_06284_),
    .o1(_08422_));
 b15nor002an1n04x5 _33839_ (.a(net557),
    .b(_06133_),
    .o1(_08423_));
 b15aoi022aq1n04x5 _33840_ (.a(_06158_),
    .b(_07062_),
    .c(_08423_),
    .d(net565),
    .o1(_08424_));
 b15aoi012an1n02x5 _33841_ (.a(net554),
    .b(_08417_),
    .c(_07062_),
    .o1(_08425_));
 b15aoi013al1n04x5 _33842_ (.a(_08419_),
    .b(_08422_),
    .c(_08424_),
    .d(_08425_),
    .o1(_08426_));
 b15nandp2al1n04x5 _33843_ (.a(\us33.a[7] ),
    .b(_06118_),
    .o1(_08427_));
 b15nanb02an1n04x5 _33844_ (.a(net553),
    .b(net545),
    .out0(_08428_));
 b15oai012an1n02x5 _33845_ (.a(_08428_),
    .b(_07097_),
    .c(_07865_),
    .o1(_08429_));
 b15nona23an1n04x5 _33846_ (.a(_07067_),
    .b(_08427_),
    .c(_08429_),
    .d(_06089_),
    .out0(_08430_));
 b15aoi012ar1n02x5 _33847_ (.a(_07084_),
    .b(_06220_),
    .c(\us33.a[5] ),
    .o1(_08431_));
 b15orn003al1n02x5 _33848_ (.a(_06179_),
    .b(_06306_),
    .c(_08431_),
    .o(_08433_));
 b15nonb03ar1n02x5 _33849_ (.a(\us33.a[7] ),
    .b(\us33.a[5] ),
    .c(net560),
    .out0(_08434_));
 b15nonb02as1n04x5 _33850_ (.a(\us33.a[6] ),
    .b(net551),
    .out0(_08435_));
 b15and003ar1n02x5 _33851_ (.a(_06264_),
    .b(_08434_),
    .c(_08435_),
    .o(_08436_));
 b15norp03ar1n02x5 _33852_ (.a(net551),
    .b(_06100_),
    .c(_06287_),
    .o1(_08437_));
 b15mdn022ar1n03x5 _33853_ (.a(_06235_),
    .b(_06274_),
    .o1(_08438_),
    .sa(net560));
 b15aoi012ah1n02x5 _33854_ (.a(_08436_),
    .b(_08437_),
    .c(_08438_),
    .o1(_08439_));
 b15nand04ar1n03x5 _33855_ (.a(net565),
    .b(net553),
    .c(\us33.a[5] ),
    .d(\us33.a[6] ),
    .o1(_08440_));
 b15orn002al1n04x5 _33856_ (.a(net551),
    .b(\us33.a[7] ),
    .o(_08441_));
 b15oaoi13an1n03x5 _33857_ (.a(_08440_),
    .b(_08441_),
    .c(_06269_),
    .d(net558),
    .o1(_08442_));
 b15aob012aq1n04x5 _33858_ (.a(_06103_),
    .b(_07845_),
    .c(net553),
    .out0(_08444_));
 b15aoi013an1n03x5 _33859_ (.a(_08442_),
    .b(_08444_),
    .c(_08227_),
    .d(_07067_),
    .o1(_08445_));
 b15nand04as1n08x5 _33860_ (.a(_08430_),
    .b(_08433_),
    .c(_08439_),
    .d(_08445_),
    .o1(_08446_));
 b15aoi012ar1n04x5 _33861_ (.a(_07080_),
    .b(_07867_),
    .c(_06158_),
    .o1(_08447_));
 b15aoai13al1n06x5 _33862_ (.a(_06219_),
    .b(_06215_),
    .c(_07791_),
    .d(_07010_),
    .o1(_08448_));
 b15norp02aq1n02x5 _33863_ (.a(net561),
    .b(_07012_),
    .o1(_08449_));
 b15aoi013al1n06x5 _33864_ (.a(_08449_),
    .b(_06341_),
    .c(_06111_),
    .d(net561),
    .o1(_08450_));
 b15oai022an1n12x5 _33865_ (.a(_06179_),
    .b(_08447_),
    .c(_08448_),
    .d(_08450_),
    .o1(_08451_));
 b15nor002al1n02x5 _33866_ (.a(net551),
    .b(_06145_),
    .o1(_08452_));
 b15oaoi13aq1n03x5 _33867_ (.a(_07846_),
    .b(_07822_),
    .c(net563),
    .d(_07845_),
    .o1(_08453_));
 b15and003ar1n02x5 _33868_ (.a(_06089_),
    .b(_06211_),
    .c(net544),
    .o(_08455_));
 b15oai012aq1n08x5 _33869_ (.a(_08452_),
    .b(_08453_),
    .c(_08455_),
    .o1(_08456_));
 b15nor002ah1n02x5 _33870_ (.a(_06253_),
    .b(_06287_),
    .o1(_08457_));
 b15oai022an1n06x5 _33871_ (.a(_06201_),
    .b(_06091_),
    .c(_06244_),
    .d(net562),
    .o1(_08458_));
 b15nor003al1n08x5 _33872_ (.a(_06091_),
    .b(_06096_),
    .c(_06127_),
    .o1(_08459_));
 b15aoi022ar1n12x5 _33873_ (.a(_08457_),
    .b(_08458_),
    .c(_08459_),
    .d(_06111_),
    .o1(_08460_));
 b15norp03ar1n02x5 _33874_ (.a(net553),
    .b(_06298_),
    .c(_07797_),
    .o1(_08461_));
 b15aoi012an1n02x5 _33875_ (.a(_08461_),
    .b(_06243_),
    .c(net553),
    .o1(_08462_));
 b15oai112al1n08x5 _33876_ (.a(_08456_),
    .b(_08460_),
    .c(_08462_),
    .d(_06089_),
    .o1(_08463_));
 b15nor004ah1n04x5 _33877_ (.a(_08426_),
    .b(_08446_),
    .c(_08451_),
    .d(_08463_),
    .o1(_08464_));
 b15andc04as1n16x5 _33878_ (.a(_08389_),
    .b(_08395_),
    .c(_08416_),
    .d(_08464_),
    .o(_08466_));
 b15xor002an1n16x5 _33879_ (.a(_08166_),
    .b(_08466_),
    .out0(_08467_));
 b15nandp2al1n02x5 _33880_ (.a(_06786_),
    .b(net680),
    .o1(_08468_));
 b15norp03an1n02x5 _33881_ (.a(net677),
    .b(_08468_),
    .c(_06854_),
    .o1(_08469_));
 b15oai112ah1n04x5 _33882_ (.a(_06822_),
    .b(_06839_),
    .c(_06966_),
    .d(net684),
    .o1(_08470_));
 b15aoai13al1n08x5 _33883_ (.a(_08470_),
    .b(_07282_),
    .c(_06792_),
    .d(_07279_),
    .o1(_08471_));
 b15aoi012al1n04x5 _33884_ (.a(_08469_),
    .b(_08471_),
    .c(net677),
    .o1(_08472_));
 b15nandp2al1n05x5 _33885_ (.a(_06813_),
    .b(_07372_),
    .o1(_08473_));
 b15nandp3al1n03x5 _33886_ (.a(_06852_),
    .b(_06839_),
    .c(_07363_),
    .o1(_08474_));
 b15aoi012al1n06x5 _33887_ (.a(_06786_),
    .b(_08473_),
    .c(_08474_),
    .o1(_08475_));
 b15nandp3al1n04x5 _33888_ (.a(_06999_),
    .b(_06777_),
    .c(_06911_),
    .o1(_08477_));
 b15nand02an1n04x5 _33889_ (.a(_06839_),
    .b(_07928_),
    .o1(_08478_));
 b15aoi112ah1n06x5 _33890_ (.a(_06882_),
    .b(_06869_),
    .c(_08477_),
    .d(_08478_),
    .o1(_08479_));
 b15oai112al1n02x5 _33891_ (.a(_06999_),
    .b(_06768_),
    .c(_07348_),
    .d(_06882_),
    .o1(_08480_));
 b15norp03as1n04x5 _33892_ (.a(net678),
    .b(_07306_),
    .c(_08480_),
    .o1(_08481_));
 b15nor004as1n12x5 _33893_ (.a(_06983_),
    .b(_08475_),
    .c(_08479_),
    .d(_08481_),
    .o1(_08482_));
 b15nandp2al1n02x5 _33894_ (.a(_06912_),
    .b(_06844_),
    .o1(_08483_));
 b15nanb02aq1n04x5 _33895_ (.a(net675),
    .b(net669),
    .out0(_08484_));
 b15oa0022al1n04x5 _33896_ (.a(_06826_),
    .b(_07512_),
    .c(_06838_),
    .d(_08484_),
    .o(_08485_));
 b15oai013an1n08x5 _33897_ (.a(_08483_),
    .b(_08485_),
    .c(_07531_),
    .d(_06758_),
    .o1(_08486_));
 b15norp03ar1n02x5 _33898_ (.a(net670),
    .b(net671),
    .c(\us22.a[3] ),
    .o1(_08488_));
 b15aoai13ar1n02x5 _33899_ (.a(_06839_),
    .b(_08488_),
    .c(_06927_),
    .d(net670),
    .o1(_08489_));
 b15nor002aq1n12x5 _33900_ (.a(_06933_),
    .b(_07302_),
    .o1(_08490_));
 b15aob012ar1n02x5 _33901_ (.a(_08489_),
    .b(_06955_),
    .c(_08490_),
    .out0(_08491_));
 b15aoi112aq1n03x5 _33902_ (.a(_06792_),
    .b(_08486_),
    .c(_08491_),
    .d(_06758_),
    .o1(_08492_));
 b15norp02ar1n02x5 _33903_ (.a(_06786_),
    .b(_06945_),
    .o1(_08493_));
 b15nonb02an1n04x5 _33904_ (.a(net690),
    .b(net676),
    .out0(_08494_));
 b15nor002ar1n12x5 _33905_ (.a(\us22.a[5] ),
    .b(net670),
    .o1(_08495_));
 b15nona23al1n08x5 _33906_ (.a(_06869_),
    .b(_08494_),
    .c(_08495_),
    .d(_06999_),
    .out0(_08496_));
 b15oai012al1n06x5 _33907_ (.a(_08496_),
    .b(_06973_),
    .c(_07356_),
    .o1(_08497_));
 b15nor004as1n03x5 _33908_ (.a(net685),
    .b(_06940_),
    .c(_08493_),
    .d(_08497_),
    .o1(_08499_));
 b15oai112aq1n12x5 _33909_ (.a(_08472_),
    .b(_08482_),
    .c(_08492_),
    .d(_08499_),
    .o1(_08500_));
 b15aoi013ah1n06x5 _33910_ (.a(net678),
    .b(_06777_),
    .c(_06852_),
    .d(net683),
    .o1(_08501_));
 b15oai013ar1n04x5 _33911_ (.a(_08501_),
    .b(_06824_),
    .c(_06748_),
    .d(net683),
    .o1(_08502_));
 b15nanb02as1n06x5 _33912_ (.a(net669),
    .b(\us22.a[5] ),
    .out0(_08503_));
 b15nandp2ar1n03x5 _33913_ (.a(net683),
    .b(_07309_),
    .o1(_08504_));
 b15oai022al1n08x5 _33914_ (.a(_06954_),
    .b(_08503_),
    .c(_08504_),
    .d(_06922_),
    .o1(_08505_));
 b15nonb02ah1n06x5 _33915_ (.a(net676),
    .b(net690),
    .out0(_08506_));
 b15aoi012al1n06x5 _33916_ (.a(_08502_),
    .b(_08505_),
    .c(_08506_),
    .o1(_08507_));
 b15nor002aq1n06x5 _33917_ (.a(_06758_),
    .b(_07387_),
    .o1(_08508_));
 b15aoai13al1n04x5 _33918_ (.a(net690),
    .b(_08508_),
    .c(_06986_),
    .d(_07546_),
    .o1(_08510_));
 b15nor002ah1n04x5 _33919_ (.a(_06981_),
    .b(_06790_),
    .o1(_08511_));
 b15nand02ar1n02x5 _33920_ (.a(_06761_),
    .b(_07329_),
    .o1(_08512_));
 b15oai022al1n02x5 _33921_ (.a(_06769_),
    .b(_06748_),
    .c(_08512_),
    .d(net671),
    .o1(_08513_));
 b15nor003al1n02x5 _33922_ (.a(_06792_),
    .b(_07277_),
    .c(_06824_),
    .o1(_08514_));
 b15nor004ah1n03x5 _33923_ (.a(_06826_),
    .b(_08511_),
    .c(_08513_),
    .d(_08514_),
    .o1(_08515_));
 b15norp03al1n02x5 _33924_ (.a(\us22.a[7] ),
    .b(_06783_),
    .c(_07306_),
    .o1(_08516_));
 b15nand02ar1n02x5 _33925_ (.a(net674),
    .b(_07329_),
    .o1(_08517_));
 b15aoi012ar1n02x5 _33926_ (.a(_07365_),
    .b(_06786_),
    .c(_06882_),
    .o1(_08518_));
 b15oaoi13ar1n02x5 _33927_ (.a(net671),
    .b(_08517_),
    .c(_08518_),
    .d(_06984_),
    .o1(_08519_));
 b15oai012aq1n04x5 _33928_ (.a(net680),
    .b(_08516_),
    .c(_08519_),
    .o1(_08521_));
 b15aoi013ah1n04x5 _33929_ (.a(_08507_),
    .b(_08510_),
    .c(_08515_),
    .d(_08521_),
    .o1(_08522_));
 b15mdn022al1n03x5 _33930_ (.a(_06924_),
    .b(_06844_),
    .o1(_08523_),
    .sa(_06792_));
 b15oai112al1n02x5 _33931_ (.a(net680),
    .b(_06945_),
    .c(_08523_),
    .d(net690),
    .o1(_08524_));
 b15xor002al1n02x5 _33932_ (.a(net670),
    .b(\us22.a[3] ),
    .out0(_08525_));
 b15nand03aq1n04x5 _33933_ (.a(_06872_),
    .b(_06768_),
    .c(_08525_),
    .o1(_08526_));
 b15nonb03ah1n02x5 _33934_ (.a(\us22.a[3] ),
    .b(net670),
    .c(net676),
    .out0(_08527_));
 b15aoi012ah1n04x5 _33935_ (.a(_08527_),
    .b(_07361_),
    .c(_07523_),
    .o1(_08528_));
 b15nand02an1n03x5 _33936_ (.a(_07319_),
    .b(net671),
    .o1(_08529_));
 b15oai122aq1n12x5 _33937_ (.a(_08526_),
    .b(_08528_),
    .c(_08529_),
    .d(_06981_),
    .e(_06990_),
    .o1(_08530_));
 b15nor004aq1n02x5 _33938_ (.a(_06826_),
    .b(_06933_),
    .c(_06850_),
    .d(_06781_),
    .o1(_08532_));
 b15oai013as1n02x5 _33939_ (.a(_08524_),
    .b(_08530_),
    .c(_08532_),
    .d(net680),
    .o1(_08533_));
 b15aoi012ar1n02x5 _33940_ (.a(_06852_),
    .b(_06904_),
    .c(_06822_),
    .o1(_08534_));
 b15norp03ar1n02x5 _33941_ (.a(net690),
    .b(_06933_),
    .c(_08534_),
    .o1(_08535_));
 b15oai012ar1n02x5 _33942_ (.a(\us22.a[3] ),
    .b(_07545_),
    .c(_06758_),
    .o1(_08536_));
 b15aoi112aq1n02x5 _33943_ (.a(_08535_),
    .b(_08536_),
    .c(_08490_),
    .d(_06911_),
    .o1(_08537_));
 b15nano22an1n02x5 _33944_ (.a(net670),
    .b(net671),
    .c(net690),
    .out0(_08538_));
 b15nonb03an1n02x5 _33945_ (.a(net690),
    .b(net671),
    .c(net670),
    .out0(_08539_));
 b15oai112ah1n06x5 _33946_ (.a(\us22.a[1] ),
    .b(_06823_),
    .c(_08538_),
    .d(_08539_),
    .o1(_08540_));
 b15nand02ar1n02x5 _33947_ (.a(net680),
    .b(_06915_),
    .o1(_08541_));
 b15aoai13ar1n02x5 _33948_ (.a(_08540_),
    .b(_08541_),
    .c(_06878_),
    .d(_06778_),
    .o1(_08543_));
 b15oai013ar1n02x5 _33949_ (.a(_06826_),
    .b(_06775_),
    .c(_06904_),
    .d(_06821_),
    .o1(_08544_));
 b15nonb02as1n04x5 _33950_ (.a(net683),
    .b(net673),
    .out0(_08545_));
 b15aoi022ar1n08x5 _33951_ (.a(_06904_),
    .b(_06768_),
    .c(_08545_),
    .d(\us22.a[4] ),
    .o1(_08546_));
 b15aoi022ah1n06x5 _33952_ (.a(_06960_),
    .b(_08495_),
    .c(_07979_),
    .d(_06896_),
    .o1(_08547_));
 b15oai022as1n06x5 _33953_ (.a(_06969_),
    .b(_08546_),
    .c(_08547_),
    .d(\us22.a[4] ),
    .o1(_08548_));
 b15aoi112aq1n02x5 _33954_ (.a(_08543_),
    .b(_08544_),
    .c(net690),
    .d(_08548_),
    .o1(_08549_));
 b15norp03ar1n02x5 _33955_ (.a(net690),
    .b(_06792_),
    .c(_06878_),
    .o1(_08550_));
 b15aoai13as1n02x5 _33956_ (.a(_06758_),
    .b(_08550_),
    .c(_06844_),
    .d(_06792_),
    .o1(_08551_));
 b15aoai13aq1n04x5 _33957_ (.a(_08533_),
    .b(_08537_),
    .c(_08549_),
    .d(_08551_),
    .o1(_08552_));
 b15orn003aq1n24x5 _33958_ (.a(_08500_),
    .b(_08522_),
    .c(_08552_),
    .o(_08554_));
 b15xor002ar1n03x5 _33959_ (.a(_08467_),
    .b(_08554_),
    .out0(_08555_));
 b15xor003an1n02x5 _33960_ (.a(_06354_),
    .b(_08384_),
    .c(_08555_),
    .out0(_08556_));
 b15cmbn22ah1n04x5 _33961_ (.clk1(\text_in_r[100] ),
    .clk2(_08556_),
    .clkout(_08557_),
    .s(net535));
 b15xor002as1n02x5 _33962_ (.a(\u0.w[0][4] ),
    .b(_08557_),
    .out0(_00101_));
 b15nor004ar1n02x5 _33963_ (.a(_05821_),
    .b(_05883_),
    .c(_05854_),
    .d(_08368_),
    .o1(_08558_));
 b15oaoi13ar1n02x5 _33964_ (.a(net930),
    .b(_06034_),
    .c(_05854_),
    .d(_05883_),
    .o1(_08559_));
 b15aoai13aq1n02x5 _33965_ (.a(net924),
    .b(_08558_),
    .c(_08559_),
    .d(_08368_),
    .o1(_08560_));
 b15aob012ar1n02x5 _33966_ (.a(_05924_),
    .b(_06019_),
    .c(_05969_),
    .out0(_08561_));
 b15aoi012ah1n02x5 _33967_ (.a(_08126_),
    .b(_08561_),
    .c(_05911_),
    .o1(_08562_));
 b15oai012al1n06x5 _33968_ (.a(_08560_),
    .b(_08562_),
    .c(_06037_),
    .o1(_08564_));
 b15norp03ar1n03x5 _33969_ (.a(_05911_),
    .b(_05966_),
    .c(_05967_),
    .o1(_08565_));
 b15norp02aq1n03x5 _33970_ (.a(\us00.a[3] ),
    .b(_07405_),
    .o1(_08566_));
 b15oaoi13aq1n03x5 _33971_ (.a(_05918_),
    .b(_05917_),
    .c(_08565_),
    .d(_08566_),
    .o1(_08567_));
 b15nor004ah1n03x5 _33972_ (.a(net915),
    .b(_05911_),
    .c(_05883_),
    .d(_05894_),
    .o1(_08568_));
 b15oai022aq1n04x5 _33973_ (.a(_05883_),
    .b(_05929_),
    .c(_05997_),
    .d(net933),
    .o1(_08569_));
 b15aoi112ar1n06x5 _33974_ (.a(_08148_),
    .b(_08568_),
    .c(_08569_),
    .d(_07634_),
    .o1(_08570_));
 b15norp03al1n02x5 _33975_ (.a(_05911_),
    .b(_05894_),
    .c(_05854_),
    .o1(_08571_));
 b15aoai13ah1n03x5 _33976_ (.a(_05975_),
    .b(_08571_),
    .c(_06388_),
    .d(net915),
    .o1(_08572_));
 b15aoi013ah1n06x5 _33977_ (.a(_08567_),
    .b(_08570_),
    .c(_08572_),
    .d(_05918_),
    .o1(_08573_));
 b15aoi122aq1n02x5 _33978_ (.a(net930),
    .b(_07636_),
    .c(_05895_),
    .d(_06006_),
    .e(_05827_),
    .o1(_08575_));
 b15aob012ar1n02x5 _33979_ (.a(net924),
    .b(_05972_),
    .c(_06033_),
    .out0(_08576_));
 b15oai022ar1n02x5 _33980_ (.a(net924),
    .b(_06078_),
    .c(_05972_),
    .d(_05918_),
    .o1(_08577_));
 b15aoi022ar1n02x5 _33981_ (.a(_05968_),
    .b(_06006_),
    .c(_08577_),
    .d(_05969_),
    .o1(_08578_));
 b15aoi013aq1n02x5 _33982_ (.a(_08575_),
    .b(_08576_),
    .c(_08578_),
    .d(net930),
    .o1(_08579_));
 b15oai012ah1n04x5 _33983_ (.a(_05921_),
    .b(_06037_),
    .c(net930),
    .o1(_08580_));
 b15nor002ar1n04x5 _33984_ (.a(net933),
    .b(_05942_),
    .o1(_08581_));
 b15nor002al1n03x5 _33985_ (.a(_05882_),
    .b(_05846_),
    .o1(_08582_));
 b15oai012ah1n04x5 _33986_ (.a(_05891_),
    .b(_05929_),
    .c(_05883_),
    .o1(_08583_));
 b15nandp2al1n03x5 _33987_ (.a(net927),
    .b(_05894_),
    .o1(_08584_));
 b15norp03aq1n08x5 _33988_ (.a(_05911_),
    .b(_05928_),
    .c(_05854_),
    .o1(_08586_));
 b15aoi222as1n08x5 _33989_ (.a(_08580_),
    .b(_08581_),
    .c(_08582_),
    .d(_08583_),
    .e(_08584_),
    .f(_08586_),
    .o1(_08587_));
 b15nonb03ar1n02x5 _33990_ (.a(net933),
    .b(net914),
    .c(net921),
    .out0(_08588_));
 b15aoi012ah1n02x5 _33991_ (.a(_08588_),
    .b(_05969_),
    .c(net921),
    .o1(_08589_));
 b15nandp3ar1n02x5 _33992_ (.a(net930),
    .b(_05906_),
    .c(_06020_),
    .o1(_08590_));
 b15oa0022aq1n03x5 _33993_ (.a(_05911_),
    .b(_06435_),
    .c(_08589_),
    .d(_08590_),
    .o(_08591_));
 b15oab012ar1n02x5 _33994_ (.a(net934),
    .b(net931),
    .c(net917),
    .out0(_08592_));
 b15nor004ah1n04x5 _33995_ (.a(net915),
    .b(_05928_),
    .c(_05884_),
    .d(_08592_),
    .o1(_08593_));
 b15oai112ar1n02x5 _33996_ (.a(_06003_),
    .b(_05895_),
    .c(_06378_),
    .d(net921),
    .o1(_08594_));
 b15oab012al1n04x5 _33997_ (.a(_08593_),
    .b(_08594_),
    .c(_07605_),
    .out0(_08595_));
 b15nand04ar1n12x5 _33998_ (.a(_07672_),
    .b(_08587_),
    .c(_08591_),
    .d(_08595_),
    .o1(_08597_));
 b15ornc04as1n04x5 _33999_ (.a(_08564_),
    .b(_08573_),
    .c(_08579_),
    .d(_08597_),
    .o(_08598_));
 b15and002ar1n02x5 _34000_ (.a(\us00.a[1] ),
    .b(_07411_),
    .o(_08599_));
 b15oai012ar1n02x5 _34001_ (.a(net927),
    .b(_05827_),
    .c(_06046_),
    .o1(_08600_));
 b15aob012ar1n02x5 _34002_ (.a(_08600_),
    .b(_08157_),
    .c(\us00.a[0] ),
    .out0(_08601_));
 b15aoi112aq1n02x5 _34003_ (.a(net924),
    .b(_08599_),
    .c(_08601_),
    .d(_05821_),
    .o1(_08602_));
 b15nandp3ar1n02x5 _34004_ (.a(net931),
    .b(_05898_),
    .c(_05840_),
    .o1(_08603_));
 b15oaoi13an1n03x5 _34005_ (.a(\us00.a[0] ),
    .b(_08603_),
    .c(_06405_),
    .d(net931),
    .o1(_08604_));
 b15aoai13an1n08x5 _34006_ (.a(\us00.a[2] ),
    .b(_08604_),
    .c(_05915_),
    .d(net933),
    .o1(_08605_));
 b15aoi012ar1n02x5 _34007_ (.a(net930),
    .b(_05899_),
    .c(_05977_),
    .o1(_08606_));
 b15oaoi13aq1n02x5 _34008_ (.a(_07394_),
    .b(\us00.a[0] ),
    .c(_08157_),
    .d(_08606_),
    .o1(_08608_));
 b15aoi013aq1n04x5 _34009_ (.a(_08602_),
    .b(_08605_),
    .c(_08608_),
    .d(net924),
    .o1(_08609_));
 b15nona22an1n02x5 _34010_ (.a(net933),
    .b(net924),
    .c(net930),
    .out0(_08610_));
 b15oai012ar1n03x5 _34011_ (.a(net928),
    .b(_06034_),
    .c(_08610_),
    .o1(_08611_));
 b15norp03as1n03x5 _34012_ (.a(_05928_),
    .b(_05929_),
    .c(_06050_),
    .o1(_08612_));
 b15oaoi13ah1n02x5 _34013_ (.a(_08095_),
    .b(_05959_),
    .c(_05928_),
    .d(_05929_),
    .o1(_08613_));
 b15oaoi13as1n03x5 _34014_ (.a(_08611_),
    .b(_05969_),
    .c(_08612_),
    .d(_08613_),
    .o1(_08614_));
 b15aoai13ar1n02x5 _34015_ (.a(_05918_),
    .b(_08610_),
    .c(_05891_),
    .d(_05972_),
    .o1(_08615_));
 b15norp02an1n02x5 _34016_ (.a(_05972_),
    .b(_08095_),
    .o1(_08616_));
 b15oaoi13an1n03x5 _34017_ (.a(_08615_),
    .b(net933),
    .c(_08616_),
    .d(_08612_),
    .o1(_08617_));
 b15nanb02ar1n12x5 _34018_ (.a(\us00.a[5] ),
    .b(net917),
    .out0(_08619_));
 b15aoi012ah1n02x5 _34019_ (.a(_08619_),
    .b(_08115_),
    .c(_06449_),
    .o1(_08620_));
 b15norp03aq1n03x5 _34020_ (.a(net917),
    .b(_05894_),
    .c(_05935_),
    .o1(_08621_));
 b15oaoi13an1n04x5 _34021_ (.a(_05964_),
    .b(net914),
    .c(_08620_),
    .d(_08621_),
    .o1(_08622_));
 b15oaoi13as1n08x5 _34022_ (.a(_08614_),
    .b(_08617_),
    .c(_05911_),
    .d(_08622_),
    .o1(_08623_));
 b15norp03as1n08x5 _34023_ (.a(_06054_),
    .b(_06065_),
    .c(_08623_),
    .o1(_08624_));
 b15nona23as1n32x5 _34024_ (.a(_08598_),
    .b(_08609_),
    .c(_08624_),
    .d(_08328_),
    .out0(_08625_));
 b15nor003ah1n03x5 _34025_ (.a(_06201_),
    .b(_06089_),
    .c(_06125_),
    .o1(_08626_));
 b15oai013as1n08x5 _34026_ (.a(_06179_),
    .b(_06235_),
    .c(_06318_),
    .d(_08428_),
    .o1(_08627_));
 b15oai022aq1n06x5 _34027_ (.a(\us33.a[2] ),
    .b(_06125_),
    .c(_06197_),
    .d(net554),
    .o1(_08628_));
 b15aoi112an1n08x5 _34028_ (.a(_08626_),
    .b(_08627_),
    .c(_08628_),
    .d(net567),
    .o1(_08630_));
 b15xnr002aq1n12x5 _34029_ (.a(\us33.a[3] ),
    .b(net559),
    .out0(_08631_));
 b15oai022ar1n02x5 _34030_ (.a(_06125_),
    .b(_07010_),
    .c(_08631_),
    .d(_06197_),
    .o1(_08632_));
 b15norp02ar1n03x5 _34031_ (.a(_06179_),
    .b(_08632_),
    .o1(_08633_));
 b15aoi022as1n04x5 _34032_ (.a(_08417_),
    .b(_06221_),
    .c(_07025_),
    .d(net554),
    .o1(_08634_));
 b15oaoi13al1n08x5 _34033_ (.a(_08630_),
    .b(_08633_),
    .c(net566),
    .d(_08634_),
    .o1(_08635_));
 b15aoi012ar1n04x5 _34034_ (.a(_06158_),
    .b(_06313_),
    .c(net566),
    .o1(_08636_));
 b15aoi012ar1n04x5 _34035_ (.a(_08189_),
    .b(_06245_),
    .c(_06089_),
    .o1(_08637_));
 b15norp03ar1n24x5 _34036_ (.a(_06089_),
    .b(_06096_),
    .c(_06244_),
    .o1(_08638_));
 b15oab012ah1n03x5 _34037_ (.a(_08638_),
    .b(_07817_),
    .c(net566),
    .out0(_08639_));
 b15oai222aq1n16x5 _34038_ (.a(_06105_),
    .b(_08636_),
    .c(_08637_),
    .d(_07057_),
    .e(_08639_),
    .f(net555),
    .o1(_08641_));
 b15nandp3ah1n03x5 _34039_ (.a(net565),
    .b(net551),
    .c(\us33.a[7] ),
    .o1(_08642_));
 b15aoi112aq1n08x5 _34040_ (.a(_06108_),
    .b(_06235_),
    .c(_08441_),
    .d(_08642_),
    .o1(_08643_));
 b15oai013ah1n04x5 _34041_ (.a(net555),
    .b(_06174_),
    .c(_06287_),
    .d(_07813_),
    .o1(_08644_));
 b15oai022aq1n04x5 _34042_ (.a(_06218_),
    .b(_06135_),
    .c(_07828_),
    .d(_07823_),
    .o1(_08645_));
 b15aoi112ah1n04x5 _34043_ (.a(_08643_),
    .b(_08644_),
    .c(net560),
    .d(_08645_),
    .o1(_08646_));
 b15nano23an1n03x5 _34044_ (.a(net564),
    .b(_06206_),
    .c(_07780_),
    .d(net547),
    .out0(_08647_));
 b15aoi012as1n02x5 _34045_ (.a(_08647_),
    .b(_06333_),
    .c(_06313_),
    .o1(_08648_));
 b15aoi012an1n08x5 _34046_ (.a(_08646_),
    .b(_08648_),
    .c(_06201_),
    .o1(_08649_));
 b15nandp2aq1n02x5 _34047_ (.a(net560),
    .b(_06295_),
    .o1(_08650_));
 b15nor002ar1n02x5 _34048_ (.a(_07090_),
    .b(_06345_),
    .o1(_08652_));
 b15aoi013al1n04x5 _34049_ (.a(_08652_),
    .b(_07048_),
    .c(_06207_),
    .d(net547),
    .o1(_08653_));
 b15oaoi13as1n08x5 _34050_ (.a(_06201_),
    .b(_08650_),
    .c(_08653_),
    .d(_07828_),
    .o1(_08654_));
 b15nor004ah1n08x5 _34051_ (.a(_08635_),
    .b(_08641_),
    .c(_08649_),
    .d(_08654_),
    .o1(_08655_));
 b15aoi022an1n08x5 _34052_ (.a(_06220_),
    .b(_06243_),
    .c(_08423_),
    .d(_06264_),
    .o1(_08656_));
 b15norp02ar1n02x5 _34053_ (.a(_06243_),
    .b(_07024_),
    .o1(_08657_));
 b15nand02ar1n02x5 _34054_ (.a(_06111_),
    .b(_08631_),
    .o1(_08658_));
 b15oai112ar1n02x5 _34055_ (.a(net562),
    .b(_08658_),
    .c(_07804_),
    .d(_06111_),
    .o1(_08659_));
 b15oa0022aq1n03x5 _34056_ (.a(net562),
    .b(_08656_),
    .c(_08657_),
    .d(_08659_),
    .o(_08660_));
 b15nand02ar1n02x5 _34057_ (.a(\us33.a[3] ),
    .b(_06313_),
    .o1(_08661_));
 b15oaoi13ar1n03x5 _34058_ (.a(\us33.a[0] ),
    .b(_08661_),
    .c(_06195_),
    .d(\us33.a[3] ),
    .o1(_08663_));
 b15nanb03ar1n06x5 _34059_ (.a(net552),
    .b(net548),
    .c(net554),
    .out0(_08664_));
 b15oai012aq1n06x5 _34060_ (.a(_08664_),
    .b(_06135_),
    .c(net554),
    .o1(_08665_));
 b15aoi122ar1n04x5 _34061_ (.a(_08663_),
    .b(_08665_),
    .c(_07069_),
    .d(_06240_),
    .e(_06221_),
    .o1(_08666_));
 b15aoi022ah1n04x5 _34062_ (.a(\us33.a[3] ),
    .b(_06240_),
    .c(_06245_),
    .d(_06127_),
    .o1(_08667_));
 b15oaoi13as1n08x5 _34063_ (.a(net562),
    .b(_08666_),
    .c(_08667_),
    .d(_06111_),
    .o1(_08668_));
 b15nor003ar1n02x5 _34064_ (.a(\us33.a[0] ),
    .b(net557),
    .c(net550),
    .o1(_08669_));
 b15nor003aq1n04x5 _34065_ (.a(_06096_),
    .b(_07020_),
    .c(_08669_),
    .o1(_08670_));
 b15orn003al1n03x5 _34066_ (.a(_07797_),
    .b(_08423_),
    .c(_08638_),
    .o(_08671_));
 b15oai022aq1n04x5 _34067_ (.a(_06230_),
    .b(_07856_),
    .c(_06339_),
    .d(_07030_),
    .o1(_08672_));
 b15aoi022an1n12x5 _34068_ (.a(_08670_),
    .b(_08671_),
    .c(_08672_),
    .d(_06201_),
    .o1(_08674_));
 b15nonb02al1n08x5 _34069_ (.a(net558),
    .b(\us33.a[5] ),
    .out0(_08675_));
 b15nand04ah1n08x5 _34070_ (.a(\us33.a[7] ),
    .b(_06264_),
    .c(_08675_),
    .d(_08435_),
    .o1(_08676_));
 b15orn003al1n02x5 _34071_ (.a(_06089_),
    .b(_06298_),
    .c(_06300_),
    .o(_08677_));
 b15nandp3aq1n03x5 _34072_ (.a(_06324_),
    .b(_06193_),
    .c(_06242_),
    .o1(_08678_));
 b15oai112aq1n08x5 _34073_ (.a(_08676_),
    .b(_08677_),
    .c(_08397_),
    .d(_08678_),
    .o1(_08679_));
 b15nor004al1n02x5 _34074_ (.a(net555),
    .b(net547),
    .c(net551),
    .d(\us33.a[6] ),
    .o1(_08680_));
 b15aoi013ah1n02x5 _34075_ (.a(_08680_),
    .b(_08201_),
    .c(net547),
    .d(_06111_),
    .o1(_08681_));
 b15nano23aq1n06x5 _34076_ (.a(net558),
    .b(net544),
    .c(_08681_),
    .d(net563),
    .out0(_08682_));
 b15oai022ar1n02x5 _34077_ (.a(net551),
    .b(_06218_),
    .c(_06103_),
    .d(_06318_),
    .o1(_08683_));
 b15and003as1n02x5 _34078_ (.a(net547),
    .b(_07033_),
    .c(_08683_),
    .o(_08685_));
 b15nonb03ar1n03x5 _34079_ (.a(net558),
    .b(\us33.a[7] ),
    .c(net553),
    .out0(_08686_));
 b15nano23al1n03x5 _34080_ (.a(\us33.a[5] ),
    .b(net551),
    .c(\us33.a[6] ),
    .d(net560),
    .out0(_08687_));
 b15aoai13an1n08x5 _34081_ (.a(_08686_),
    .b(_08687_),
    .c(_08435_),
    .d(_06257_),
    .o1(_08688_));
 b15nandp3an1n08x5 _34082_ (.a(net544),
    .b(_06324_),
    .c(_06333_),
    .o1(_08689_));
 b15nandp2aq1n03x5 _34083_ (.a(net555),
    .b(net545),
    .o1(_08690_));
 b15oai122ar1n16x5 _34084_ (.a(_08688_),
    .b(_08689_),
    .c(_08690_),
    .d(_07063_),
    .e(net560),
    .o1(_08691_));
 b15nor004as1n08x5 _34085_ (.a(_08679_),
    .b(_08682_),
    .c(_08685_),
    .d(_08691_),
    .o1(_08692_));
 b15oai022aq1n02x5 _34086_ (.a(net564),
    .b(_06105_),
    .c(_07797_),
    .d(net555),
    .o1(_08693_));
 b15oai022an1n02x5 _34087_ (.a(net560),
    .b(_07804_),
    .c(_07093_),
    .d(_06155_),
    .o1(_08694_));
 b15oai012as1n06x5 _34088_ (.a(_06302_),
    .b(_08693_),
    .c(_08694_),
    .o1(_08696_));
 b15oai022as1n02x5 _34089_ (.a(_06127_),
    .b(_06230_),
    .c(_07100_),
    .d(_06310_),
    .o1(_08697_));
 b15oai022ah1n02x5 _34090_ (.a(net557),
    .b(_07838_),
    .c(_08689_),
    .d(net545),
    .o1(_08698_));
 b15aoi022an1n08x5 _34091_ (.a(net564),
    .b(_08697_),
    .c(_08698_),
    .d(_06264_),
    .o1(_08699_));
 b15nand04as1n16x5 _34092_ (.a(_08674_),
    .b(_08692_),
    .c(_08696_),
    .d(_08699_),
    .o1(_08700_));
 b15nano23as1n24x5 _34093_ (.a(_08655_),
    .b(_08660_),
    .c(_08668_),
    .d(_08700_),
    .out0(_08701_));
 b15xnr002ar1n03x5 _34094_ (.a(_08383_),
    .b(_08701_),
    .out0(_08702_));
 b15xor002al1n02x5 _34095_ (.a(_08625_),
    .b(_08702_),
    .out0(_08703_));
 b15nor002ah1n02x5 _34096_ (.a(net681),
    .b(_07282_),
    .o1(_08704_));
 b15nandp2ar1n08x5 _34097_ (.a(net688),
    .b(_07372_),
    .o1(_08705_));
 b15aoi013al1n03x5 _34098_ (.a(net679),
    .b(_06769_),
    .c(_07984_),
    .d(_08705_),
    .o1(_08707_));
 b15oai012ah1n08x5 _34099_ (.a(_06792_),
    .b(_08704_),
    .c(_08707_),
    .o1(_08708_));
 b15nandp3ah1n03x5 _34100_ (.a(net669),
    .b(_06777_),
    .c(_07928_),
    .o1(_08709_));
 b15aoi013ah1n02x5 _34101_ (.a(_06792_),
    .b(net678),
    .c(_07387_),
    .d(_08709_),
    .o1(_08710_));
 b15oai012ar1n03x5 _34102_ (.a(_08501_),
    .b(_07269_),
    .c(_06786_),
    .o1(_08711_));
 b15oai022al1n04x5 _34103_ (.a(_06858_),
    .b(_06778_),
    .c(_06980_),
    .d(_06906_),
    .o1(_08712_));
 b15aoi022ah1n04x5 _34104_ (.a(_08710_),
    .b(_08711_),
    .c(_08712_),
    .d(_07901_),
    .o1(_08713_));
 b15nand04ar1n02x5 _34105_ (.a(_06792_),
    .b(_06896_),
    .c(_06768_),
    .d(_06980_),
    .o1(_08714_));
 b15nand02ar1n02x5 _34106_ (.a(_06866_),
    .b(_07348_),
    .o1(_08715_));
 b15aoi012ah1n02x5 _34107_ (.a(net678),
    .b(_08714_),
    .c(_08715_),
    .o1(_08716_));
 b15aoi012ar1n02x5 _34108_ (.a(_06786_),
    .b(_06977_),
    .c(_07906_),
    .o1(_08718_));
 b15nano23aq1n03x5 _34109_ (.a(_06999_),
    .b(_07366_),
    .c(_08718_),
    .d(_06849_),
    .out0(_08719_));
 b15nandp2ar1n02x5 _34110_ (.a(net679),
    .b(_06748_),
    .o1(_08720_));
 b15nandp2ar1n02x5 _34111_ (.a(_07364_),
    .b(_07348_),
    .o1(_08721_));
 b15oaoi13an1n04x5 _34112_ (.a(_08720_),
    .b(_08721_),
    .c(_06758_),
    .d(_06906_),
    .o1(_08722_));
 b15nor004aq1n08x5 _34113_ (.a(_06861_),
    .b(_08716_),
    .c(_08719_),
    .d(_08722_),
    .o1(_08723_));
 b15norp02aq1n02x5 _34114_ (.a(_06915_),
    .b(_07344_),
    .o1(_08724_));
 b15aoai13an1n02x5 _34115_ (.a(_06914_),
    .b(_08724_),
    .c(_06924_),
    .d(_06915_),
    .o1(_08725_));
 b15oai112an1n04x5 _34116_ (.a(_06758_),
    .b(_06915_),
    .c(_06940_),
    .d(_06993_),
    .o1(_08726_));
 b15oai022aq1n06x5 _34117_ (.a(net680),
    .b(_06783_),
    .c(_07899_),
    .d(_06984_),
    .o1(_08727_));
 b15nandp3as1n03x5 _34118_ (.a(_06822_),
    .b(_07361_),
    .c(_08727_),
    .o1(_08729_));
 b15andc04ah1n03x5 _34119_ (.a(_07349_),
    .b(_08725_),
    .c(_08726_),
    .d(_08729_),
    .o(_08730_));
 b15nand04an1n16x5 _34120_ (.a(_08708_),
    .b(_08713_),
    .c(_08723_),
    .d(_08730_),
    .o1(_08731_));
 b15nand02an1n08x5 _34121_ (.a(_07372_),
    .b(_07901_),
    .o1(_08732_));
 b15nand04as1n03x5 _34122_ (.a(net678),
    .b(_06822_),
    .c(_06839_),
    .d(_06775_),
    .o1(_08733_));
 b15oai112ar1n12x5 _34123_ (.a(_08732_),
    .b(_08733_),
    .c(_07377_),
    .d(_07269_),
    .o1(_08734_));
 b15oai012an1n02x5 _34124_ (.a(_06786_),
    .b(_07356_),
    .c(_07910_),
    .o1(_08735_));
 b15nor003ah1n06x5 _34125_ (.a(net686),
    .b(net682),
    .c(net679),
    .o1(_08736_));
 b15aoi012an1n04x5 _34126_ (.a(_06786_),
    .b(_06924_),
    .c(_08736_),
    .o1(_08737_));
 b15oai112al1n12x5 _34127_ (.a(_07576_),
    .b(_08737_),
    .c(net681),
    .d(_07282_),
    .o1(_08738_));
 b15aoi012ar1n02x5 _34128_ (.a(_07338_),
    .b(_06841_),
    .c(_06778_),
    .o1(_08740_));
 b15oai022aq1n06x5 _34129_ (.a(_08734_),
    .b(_08735_),
    .c(_08738_),
    .d(_08740_),
    .o1(_08741_));
 b15aoi022an1n06x5 _34130_ (.a(_06927_),
    .b(_07943_),
    .c(_07907_),
    .d(_08495_),
    .o1(_08742_));
 b15nano22ar1n05x5 _34131_ (.a(net672),
    .b(\us22.a[0] ),
    .c(net679),
    .out0(_08743_));
 b15aoi022al1n12x5 _34132_ (.a(_06777_),
    .b(_06950_),
    .c(_08743_),
    .d(_06839_),
    .o1(_08744_));
 b15obai22ar1n12x5 _34133_ (.a(_08506_),
    .b(_08742_),
    .c(_08744_),
    .d(net669),
    .out0(_08745_));
 b15oai112an1n12x5 _34134_ (.a(_06826_),
    .b(_07984_),
    .c(_07282_),
    .d(_06792_),
    .o1(_08746_));
 b15aoi012ar1n02x5 _34135_ (.a(net689),
    .b(net678),
    .c(_07387_),
    .o1(_08747_));
 b15aoi022as1n04x5 _34136_ (.a(net683),
    .b(_08745_),
    .c(_08746_),
    .d(_08747_),
    .o1(_08748_));
 b15aoi013ar1n02x5 _34137_ (.a(net677),
    .b(_06767_),
    .c(_06768_),
    .d(net689),
    .o1(_08749_));
 b15oaoi13ar1n03x5 _34138_ (.a(_08749_),
    .b(_06769_),
    .c(_07269_),
    .d(_06792_),
    .o1(_08751_));
 b15nano22aq1n02x5 _34139_ (.a(\us22.a[4] ),
    .b(\us22.a[6] ),
    .c(net670),
    .out0(_08752_));
 b15aoai13an1n06x5 _34140_ (.a(_07906_),
    .b(_08752_),
    .c(_07948_),
    .d(_06822_),
    .o1(_08753_));
 b15oaoi13aq1n08x5 _34141_ (.a(\us22.a[5] ),
    .b(_08753_),
    .c(_06965_),
    .d(_06936_),
    .o1(_08754_));
 b15oai122ar1n12x5 _34142_ (.a(_06786_),
    .b(_06826_),
    .c(_06901_),
    .d(_06990_),
    .e(_06854_),
    .o1(_08755_));
 b15nandp3an1n02x5 _34143_ (.a(_06777_),
    .b(_06852_),
    .c(_07361_),
    .o1(_08756_));
 b15oai112ar1n08x5 _34144_ (.a(net689),
    .b(_08756_),
    .c(_07361_),
    .d(_06878_),
    .o1(_08757_));
 b15aoi112an1n04x5 _34145_ (.a(_08751_),
    .b(_08754_),
    .c(_08755_),
    .d(_08757_),
    .o1(_08758_));
 b15oai112al1n12x5 _34146_ (.a(_08741_),
    .b(_08748_),
    .c(net683),
    .d(_08758_),
    .o1(_08759_));
 b15nandp3ar1n02x5 _34147_ (.a(net671),
    .b(_07277_),
    .c(_07288_),
    .o1(_08760_));
 b15aoi022al1n02x5 _34148_ (.a(_07277_),
    .b(_06852_),
    .c(_06960_),
    .d(\us22.a[7] ),
    .o1(_08761_));
 b15oaoi13ar1n02x5 _34149_ (.a(_07319_),
    .b(_08760_),
    .c(_08761_),
    .d(_07948_),
    .o1(_08762_));
 b15norp02ar1n02x5 _34150_ (.a(_08468_),
    .b(_07269_),
    .o1(_08763_));
 b15oab012al1n04x5 _34151_ (.a(_06792_),
    .b(_08762_),
    .c(_08763_),
    .out0(_08764_));
 b15norp03al1n03x5 _34152_ (.a(_06882_),
    .b(_06921_),
    .c(_06800_),
    .o1(_08765_));
 b15oai022aq1n02x5 _34153_ (.a(_06800_),
    .b(_07512_),
    .c(_08484_),
    .d(_06863_),
    .o1(_08766_));
 b15aoai13as1n04x5 _34154_ (.a(\us22.a[6] ),
    .b(_08765_),
    .c(_08766_),
    .d(net673),
    .o1(_08767_));
 b15oaoi13aq1n04x5 _34155_ (.a(_06786_),
    .b(_08767_),
    .c(_07269_),
    .d(_06800_),
    .o1(_08768_));
 b15aoi112an1n04x5 _34156_ (.a(net689),
    .b(net683),
    .c(_06906_),
    .d(_06973_),
    .o1(_08769_));
 b15oai013aq1n12x5 _34157_ (.a(net677),
    .b(_08764_),
    .c(_08768_),
    .d(_08769_),
    .o1(_08770_));
 b15nona22as1n32x5 _34158_ (.a(_08731_),
    .b(_08759_),
    .c(_08770_),
    .out0(_08772_));
 b15aoi022ar1n02x5 _34159_ (.a(_06574_),
    .b(_07250_),
    .c(_07251_),
    .d(_06631_),
    .o1(_08773_));
 b15oai022ah1n04x5 _34160_ (.a(_06605_),
    .b(_06627_),
    .c(_08773_),
    .d(net820),
    .o1(_08774_));
 b15nandp3as1n08x5 _34161_ (.a(net804),
    .b(_07249_),
    .c(_08774_),
    .o1(_08775_));
 b15aoi112ar1n02x5 _34162_ (.a(\us11.a[0] ),
    .b(_06632_),
    .c(_06587_),
    .d(_06686_),
    .o1(_08776_));
 b15aoai13ar1n04x5 _34163_ (.a(_06650_),
    .b(_08776_),
    .c(_08255_),
    .d(\us11.a[0] ),
    .o1(_08777_));
 b15aoi112ar1n02x5 _34164_ (.a(\us11.a[3] ),
    .b(_06624_),
    .c(_06600_),
    .d(_06661_),
    .o1(_08778_));
 b15aoai13an1n03x5 _34165_ (.a(net813),
    .b(_08778_),
    .c(_07996_),
    .d(_06624_),
    .o1(_08779_));
 b15nand03as1n08x5 _34166_ (.a(_08775_),
    .b(_08777_),
    .c(_08779_),
    .o1(_08780_));
 b15aoai13ar1n03x5 _34167_ (.a(_06567_),
    .b(_06606_),
    .c(\us11.a[0] ),
    .d(_07206_),
    .o1(_08781_));
 b15aoi022an1n04x5 _34168_ (.a(net813),
    .b(_07206_),
    .c(_06606_),
    .d(_06476_),
    .o1(_08783_));
 b15oaoi13ah1n04x5 _34169_ (.a(\us11.a[3] ),
    .b(_08781_),
    .c(_08783_),
    .d(_06632_),
    .o1(_08784_));
 b15oai112ar1n04x5 _34170_ (.a(\us11.a[3] ),
    .b(_06593_),
    .c(_06631_),
    .d(_06709_),
    .o1(_08785_));
 b15oai013ar1n02x5 _34171_ (.a(_08785_),
    .b(_08254_),
    .c(_07169_),
    .d(\us11.a[3] ),
    .o1(_08786_));
 b15oai022an1n02x5 _34172_ (.a(net805),
    .b(net811),
    .c(_06525_),
    .d(_07155_),
    .o1(_08787_));
 b15aoi012as1n04x5 _34173_ (.a(_06476_),
    .b(_06533_),
    .c(_08787_),
    .o1(_08788_));
 b15and002aq1n02x5 _34174_ (.a(_08786_),
    .b(_08788_),
    .o(_08789_));
 b15aoi122al1n06x5 _34175_ (.a(net819),
    .b(net810),
    .c(_06509_),
    .d(_06676_),
    .e(_06548_),
    .o1(_08790_));
 b15oai012ah1n04x5 _34176_ (.a(_06558_),
    .b(_06709_),
    .c(_07155_),
    .o1(_08791_));
 b15aoi012an1n02x5 _34177_ (.a(_07169_),
    .b(_08791_),
    .c(_06476_),
    .o1(_08792_));
 b15oai022aq1n08x5 _34178_ (.a(_08789_),
    .b(_08790_),
    .c(_08792_),
    .d(net813),
    .o1(_08794_));
 b15oai112ar1n02x5 _34179_ (.a(_06545_),
    .b(_06682_),
    .c(_06565_),
    .d(net797),
    .o1(_08795_));
 b15oai022as1n02x5 _34180_ (.a(_06703_),
    .b(_06639_),
    .c(_06698_),
    .d(_08795_),
    .o1(_08796_));
 b15aoai13ar1n02x5 _34181_ (.a(_07232_),
    .b(_06682_),
    .c(_06577_),
    .d(net799),
    .o1(_08797_));
 b15oai112ar1n04x5 _34182_ (.a(_06605_),
    .b(_06700_),
    .c(net820),
    .d(_06514_),
    .o1(_08798_));
 b15nandp2ar1n04x5 _34183_ (.a(_08797_),
    .b(_08798_),
    .o1(_08799_));
 b15oai012ah1n08x5 _34184_ (.a(_06536_),
    .b(_08796_),
    .c(_08799_),
    .o1(_08800_));
 b15oai012ar1n02x5 _34185_ (.a(net809),
    .b(_06645_),
    .c(_06722_),
    .o1(_08801_));
 b15oai012an1n02x5 _34186_ (.a(net820),
    .b(_06518_),
    .c(_07245_),
    .o1(_08802_));
 b15oai022ar1n02x5 _34187_ (.a(net809),
    .b(_06580_),
    .c(_06705_),
    .d(_06574_),
    .o1(_08803_));
 b15nano22ar1n03x5 _34188_ (.a(_08801_),
    .b(_08802_),
    .c(_08803_),
    .out0(_08805_));
 b15aoi012ar1n02x5 _34189_ (.a(_06659_),
    .b(_06610_),
    .c(_06587_),
    .o1(_08806_));
 b15nand03ah1n03x5 _34190_ (.a(_06632_),
    .b(_06586_),
    .c(_06555_),
    .o1(_08807_));
 b15oai012ar1n12x5 _34191_ (.a(_08807_),
    .b(_06610_),
    .c(_06632_),
    .o1(_08808_));
 b15oaoi13ah1n04x5 _34192_ (.a(_08805_),
    .b(_08806_),
    .c(_08808_),
    .d(net820),
    .o1(_08809_));
 b15oaoi13aq1n02x5 _34193_ (.a(_06628_),
    .b(_06589_),
    .c(_06610_),
    .d(_06703_),
    .o1(_08810_));
 b15oai012ar1n02x5 _34194_ (.a(net808),
    .b(_06514_),
    .c(_06476_),
    .o1(_08811_));
 b15oaoi13al1n02x5 _34195_ (.a(_08811_),
    .b(_06558_),
    .c(_06728_),
    .d(_06565_),
    .o1(_08812_));
 b15orn003ar1n02x5 _34196_ (.a(_07749_),
    .b(_06645_),
    .c(_07754_),
    .o(_08813_));
 b15oaoi13ar1n03x5 _34197_ (.a(_07210_),
    .b(_08813_),
    .c(_06675_),
    .d(_08049_),
    .o1(_08814_));
 b15norp03as1n04x5 _34198_ (.a(_08810_),
    .b(_08812_),
    .c(_08814_),
    .o1(_08816_));
 b15nandp2ar1n03x5 _34199_ (.a(_06538_),
    .b(_06499_),
    .o1(_08817_));
 b15aoi022al1n04x5 _34200_ (.a(_06527_),
    .b(_06545_),
    .c(_06539_),
    .d(_06624_),
    .o1(_08818_));
 b15nandp2ar1n03x5 _34201_ (.a(_06577_),
    .b(_07173_),
    .o1(_08819_));
 b15aoi012an1n02x5 _34202_ (.a(_06652_),
    .b(_06553_),
    .c(_06552_),
    .o1(_08820_));
 b15oai022ah1n06x5 _34203_ (.a(_08817_),
    .b(_08818_),
    .c(_08819_),
    .d(_08820_),
    .o1(_08821_));
 b15nand04as1n02x5 _34204_ (.a(_06476_),
    .b(_06539_),
    .c(_06638_),
    .d(_06628_),
    .o1(_08822_));
 b15aob012ar1n03x5 _34205_ (.a(_08008_),
    .b(_07225_),
    .c(_06632_),
    .out0(_08823_));
 b15oai112ah1n06x5 _34206_ (.a(_06653_),
    .b(_08822_),
    .c(_08823_),
    .d(_06661_),
    .o1(_08824_));
 b15nand04ar1n02x5 _34207_ (.a(_06476_),
    .b(_06501_),
    .c(_06556_),
    .d(_06650_),
    .o1(_08825_));
 b15oaoi13aq1n03x5 _34208_ (.a(net815),
    .b(_08825_),
    .c(_06628_),
    .d(_06686_),
    .o1(_08827_));
 b15nor004an1n08x5 _34209_ (.a(_06630_),
    .b(_08821_),
    .c(_08824_),
    .d(_08827_),
    .o1(_08828_));
 b15nand04as1n16x5 _34210_ (.a(_08800_),
    .b(_08809_),
    .c(_08816_),
    .d(_08828_),
    .o1(_08829_));
 b15nor004as1n12x5 _34211_ (.a(_08780_),
    .b(_08784_),
    .c(_08794_),
    .d(_08829_),
    .o1(_08830_));
 b15xor002an1n16x5 _34212_ (.a(_08772_),
    .b(_08830_),
    .out0(_08831_));
 b15xor002ar1n02x5 _34213_ (.a(_08703_),
    .b(_08831_),
    .out0(_08832_));
 b15cmbn22an1n04x5 _34214_ (.clk1(\text_in_r[101] ),
    .clk2(_08832_),
    .clkout(_08833_),
    .s(net535));
 b15xor002al1n02x5 _34215_ (.a(\u0.w[0][5] ),
    .b(_08833_),
    .out0(_00102_));
 b15nand02ar1n02x5 _34216_ (.a(net538),
    .b(\text_in_r[102] ),
    .o1(_08834_));
 b15oaoi13aq1n03x5 _34217_ (.a(_07378_),
    .b(_07576_),
    .c(net689),
    .d(_06867_),
    .o1(_08835_));
 b15oaoi13ar1n02x5 _34218_ (.a(_07580_),
    .b(_06945_),
    .c(_07282_),
    .d(net678),
    .o1(_08837_));
 b15norp03ar1n02x5 _34219_ (.a(net678),
    .b(_07282_),
    .c(_06748_),
    .o1(_08838_));
 b15nor004al1n02x5 _34220_ (.a(net681),
    .b(_08835_),
    .c(_08837_),
    .d(_08838_),
    .o1(_08839_));
 b15norp02ar1n02x5 _34221_ (.a(_06862_),
    .b(_07580_),
    .o1(_08840_));
 b15oaoi13ar1n02x5 _34222_ (.a(_06786_),
    .b(_08732_),
    .c(_06906_),
    .d(net684),
    .o1(_08841_));
 b15aoi112ar1n02x5 _34223_ (.a(_08840_),
    .b(_08841_),
    .c(net678),
    .d(_06844_),
    .o1(_08842_));
 b15aoi012ar1n02x5 _34224_ (.a(_08839_),
    .b(_08842_),
    .c(net681),
    .o1(_08843_));
 b15nand02ar1n02x5 _34225_ (.a(net679),
    .b(_06859_),
    .o1(_08844_));
 b15oai012ar1n02x5 _34226_ (.a(_07372_),
    .b(_07546_),
    .c(_06786_),
    .o1(_08845_));
 b15oaoi13an1n03x5 _34227_ (.a(_08844_),
    .b(_08845_),
    .c(_07546_),
    .d(_06769_),
    .o1(_08846_));
 b15nand02ar1n02x5 _34228_ (.a(_06792_),
    .b(_07364_),
    .o1(_08848_));
 b15oaoi13ah1n02x5 _34229_ (.a(_06858_),
    .b(_08848_),
    .c(_07282_),
    .d(_06826_),
    .o1(_08849_));
 b15oai112al1n12x5 _34230_ (.a(_06823_),
    .b(_07365_),
    .c(_06966_),
    .d(_06999_),
    .o1(_08850_));
 b15nandp2ah1n03x5 _34231_ (.a(_07942_),
    .b(_08495_),
    .o1(_08851_));
 b15nor003as1n04x5 _34232_ (.a(_06790_),
    .b(_08494_),
    .c(_08506_),
    .o1(_08852_));
 b15oai022aq1n16x5 _34233_ (.a(_06826_),
    .b(_08850_),
    .c(_08851_),
    .d(_08852_),
    .o1(_08853_));
 b15nor004al1n06x5 _34234_ (.a(_06962_),
    .b(_08846_),
    .c(_08849_),
    .d(_08853_),
    .o1(_08854_));
 b15nand02ar1n02x5 _34235_ (.a(net681),
    .b(_07364_),
    .o1(_08855_));
 b15oaoi13al1n02x5 _34236_ (.a(_06826_),
    .b(_08855_),
    .c(_06981_),
    .d(_06792_),
    .o1(_08856_));
 b15aoai13al1n04x5 _34237_ (.a(net688),
    .b(_08856_),
    .c(_06849_),
    .d(_08490_),
    .o1(_08857_));
 b15oai112as1n04x5 _34238_ (.a(_06826_),
    .b(_07278_),
    .c(_06981_),
    .d(net684),
    .o1(_08859_));
 b15oai022al1n04x5 _34239_ (.a(net681),
    .b(_06906_),
    .c(_07344_),
    .d(_07508_),
    .o1(_08860_));
 b15oai012ah1n03x5 _34240_ (.a(_08859_),
    .b(_08860_),
    .c(_06826_),
    .o1(_08861_));
 b15nandp3al1n08x5 _34241_ (.a(_06822_),
    .b(_06839_),
    .c(_08736_),
    .o1(_08862_));
 b15aoi013as1n06x5 _34242_ (.a(net688),
    .b(_06777_),
    .c(_06852_),
    .d(_07906_),
    .o1(_08863_));
 b15aoi013aq1n06x5 _34243_ (.a(_06786_),
    .b(_06822_),
    .c(_06839_),
    .d(_07363_),
    .o1(_08864_));
 b15norp03ar1n04x5 _34244_ (.a(net672),
    .b(net682),
    .c(net679),
    .o1(_08865_));
 b15aoai13an1n08x5 _34245_ (.a(_06876_),
    .b(_08865_),
    .c(_06889_),
    .d(net672),
    .o1(_08866_));
 b15aoi022an1n24x5 _34246_ (.a(_08862_),
    .b(_08863_),
    .c(_08864_),
    .d(_08866_),
    .o1(_08867_));
 b15norp03ar1n04x5 _34247_ (.a(net675),
    .b(_06826_),
    .c(_07302_),
    .o1(_08868_));
 b15oai012ar1n02x5 _34248_ (.a(_06800_),
    .b(_06863_),
    .c(net689),
    .o1(_08870_));
 b15oai012ar1n02x5 _34249_ (.a(_07279_),
    .b(_06859_),
    .c(net689),
    .o1(_08871_));
 b15aoi022aq1n04x5 _34250_ (.a(net674),
    .b(_08870_),
    .c(_08871_),
    .d(_07910_),
    .o1(_08872_));
 b15aoi112ah1n04x5 _34251_ (.a(_07541_),
    .b(_08867_),
    .c(_08868_),
    .d(_08872_),
    .o1(_08873_));
 b15nand04al1n12x5 _34252_ (.a(_08854_),
    .b(_08857_),
    .c(_08861_),
    .d(_08873_),
    .o1(_08874_));
 b15orn002ar1n08x5 _34253_ (.a(_08843_),
    .b(_08874_),
    .o(_08875_));
 b15oai012ah1n03x5 _34254_ (.a(_07332_),
    .b(_07545_),
    .c(_06792_),
    .o1(_08876_));
 b15aoai13an1n06x5 _34255_ (.a(net681),
    .b(_07582_),
    .c(_08876_),
    .d(net689),
    .o1(_08877_));
 b15aoi012ah1n02x5 _34256_ (.a(net677),
    .b(_06784_),
    .c(net684),
    .o1(_08878_));
 b15oai122as1n08x5 _34257_ (.a(_08878_),
    .b(_06915_),
    .c(_06906_),
    .d(net689),
    .e(_06878_),
    .o1(_08879_));
 b15oai012al1n06x5 _34258_ (.a(_07384_),
    .b(_07910_),
    .c(_06786_),
    .o1(_08881_));
 b15oai022as1n02x5 _34259_ (.a(net681),
    .b(_07545_),
    .c(_07910_),
    .d(net684),
    .o1(_08882_));
 b15aoi222as1n08x5 _34260_ (.a(net681),
    .b(_08879_),
    .c(_08881_),
    .d(_07291_),
    .e(_08882_),
    .f(_06786_),
    .o1(_08883_));
 b15aoi012al1n08x5 _34261_ (.a(net677),
    .b(_08877_),
    .c(_08883_),
    .o1(_08884_));
 b15aoai13al1n02x5 _34262_ (.a(net689),
    .b(_06844_),
    .c(_06807_),
    .d(_06758_),
    .o1(_08885_));
 b15oai112ar1n06x5 _34263_ (.a(_06826_),
    .b(_08885_),
    .c(_07344_),
    .d(net684),
    .o1(_08886_));
 b15nand04ah1n03x5 _34264_ (.a(_06786_),
    .b(_06758_),
    .c(_06852_),
    .d(_06839_),
    .o1(_08887_));
 b15oai012as1n03x5 _34265_ (.a(_08887_),
    .b(_07273_),
    .c(_06792_),
    .o1(_08888_));
 b15nand03as1n08x5 _34266_ (.a(net682),
    .b(_06852_),
    .c(_06839_),
    .o1(_08889_));
 b15oaoi13aq1n08x5 _34267_ (.a(_06850_),
    .b(_08889_),
    .c(_07269_),
    .d(net681),
    .o1(_08890_));
 b15oai013ah1n06x5 _34268_ (.a(_08886_),
    .b(_08888_),
    .c(_08890_),
    .d(_06826_),
    .o1(_08892_));
 b15nand02al1n03x5 _34269_ (.a(net685),
    .b(_06862_),
    .o1(_08893_));
 b15nand02ar1n02x5 _34270_ (.a(net681),
    .b(_06924_),
    .o1(_08894_));
 b15oai013ah1n03x5 _34271_ (.a(_08894_),
    .b(_06769_),
    .c(net677),
    .d(net681),
    .o1(_08895_));
 b15oai112ar1n12x5 _34272_ (.a(net689),
    .b(_08893_),
    .c(_08895_),
    .d(net685),
    .o1(_08896_));
 b15oai012ar1n03x5 _34273_ (.a(_06906_),
    .b(_08705_),
    .c(net678),
    .o1(_08897_));
 b15oai012ar1n02x5 _34274_ (.a(_06906_),
    .b(_06981_),
    .c(_06758_),
    .o1(_08898_));
 b15aoi022as1n04x5 _34275_ (.a(_06758_),
    .b(_08897_),
    .c(_08898_),
    .d(net678),
    .o1(_08899_));
 b15oai112an1n16x5 _34276_ (.a(_08892_),
    .b(_08896_),
    .c(_08899_),
    .d(net685),
    .o1(_08900_));
 b15norp03as1n24x5 _34277_ (.a(_08875_),
    .b(_08884_),
    .c(_08900_),
    .o1(_08901_));
 b15norp03aq1n02x5 _34278_ (.a(_06096_),
    .b(_06244_),
    .c(_07804_),
    .o1(_08903_));
 b15norp03as1n04x5 _34279_ (.a(_06171_),
    .b(_06287_),
    .c(_07011_),
    .o1(_08904_));
 b15nor003al1n02x5 _34280_ (.a(_06145_),
    .b(_06135_),
    .c(_06287_),
    .o1(_08905_));
 b15nanb03ar1n04x5 _34281_ (.a(\us33.a[6] ),
    .b(\us33.a[7] ),
    .c(net554),
    .out0(_08906_));
 b15oaoi13aq1n08x5 _34282_ (.a(_08906_),
    .b(_06187_),
    .c(\us33.a[4] ),
    .d(_08675_),
    .o1(_08907_));
 b15nor004al1n04x5 _34283_ (.a(_08903_),
    .b(_08904_),
    .c(_08905_),
    .d(_08907_),
    .o1(_08908_));
 b15aoai13an1n03x5 _34284_ (.a(_06111_),
    .b(_08459_),
    .c(_08638_),
    .d(net554),
    .o1(_08909_));
 b15aoai13al1n03x5 _34285_ (.a(_06111_),
    .b(_08189_),
    .c(_08417_),
    .d(net559),
    .o1(_08910_));
 b15aoi013an1n04x5 _34286_ (.a(_06179_),
    .b(_08908_),
    .c(_08909_),
    .d(_08910_),
    .o1(_08911_));
 b15oaoi13as1n02x5 _34287_ (.a(_06197_),
    .b(_07045_),
    .c(_08631_),
    .d(\us33.a[0] ),
    .o1(_08912_));
 b15norp03al1n02x5 _34288_ (.a(_06096_),
    .b(_06244_),
    .c(_06155_),
    .o1(_08914_));
 b15norp02ar1n02x5 _34289_ (.a(_07804_),
    .b(_06197_),
    .o1(_08915_));
 b15oaoi13as1n02x5 _34290_ (.a(_08912_),
    .b(_06179_),
    .c(_08914_),
    .d(_08915_),
    .o1(_08916_));
 b15nand02ar1n02x5 _34291_ (.a(net559),
    .b(_06312_),
    .o1(_08917_));
 b15oai013al1n03x5 _34292_ (.a(_08664_),
    .b(_07804_),
    .c(_06135_),
    .d(net562),
    .o1(_08918_));
 b15norp02ar1n02x5 _34293_ (.a(\us33.a[0] ),
    .b(_06287_),
    .o1(_08919_));
 b15aoi022aq1n02x5 _34294_ (.a(_07014_),
    .b(_08917_),
    .c(_08918_),
    .d(_08919_),
    .o1(_08920_));
 b15oai022al1n06x5 _34295_ (.a(_06179_),
    .b(_06133_),
    .c(_06287_),
    .d(_06174_),
    .o1(_08921_));
 b15nandp2al1n03x5 _34296_ (.a(net559),
    .b(_07075_),
    .o1(_08922_));
 b15aoi222as1n08x5 _34297_ (.a(_06158_),
    .b(_08231_),
    .c(_07118_),
    .d(_08921_),
    .e(_08922_),
    .f(_06240_),
    .o1(_08923_));
 b15oai112as1n08x5 _34298_ (.a(_08916_),
    .b(_08920_),
    .c(net554),
    .d(_08923_),
    .o1(_08925_));
 b15aoai13an1n03x5 _34299_ (.a(net563),
    .b(_07867_),
    .c(_06140_),
    .d(net565),
    .o1(_08926_));
 b15oaoi13al1n08x5 _34300_ (.a(_08427_),
    .b(_08926_),
    .c(net565),
    .d(_07865_),
    .o1(_08927_));
 b15oai022ar1n02x5 _34301_ (.a(net555),
    .b(_07040_),
    .c(_07100_),
    .d(_06195_),
    .o1(_08928_));
 b15ao0012al1n06x5 _34302_ (.a(_08927_),
    .b(_08928_),
    .c(_07033_),
    .o(_08929_));
 b15oai112al1n02x5 _34303_ (.a(_06197_),
    .b(_06312_),
    .c(_06236_),
    .d(_06091_),
    .o1(_08930_));
 b15oai112ah1n04x5 _34304_ (.a(_06221_),
    .b(_08930_),
    .c(_06312_),
    .d(_08417_),
    .o1(_08931_));
 b15orn003ar1n02x5 _34305_ (.a(_07108_),
    .b(_06195_),
    .c(_07016_),
    .o(_08932_));
 b15oai022ar1n12x5 _34306_ (.a(_06201_),
    .b(_07784_),
    .c(_06127_),
    .d(net545),
    .o1(_08933_));
 b15aoi013aq1n02x5 _34307_ (.a(_08904_),
    .b(_08933_),
    .c(net543),
    .d(_06118_),
    .o1(_08934_));
 b15oai112aq1n08x5 _34308_ (.a(_08931_),
    .b(_08932_),
    .c(_08934_),
    .d(\us33.a[0] ),
    .o1(_08936_));
 b15nor004an1n12x5 _34309_ (.a(_08911_),
    .b(_08925_),
    .c(_08929_),
    .d(_08936_),
    .o1(_08937_));
 b15norp02ar1n02x5 _34310_ (.a(net556),
    .b(_07839_),
    .o1(_08938_));
 b15aoai13as1n02x5 _34311_ (.a(_06179_),
    .b(_08938_),
    .c(_06245_),
    .d(net556),
    .o1(_08939_));
 b15norp03aq1n02x5 _34312_ (.a(_06135_),
    .b(_06287_),
    .c(_07075_),
    .o1(_08940_));
 b15aoi012al1n04x5 _34313_ (.a(_08940_),
    .b(_07075_),
    .c(_06295_),
    .o1(_08941_));
 b15oai112ah1n06x5 _34314_ (.a(net559),
    .b(_08939_),
    .c(_08941_),
    .d(_06201_),
    .o1(_08942_));
 b15oaoi13al1n03x5 _34315_ (.a(net556),
    .b(_07838_),
    .c(_06327_),
    .d(_07032_),
    .o1(_08943_));
 b15aoi012an1n02x5 _34316_ (.a(_06201_),
    .b(_07817_),
    .c(_08396_),
    .o1(_08944_));
 b15oai013al1n06x5 _34317_ (.a(_08942_),
    .b(_08943_),
    .c(_08944_),
    .d(net559),
    .o1(_08945_));
 b15oaoi13ar1n02x5 _34318_ (.a(_06179_),
    .b(_06100_),
    .c(_06127_),
    .d(net566),
    .o1(_08947_));
 b15oab012an1n03x5 _34319_ (.a(_06298_),
    .b(_08947_),
    .c(_06220_),
    .out0(_08948_));
 b15oai022aq1n06x5 _34320_ (.a(_07839_),
    .b(_06100_),
    .c(_06230_),
    .d(net556),
    .o1(_08949_));
 b15aoi112al1n08x5 _34321_ (.a(_07816_),
    .b(_08948_),
    .c(_08949_),
    .d(_06207_),
    .o1(_08950_));
 b15aoi022aq1n02x5 _34322_ (.a(_06242_),
    .b(_06295_),
    .c(_07835_),
    .d(_08418_),
    .o1(_08951_));
 b15oai112aq1n08x5 _34323_ (.a(net561),
    .b(_06341_),
    .c(_07110_),
    .d(_06242_),
    .o1(_08952_));
 b15aoi012al1n06x5 _34324_ (.a(_06201_),
    .b(_08951_),
    .c(_08952_),
    .o1(_08953_));
 b15oab012ar1n02x5 _34325_ (.a(_07812_),
    .b(_07026_),
    .c(_06325_),
    .out0(_08954_));
 b15oai122al1n08x5 _34326_ (.a(net566),
    .b(_06127_),
    .c(_07817_),
    .d(_08954_),
    .e(_06201_),
    .o1(_08955_));
 b15aoai13an1n02x5 _34327_ (.a(_06294_),
    .b(_06240_),
    .c(net562),
    .d(_06243_),
    .o1(_08956_));
 b15aoai13an1n06x5 _34328_ (.a(_08956_),
    .b(_07016_),
    .c(_06230_),
    .d(_07839_),
    .o1(_08958_));
 b15oaoi13ar1n08x5 _34329_ (.a(_08953_),
    .b(_08955_),
    .c(_08958_),
    .d(net566),
    .o1(_08959_));
 b15andc04as1n16x5 _34330_ (.a(_08937_),
    .b(_08945_),
    .c(_08950_),
    .d(_08959_),
    .o(_08960_));
 b15xor002ah1n16x5 _34331_ (.a(_08625_),
    .b(_08960_),
    .out0(_08961_));
 b15xor002as1n04x5 _34332_ (.a(_08901_),
    .b(_08961_),
    .out0(_08962_));
 b15oaoi13al1n02x5 _34333_ (.a(_06574_),
    .b(_07198_),
    .c(_06554_),
    .d(net819),
    .o1(_08963_));
 b15oai012as1n03x5 _34334_ (.a(net817),
    .b(_06509_),
    .c(_08963_),
    .o1(_08964_));
 b15oai012ar1n02x5 _34335_ (.a(_06661_),
    .b(_06589_),
    .c(net819),
    .o1(_08965_));
 b15aoi022as1n02x5 _34336_ (.a(_06567_),
    .b(_07142_),
    .c(_08965_),
    .d(net813),
    .o1(_08966_));
 b15norp03ar1n02x5 _34337_ (.a(net797),
    .b(net799),
    .c(net811),
    .o1(_08967_));
 b15aoai13ar1n02x5 _34338_ (.a(net805),
    .b(_08967_),
    .c(_07202_),
    .d(net797),
    .o1(_08969_));
 b15oaoi13an1n03x5 _34339_ (.a(_07188_),
    .b(_08969_),
    .c(_06631_),
    .d(_06722_),
    .o1(_08970_));
 b15oai012as1n08x5 _34340_ (.a(net819),
    .b(_06509_),
    .c(_08970_),
    .o1(_08971_));
 b15aoi013as1n06x5 _34341_ (.a(net810),
    .b(_08964_),
    .c(_08966_),
    .d(_08971_),
    .o1(_08972_));
 b15nandp2an1n05x5 _34342_ (.a(net818),
    .b(net813),
    .o1(_08973_));
 b15oai012ar1n02x5 _34343_ (.a(\us11.a[3] ),
    .b(_08973_),
    .c(\us11.a[0] ),
    .o1(_08974_));
 b15oai012ar1n02x5 _34344_ (.a(_06580_),
    .b(_06567_),
    .c(_06476_),
    .o1(_08975_));
 b15oaoi13an1n02x5 _34345_ (.a(_08974_),
    .b(_08975_),
    .c(_06574_),
    .d(_06709_),
    .o1(_08976_));
 b15aoi112ar1n02x5 _34346_ (.a(_06593_),
    .b(_06616_),
    .c(_06628_),
    .d(\us11.a[0] ),
    .o1(_08977_));
 b15oai122as1n02x5 _34347_ (.a(_08973_),
    .b(_07754_),
    .c(_06567_),
    .d(_08977_),
    .e(_07725_),
    .o1(_08978_));
 b15oaoi13ar1n02x5 _34348_ (.a(_06536_),
    .b(_06600_),
    .c(_07258_),
    .d(_06514_),
    .o1(_08980_));
 b15aoai13al1n02x5 _34349_ (.a(_08980_),
    .b(net811),
    .c(_06527_),
    .d(_06606_),
    .o1(_08981_));
 b15nona23an1n05x5 _34350_ (.a(_07178_),
    .b(_08976_),
    .c(_08978_),
    .d(_08981_),
    .out0(_08982_));
 b15norp02ar1n02x5 _34351_ (.a(net805),
    .b(_07212_),
    .o1(_08983_));
 b15aoi012ar1n02x5 _34352_ (.a(_08983_),
    .b(_06714_),
    .c(net805),
    .o1(_08984_));
 b15nandp3ar1n02x5 _34353_ (.a(net810),
    .b(_07250_),
    .c(_07263_),
    .o1(_08985_));
 b15aoi022ar1n02x5 _34354_ (.a(net819),
    .b(_07240_),
    .c(_07137_),
    .d(net817),
    .o1(_08986_));
 b15oai022ar1n02x5 _34355_ (.a(_08984_),
    .b(_08985_),
    .c(_08986_),
    .d(_07161_),
    .o1(_08987_));
 b15norp02ar1n02x5 _34356_ (.a(net819),
    .b(_06659_),
    .o1(_08988_));
 b15aoai13ar1n02x5 _34357_ (.a(_08988_),
    .b(_06647_),
    .c(_07206_),
    .d(net816),
    .o1(_08989_));
 b15aoi022ar1n02x5 _34358_ (.a(net810),
    .b(_07191_),
    .c(_06642_),
    .d(_08035_),
    .o1(_08991_));
 b15oai012al1n02x5 _34359_ (.a(_08989_),
    .b(_08991_),
    .c(_07729_),
    .o1(_08992_));
 b15orn003an1n03x5 _34360_ (.a(_08982_),
    .b(_08987_),
    .c(_08992_),
    .o(_08993_));
 b15and003ar1n02x5 _34361_ (.a(net803),
    .b(_07132_),
    .c(_07218_),
    .o(_08994_));
 b15nor003as1n02x5 _34362_ (.a(net803),
    .b(_07148_),
    .c(_07161_),
    .o1(_08995_));
 b15oai012al1n06x5 _34363_ (.a(_06654_),
    .b(_08994_),
    .c(_08995_),
    .o1(_08996_));
 b15norp02as1n02x5 _34364_ (.a(_07229_),
    .b(_08294_),
    .o1(_08997_));
 b15oai112ah1n08x5 _34365_ (.a(_07680_),
    .b(_08996_),
    .c(_08997_),
    .d(_07130_),
    .o1(_08998_));
 b15nand03ar1n03x5 _34366_ (.a(_06476_),
    .b(_06574_),
    .c(_06700_),
    .o1(_08999_));
 b15oai012ah1n04x5 _34367_ (.a(_08999_),
    .b(_07130_),
    .c(_06589_),
    .o1(_09000_));
 b15aoai13as1n08x5 _34368_ (.a(_06632_),
    .b(_08998_),
    .c(_09000_),
    .d(net810),
    .o1(_09002_));
 b15oai012ar1n03x5 _34369_ (.a(_06499_),
    .b(_07223_),
    .c(_07240_),
    .o1(_09003_));
 b15aoi022ar1n06x5 _34370_ (.a(_07725_),
    .b(_06518_),
    .c(_06606_),
    .d(_06567_),
    .o1(_09004_));
 b15oaoi13aq1n04x5 _34371_ (.a(\us11.a[0] ),
    .b(_09003_),
    .c(_09004_),
    .d(\us11.a[3] ),
    .o1(_09005_));
 b15aoai13al1n08x5 _34372_ (.a(net816),
    .b(_07150_),
    .c(_06726_),
    .d(net811),
    .o1(_09006_));
 b15nand03an1n08x5 _34373_ (.a(_06574_),
    .b(_07240_),
    .c(_06609_),
    .o1(_09007_));
 b15aoai13ar1n08x5 _34374_ (.a(_08010_),
    .b(net809),
    .c(_09006_),
    .d(_09007_),
    .o1(_09008_));
 b15norp03ar1n03x5 _34375_ (.a(net814),
    .b(_06527_),
    .c(_06661_),
    .o1(_09009_));
 b15oai013aq1n02x5 _34376_ (.a(net809),
    .b(_06722_),
    .c(_06542_),
    .d(_07703_),
    .o1(_09010_));
 b15nandp3ar1n02x5 _34377_ (.a(_06574_),
    .b(_06539_),
    .c(_06638_),
    .o1(_09011_));
 b15nandp2aq1n02x5 _34378_ (.a(net821),
    .b(_06652_),
    .o1(_09013_));
 b15aob012al1n06x5 _34379_ (.a(net815),
    .b(_09011_),
    .c(_09013_),
    .out0(_09014_));
 b15oai112al1n08x5 _34380_ (.a(net814),
    .b(_06527_),
    .c(_06509_),
    .d(_06676_),
    .o1(_09015_));
 b15nona23an1n12x5 _34381_ (.a(_09009_),
    .b(_09010_),
    .c(_09014_),
    .d(_09015_),
    .out0(_09016_));
 b15oai013al1n02x5 _34382_ (.a(_06536_),
    .b(_07263_),
    .c(_06709_),
    .d(net813),
    .o1(_09017_));
 b15aoi012as1n02x5 _34383_ (.a(_09017_),
    .b(_07137_),
    .c(_06631_),
    .o1(_09018_));
 b15nor003ah1n02x5 _34384_ (.a(_06728_),
    .b(_06514_),
    .c(_06602_),
    .o1(_09019_));
 b15aoi022ar1n08x5 _34385_ (.a(_07206_),
    .b(_06616_),
    .c(_09019_),
    .d(net819),
    .o1(_09020_));
 b15norp02aq1n02x5 _34386_ (.a(net818),
    .b(_06593_),
    .o1(_09021_));
 b15aoai13an1n06x5 _34387_ (.a(net813),
    .b(_09021_),
    .c(_06624_),
    .d(_07206_),
    .o1(_09022_));
 b15aoai13an1n06x5 _34388_ (.a(_06476_),
    .b(_07137_),
    .c(_07240_),
    .d(net813),
    .o1(_09024_));
 b15nand04ah1n12x5 _34389_ (.a(_09018_),
    .b(_09020_),
    .c(_09022_),
    .d(_09024_),
    .o1(_09025_));
 b15aoi112as1n08x5 _34390_ (.a(_09005_),
    .b(_09008_),
    .c(_09016_),
    .d(_09025_),
    .o1(_09026_));
 b15nona23as1n32x5 _34391_ (.a(_08972_),
    .b(_08993_),
    .c(_09002_),
    .d(_09026_),
    .out0(_09027_));
 b15aoai13an1n03x5 _34392_ (.a(\us00.a[0] ),
    .b(_06076_),
    .c(_05997_),
    .d(net927),
    .o1(_09028_));
 b15oai013ah1n02x5 _34393_ (.a(_09028_),
    .b(_06046_),
    .c(_06024_),
    .d(net930),
    .o1(_09029_));
 b15nor002ar1n03x5 _34394_ (.a(_05899_),
    .b(_09029_),
    .o1(_09030_));
 b15aoi022ar1n02x5 _34395_ (.a(_06032_),
    .b(_06378_),
    .c(_06024_),
    .d(_09028_),
    .o1(_09031_));
 b15nor002aq1n02x5 _34396_ (.a(net927),
    .b(_09031_),
    .o1(_09032_));
 b15aoi012an1n02x5 _34397_ (.a(_06378_),
    .b(_06033_),
    .c(_09029_),
    .o1(_09033_));
 b15oai013ah1n06x5 _34398_ (.a(net924),
    .b(_09030_),
    .c(_09032_),
    .d(_09033_),
    .o1(_09035_));
 b15aoi012an1n02x5 _34399_ (.a(net934),
    .b(_06046_),
    .c(_06049_),
    .o1(_09036_));
 b15oai013ar1n02x5 _34400_ (.a(net928),
    .b(_05934_),
    .c(_05966_),
    .d(net931),
    .o1(_09037_));
 b15oai012aq1n04x5 _34401_ (.a(_09037_),
    .b(_07475_),
    .c(net928),
    .o1(_09038_));
 b15aoi013ar1n06x5 _34402_ (.a(_09036_),
    .b(_09038_),
    .c(net934),
    .d(_07427_),
    .o1(_09039_));
 b15aoi012al1n04x5 _34403_ (.a(_05984_),
    .b(_07594_),
    .c(_05841_),
    .o1(_09040_));
 b15aoai13ar1n03x5 _34404_ (.a(net928),
    .b(_08586_),
    .c(_05827_),
    .d(net934),
    .o1(_09041_));
 b15aoi022al1n06x5 _34405_ (.a(net925),
    .b(_07636_),
    .c(_06453_),
    .d(_06000_),
    .o1(_09042_));
 b15oai112aq1n08x5 _34406_ (.a(_09041_),
    .b(_09042_),
    .c(net925),
    .d(_06465_),
    .o1(_09043_));
 b15oaoi13as1n08x5 _34407_ (.a(_09039_),
    .b(_05821_),
    .c(_09040_),
    .d(_09043_),
    .o1(_09044_));
 b15oai012aq1n04x5 _34408_ (.a(\us00.a[2] ),
    .b(_05899_),
    .c(_07634_),
    .o1(_09046_));
 b15oai022an1n08x5 _34409_ (.a(_06364_),
    .b(_07646_),
    .c(_06078_),
    .d(net926),
    .o1(_09047_));
 b15oai112ah1n12x5 _34410_ (.a(\us00.a[0] ),
    .b(_09046_),
    .c(_09047_),
    .d(\us00.a[2] ),
    .o1(_09048_));
 b15oai112al1n06x5 _34411_ (.a(\us00.a[5] ),
    .b(net927),
    .c(_05969_),
    .d(\us00.a[6] ),
    .o1(_09049_));
 b15oaoi13ah1n08x5 _34412_ (.a(_07668_),
    .b(_09049_),
    .c(_06382_),
    .d(_08619_),
    .o1(_09050_));
 b15oai012ar1n12x5 _34413_ (.a(net930),
    .b(_06032_),
    .c(_09050_),
    .o1(_09051_));
 b15aoai13an1n06x5 _34414_ (.a(_05821_),
    .b(_07410_),
    .c(_06032_),
    .d(\us00.a[0] ),
    .o1(_09052_));
 b15aoai13as1n08x5 _34415_ (.a(_09048_),
    .b(net924),
    .c(_09051_),
    .d(_09052_),
    .o1(_09053_));
 b15aoi122ar1n08x5 _34416_ (.a(net930),
    .b(net924),
    .c(_06026_),
    .d(_05947_),
    .e(_07636_),
    .o1(_09054_));
 b15norp03al1n02x5 _34417_ (.a(_05918_),
    .b(net924),
    .c(_05972_),
    .o1(_09055_));
 b15aoai13as1n03x5 _34418_ (.a(net933),
    .b(_09055_),
    .c(_05932_),
    .d(net924),
    .o1(_09057_));
 b15norp03aq1n02x5 _34419_ (.a(_05928_),
    .b(_05854_),
    .c(_05846_),
    .o1(_09058_));
 b15aoi012ar1n04x5 _34420_ (.a(_09058_),
    .b(_05971_),
    .c(_06024_),
    .o1(_09059_));
 b15aoi013aq1n08x5 _34421_ (.a(_09054_),
    .b(_09057_),
    .c(_09059_),
    .d(net930),
    .o1(_09060_));
 b15nand02ar1n02x5 _34422_ (.a(_05827_),
    .b(_07656_),
    .o1(_09061_));
 b15nandp3ar1n02x5 _34423_ (.a(net931),
    .b(net928),
    .c(_07637_),
    .o1(_09062_));
 b15aoi012ar1n02x5 _34424_ (.a(_05911_),
    .b(_09061_),
    .c(_09062_),
    .o1(_09063_));
 b15aoai13ar1n02x5 _34425_ (.a(_05969_),
    .b(_05911_),
    .c(_05955_),
    .d(_05844_),
    .o1(_09064_));
 b15aoi122an1n02x5 _34426_ (.a(net928),
    .b(_05899_),
    .c(_07451_),
    .d(_09064_),
    .e(_05841_),
    .o1(_09065_));
 b15nona23al1n04x5 _34427_ (.a(_09063_),
    .b(_09065_),
    .c(_06016_),
    .d(_08102_),
    .out0(_09066_));
 b15nandp2ar1n02x5 _34428_ (.a(_05851_),
    .b(_05915_),
    .o1(_09068_));
 b15nandp2ar1n03x5 _34429_ (.a(net935),
    .b(_05947_),
    .o1(_09069_));
 b15oaoi13aq1n04x5 _34430_ (.a(net932),
    .b(_09068_),
    .c(_07448_),
    .d(_09069_),
    .o1(_09070_));
 b15oai112as1n02x5 _34431_ (.a(\us00.a[3] ),
    .b(_07463_),
    .c(_05917_),
    .d(_06432_),
    .o1(_09071_));
 b15oai013aq1n06x5 _34432_ (.a(_09071_),
    .b(_05851_),
    .c(_05882_),
    .d(_06405_),
    .o1(_09072_));
 b15aoi012al1n02x5 _34433_ (.a(_06003_),
    .b(_05844_),
    .c(_05969_),
    .o1(_09073_));
 b15oai013aq1n06x5 _34434_ (.a(_07458_),
    .b(_09073_),
    .c(_05883_),
    .d(_05835_),
    .o1(_09074_));
 b15oai112an1n12x5 _34435_ (.a(net929),
    .b(_06368_),
    .c(_08342_),
    .d(_08343_),
    .o1(_09075_));
 b15nandp2ar1n02x5 _34436_ (.a(_05898_),
    .b(_05975_),
    .o1(_09076_));
 b15oai013ah1n04x5 _34437_ (.a(_09075_),
    .b(_08141_),
    .c(_09076_),
    .d(net935),
    .o1(_09077_));
 b15nor004aq1n12x5 _34438_ (.a(_09070_),
    .b(_09072_),
    .c(_09074_),
    .d(_09077_),
    .o1(_09079_));
 b15nandp2al1n02x5 _34439_ (.a(_06056_),
    .b(_05915_),
    .o1(_09080_));
 b15oaoi13al1n04x5 _34440_ (.a(_05851_),
    .b(_09080_),
    .c(_05821_),
    .d(_07646_),
    .o1(_09081_));
 b15nandp2ar1n02x5 _34441_ (.a(_07637_),
    .b(_07451_),
    .o1(_09082_));
 b15oaoi13an1n04x5 _34442_ (.a(net932),
    .b(_09082_),
    .c(_06465_),
    .d(_05851_),
    .o1(_09083_));
 b15aoi012ar1n02x5 _34443_ (.a(net935),
    .b(_05835_),
    .c(_05846_),
    .o1(_09084_));
 b15oab012ar1n04x5 _34444_ (.a(_06405_),
    .b(_07666_),
    .c(_09084_),
    .out0(_09085_));
 b15norp03al1n12x5 _34445_ (.a(_09081_),
    .b(_09083_),
    .c(_09085_),
    .o1(_09086_));
 b15nona23ah1n16x5 _34446_ (.a(_09060_),
    .b(_09066_),
    .c(_09079_),
    .d(_09086_),
    .out0(_09087_));
 b15nano23as1n24x5 _34447_ (.a(_09035_),
    .b(_09044_),
    .c(_09053_),
    .d(_09087_),
    .out0(_09088_));
 b15xor002ah1n16x5 _34448_ (.a(_09027_),
    .b(_09088_),
    .out0(_09090_));
 b15xor002as1n08x5 _34449_ (.a(_08962_),
    .b(_09090_),
    .out0(_09091_));
 b15oai012ar1n02x5 _34450_ (.a(_08834_),
    .b(_09091_),
    .c(net538),
    .o1(_09092_));
 b15xor002ar1n02x5 _34451_ (.a(\u0.w[0][6] ),
    .b(_09092_),
    .out0(_00103_));
 b15inv040as1n06x5 _34452_ (.a(\text_in_r[103] ),
    .o1(_09093_));
 b15aoi012as1n06x5 _34453_ (.a(net809),
    .b(_09007_),
    .c(_09006_),
    .o1(_09094_));
 b15nand02as1n03x5 _34454_ (.a(_07173_),
    .b(_06700_),
    .o1(_09095_));
 b15oaoi13aq1n03x5 _34455_ (.a(net821),
    .b(_09095_),
    .c(_06542_),
    .d(_06661_),
    .o1(_09096_));
 b15nor002ar1n02x5 _34456_ (.a(net804),
    .b(net815),
    .o1(_09097_));
 b15oai112as1n06x5 _34457_ (.a(_07249_),
    .b(_07747_),
    .c(_09097_),
    .d(net814),
    .o1(_09098_));
 b15aoi122al1n06x5 _34458_ (.a(_09098_),
    .b(_06706_),
    .c(_06589_),
    .d(_06577_),
    .e(_06728_),
    .o1(_09100_));
 b15nor003ar1n02x5 _34459_ (.a(net803),
    .b(net800),
    .c(net817),
    .o1(_09101_));
 b15aoi013ah1n03x5 _34460_ (.a(_09101_),
    .b(_06705_),
    .c(net800),
    .d(net803),
    .o1(_09102_));
 b15nor003an1n12x5 _34461_ (.a(_07161_),
    .b(_07737_),
    .c(_09102_),
    .o1(_09103_));
 b15aoi112aq1n02x5 _34462_ (.a(_06577_),
    .b(_08008_),
    .c(_07764_),
    .d(_06587_),
    .o1(_09104_));
 b15nor004ah1n04x5 _34463_ (.a(_09096_),
    .b(_09100_),
    .c(_09103_),
    .d(_09104_),
    .o1(_09105_));
 b15aoi022ar1n16x5 _34464_ (.a(_06691_),
    .b(_07230_),
    .c(_07218_),
    .d(_07209_),
    .o1(_09106_));
 b15nor004al1n06x5 _34465_ (.a(net802),
    .b(net814),
    .c(_06642_),
    .d(_09106_),
    .o1(_09107_));
 b15oai013aq1n03x5 _34466_ (.a(_09013_),
    .b(_06624_),
    .c(_06686_),
    .d(net814),
    .o1(_09108_));
 b15aoi122an1n04x5 _34467_ (.a(_09107_),
    .b(_08023_),
    .c(_06606_),
    .d(_06536_),
    .e(_09108_),
    .o1(_09109_));
 b15aoi112aq1n02x5 _34468_ (.a(_06587_),
    .b(_06659_),
    .c(_07157_),
    .d(net815),
    .o1(_09111_));
 b15nor002an1n02x5 _34469_ (.a(net804),
    .b(_06705_),
    .o1(_09112_));
 b15nand03ar1n06x5 _34470_ (.a(net799),
    .b(_06530_),
    .c(_07251_),
    .o1(_09113_));
 b15aoi112aq1n06x5 _34471_ (.a(_09112_),
    .b(_09113_),
    .c(net804),
    .d(net815),
    .o1(_09114_));
 b15oai012ah1n02x5 _34472_ (.a(_08047_),
    .b(_06704_),
    .c(_06628_),
    .o1(_09115_));
 b15nor003al1n06x5 _34473_ (.a(_09111_),
    .b(_09114_),
    .c(_09115_),
    .o1(_09116_));
 b15aoi012al1n02x5 _34474_ (.a(_06632_),
    .b(_07156_),
    .c(_06628_),
    .o1(_09117_));
 b15nand04aq1n02x5 _34475_ (.a(net809),
    .b(_06538_),
    .c(_06539_),
    .d(_06642_),
    .o1(_09118_));
 b15oaoi13an1n04x5 _34476_ (.a(_09117_),
    .b(_09118_),
    .c(_06558_),
    .d(net809),
    .o1(_09119_));
 b15nand03ar1n03x5 _34477_ (.a(_06536_),
    .b(_06698_),
    .c(_07721_),
    .o1(_09120_));
 b15aoi012ar1n02x5 _34478_ (.a(_06602_),
    .b(_06565_),
    .c(_06638_),
    .o1(_09122_));
 b15oai013as1n03x5 _34479_ (.a(_09120_),
    .b(_09122_),
    .c(_08049_),
    .d(_06488_),
    .o1(_09123_));
 b15oai012ar1n02x5 _34480_ (.a(_06606_),
    .b(_06616_),
    .c(net809),
    .o1(_09124_));
 b15aoi012ar1n02x5 _34481_ (.a(_06499_),
    .b(_06530_),
    .c(net820),
    .o1(_09125_));
 b15oaoi13as1n03x5 _34482_ (.a(net815),
    .b(_09124_),
    .c(_09125_),
    .d(_06610_),
    .o1(_09126_));
 b15nand03aq1n03x5 _34483_ (.a(net804),
    .b(net799),
    .c(_06698_),
    .o1(_09127_));
 b15aoai13ah1n02x5 _34484_ (.a(net802),
    .b(_08027_),
    .c(_07147_),
    .d(net797),
    .o1(_09128_));
 b15nand03aq1n03x5 _34485_ (.a(net815),
    .b(net808),
    .c(_07747_),
    .o1(_09129_));
 b15aoi012aq1n06x5 _34486_ (.a(_09127_),
    .b(_09128_),
    .c(_09129_),
    .o1(_09130_));
 b15nor004an1n06x5 _34487_ (.a(_09119_),
    .b(_09123_),
    .c(_09126_),
    .d(_09130_),
    .o1(_09131_));
 b15nand04ah1n12x5 _34488_ (.a(_09105_),
    .b(_09109_),
    .c(_09116_),
    .d(_09131_),
    .o1(_09133_));
 b15nor003al1n02x5 _34489_ (.a(net821),
    .b(_06499_),
    .c(_06530_),
    .o1(_09134_));
 b15aoi012ar1n02x5 _34490_ (.a(net815),
    .b(_07161_),
    .c(net821),
    .o1(_09135_));
 b15aoi012al1n02x5 _34491_ (.a(_06703_),
    .b(_08008_),
    .c(_06659_),
    .o1(_09136_));
 b15nor004ar1n04x5 _34492_ (.a(_06600_),
    .b(_09134_),
    .c(_09135_),
    .d(_09136_),
    .o1(_09137_));
 b15nand04ar1n02x5 _34493_ (.a(_06574_),
    .b(net809),
    .c(_06577_),
    .d(_07721_),
    .o1(_09138_));
 b15aoi022ar1n02x5 _34494_ (.a(_06580_),
    .b(_06673_),
    .c(_08023_),
    .d(_06509_),
    .o1(_09139_));
 b15oai012al1n02x5 _34495_ (.a(_09138_),
    .b(_09139_),
    .c(_06574_),
    .o1(_09140_));
 b15aob012ar1n02x5 _34496_ (.a(net809),
    .b(_06554_),
    .c(_06704_),
    .out0(_09141_));
 b15oaoi13as1n02x5 _34497_ (.a(_07130_),
    .b(_09141_),
    .c(net809),
    .d(_06728_),
    .o1(_09142_));
 b15orn003ah1n04x5 _34498_ (.a(_09137_),
    .b(_09140_),
    .c(_09142_),
    .o(_09144_));
 b15oai013ar1n02x5 _34499_ (.a(_06542_),
    .b(_06628_),
    .c(_06632_),
    .d(_07191_),
    .o1(_09145_));
 b15nandp3ar1n02x5 _34500_ (.a(_06536_),
    .b(_07191_),
    .c(_07156_),
    .o1(_09146_));
 b15oai112ar1n04x5 _34501_ (.a(_06545_),
    .b(_06638_),
    .c(_07156_),
    .d(_06548_),
    .o1(_09147_));
 b15aoi022ar1n02x5 _34502_ (.a(net821),
    .b(_09145_),
    .c(_09146_),
    .d(_09147_),
    .o1(_09148_));
 b15aoi013ar1n02x5 _34503_ (.a(_06476_),
    .b(net818),
    .c(_06509_),
    .d(_06530_),
    .o1(_09149_));
 b15oai012ar1n02x5 _34504_ (.a(_09149_),
    .b(_07177_),
    .c(_06593_),
    .o1(_09150_));
 b15aoi012ar1n02x5 _34505_ (.a(net818),
    .b(_06580_),
    .c(_07173_),
    .o1(_09151_));
 b15nandp3al1n02x5 _34506_ (.a(_06536_),
    .b(_06538_),
    .c(_06545_),
    .o1(_09152_));
 b15aoi013ar1n03x5 _34507_ (.a(_09151_),
    .b(_07989_),
    .c(_09152_),
    .d(net818),
    .o1(_09153_));
 b15oai012ar1n03x5 _34508_ (.a(_06476_),
    .b(_07161_),
    .c(_07198_),
    .o1(_09155_));
 b15oaoi13an1n03x5 _34509_ (.a(_09148_),
    .b(_09150_),
    .c(_09153_),
    .d(_09155_),
    .o1(_09156_));
 b15nor003ah1n02x5 _34510_ (.a(net813),
    .b(_06615_),
    .c(_06637_),
    .o1(_09157_));
 b15norp03as1n02x5 _34511_ (.a(_06574_),
    .b(\us11.a[3] ),
    .c(_06709_),
    .o1(_09158_));
 b15oai012ar1n08x5 _34512_ (.a(net818),
    .b(_09157_),
    .c(_09158_),
    .o1(_09159_));
 b15nandp3ar1n02x5 _34513_ (.a(net814),
    .b(net809),
    .c(_06509_),
    .o1(_09160_));
 b15aob012ar1n02x5 _34514_ (.a(_06632_),
    .b(_09095_),
    .c(_09160_),
    .out0(_09161_));
 b15nor003ar1n02x5 _34515_ (.a(\us11.a[7] ),
    .b(net811),
    .c(_06675_),
    .o1(_09162_));
 b15norp03al1n02x5 _34516_ (.a(_06552_),
    .b(_06645_),
    .c(_08973_),
    .o1(_09163_));
 b15oai112ah1n04x5 _34517_ (.a(_07749_),
    .b(net820),
    .c(_09162_),
    .d(_09163_),
    .o1(_09164_));
 b15aoi012ar1n02x5 _34518_ (.a(_07135_),
    .b(_07721_),
    .c(_06706_),
    .o1(_09166_));
 b15aob012ah1n02x5 _34519_ (.a(net809),
    .b(_09164_),
    .c(_09166_),
    .out0(_09167_));
 b15nand04as1n06x5 _34520_ (.a(_09156_),
    .b(_09159_),
    .c(_09161_),
    .d(_09167_),
    .o1(_09168_));
 b15nor004as1n12x5 _34521_ (.a(_09094_),
    .b(_09133_),
    .c(_09144_),
    .d(_09168_),
    .o1(_09169_));
 b15xor002as1n16x5 _34522_ (.a(_06088_),
    .b(_09169_),
    .out0(_09170_));
 b15nand04al1n08x5 _34523_ (.a(net678),
    .b(_06800_),
    .c(_06863_),
    .d(_06844_),
    .o1(_09171_));
 b15nor004al1n03x5 _34524_ (.a(\us22.a[4] ),
    .b(_06999_),
    .c(_07906_),
    .d(_07361_),
    .o1(_09172_));
 b15norp03ar1n02x5 _34525_ (.a(_07948_),
    .b(\us22.a[6] ),
    .c(_06990_),
    .o1(_09173_));
 b15oai112ar1n04x5 _34526_ (.a(net680),
    .b(_08495_),
    .c(_09172_),
    .d(_09173_),
    .o1(_09174_));
 b15aoi013ar1n02x5 _34527_ (.a(_06959_),
    .b(_06777_),
    .c(\us22.a[3] ),
    .d(net669),
    .o1(_09175_));
 b15nand02ar1n02x5 _34528_ (.a(\us22.a[6] ),
    .b(_07546_),
    .o1(_09177_));
 b15oai112an1n02x5 _34529_ (.a(_09171_),
    .b(_09174_),
    .c(_09175_),
    .d(_09177_),
    .o1(_09178_));
 b15and002ah1n03x5 _34530_ (.a(net690),
    .b(_09178_),
    .o(_09179_));
 b15norp03ar1n02x5 _34531_ (.a(_06792_),
    .b(net680),
    .c(_06981_),
    .o1(_09180_));
 b15aoai13al1n02x5 _34532_ (.a(_06826_),
    .b(_09180_),
    .c(_08508_),
    .d(_06792_),
    .o1(_09181_));
 b15norp02ah1n04x5 _34533_ (.a(net690),
    .b(_09181_),
    .o1(_09182_));
 b15nanb02as1n02x5 _34534_ (.a(net683),
    .b(\us22.a[4] ),
    .out0(_09183_));
 b15orn003ar1n02x5 _34535_ (.a(_06826_),
    .b(_06922_),
    .c(_08503_),
    .o(_09184_));
 b15nand03ar1n06x5 _34536_ (.a(net687),
    .b(_06927_),
    .c(_07309_),
    .o1(_09185_));
 b15oaoi13aq1n02x5 _34537_ (.a(_09183_),
    .b(_09184_),
    .c(_09185_),
    .d(_06786_),
    .o1(_09186_));
 b15oai013ah1n02x5 _34538_ (.a(_09185_),
    .b(_08503_),
    .c(_06922_),
    .d(net678),
    .o1(_09188_));
 b15aoi013al1n04x5 _34539_ (.a(_09186_),
    .b(_09188_),
    .c(_07948_),
    .d(net683),
    .o1(_09189_));
 b15aoi012ar1n02x5 _34540_ (.a(_06786_),
    .b(_06790_),
    .c(_07354_),
    .o1(_09190_));
 b15oai012ar1n03x5 _34541_ (.a(_07364_),
    .b(_07937_),
    .c(_09190_),
    .o1(_09191_));
 b15nand04aq1n02x5 _34542_ (.a(\us22.a[0] ),
    .b(_06792_),
    .c(_06822_),
    .d(_06839_),
    .o1(_09192_));
 b15nand04an1n06x5 _34543_ (.a(_06882_),
    .b(_06823_),
    .c(_06922_),
    .d(_06954_),
    .o1(_09193_));
 b15oaoi13ar1n04x5 _34544_ (.a(_06869_),
    .b(_09192_),
    .c(_09193_),
    .d(\us22.a[0] ),
    .o1(_09194_));
 b15nano23an1n03x5 _34545_ (.a(_09191_),
    .b(_07359_),
    .c(_08867_),
    .d(_09194_),
    .out0(_09195_));
 b15nandp2ah1n03x5 _34546_ (.a(_06844_),
    .b(_07504_),
    .o1(_09196_));
 b15nandp2ar1n03x5 _34547_ (.a(_09196_),
    .b(_07553_),
    .o1(_09197_));
 b15oai022ar1n02x5 _34548_ (.a(net678),
    .b(_06936_),
    .c(_06837_),
    .d(_06781_),
    .o1(_09199_));
 b15aoai13an1n03x5 _34549_ (.a(_06775_),
    .b(_09197_),
    .c(_09199_),
    .d(_06777_),
    .o1(_09200_));
 b15nand02ar1n02x5 _34550_ (.a(\us22.a[5] ),
    .b(net688),
    .o1(_09201_));
 b15nand04as1n04x5 _34551_ (.a(_07523_),
    .b(_06927_),
    .c(_07521_),
    .d(_09201_),
    .o1(_09202_));
 b15oai112as1n02x5 _34552_ (.a(net683),
    .b(_09202_),
    .c(_06824_),
    .d(_06990_),
    .o1(_09203_));
 b15nand04ar1n02x5 _34553_ (.a(_06882_),
    .b(_07942_),
    .c(_06768_),
    .d(_06748_),
    .o1(_09204_));
 b15oai013aq1n02x5 _34554_ (.a(_09204_),
    .b(_06748_),
    .c(_06934_),
    .d(_06921_),
    .o1(_09205_));
 b15nandp2ar1n02x5 _34555_ (.a(_07319_),
    .b(_06882_),
    .o1(_09206_));
 b15oai013ah1n04x5 _34556_ (.a(_09196_),
    .b(_07970_),
    .c(_09206_),
    .d(_07338_),
    .o1(_09207_));
 b15oai013as1n03x5 _34557_ (.a(_09203_),
    .b(_09205_),
    .c(_09207_),
    .d(net680),
    .o1(_09208_));
 b15nand04ah1n08x5 _34558_ (.a(_09189_),
    .b(_09195_),
    .c(_09200_),
    .d(_09208_),
    .o1(_09210_));
 b15aoi012al1n02x5 _34559_ (.a(net678),
    .b(_07372_),
    .c(_07535_),
    .o1(_09211_));
 b15oai012ar1n08x5 _34560_ (.a(_09211_),
    .b(_06748_),
    .c(_06975_),
    .o1(_09212_));
 b15nand04as1n08x5 _34561_ (.a(net689),
    .b(net681),
    .c(_06767_),
    .d(_06823_),
    .o1(_09213_));
 b15aoi022ar1n24x5 _34562_ (.a(_07910_),
    .b(_07273_),
    .c(_09213_),
    .d(net684),
    .o1(_09214_));
 b15nano22ar1n02x5 _34563_ (.a(net675),
    .b(\us22.a[6] ),
    .c(net683),
    .out0(_09215_));
 b15aoi013ar1n03x5 _34564_ (.a(_09215_),
    .b(_06966_),
    .c(_06999_),
    .d(_07948_),
    .o1(_09216_));
 b15nandp2ah1n02x5 _34565_ (.a(_06792_),
    .b(_07310_),
    .o1(_09217_));
 b15oai122an1n08x5 _34566_ (.a(net678),
    .b(_06748_),
    .c(_08889_),
    .d(_09216_),
    .e(_09217_),
    .o1(_09218_));
 b15nor004al1n02x5 _34567_ (.a(net675),
    .b(net669),
    .c(\us22.a[6] ),
    .d(net687),
    .o1(_09219_));
 b15aoai13ah1n02x5 _34568_ (.a(_08545_),
    .b(_09219_),
    .c(_07306_),
    .d(_06836_),
    .o1(_09221_));
 b15nand03aq1n06x5 _34569_ (.a(_06999_),
    .b(_07546_),
    .c(_07309_),
    .o1(_09222_));
 b15nand04an1n06x5 _34570_ (.a(net673),
    .b(_06882_),
    .c(\us22.a[6] ),
    .d(_07291_),
    .o1(_09223_));
 b15aoai13ah1n06x5 _34571_ (.a(_09221_),
    .b(net675),
    .c(_09222_),
    .d(_09223_),
    .o1(_09224_));
 b15oai013al1n08x5 _34572_ (.a(_09212_),
    .b(_09214_),
    .c(_09218_),
    .d(_09224_),
    .o1(_09225_));
 b15oai012ar1n04x5 _34573_ (.a(_07512_),
    .b(_08484_),
    .c(_06786_),
    .o1(_09226_));
 b15norp03ar1n03x5 _34574_ (.a(_07319_),
    .b(_06800_),
    .c(_07287_),
    .o1(_09227_));
 b15obai22an1n02x5 _34575_ (.a(_07943_),
    .b(_07287_),
    .c(net673),
    .d(_06781_),
    .out0(_09228_));
 b15aoi012ar1n02x5 _34576_ (.a(_09183_),
    .b(_06915_),
    .c(_06826_),
    .o1(_09229_));
 b15aoi022ar1n02x5 _34577_ (.a(_09226_),
    .b(_09227_),
    .c(_09228_),
    .d(_09229_),
    .o1(_09230_));
 b15nor004aq1n03x5 _34578_ (.a(_06933_),
    .b(_07302_),
    .c(_06966_),
    .d(_07338_),
    .o1(_09232_));
 b15oai022aq1n02x5 _34579_ (.a(_06980_),
    .b(_08503_),
    .c(_07904_),
    .d(_06984_),
    .o1(_09233_));
 b15aoi013ar1n02x5 _34580_ (.a(_09232_),
    .b(_09233_),
    .c(\us22.a[6] ),
    .d(_07901_),
    .o1(_09234_));
 b15oai112ah1n02x5 _34581_ (.a(_06758_),
    .b(_06807_),
    .c(_06911_),
    .d(_06826_),
    .o1(_09235_));
 b15aoi022an1n04x5 _34582_ (.a(_06927_),
    .b(_07288_),
    .c(_07339_),
    .d(_06767_),
    .o1(_09236_));
 b15oai013aq1n08x5 _34583_ (.a(_09235_),
    .b(_09236_),
    .c(_06790_),
    .d(net674),
    .o1(_09237_));
 b15nandp3ah1n03x5 _34584_ (.a(_06866_),
    .b(_06889_),
    .c(_07378_),
    .o1(_09238_));
 b15aoi022ar1n02x5 _34585_ (.a(_06775_),
    .b(_06823_),
    .c(_06768_),
    .d(net686),
    .o1(_09239_));
 b15oai013ar1n03x5 _34586_ (.a(_09238_),
    .b(_09239_),
    .c(_06837_),
    .d(_07302_),
    .o1(_09240_));
 b15nano23ah1n03x5 _34587_ (.a(_09230_),
    .b(_09234_),
    .c(_09237_),
    .d(_09240_),
    .out0(_09241_));
 b15nano23aq1n05x5 _34588_ (.a(_06823_),
    .b(_06926_),
    .c(_06748_),
    .d(net671),
    .out0(_09243_));
 b15orn003al1n03x5 _34589_ (.a(_06790_),
    .b(_06995_),
    .c(_08494_),
    .o(_09244_));
 b15oai012as1n03x5 _34590_ (.a(_09244_),
    .b(_06981_),
    .c(_06859_),
    .o1(_09245_));
 b15oai013ah1n08x5 _34591_ (.a(_06826_),
    .b(_08511_),
    .c(_09243_),
    .d(_09245_),
    .o1(_09246_));
 b15aoi022ar1n04x5 _34592_ (.a(_07309_),
    .b(_07367_),
    .c(_07931_),
    .d(_06912_),
    .o1(_09247_));
 b15nor003as1n04x5 _34593_ (.a(net675),
    .b(_06761_),
    .c(_09247_),
    .o1(_09248_));
 b15oai022aq1n06x5 _34594_ (.a(_07384_),
    .b(_06790_),
    .c(_06980_),
    .d(_06778_),
    .o1(_09249_));
 b15aoi112ar1n06x5 _34595_ (.a(_06918_),
    .b(_09248_),
    .c(_09249_),
    .d(_06826_),
    .o1(_09250_));
 b15nand04ah1n12x5 _34596_ (.a(_09225_),
    .b(_09241_),
    .c(_09246_),
    .d(_09250_),
    .o1(_09251_));
 b15nor004as1n12x5 _34597_ (.a(_09179_),
    .b(_09182_),
    .c(_09210_),
    .d(_09251_),
    .o1(_09252_));
 b15norp02as1n02x5 _34598_ (.a(_06207_),
    .b(_07058_),
    .o1(_09254_));
 b15oai012ah1n02x5 _34599_ (.a(_06133_),
    .b(_06197_),
    .c(net554),
    .o1(_09255_));
 b15aboi22ah1n06x5 _34600_ (.a(_07092_),
    .b(_09254_),
    .c(_09255_),
    .d(_08418_),
    .out0(_09256_));
 b15norp03ah1n08x5 _34601_ (.a(net556),
    .b(_06345_),
    .c(_07079_),
    .o1(_09257_));
 b15oaoi13ar1n03x5 _34602_ (.a(_09257_),
    .b(_06295_),
    .c(_06163_),
    .d(_06294_),
    .o1(_09258_));
 b15aoi022ar1n02x5 _34603_ (.a(_06220_),
    .b(_07812_),
    .c(_06221_),
    .d(_06313_),
    .o1(_09259_));
 b15oai022an1n02x5 _34604_ (.a(\us33.a[0] ),
    .b(_09258_),
    .c(_09259_),
    .d(_07030_),
    .o1(_09260_));
 b15nand03ar1n03x5 _34605_ (.a(net559),
    .b(net552),
    .c(net543),
    .o1(_09261_));
 b15nona22ar1n02x5 _34606_ (.a(net548),
    .b(net546),
    .c(net554),
    .out0(_09262_));
 b15oaoi13ah1n03x5 _34607_ (.a(_09261_),
    .b(_09262_),
    .c(_07052_),
    .d(net562),
    .o1(_09263_));
 b15oai013as1n02x5 _34608_ (.a(net567),
    .b(net546),
    .c(_06244_),
    .d(_06127_),
    .o1(_09265_));
 b15oai013as1n02x5 _34609_ (.a(_06197_),
    .b(_06306_),
    .c(_07011_),
    .d(net562),
    .o1(_09266_));
 b15aoi112aq1n06x5 _34610_ (.a(_09263_),
    .b(_09265_),
    .c(_09266_),
    .d(\us33.a[2] ),
    .o1(_09267_));
 b15oai022ar1n04x5 _34611_ (.a(_06272_),
    .b(_06199_),
    .c(_07838_),
    .d(_06155_),
    .o1(_09268_));
 b15oab012al1n02x5 _34612_ (.a(_09267_),
    .b(_09268_),
    .c(\us33.a[0] ),
    .out0(_09269_));
 b15nonb03aq1n06x5 _34613_ (.a(_09256_),
    .b(_09260_),
    .c(_09269_),
    .out0(_09270_));
 b15nor003an1n02x5 _34614_ (.a(net559),
    .b(_06091_),
    .c(_06096_),
    .o1(_09271_));
 b15oai012aq1n06x5 _34615_ (.a(_06111_),
    .b(_07834_),
    .c(_09271_),
    .o1(_09272_));
 b15aoi012ar1n02x5 _34616_ (.a(_06201_),
    .b(_08417_),
    .c(_06207_),
    .o1(_09273_));
 b15aoi012al1n02x5 _34617_ (.a(_08638_),
    .b(_08417_),
    .c(net562),
    .o1(_09274_));
 b15oai112al1n06x5 _34618_ (.a(_09272_),
    .b(_09273_),
    .c(_06111_),
    .d(_09274_),
    .o1(_09276_));
 b15oai022aq1n04x5 _34619_ (.a(net562),
    .b(_06230_),
    .c(_07026_),
    .d(_06133_),
    .o1(_09277_));
 b15aoi012an1n02x5 _34620_ (.a(_06111_),
    .b(_06243_),
    .c(net562),
    .o1(_09278_));
 b15aoi112ah1n04x5 _34621_ (.a(net559),
    .b(_09278_),
    .c(_06195_),
    .d(_07839_),
    .o1(_09279_));
 b15oai013ah1n06x5 _34622_ (.a(_09276_),
    .b(_09277_),
    .c(_09279_),
    .d(net556),
    .o1(_09280_));
 b15aoi012ar1n02x5 _34623_ (.a(net556),
    .b(_08417_),
    .c(_06327_),
    .o1(_09281_));
 b15aoai13ar1n02x5 _34624_ (.a(net562),
    .b(_06313_),
    .c(_07033_),
    .d(_08417_),
    .o1(_09282_));
 b15oai112an1n04x5 _34625_ (.a(_09281_),
    .b(_09282_),
    .c(_07032_),
    .d(_07012_),
    .o1(_09283_));
 b15nandp2ar1n05x5 _34626_ (.a(_08239_),
    .b(_09283_),
    .o1(_09284_));
 b15oai022ah1n06x5 _34627_ (.a(_06135_),
    .b(_06294_),
    .c(_08631_),
    .d(_06174_),
    .o1(_09285_));
 b15nand03ar1n08x5 _34628_ (.a(net562),
    .b(_06217_),
    .c(_09285_),
    .o1(_09287_));
 b15oai022ah1n06x5 _34629_ (.a(_06100_),
    .b(_07074_),
    .c(_07817_),
    .d(_06223_),
    .o1(_09288_));
 b15aob012ah1n02x5 _34630_ (.a(_06272_),
    .b(_07835_),
    .c(_06264_),
    .out0(_09289_));
 b15aoi012as1n06x5 _34631_ (.a(_09288_),
    .b(_09289_),
    .c(_07804_),
    .o1(_09290_));
 b15oai112as1n16x5 _34632_ (.a(_09284_),
    .b(_09287_),
    .c(_09290_),
    .d(net562),
    .o1(_09291_));
 b15aoi013an1n03x5 _34633_ (.a(net555),
    .b(_06266_),
    .c(_06265_),
    .d(_07075_),
    .o1(_09292_));
 b15aoi022as1n06x5 _34634_ (.a(_06158_),
    .b(_06143_),
    .c(_06217_),
    .d(_07791_),
    .o1(_09293_));
 b15oai012ar1n08x5 _34635_ (.a(_09292_),
    .b(_09293_),
    .c(_06242_),
    .o1(_09294_));
 b15aoi012ar1n02x5 _34636_ (.a(_07012_),
    .b(_07010_),
    .c(_06179_),
    .o1(_09295_));
 b15oai012an1n02x5 _34637_ (.a(net556),
    .b(_06325_),
    .c(_09295_),
    .o1(_09296_));
 b15aoi022ar1n02x5 _34638_ (.a(net559),
    .b(_08417_),
    .c(_07036_),
    .d(net566),
    .o1(_09298_));
 b15oaoi13an1n02x5 _34639_ (.a(_06179_),
    .b(_09298_),
    .c(_06195_),
    .d(net566),
    .o1(_09299_));
 b15aoi112ar1n02x5 _34640_ (.a(net559),
    .b(_07025_),
    .c(_06158_),
    .d(_06111_),
    .o1(_09300_));
 b15aoi112an1n02x5 _34641_ (.a(net561),
    .b(_09300_),
    .c(_07839_),
    .d(net559),
    .o1(_09301_));
 b15oai013aq1n04x5 _34642_ (.a(_09294_),
    .b(_09296_),
    .c(_09299_),
    .d(_09301_),
    .o1(_09302_));
 b15norp02aq1n02x5 _34643_ (.a(_06325_),
    .b(_06199_),
    .o1(_09303_));
 b15oai022as1n02x5 _34644_ (.a(_06325_),
    .b(_06127_),
    .c(_07838_),
    .d(_06105_),
    .o1(_09304_));
 b15aoai13an1n06x5 _34645_ (.a(net566),
    .b(_09303_),
    .c(_09304_),
    .d(_06179_),
    .o1(_09305_));
 b15norp02ar1n03x5 _34646_ (.a(_07040_),
    .b(_07093_),
    .o1(_09306_));
 b15oaoi13as1n02x5 _34647_ (.a(_06179_),
    .b(_08396_),
    .c(_07040_),
    .d(net566),
    .o1(_09307_));
 b15oai012al1n08x5 _34648_ (.a(_06163_),
    .b(_09306_),
    .c(_09307_),
    .o1(_09309_));
 b15aoi122ar1n06x5 _34649_ (.a(net557),
    .b(_06312_),
    .c(_08189_),
    .d(_06245_),
    .e(net555),
    .o1(_09310_));
 b15aoi022ar1n02x5 _34650_ (.a(net556),
    .b(_07025_),
    .c(_07103_),
    .d(_06245_),
    .o1(_09311_));
 b15ao0012an1n03x5 _34651_ (.a(_09310_),
    .b(_09311_),
    .c(net559),
    .o(_09312_));
 b15nand04an1n16x5 _34652_ (.a(_09302_),
    .b(_09305_),
    .c(_09309_),
    .d(_09312_),
    .o1(_09313_));
 b15nano23as1n24x5 _34653_ (.a(_09270_),
    .b(_09280_),
    .c(_09291_),
    .d(_09313_),
    .out0(_09314_));
 b15xnr002aq1n02x5 _34654_ (.a(_09088_),
    .b(_09314_),
    .out0(_09315_));
 b15xor002ar1n03x5 _34655_ (.a(_09252_),
    .b(_09315_),
    .out0(_09316_));
 b15xor002aq1n03x5 _34656_ (.a(_09170_),
    .b(_09316_),
    .out0(_09317_));
 b15mdn022ar1n08x5 _34657_ (.a(_09093_),
    .b(_09317_),
    .o1(_09318_),
    .sa(net535));
 b15xor002ar1n02x5 _34658_ (.a(\u0.w[0][7] ),
    .b(_09318_),
    .out0(_00104_));
 b15inv000an1n05x5 _34659_ (.a(\text_in_r[104] ),
    .o1(_09320_));
 b15xnr002as1n16x5 _34660_ (.a(_06353_),
    .b(_09252_),
    .out0(_09321_));
 b15xor002ar1n12x5 _34661_ (.a(_06741_),
    .b(_07126_),
    .out0(_09322_));
 b15xor002aq1n06x5 _34662_ (.a(_09321_),
    .b(_09322_),
    .out0(_09323_));
 b15mdn022al1n12x5 _34663_ (.a(_09320_),
    .b(_09323_),
    .o1(_09324_),
    .sa(net535));
 b15xor002an1n16x5 _34664_ (.a(\u0.w[0][8] ),
    .b(_09324_),
    .out0(_00065_));
 b15xor002ar1n03x5 _34665_ (.a(_07267_),
    .b(_07125_),
    .out0(_09325_));
 b15xor003aq1n06x5 _34666_ (.a(_07004_),
    .b(_07887_),
    .c(_09325_),
    .out0(_09326_));
 b15xor002ar1n02x5 _34667_ (.a(_09321_),
    .b(_09326_),
    .out0(_09327_));
 b15cmbn22as1n03x5 _34668_ (.clk1(\text_in_r[105] ),
    .clk2(_09327_),
    .clkout(_09329_),
    .s(net535));
 b15xor002an1n06x5 _34669_ (.a(\u0.w[0][9] ),
    .b(_09329_),
    .out0(_00066_));
 b15inv040an1n05x5 _34670_ (.a(\text_in_r[106] ),
    .o1(_09330_));
 b15xor002ah1n04x5 _34671_ (.a(_07886_),
    .b(_08244_),
    .out0(_09331_));
 b15xor002as1n08x5 _34672_ (.a(_07392_),
    .b(_09331_),
    .out0(_09332_));
 b15xor002ah1n12x5 _34673_ (.a(_07776_),
    .b(_09332_),
    .out0(_09333_));
 b15mdn022ar1n03x5 _34674_ (.a(_09330_),
    .b(_09333_),
    .o1(_09334_),
    .sa(net538));
 b15xor002al1n02x5 _34675_ (.a(\u0.w[0][10] ),
    .b(_09334_),
    .out0(_00067_));
 b15xor002ah1n16x5 _34676_ (.a(_07586_),
    .b(_08244_),
    .out0(_09335_));
 b15xor003aq1n16x5 _34677_ (.a(_08077_),
    .b(_08467_),
    .c(_09335_),
    .out0(_09336_));
 b15xor002ah1n16x5 _34678_ (.a(_09321_),
    .b(_09336_),
    .out0(_09338_));
 b15cmbn22ar1n02x5 _34679_ (.clk1(\text_in_r[107] ),
    .clk2(_09338_),
    .clkout(_09339_),
    .s(net538));
 b15xor002ar1n02x5 _34680_ (.a(\u0.w[0][11] ),
    .b(_09339_),
    .out0(_00068_));
 b15xor003an1n08x5 _34681_ (.a(_07988_),
    .b(_08466_),
    .c(_08701_),
    .out0(_09340_));
 b15xor002as1n06x5 _34682_ (.a(_08384_),
    .b(_09340_),
    .out0(_09341_));
 b15xor002an1n16x5 _34683_ (.a(_09321_),
    .b(_09341_),
    .out0(_09342_));
 b15cmbn22ar1n02x5 _34684_ (.clk1(\text_in_r[108] ),
    .clk2(_09342_),
    .clkout(_09343_),
    .s(net538));
 b15xor002ar1n02x5 _34685_ (.a(\u0.w[0][12] ),
    .b(_09343_),
    .out0(_00069_));
 b15inv040ah1n02x5 _34686_ (.a(\text_in_r[109] ),
    .o1(_09344_));
 b15xor002as1n12x5 _34687_ (.a(_08554_),
    .b(_08701_),
    .out0(_09345_));
 b15xor002as1n06x5 _34688_ (.a(_08830_),
    .b(_09345_),
    .out0(_09347_));
 b15xor002as1n08x5 _34689_ (.a(_08961_),
    .b(_09347_),
    .out0(_09348_));
 b15mdn022an1n03x5 _34690_ (.a(_09344_),
    .b(_09348_),
    .o1(_09349_),
    .sa(net538));
 b15xor002ar1n02x5 _34691_ (.a(\u0.w[0][13] ),
    .b(_09349_),
    .out0(_00070_));
 b15inv040ah1n02x5 _34692_ (.a(\text_in_r[110] ),
    .o1(_09350_));
 b15xor002ar1n02x5 _34693_ (.a(_08960_),
    .b(_09314_),
    .out0(_09351_));
 b15xor002al1n02x5 _34694_ (.a(_08772_),
    .b(_09351_),
    .out0(_09352_));
 b15xor002as1n02x5 _34695_ (.a(_09090_),
    .b(_09352_),
    .out0(_09353_));
 b15mdn022ar1n03x5 _34696_ (.a(_09350_),
    .b(_09353_),
    .o1(_09354_),
    .sa(net538));
 b15xor002aq1n02x5 _34697_ (.a(\u0.w[0][14] ),
    .b(_09354_),
    .out0(_00071_));
 b15inv020as1n05x5 _34698_ (.a(\text_in_r[111] ),
    .o1(_09356_));
 b15xnr002ah1n12x5 _34699_ (.a(_08901_),
    .b(_09314_),
    .out0(_09357_));
 b15xor003an1n16x5 _34700_ (.a(_06353_),
    .b(_09170_),
    .c(_09357_),
    .out0(_09358_));
 b15mdn022al1n03x5 _34701_ (.a(_09356_),
    .b(_09358_),
    .o1(_09359_),
    .sa(net538));
 b15xor002ar1n02x5 _34702_ (.a(\u0.w[0][15] ),
    .b(_09359_),
    .out0(_00072_));
 b15xnr002as1n12x5 _34703_ (.a(_09169_),
    .b(_09252_),
    .out0(_09360_));
 b15xor003as1n06x5 _34704_ (.a(_07004_),
    .b(_07126_),
    .c(_09360_),
    .out0(_09361_));
 b15norp02ar1n02x5 _34705_ (.a(net536),
    .b(_09361_),
    .o1(_09362_));
 b15inv040as1n02x5 _34706_ (.a(\text_in_r[112] ),
    .o1(_09363_));
 b15aoi012ar1n02x5 _34707_ (.a(_09362_),
    .b(_09363_),
    .c(net536),
    .o1(_09364_));
 b15xor002ar1n02x5 _34708_ (.a(\u0.w[0][16] ),
    .b(_09364_),
    .out0(_00033_));
 b15inv040ah1n02x5 _34709_ (.a(\text_in_r[113] ),
    .o1(_09366_));
 b15qgbxo2an1n05x5 _34710_ (.a(_07887_),
    .b(_09360_),
    .out0(_09367_));
 b15xor002ah1n03x5 _34711_ (.a(_07005_),
    .b(_07392_),
    .out0(_09368_));
 b15xor002aq1n08x5 _34712_ (.a(_09367_),
    .b(_09368_),
    .out0(_09369_));
 b15mdn022aq1n02x5 _34713_ (.a(_09366_),
    .b(_09369_),
    .o1(_09370_),
    .sa(net536));
 b15xor002al1n02x5 _34714_ (.a(\u0.w[0][17] ),
    .b(_09370_),
    .out0(_00034_));
 b15xor002ar1n08x5 _34715_ (.a(_07679_),
    .b(_09335_),
    .out0(_09371_));
 b15xor002as1n03x5 _34716_ (.a(_07393_),
    .b(_09371_),
    .out0(_09372_));
 b15cmbn22al1n08x5 _34717_ (.clk1(\text_in_r[114] ),
    .clk2(_09372_),
    .clkout(_09373_),
    .s(net536));
 b15xor002ah1n08x5 _34718_ (.a(\u0.w[0][18] ),
    .b(_09373_),
    .out0(_00035_));
 b15xor002an1n02x5 _34719_ (.a(_08467_),
    .b(_09360_),
    .out0(_09375_));
 b15xnr002al1n03x5 _34720_ (.a(_07586_),
    .b(_07988_),
    .out0(_09376_));
 b15xor002al1n03x5 _34721_ (.a(_07775_),
    .b(_09376_),
    .out0(_09377_));
 b15xor002an1n04x5 _34722_ (.a(_09375_),
    .b(_09377_),
    .out0(_09378_));
 b15cmbn22ah1n04x5 _34723_ (.clk1(\text_in_r[115] ),
    .clk2(_09378_),
    .clkout(_09379_),
    .s(net536));
 b15xor002an1n06x5 _34724_ (.a(\u0.w[0][19] ),
    .b(_09379_),
    .out0(_00036_));
 b15inv040ah1n02x5 _34725_ (.a(\text_in_r[116] ),
    .o1(_09380_));
 b15qgbxo2an1n10x5 _34726_ (.a(_08078_),
    .b(_09345_),
    .out0(_09381_));
 b15xor002ah1n04x5 _34727_ (.a(_08383_),
    .b(_09360_),
    .out0(_09382_));
 b15xor002as1n08x5 _34728_ (.a(_09381_),
    .b(_09382_),
    .out0(_09384_));
 b15mdn022aq1n06x5 _34729_ (.a(_09380_),
    .b(_09384_),
    .o1(_09385_),
    .sa(net536));
 b15xor002al1n04x5 _34730_ (.a(\u0.w[0][20] ),
    .b(_09385_),
    .out0(_00037_));
 b15xor003al1n12x5 _34731_ (.a(net394),
    .b(_08554_),
    .c(_08772_),
    .out0(_09386_));
 b15xor002an1n12x5 _34732_ (.a(_08961_),
    .b(_09386_),
    .out0(_09387_));
 b15nor002an1n04x5 _34733_ (.a(net536),
    .b(_09387_),
    .o1(_09388_));
 b15inv000ah1n04x5 _34734_ (.a(\text_in_r[117] ),
    .o1(_09389_));
 b15aoi012ah1n12x5 _34735_ (.a(_09388_),
    .b(_09389_),
    .c(net536),
    .o1(_09390_));
 b15xor002as1n16x5 _34736_ (.a(\u0.w[0][21] ),
    .b(_09390_),
    .out0(_00038_));
 b15inv020as1n10x5 _34737_ (.a(\text_in_r[118] ),
    .o1(_09391_));
 b15xor003aq1n12x5 _34738_ (.a(_08831_),
    .b(_09088_),
    .c(_09357_),
    .out0(_09393_));
 b15mdn022as1n12x5 _34739_ (.a(_09391_),
    .b(_09393_),
    .o1(_09394_),
    .sa(net537));
 b15xor002as1n16x5 _34740_ (.a(\u0.w[0][22] ),
    .b(_09394_),
    .out0(_00039_));
 b15xor003aq1n08x5 _34741_ (.a(_06088_),
    .b(_08901_),
    .c(_09027_),
    .out0(_09395_));
 b15xor002as1n08x5 _34742_ (.a(_09321_),
    .b(_09395_),
    .out0(_09396_));
 b15cmbn22al1n04x5 _34743_ (.clk1(\text_in_r[119] ),
    .clk2(_09396_),
    .clkout(_09397_),
    .s(net536));
 b15xor002as1n03x5 _34744_ (.a(\u0.w[0][23] ),
    .b(_09397_),
    .out0(_00040_));
 b15inv000ah1n05x5 _34745_ (.a(\text_in_r[120] ),
    .o1(_09398_));
 b15xor003ah1n04x5 _34746_ (.a(_07005_),
    .b(_07125_),
    .c(_09170_),
    .out0(_09399_));
 b15mdn022ar1n02x5 _34747_ (.a(_09398_),
    .b(_09399_),
    .o1(_09400_),
    .sa(net535));
 b15xor002ar1n02x5 _34748_ (.a(\u0.w[0][24] ),
    .b(_09400_),
    .out0(_00001_));
 b15xor002ar1n03x5 _34749_ (.a(_06741_),
    .b(_07886_),
    .out0(_09402_));
 b15xor002aq1n03x5 _34750_ (.a(_06474_),
    .b(_09402_),
    .out0(_09403_));
 b15xor003aq1n06x5 _34751_ (.a(_07393_),
    .b(_09170_),
    .c(_09403_),
    .out0(_09404_));
 b15cmbn22ar1n02x5 _34752_ (.clk1(\text_in_r[121] ),
    .clk2(_09404_),
    .clkout(_09405_),
    .s(net535));
 b15xor002ar1n02x5 _34753_ (.a(\u0.w[0][25] ),
    .b(_09405_),
    .out0(_00002_));
 b15xor003aq1n06x5 _34754_ (.a(_07267_),
    .b(_07492_),
    .c(_07775_),
    .out0(_09406_));
 b15xor002ar1n08x5 _34755_ (.a(_09335_),
    .b(_09406_),
    .out0(_09407_));
 b15nor002aq1n04x5 _34756_ (.a(net535),
    .b(_09407_),
    .o1(_09408_));
 b15inv040ah1n02x5 _34757_ (.a(\text_in_r[122] ),
    .o1(_09409_));
 b15aoi012ar1n02x5 _34758_ (.a(_09408_),
    .b(_09409_),
    .c(net535),
    .o1(_09411_));
 b15xor002ar1n02x5 _34759_ (.a(\u0.w[0][26] ),
    .b(_09411_),
    .out0(_00003_));
 b15inv000an1n06x5 _34760_ (.a(\text_in_r[123] ),
    .o1(_09412_));
 b15xor002al1n04x5 _34761_ (.a(_07776_),
    .b(_08078_),
    .out0(_09413_));
 b15xor003al1n06x5 _34762_ (.a(_08466_),
    .b(_09170_),
    .c(_09413_),
    .out0(_09414_));
 b15mdn022ar1n03x5 _34763_ (.a(_09412_),
    .b(_09414_),
    .o1(_09415_),
    .sa(net535));
 b15xor002ar1n02x5 _34764_ (.a(\u0.w[0][27] ),
    .b(_09415_),
    .out0(_00004_));
 b15xnr002aq1n04x5 _34765_ (.a(_08077_),
    .b(_08166_),
    .out0(_09416_));
 b15xor002al1n03x5 _34766_ (.a(net394),
    .b(_09416_),
    .out0(_09417_));
 b15xor003ah1n03x5 _34767_ (.a(_09170_),
    .b(_09345_),
    .c(_09417_),
    .out0(_09418_));
 b15cmbn22ar1n02x5 _34768_ (.clk1(\text_in_r[124] ),
    .clk2(_09418_),
    .clkout(_09420_),
    .s(net535));
 b15xor002ar1n02x5 _34769_ (.a(\u0.w[0][28] ),
    .b(_09420_),
    .out0(_00005_));
 b15xor002ar1n02x5 _34770_ (.a(_08831_),
    .b(_08960_),
    .out0(_09421_));
 b15xor002ar1n02x5 _34771_ (.a(_08384_),
    .b(_09421_),
    .out0(_09422_));
 b15cmbn22ar1n02x5 _34772_ (.clk1(\text_in_r[125] ),
    .clk2(_09422_),
    .clkout(_09423_),
    .s(net535));
 b15xor002ar1n02x5 _34773_ (.a(\u0.w[0][29] ),
    .b(_09423_),
    .out0(_00006_));
 b15inv000ah1n10x5 _34774_ (.a(\text_in_r[126] ),
    .o1(_09424_));
 b15xor002as1n02x5 _34775_ (.a(_08830_),
    .b(_09027_),
    .out0(_09425_));
 b15xor002an1n02x5 _34776_ (.a(_08625_),
    .b(_09425_),
    .out0(_09426_));
 b15xnr002ar1n03x5 _34777_ (.a(_09357_),
    .b(_09426_),
    .out0(_09427_));
 b15mdn022ar1n03x5 _34778_ (.a(_09424_),
    .b(_09427_),
    .o1(_09429_),
    .sa(net535));
 b15xor002al1n02x5 _34779_ (.a(\u0.w[0][30] ),
    .b(_09429_),
    .out0(_00007_));
 b15inv040ah1n02x5 _34780_ (.a(\text_in_r[127] ),
    .o1(_09430_));
 b15xor002al1n02x5 _34781_ (.a(_09090_),
    .b(_09169_),
    .out0(_09431_));
 b15xor002ar1n02x5 _34782_ (.a(_09321_),
    .b(_09431_),
    .out0(_09432_));
 b15mdn022ar1n02x5 _34783_ (.a(_09430_),
    .b(_09432_),
    .o1(_09433_),
    .sa(net535));
 b15xor002al1n02x5 _34784_ (.a(\u0.w[0][31] ),
    .b(_09433_),
    .out0(_00008_));
 b15xnr002al1n12x5 _34785_ (.a(\u0.w[0][24] ),
    .b(_06474_),
    .out0(_00153_));
 b15xnr002ah1n03x5 _34786_ (.a(\u0.w[0][25] ),
    .b(_07492_),
    .out0(_00154_));
 b15xnr002as1n02x5 _34787_ (.a(\u0.w[0][26] ),
    .b(_07679_),
    .out0(_00155_));
 b15xor002aq1n08x5 _34788_ (.a(\u0.w[0][27] ),
    .b(_08166_),
    .out0(_00156_));
 b15xnr002al1n12x5 _34789_ (.a(\u0.w[0][28] ),
    .b(_08383_),
    .out0(_00157_));
 b15xor002ah1n16x5 _34790_ (.a(\u0.w[0][29] ),
    .b(_08625_),
    .out0(_00158_));
 b15xnr002ah1n12x5 _34791_ (.a(\u0.w[0][30] ),
    .b(_09088_),
    .out0(_00159_));
 b15xor002aq1n02x5 _34792_ (.a(\u0.w[0][31] ),
    .b(_06088_),
    .out0(_00160_));
 b15xor002ar1n02x5 _34793_ (.a(\u0.w[1][24] ),
    .b(_02771_),
    .out0(_00249_));
 b15xor002as1n02x5 _34794_ (.a(\u0.w[1][25] ),
    .b(_03633_),
    .out0(_00250_));
 b15xnr002ar1n08x5 _34795_ (.a(\u0.w[1][26] ),
    .b(_04217_),
    .out0(_00251_));
 b15xor002as1n12x5 _34796_ (.a(\u0.w[1][27] ),
    .b(_04478_),
    .out0(_00252_));
 b15xor002an1n04x5 _34797_ (.a(\u0.w[1][28] ),
    .b(_04955_),
    .out0(_00253_));
 b15xor002ar1n02x5 _34798_ (.a(\u0.w[1][29] ),
    .b(_05229_),
    .out0(_00254_));
 b15xnr002al1n04x5 _34799_ (.a(\u0.w[1][30] ),
    .b(_05361_),
    .out0(_00255_));
 b15xnr002an1n12x5 _34800_ (.a(\u0.w[1][31] ),
    .b(_03413_),
    .out0(_00256_));
 b15xnr002ah1n12x5 _34801_ (.a(net523),
    .b(_16424_),
    .out0(_00209_));
 b15xnr002an1n08x5 _34802_ (.a(net522),
    .b(_17281_),
    .out0(_00210_));
 b15xor002as1n06x5 _34803_ (.a(net521),
    .b(_00706_),
    .out0(_00211_));
 b15xnr002an1n16x5 _34804_ (.a(\u0.w[2][27] ),
    .b(_00973_),
    .out0(_00212_));
 b15xnr002ar1n08x5 _34805_ (.a(\u0.w[2][28] ),
    .b(_01209_),
    .out0(_00213_));
 b15xnr002ah1n03x5 _34806_ (.a(\u0.w[2][29] ),
    .b(_01689_),
    .out0(_00214_));
 b15xor002al1n02x5 _34807_ (.a(\u0.w[2][30] ),
    .b(_01871_),
    .out0(_00215_));
 b15xor002ar1n02x5 _34808_ (.a(\u0.w[2][31] ),
    .b(_17068_),
    .out0(_00216_));
 b15xor002al1n02x5 _34809_ (.a(net432),
    .b(_12776_),
    .out0(_00177_));
 b15xor002ar1n02x5 _34810_ (.a(net425),
    .b(_13768_),
    .out0(_00178_));
 b15xor002ar1n02x5 _34811_ (.a(_04168_),
    .b(_14493_),
    .out0(_00179_));
 b15xor002ar1n02x5 _34812_ (.a(net417),
    .b(_14826_),
    .out0(_00180_));
 b15xor002ar1n02x5 _34813_ (.a(\u0.tmp_w[28] ),
    .b(_15034_),
    .out0(_00181_));
 b15xor002ar1n02x5 _34814_ (.a(net411),
    .b(_15231_),
    .out0(_00182_));
 b15xor002ar1n02x5 _34815_ (.a(net408),
    .b(_15491_),
    .out0(_00183_));
 b15xnr002ar1n02x5 _34816_ (.a(net406),
    .b(_13663_),
    .out0(_00184_));
 b15xnr002al1n02x5 _34817_ (.a(\u0.w[0][16] ),
    .b(_06741_),
    .out0(_00145_));
 b15xor002ar1n03x5 _34818_ (.a(\u0.w[0][17] ),
    .b(_07267_),
    .out0(_00146_));
 b15xnr002al1n02x5 _34819_ (.a(\u0.w[0][18] ),
    .b(_07775_),
    .out0(_00147_));
 b15xor002ar1n02x5 _34820_ (.a(\u0.w[0][19] ),
    .b(_08077_),
    .out0(_00148_));
 b15xnr002al1n16x5 _34821_ (.a(\u0.w[0][20] ),
    .b(net394),
    .out0(_00149_));
 b15xnr002ah1n08x5 _34822_ (.a(\u0.w[0][21] ),
    .b(_08830_),
    .out0(_00150_));
 b15xor002al1n08x5 _34823_ (.a(\u0.w[0][22] ),
    .b(_09027_),
    .out0(_00151_));
 b15xnr002aq1n08x5 _34824_ (.a(\u0.w[0][23] ),
    .b(_09169_),
    .out0(_00152_));
 b15xnr002ar1n03x5 _34825_ (.a(\u0.w[1][16] ),
    .b(net401),
    .out0(_00241_));
 b15xor002ar1n02x5 _34826_ (.a(\u0.w[1][17] ),
    .b(_03769_),
    .out0(_00242_));
 b15xnr002ar1n08x5 _34827_ (.a(\u0.w[1][18] ),
    .b(net399),
    .out0(_00243_));
 b15xor002ar1n02x5 _34828_ (.a(\u0.w[1][19] ),
    .b(net398),
    .out0(_00244_));
 b15xnr002aq1n08x5 _34829_ (.a(\u0.w[1][20] ),
    .b(_04721_),
    .out0(_00245_));
 b15xnr002ar1n02x5 _34830_ (.a(\u0.w[1][21] ),
    .b(_05102_),
    .out0(_00246_));
 b15xor002al1n03x5 _34831_ (.a(\u0.w[1][22] ),
    .b(_05418_),
    .out0(_00247_));
 b15xor002ah1n12x5 _34832_ (.a(\u0.w[1][23] ),
    .b(net396),
    .out0(_00248_));
 b15xnr002ah1n12x5 _34833_ (.a(net527),
    .b(_16689_),
    .out0(_00201_));
 b15xnr002an1n16x5 _34834_ (.a(net526),
    .b(_17196_),
    .out0(_00202_));
 b15xor002al1n16x5 _34835_ (.a(net525),
    .b(_17615_),
    .out0(_00203_));
 b15xnr002al1n16x5 _34836_ (.a(net524),
    .b(_00905_),
    .out0(_00204_));
 b15xnr002an1n12x5 _34837_ (.a(\u0.w[2][20] ),
    .b(_01285_),
    .out0(_00205_));
 b15xnr002ar1n08x5 _34838_ (.a(\u0.w[2][21] ),
    .b(_01620_),
    .out0(_00206_));
 b15qgbxo2an1n05x5 _34839_ (.a(\u0.w[2][22] ),
    .b(_01940_),
    .out0(_00207_));
 b15xnr002as1n06x5 _34840_ (.a(\u0.w[2][23] ),
    .b(_02121_),
    .out0(_00208_));
 b15xor002al1n03x5 _34841_ (.a(_11579_),
    .b(_13019_),
    .out0(_00169_));
 b15xor002as1n02x5 _34842_ (.a(_11696_),
    .b(_13891_),
    .out0(_00170_));
 b15xor002al1n04x5 _34843_ (.a(_11603_),
    .b(_14247_),
    .out0(_00171_));
 b15xor002al1n02x5 _34844_ (.a(_11666_),
    .b(_14673_),
    .out0(_00172_));
 b15xor002ar1n02x5 _34845_ (.a(net447),
    .b(_14973_),
    .out0(_00173_));
 b15xor002as1n16x5 _34846_ (.a(_11689_),
    .b(_15173_),
    .out0(_00174_));
 b15xor002as1n16x5 _34847_ (.a(_11939_),
    .b(_15428_),
    .out0(_00175_));
 b15xor002ar1n02x5 _34848_ (.a(net433),
    .b(_15797_),
    .out0(_00176_));
 b15xor002ar1n08x5 _34849_ (.a(\u0.w[0][8] ),
    .b(_07004_),
    .out0(_00137_));
 b15xnr002ah1n02x5 _34850_ (.a(\u0.w[0][9] ),
    .b(_07392_),
    .out0(_00138_));
 b15xnr002as1n04x5 _34851_ (.a(\u0.w[0][10] ),
    .b(_07586_),
    .out0(_00139_));
 b15xnr002as1n12x5 _34852_ (.a(\u0.w[0][11] ),
    .b(_07988_),
    .out0(_00140_));
 b15xor002as1n08x5 _34853_ (.a(\u0.w[0][12] ),
    .b(_08554_),
    .out0(_00141_));
 b15xor002as1n12x5 _34854_ (.a(\u0.w[0][13] ),
    .b(_08772_),
    .out0(_00142_));
 b15xnr002an1n16x5 _34855_ (.a(\u0.w[0][14] ),
    .b(_08901_),
    .out0(_00143_));
 b15xnr002as1n12x5 _34856_ (.a(\u0.w[0][15] ),
    .b(_09252_),
    .out0(_00144_));
 b15xnr002ar1n02x5 _34857_ (.a(\u0.w[1][8] ),
    .b(net400),
    .out0(_00225_));
 b15xnr002an1n06x5 _34858_ (.a(\u0.w[1][9] ),
    .b(net393),
    .out0(_00226_));
 b15xor002an1n12x5 _34859_ (.a(\u0.w[1][10] ),
    .b(net392),
    .out0(_00227_));
 b15xnr002ah1n12x5 _34860_ (.a(\u0.w[1][11] ),
    .b(net397),
    .out0(_00228_));
 b15xnr002al1n08x5 _34861_ (.a(\u0.w[1][12] ),
    .b(_04800_),
    .out0(_00229_));
 b15xnr002ar1n04x5 _34862_ (.a(\u0.w[1][13] ),
    .b(_05030_),
    .out0(_00230_));
 b15xor002as1n12x5 _34863_ (.a(\u0.w[1][14] ),
    .b(_05300_),
    .out0(_00231_));
 b15xnr002ar1n02x5 _34864_ (.a(\u0.w[1][15] ),
    .b(net395),
    .out0(_00232_));
 b15xor002al1n02x5 _34865_ (.a(net529),
    .b(_16168_),
    .out0(_00193_));
 b15xnr002al1n02x5 _34866_ (.a(net528),
    .b(_17526_),
    .out0(_00194_));
 b15xor002ar1n02x5 _34867_ (.a(\u0.w[2][10] ),
    .b(_00618_),
    .out0(_00195_));
 b15xnr002aq1n02x5 _34868_ (.a(\u0.w[2][11] ),
    .b(_01049_),
    .out0(_00196_));
 b15xnr002al1n03x5 _34869_ (.a(\u0.w[2][12] ),
    .b(_01426_),
    .out0(_00197_));
 b15xor002ar1n02x5 _34870_ (.a(\u0.w[2][13] ),
    .b(_01500_),
    .out0(_00198_));
 b15xor002al1n02x5 _34871_ (.a(\u0.w[2][14] ),
    .b(_01813_),
    .out0(_00199_));
 b15qgbxo2an1n10x5 _34872_ (.a(\u0.w[2][15] ),
    .b(_02002_),
    .out0(_00200_));
 b15xor002al1n03x5 _34873_ (.a(_10732_),
    .b(_13297_),
    .out0(_00161_));
 b15xor002ar1n02x5 _34874_ (.a(_10893_),
    .b(_14136_),
    .out0(_00162_));
 b15xor002ar1n02x5 _34875_ (.a(_10728_),
    .b(_14337_),
    .out0(_00163_));
 b15xor002al1n03x5 _34876_ (.a(_10939_),
    .b(_14763_),
    .out0(_00164_));
 b15xor002ar1n02x5 _34877_ (.a(_11205_),
    .b(_14898_),
    .out0(_00165_));
 b15xor002aq1n16x5 _34878_ (.a(\u0.tmp_w[13] ),
    .b(_15288_),
    .out0(_00166_));
 b15xor002ar1n02x5 _34879_ (.a(_10758_),
    .b(_15614_),
    .out0(_00167_));
 b15xnr002al1n03x5 _34880_ (.a(\u0.tmp_w[15] ),
    .b(_15670_),
    .out0(_00168_));
 b15xnr002ar1n04x5 _34881_ (.a(\u0.w[0][0] ),
    .b(_07125_),
    .out0(_00129_));
 b15xor002ar1n02x5 _34882_ (.a(net532),
    .b(_07886_),
    .out0(_00130_));
 b15xnr002al1n06x5 _34883_ (.a(\u0.w[0][2] ),
    .b(_08244_),
    .out0(_00131_));
 b15xnr002ar1n08x5 _34884_ (.a(\u0.w[0][3] ),
    .b(_08466_),
    .out0(_00132_));
 b15xnr002ah1n08x5 _34885_ (.a(\u0.w[0][4] ),
    .b(_08701_),
    .out0(_00133_));
 b15xnr002aq1n16x5 _34886_ (.a(\u0.w[0][5] ),
    .b(_08960_),
    .out0(_00134_));
 b15xnr002ah1n12x5 _34887_ (.a(\u0.w[0][6] ),
    .b(_09314_),
    .out0(_00135_));
 b15xnr002ah1n06x5 _34888_ (.a(\u0.w[0][7] ),
    .b(_06353_),
    .out0(_00136_));
 b15xor002ah1n08x5 _34889_ (.a(\u0.w[1][0] ),
    .b(_03544_),
    .out0(_00217_));
 b15xor002an1n02x5 _34890_ (.a(\u0.w[1][1] ),
    .b(_04319_),
    .out0(_00218_));
 b15xnr002ah1n12x5 _34891_ (.a(\u0.w[1][2] ),
    .b(_04554_),
    .out0(_00219_));
 b15xnr002ar1n02x5 _34892_ (.a(\u0.w[1][3] ),
    .b(_04878_),
    .out0(_00220_));
 b15xnr002ah1n16x5 _34893_ (.a(\u0.w[1][4] ),
    .b(_05164_),
    .out0(_00221_));
 b15xnr002an1n16x5 _34894_ (.a(\u0.w[1][5] ),
    .b(_05485_),
    .out0(_00222_));
 b15xnr002aq1n16x5 _34895_ (.a(\u0.w[1][6] ),
    .b(_05544_),
    .out0(_00223_));
 b15xnr002ah1n16x5 _34896_ (.a(\u0.w[1][7] ),
    .b(_03034_),
    .out0(_00224_));
 b15xnr002as1n12x5 _34897_ (.a(\u0.w[2][0] ),
    .b(_17396_),
    .out0(_00185_));
 b15xnr002as1n12x5 _34898_ (.a(net531),
    .b(_00818_),
    .out0(_00186_));
 b15xnr002an1n16x5 _34899_ (.a(\u0.w[2][2] ),
    .b(_01138_),
    .out0(_00187_));
 b15xnr002as1n12x5 _34900_ (.a(net530),
    .b(_01364_),
    .out0(_00188_));
 b15xnr002an1n16x5 _34901_ (.a(\u0.w[2][4] ),
    .b(_01557_),
    .out0(_00189_));
 b15xnr002al1n03x5 _34902_ (.a(\u0.w[2][5] ),
    .b(_01754_),
    .out0(_00190_));
 b15xnr002as1n04x5 _34903_ (.a(\u0.w[2][6] ),
    .b(_02061_),
    .out0(_00191_));
 b15xnr002al1n08x5 _34904_ (.a(\u0.w[2][7] ),
    .b(_16926_),
    .out0(_00192_));
 b15xor002ar1n02x5 _34905_ (.a(_09888_),
    .b(net402),
    .out0(_00233_));
 b15xor002ar1n02x5 _34906_ (.a(_09932_),
    .b(_14424_),
    .out0(_00234_));
 b15xor002an1n03x5 _34907_ (.a(\u0.tmp_w[2] ),
    .b(_14585_),
    .out0(_00235_));
 b15xor002ar1n02x5 _34908_ (.a(_10038_),
    .b(_15106_),
    .out0(_00236_));
 b15xor002ar1n02x5 _34909_ (.a(\u0.tmp_w[4] ),
    .b(_15351_),
    .out0(_00237_));
 b15xor002ar1n02x5 _34910_ (.a(net499),
    .b(_15552_),
    .out0(_00238_));
 b15xnr002ar1n02x5 _34911_ (.a(net495),
    .b(_15727_),
    .out0(_00239_));
 b15xnr002ar1n02x5 _34912_ (.a(net491),
    .b(_13546_),
    .out0(_00240_));
 b15nand02ar1n02x5 _34913_ (.a(net947),
    .b(net131),
    .o1(_09446_));
 b15oai012ar1n02x5 _34914_ (.a(_09446_),
    .b(_12505_),
    .c(net947),
    .o1(_00393_));
 b15nanb02ar1n02x5 _34915_ (.a(net944),
    .b(\text_in_r[1] ),
    .out0(_09447_));
 b15aob012ar1n02x5 _34916_ (.a(_09447_),
    .b(net170),
    .c(net944),
    .out0(_00394_));
 b15ztpn00an1n08x5 PHY_24 ();
 b15nanb02ar1n02x5 _34918_ (.a(net944),
    .b(\text_in_r[2] ),
    .out0(_09450_));
 b15aob012ar1n02x5 _34919_ (.a(_09450_),
    .b(net181),
    .c(net944),
    .out0(_00395_));
 b15nanb02ar1n02x5 _34920_ (.a(net945),
    .b(\text_in_r[3] ),
    .out0(_09451_));
 b15aob012ar1n02x5 _34921_ (.a(_09451_),
    .b(net192),
    .c(net945),
    .out0(_00396_));
 b15nanb02ar1n02x5 _34922_ (.a(net943),
    .b(\text_in_r[4] ),
    .out0(_09452_));
 b15aob012ar1n02x5 _34923_ (.a(_09452_),
    .b(net203),
    .c(net943),
    .out0(_00397_));
 b15nand02ar1n02x5 _34924_ (.a(net936),
    .b(net214),
    .o1(_09453_));
 b15oai012ar1n02x5 _34925_ (.a(_09453_),
    .b(_15112_),
    .c(net936),
    .o1(_00398_));
 b15nand02ar1n02x5 _34926_ (.a(net944),
    .b(net225),
    .o1(_09454_));
 b15oai012ar1n02x5 _34927_ (.a(_09454_),
    .b(_15356_),
    .c(net944),
    .o1(_00399_));
 b15nanb02ar1n02x5 _34928_ (.a(net943),
    .b(\text_in_r[7] ),
    .out0(_09456_));
 b15ztpn00an1n08x5 PHY_23 ();
 b15ztpn00an1n08x5 PHY_22 ();
 b15aob012ar1n02x5 _34931_ (.a(_09456_),
    .b(net236),
    .c(net943),
    .out0(_00400_));
 b15ztpn00an1n08x5 PHY_21 ();
 b15nand02ar1n02x5 _34933_ (.a(net944),
    .b(net247),
    .o1(_09460_));
 b15oai012ar1n02x5 _34934_ (.a(_09460_),
    .b(_15807_),
    .c(net944),
    .o1(_00401_));
 b15nand02ar1n02x5 _34935_ (.a(net943),
    .b(net258),
    .o1(_09461_));
 b15oai012ar1n02x5 _34936_ (.a(_09461_),
    .b(_15810_),
    .c(net943),
    .o1(_00402_));
 b15nand02ar1n02x5 _34937_ (.a(net936),
    .b(net142),
    .o1(_09462_));
 b15oai012ar1n02x5 _34938_ (.a(_09462_),
    .b(_15816_),
    .c(net936),
    .o1(_00403_));
 b15nanb02ar1n02x5 _34939_ (.a(net943),
    .b(\text_in_r[11] ),
    .out0(_09464_));
 b15aob012ar1n02x5 _34940_ (.a(_09464_),
    .b(net153),
    .c(net943),
    .out0(_00404_));
 b15nand02ar1n02x5 _34941_ (.a(net943),
    .b(net162),
    .o1(_09465_));
 b15oai012ar1n02x5 _34942_ (.a(_09465_),
    .b(_15828_),
    .c(net943),
    .o1(_00405_));
 b15nand02ar1n02x5 _34943_ (.a(net943),
    .b(net163),
    .o1(_09466_));
 b15oai012al1n02x5 _34944_ (.a(_09466_),
    .b(_15839_),
    .c(net943),
    .o1(_00406_));
 b15nand02ar1n02x5 _34945_ (.a(net943),
    .b(net164),
    .o1(_09467_));
 b15ztpn00an1n08x5 PHY_20 ();
 b15oai012ar1n02x5 _34947_ (.a(_09467_),
    .b(_15844_),
    .c(net943),
    .o1(_00407_));
 b15nand02ar1n02x5 _34948_ (.a(net943),
    .b(net165),
    .o1(_09470_));
 b15oai012ar1n02x5 _34949_ (.a(_09470_),
    .b(_15849_),
    .c(net943),
    .o1(_00408_));
 b15nand02ar1n02x5 _34950_ (.a(net936),
    .b(net166),
    .o1(_09471_));
 b15oai012ar1n02x5 _34951_ (.a(_09471_),
    .b(_15852_),
    .c(net936),
    .o1(_00409_));
 b15nanb02ar1n02x5 _34952_ (.a(net939),
    .b(\text_in_r[17] ),
    .out0(_09472_));
 b15aob012ar1n02x5 _34953_ (.a(_09472_),
    .b(net167),
    .c(net939),
    .out0(_00410_));
 b15nand02ar1n02x5 _34954_ (.a(net939),
    .b(net168),
    .o1(_09473_));
 b15oai012ar1n02x5 _34955_ (.a(_09473_),
    .b(_15864_),
    .c(net939),
    .o1(_00411_));
 b15nanb02ar1n02x5 _34956_ (.a(net939),
    .b(\text_in_r[19] ),
    .out0(_09474_));
 b15aob012ar1n02x5 _34957_ (.a(_09474_),
    .b(net169),
    .c(net939),
    .out0(_00412_));
 b15nand02ar1n02x5 _34958_ (.a(net939),
    .b(net171),
    .o1(_09476_));
 b15oai012ar1n02x5 _34959_ (.a(_09476_),
    .b(_15876_),
    .c(net939),
    .o1(_00413_));
 b15ztpn00an1n08x5 PHY_19 ();
 b15nand02ar1n02x5 _34961_ (.a(net937),
    .b(net172),
    .o1(_09478_));
 b15oai012ar1n02x5 _34962_ (.a(_09478_),
    .b(_15883_),
    .c(net937),
    .o1(_00414_));
 b15nand02ar1n02x5 _34963_ (.a(net937),
    .b(net173),
    .o1(_09479_));
 b15oai012ar1n02x5 _34964_ (.a(_09479_),
    .b(_15885_),
    .c(net937),
    .o1(_00415_));
 b15nand02ar1n02x5 _34965_ (.a(net939),
    .b(net174),
    .o1(_09480_));
 b15oai012ar1n02x5 _34966_ (.a(_09480_),
    .b(_15893_),
    .c(net939),
    .o1(_00416_));
 b15nand02ar1n02x5 _34967_ (.a(net936),
    .b(net175),
    .o1(_09481_));
 b15oai012ar1n02x5 _34968_ (.a(_09481_),
    .b(_15895_),
    .c(net936),
    .o1(_00417_));
 b15nanb02ar1n02x5 _34969_ (.a(net943),
    .b(\text_in_r[25] ),
    .out0(_09483_));
 b15aob012ar1n02x5 _34970_ (.a(_09483_),
    .b(net176),
    .c(net943),
    .out0(_00418_));
 b15nand02ar1n02x5 _34971_ (.a(net944),
    .b(net177),
    .o1(_09484_));
 b15inv000al1n02x5 _34972_ (.a(\text_in_r[26] ),
    .o1(_09485_));
 b15oai012ar1n02x5 _34973_ (.a(_09484_),
    .b(_09485_),
    .c(net944),
    .o1(_00419_));
 b15nand02ar1n02x5 _34974_ (.a(net936),
    .b(net178),
    .o1(_09486_));
 b15ztpn00an1n08x5 PHY_18 ();
 b15oai012ar1n02x5 _34976_ (.a(_09486_),
    .b(_15909_),
    .c(net936),
    .o1(_00420_));
 b15nanb02ar1n02x5 _34977_ (.a(net943),
    .b(\text_in_r[28] ),
    .out0(_09488_));
 b15aob012ar1n02x5 _34978_ (.a(_09488_),
    .b(net179),
    .c(net943),
    .out0(_00421_));
 b15nanb02ar1n02x5 _34979_ (.a(net943),
    .b(\text_in_r[29] ),
    .out0(_09490_));
 b15aob012ar1n02x5 _34980_ (.a(_09490_),
    .b(net180),
    .c(net943),
    .out0(_00422_));
 b15nand02ar1n02x5 _34981_ (.a(net943),
    .b(net182),
    .o1(_09491_));
 b15oai012ar1n02x5 _34982_ (.a(_09491_),
    .b(_15926_),
    .c(net943),
    .o1(_00423_));
 b15nand02ar1n02x5 _34983_ (.a(net943),
    .b(net183),
    .o1(_09492_));
 b15oai012ar1n02x5 _34984_ (.a(_09492_),
    .b(_15930_),
    .c(net943),
    .o1(_00424_));
 b15nand02ar1n24x5 _34985_ (.a(net129),
    .b(net184),
    .o1(_09493_));
 b15oai012ar1n02x5 _34986_ (.a(_09493_),
    .b(_17072_),
    .c(net941),
    .o1(_00425_));
 b15ztpn00an1n08x5 PHY_17 ();
 b15nanb02ar1n02x5 _34988_ (.a(net938),
    .b(\text_in_r[33] ),
    .out0(_09496_));
 b15aob012ar1n02x5 _34989_ (.a(_09496_),
    .b(net185),
    .c(net938),
    .out0(_00426_));
 b15nand02ar1n02x5 _34990_ (.a(net938),
    .b(net186),
    .o1(_09497_));
 b15oai012ar1n02x5 _34991_ (.a(_09497_),
    .b(_17531_),
    .c(net938),
    .o1(_00427_));
 b15nanb02ar1n02x5 _34992_ (.a(net938),
    .b(\text_in_r[35] ),
    .out0(_09498_));
 b15aob012ar1n02x5 _34993_ (.a(_09498_),
    .b(net187),
    .c(net938),
    .out0(_00428_));
 b15nanb02ar1n02x5 _34994_ (.a(net937),
    .b(\text_in_r[36] ),
    .out0(_09499_));
 b15aob012ar1n02x5 _34995_ (.a(_09499_),
    .b(net188),
    .c(net937),
    .out0(_00429_));
 b15ztpn00an1n08x5 PHY_16 ();
 b15nand02ar1n02x5 _34997_ (.a(net937),
    .b(net189),
    .o1(_09501_));
 b15oai012ar1n02x5 _34998_ (.a(_09501_),
    .b(_01431_),
    .c(net937),
    .o1(_00430_));
 b15nand02ar1n02x5 _34999_ (.a(net937),
    .b(net190),
    .o1(_09503_));
 b15oai012ar1n02x5 _35000_ (.a(_09503_),
    .b(_01693_),
    .c(net937),
    .o1(_00431_));
 b15nanb02ar1n02x5 _35001_ (.a(net937),
    .b(\text_in_r[39] ),
    .out0(_09504_));
 b15ztpn00an1n08x5 PHY_15 ();
 b15aob012ar1n02x5 _35003_ (.a(_09504_),
    .b(net191),
    .c(net937),
    .out0(_00432_));
 b15nand02ar1n02x5 _35004_ (.a(net938),
    .b(net193),
    .o1(_09506_));
 b15oai012ar1n02x5 _35005_ (.a(_09506_),
    .b(_02129_),
    .c(net938),
    .o1(_00433_));
 b15nand02ar1n02x5 _35006_ (.a(net938),
    .b(net194),
    .o1(_09507_));
 b15oai012ar1n02x5 _35007_ (.a(_09507_),
    .b(_02131_),
    .c(net938),
    .o1(_00434_));
 b15nanb02ar1n02x5 _35008_ (.a(net938),
    .b(\text_in_r[42] ),
    .out0(_09509_));
 b15aob012ar1n02x5 _35009_ (.a(_09509_),
    .b(net195),
    .c(net938),
    .out0(_00435_));
 b15nand02ar1n02x5 _35010_ (.a(net938),
    .b(net196),
    .o1(_09510_));
 b15oai012ar1n02x5 _35011_ (.a(_09510_),
    .b(_02141_),
    .c(net938),
    .o1(_00436_));
 b15nanb02ar1n02x5 _35012_ (.a(net938),
    .b(\text_in_r[44] ),
    .out0(_09511_));
 b15aob012ar1n02x5 _35013_ (.a(_09511_),
    .b(net197),
    .c(net938),
    .out0(_00437_));
 b15nand02ar1n02x5 _35014_ (.a(net937),
    .b(net198),
    .o1(_09512_));
 b15ztpn00an1n08x5 PHY_14 ();
 b15oai012ar1n02x5 _35016_ (.a(_09512_),
    .b(_02152_),
    .c(net937),
    .o1(_00438_));
 b15nanb02ar1n02x5 _35017_ (.a(net938),
    .b(\text_in_r[46] ),
    .out0(_09514_));
 b15aob012ar1n02x5 _35018_ (.a(_09514_),
    .b(net199),
    .c(net938),
    .out0(_00439_));
 b15nand02ar1n02x5 _35019_ (.a(net938),
    .b(net200),
    .o1(_09516_));
 b15oai012ar1n02x5 _35020_ (.a(_09516_),
    .b(_02163_),
    .c(net938),
    .o1(_00440_));
 b15nand02ar1n02x5 _35021_ (.a(net937),
    .b(net201),
    .o1(_09517_));
 b15oai012ar1n02x5 _35022_ (.a(_09517_),
    .b(_02171_),
    .c(net937),
    .o1(_00441_));
 b15nanb02ar1n02x5 _35023_ (.a(net938),
    .b(\text_in_r[49] ),
    .out0(_09518_));
 b15aob012ar1n02x5 _35024_ (.a(_09518_),
    .b(net202),
    .c(net938),
    .out0(_00442_));
 b15nand02ar1n02x5 _35025_ (.a(net938),
    .b(net204),
    .o1(_09519_));
 b15oai012ar1n02x5 _35026_ (.a(_09519_),
    .b(_02178_),
    .c(net938),
    .o1(_00443_));
 b15nand02ar1n02x5 _35027_ (.a(net939),
    .b(net205),
    .o1(_09520_));
 b15oai012ar1n02x5 _35028_ (.a(_09520_),
    .b(_02183_),
    .c(net939),
    .o1(_00444_));
 b15ztpn00an1n08x5 PHY_13 ();
 b15nand02ar1n02x5 _35030_ (.a(net937),
    .b(net206),
    .o1(_09523_));
 b15oai012ar1n02x5 _35031_ (.a(_09523_),
    .b(_02188_),
    .c(net937),
    .o1(_00445_));
 b15nand02ar1n02x5 _35032_ (.a(net937),
    .b(net207),
    .o1(_09524_));
 b15oai012ar1n02x5 _35033_ (.a(_09524_),
    .b(_02196_),
    .c(net937),
    .o1(_00446_));
 b15nanb02ar1n02x5 _35034_ (.a(net937),
    .b(\text_in_r[54] ),
    .out0(_09525_));
 b15aob012ar1n02x5 _35035_ (.a(_09525_),
    .b(net208),
    .c(net937),
    .out0(_00447_));
 b15nand02ar1n02x5 _35036_ (.a(net937),
    .b(net209),
    .o1(_09526_));
 b15oai012ar1n02x5 _35037_ (.a(_09526_),
    .b(_02203_),
    .c(net937),
    .o1(_00448_));
 b15nand02ar1n02x5 _35038_ (.a(net938),
    .b(net210),
    .o1(_09528_));
 b15oai012ar1n02x5 _35039_ (.a(_09528_),
    .b(_02208_),
    .c(net938),
    .o1(_00449_));
 b15nandp2ar1n02x5 _35040_ (.a(net938),
    .b(net211),
    .o1(_09529_));
 b15oai012ar1n02x5 _35041_ (.a(_09529_),
    .b(_02212_),
    .c(net938),
    .o1(_00450_));
 b15nanb02ar1n02x5 _35042_ (.a(net938),
    .b(\text_in_r[58] ),
    .out0(_09530_));
 b15aob012ar1n02x5 _35043_ (.a(_09530_),
    .b(net212),
    .c(net938),
    .out0(_00451_));
 b15ztpn00an1n08x5 PHY_12 ();
 b15nanb02ar1n02x5 _35045_ (.a(net939),
    .b(\text_in_r[59] ),
    .out0(_09532_));
 b15aob012ar1n02x5 _35046_ (.a(_09532_),
    .b(net213),
    .c(net939),
    .out0(_00452_));
 b15nand02ar1n02x5 _35047_ (.a(net937),
    .b(net215),
    .o1(_09533_));
 b15ztpn00an1n08x5 PHY_11 ();
 b15oai012ar1n02x5 _35049_ (.a(_09533_),
    .b(_02225_),
    .c(net937),
    .o1(_00453_));
 b15nand02ar1n02x5 _35050_ (.a(net937),
    .b(net216),
    .o1(_09536_));
 b15oai012ar1n02x5 _35051_ (.a(_09536_),
    .b(_02232_),
    .c(net937),
    .o1(_00454_));
 b15nanb02ar1n02x5 _35052_ (.a(net937),
    .b(\text_in_r[62] ),
    .out0(_09537_));
 b15aob012ar1n02x5 _35053_ (.a(_09537_),
    .b(net217),
    .c(net937),
    .out0(_00455_));
 b15nand02ar1n02x5 _35054_ (.a(net937),
    .b(net218),
    .o1(_09538_));
 b15oai012ar1n02x5 _35055_ (.a(_09538_),
    .b(_02237_),
    .c(net937),
    .o1(_00456_));
 b15nanb02ar1n02x5 _35056_ (.a(net940),
    .b(\text_in_r[64] ),
    .out0(_09539_));
 b15aob012ar1n02x5 _35057_ (.a(_09539_),
    .b(net219),
    .c(net940),
    .out0(_00457_));
 b15nand02an1n16x5 _35058_ (.a(net947),
    .b(net220),
    .o1(_09541_));
 b15oai012ar1n02x5 _35059_ (.a(_09541_),
    .b(_03418_),
    .c(net945),
    .o1(_00458_));
 b15nanb02ar1n02x5 _35060_ (.a(net942),
    .b(\text_in_r[66] ),
    .out0(_09542_));
 b15ztpn00an1n08x5 PHY_10 ();
 b15aob012ar1n02x5 _35062_ (.a(_09542_),
    .b(net221),
    .c(net942),
    .out0(_00459_));
 b15nanb02ar1n02x5 _35063_ (.a(net940),
    .b(\text_in_r[67] ),
    .out0(_09544_));
 b15aob012ar1n02x5 _35064_ (.a(_09544_),
    .b(net222),
    .c(net940),
    .out0(_00460_));
 b15nand02ar1n02x5 _35065_ (.a(net939),
    .b(net223),
    .o1(_09545_));
 b15oai012ar1n02x5 _35066_ (.a(_09545_),
    .b(_04648_),
    .c(net939),
    .o1(_00461_));
 b15nanb02ar1n02x5 _35067_ (.a(net939),
    .b(\text_in_r[69] ),
    .out0(_09546_));
 b15aob012ar1n02x5 _35068_ (.a(_09546_),
    .b(net224),
    .c(net939),
    .out0(_00462_));
 b15ztpn00an1n08x5 PHY_9 ();
 b15nand02ar1n02x5 _35070_ (.a(net939),
    .b(net226),
    .o1(_09549_));
 b15oai012ar1n02x5 _35071_ (.a(_09549_),
    .b(_05489_),
    .c(net939),
    .o1(_00463_));
 b15nand02ar1n02x5 _35072_ (.a(net940),
    .b(net227),
    .o1(_09550_));
 b15oai012ar1n02x5 _35073_ (.a(_09550_),
    .b(_05684_),
    .c(net940),
    .o1(_00464_));
 b15nand02ar1n02x5 _35074_ (.a(net940),
    .b(net228),
    .o1(_09551_));
 b15oai012ar1n02x5 _35075_ (.a(_09551_),
    .b(_05686_),
    .c(net940),
    .o1(_00465_));
 b15nanb02ar1n02x5 _35076_ (.a(net945),
    .b(\text_in_r[73] ),
    .out0(_09552_));
 b15aob012ar1n02x5 _35077_ (.a(_09552_),
    .b(net229),
    .c(net945),
    .out0(_00466_));
 b15nanb02ar1n02x5 _35078_ (.a(net946),
    .b(\text_in_r[74] ),
    .out0(_09554_));
 b15aob012ar1n02x5 _35079_ (.a(_09554_),
    .b(net230),
    .c(net946),
    .out0(_00467_));
 b15nanb02ar1n02x5 _35080_ (.a(net946),
    .b(\text_in_r[75] ),
    .out0(_09555_));
 b15aob012ar1n02x5 _35081_ (.a(_09555_),
    .b(net231),
    .c(net946),
    .out0(_00468_));
 b15nanb02ar1n02x5 _35082_ (.a(net940),
    .b(\text_in_r[76] ),
    .out0(_09556_));
 b15aob012ar1n02x5 _35083_ (.a(_09556_),
    .b(net232),
    .c(net940),
    .out0(_00469_));
 b15nand02ar1n02x5 _35084_ (.a(net939),
    .b(net233),
    .o1(_09557_));
 b15oai012ar1n02x5 _35085_ (.a(_09557_),
    .b(_05716_),
    .c(net939),
    .o1(_00470_));
 b15nand02ar1n02x5 _35086_ (.a(net939),
    .b(net234),
    .o1(_09558_));
 b15oai012ar1n02x5 _35087_ (.a(_09558_),
    .b(_05722_),
    .c(net939),
    .o1(_00471_));
 b15nand02ar1n02x5 _35088_ (.a(net936),
    .b(net235),
    .o1(_09560_));
 b15ztpn00an1n08x5 PHY_8 ();
 b15oai012ar1n02x5 _35090_ (.a(_09560_),
    .b(_05724_),
    .c(net936),
    .o1(_00472_));
 b15nand02ar1n02x5 _35091_ (.a(net947),
    .b(net237),
    .o1(_09562_));
 b15oai012ar1n02x5 _35092_ (.a(_09562_),
    .b(_05730_),
    .c(net947),
    .o1(_00473_));
 b15nand02ar1n02x5 _35093_ (.a(net945),
    .b(net238),
    .o1(_09563_));
 b15oai012ar1n02x5 _35094_ (.a(_09563_),
    .b(_05735_),
    .c(net945),
    .o1(_00474_));
 b15nand02ar1n02x5 _35095_ (.a(net947),
    .b(net239),
    .o1(_09564_));
 b15oai012ar1n02x5 _35096_ (.a(_09564_),
    .b(_05740_),
    .c(net947),
    .o1(_00475_));
 b15ztpn00an1n08x5 PHY_7 ();
 b15nanb02ar1n02x5 _35098_ (.a(net946),
    .b(\text_in_r[83] ),
    .out0(_09567_));
 b15aob012ar1n02x5 _35099_ (.a(_09567_),
    .b(net240),
    .c(net946),
    .out0(_00476_));
 b15nand02ar1n02x5 _35100_ (.a(net944),
    .b(net241),
    .o1(_09568_));
 b15oai012ar1n02x5 _35101_ (.a(_09568_),
    .b(_05752_),
    .c(net944),
    .o1(_00477_));
 b15nanb02ar1n02x5 _35102_ (.a(net936),
    .b(\text_in_r[85] ),
    .out0(_09569_));
 b15aob012ar1n02x5 _35103_ (.a(_09569_),
    .b(net242),
    .c(net936),
    .out0(_00478_));
 b15ztpn00an1n08x5 PHY_6 ();
 b15nand02ar1n02x5 _35105_ (.a(net936),
    .b(net243),
    .o1(_09571_));
 b15oai012ar1n02x5 _35106_ (.a(_09571_),
    .b(_05765_),
    .c(net936),
    .o1(_00479_));
 b15nand02ar1n02x5 _35107_ (.a(net943),
    .b(net244),
    .o1(_09572_));
 b15oai012ar1n02x5 _35108_ (.a(_09572_),
    .b(_05772_),
    .c(net943),
    .o1(_00480_));
 b15nand02ar1n02x5 _35109_ (.a(net944),
    .b(net245),
    .o1(_09574_));
 b15oai012ar1n02x5 _35110_ (.a(_09574_),
    .b(_05775_),
    .c(net944),
    .o1(_00481_));
 b15nanb02ar1n02x5 _35111_ (.a(net945),
    .b(\text_in_r[89] ),
    .out0(_09575_));
 b15aob012ar1n02x5 _35112_ (.a(_09575_),
    .b(net246),
    .c(net945),
    .out0(_00482_));
 b15nand02ar1n02x5 _35113_ (.a(net944),
    .b(net248),
    .o1(_09576_));
 b15oai012ar1n02x5 _35114_ (.a(_09576_),
    .b(_05787_),
    .c(net944),
    .o1(_00483_));
 b15nandp2as1n08x5 _35115_ (.a(net129),
    .b(net249),
    .o1(_09577_));
 b15oai012ar1n02x5 _35116_ (.a(_09577_),
    .b(_05789_),
    .c(net945),
    .o1(_00484_));
 b15nanb02ar1n02x5 _35117_ (.a(net936),
    .b(\text_in_r[92] ),
    .out0(_09578_));
 b15ztpn00an1n08x5 PHY_5 ();
 b15aob012ar1n02x5 _35119_ (.a(_09578_),
    .b(net250),
    .c(net936),
    .out0(_00485_));
 b15nand02ar1n02x5 _35120_ (.a(net936),
    .b(net251),
    .o1(_09581_));
 b15ztpn00an1n08x5 PHY_4 ();
 b15oai012ar1n02x5 _35122_ (.a(_09581_),
    .b(_05799_),
    .c(net936),
    .o1(_00486_));
 b15nand02ar1n02x5 _35123_ (.a(net936),
    .b(net252),
    .o1(_09583_));
 b15oai012ar1n02x5 _35124_ (.a(_09583_),
    .b(_05807_),
    .c(net936),
    .o1(_00487_));
 b15nand02ar1n02x5 _35125_ (.a(net936),
    .b(net253),
    .o1(_09584_));
 b15oai012ar1n02x5 _35126_ (.a(_09584_),
    .b(_05812_),
    .c(net936),
    .o1(_00488_));
 b15nand02ar1n02x5 _35127_ (.a(net948),
    .b(net254),
    .o1(_09585_));
 b15oai012ar1n02x5 _35128_ (.a(_09585_),
    .b(_05814_),
    .c(net948),
    .o1(_00489_));
 b15nanb02ar1n02x5 _35129_ (.a(net946),
    .b(\text_in_r[97] ),
    .out0(_09587_));
 b15aob012ar1n02x5 _35130_ (.a(_09587_),
    .b(net255),
    .c(net946),
    .out0(_00490_));
 b15nandp2ar1n02x5 _35131_ (.a(net129),
    .b(net256),
    .o1(_09588_));
 b15oai012ar1n02x5 _35132_ (.a(_09588_),
    .b(_07890_),
    .c(net948),
    .o1(_00491_));
 b15ztpn00an1n08x5 PHY_3 ();
 b15nand02ah1n02x5 _35134_ (.a(net129),
    .b(net257),
    .o1(_09590_));
 b15oai012ar1n02x5 _35135_ (.a(_09590_),
    .b(_07892_),
    .c(net948),
    .o1(_00492_));
 b15nanb02ar1n02x5 _35136_ (.a(net948),
    .b(\text_in_r[100] ),
    .out0(_09591_));
 b15aob012ar1n02x5 _35137_ (.a(_09591_),
    .b(net132),
    .c(net948),
    .out0(_00493_));
 b15nanb02ar1n02x5 _35138_ (.a(net129),
    .b(\text_in_r[101] ),
    .out0(_09593_));
 b15aob012ar1n02x5 _35139_ (.a(_09593_),
    .b(net133),
    .c(net129),
    .out0(_00494_));
 b15nanb02ar1n02x5 _35140_ (.a(net941),
    .b(\text_in_r[102] ),
    .out0(_09594_));
 b15aob012ar1n02x5 _35141_ (.a(_09594_),
    .b(net134),
    .c(net941),
    .out0(_00495_));
 b15nand02ar1n02x5 _35142_ (.a(net948),
    .b(net135),
    .o1(_09595_));
 b15oai012ar1n02x5 _35143_ (.a(_09595_),
    .b(_09093_),
    .c(net948),
    .o1(_00496_));
 b15nandp2al1n02x5 _35144_ (.a(net129),
    .b(net136),
    .o1(_09596_));
 b15oai012ar1n02x5 _35145_ (.a(_09596_),
    .b(_09320_),
    .c(net948),
    .o1(_00497_));
 b15nanb02ar1n02x5 _35146_ (.a(net129),
    .b(\text_in_r[105] ),
    .out0(_09597_));
 b15aob012ar1n02x5 _35147_ (.a(_09597_),
    .b(net137),
    .c(net129),
    .out0(_00498_));
 b15nand02ar1n02x5 _35148_ (.a(net941),
    .b(net138),
    .o1(_09599_));
 b15oai012ar1n02x5 _35149_ (.a(_09599_),
    .b(_09330_),
    .c(net941),
    .o1(_00499_));
 b15nanb02ar1n02x5 _35150_ (.a(net941),
    .b(\text_in_r[107] ),
    .out0(_09600_));
 b15aob012ar1n02x5 _35151_ (.a(_09600_),
    .b(net139),
    .c(net941),
    .out0(_00500_));
 b15nanb02ar1n02x5 _35152_ (.a(net941),
    .b(\text_in_r[108] ),
    .out0(_09601_));
 b15aob012ar1n02x5 _35153_ (.a(_09601_),
    .b(net140),
    .c(net941),
    .out0(_00501_));
 b15nand02ar1n02x5 _35154_ (.a(net941),
    .b(net141),
    .o1(_09602_));
 b15oai012ar1n02x5 _35155_ (.a(_09602_),
    .b(_09344_),
    .c(net941),
    .o1(_00502_));
 b15nand02ar1n02x5 _35156_ (.a(net941),
    .b(net143),
    .o1(_09603_));
 b15ztpn00an1n08x5 PHY_2 ();
 b15oai012ar1n02x5 _35158_ (.a(_09603_),
    .b(_09350_),
    .c(net941),
    .o1(_00503_));
 b15nand02ar1n02x5 _35159_ (.a(net941),
    .b(net144),
    .o1(_09606_));
 b15oai012ar1n02x5 _35160_ (.a(_09606_),
    .b(_09356_),
    .c(net941),
    .o1(_00504_));
 b15nandp2ar1n03x5 _35161_ (.a(net947),
    .b(net145),
    .o1(_09607_));
 b15oai012ar1n02x5 _35162_ (.a(_09607_),
    .b(_09363_),
    .c(net947),
    .o1(_00505_));
 b15nand02ar1n02x5 _35163_ (.a(net946),
    .b(net146),
    .o1(_09608_));
 b15oai012ar1n02x5 _35164_ (.a(_09608_),
    .b(_09366_),
    .c(net946),
    .o1(_00506_));
 b15nanb02ar1n02x5 _35165_ (.a(net946),
    .b(\text_in_r[114] ),
    .out0(_09609_));
 b15aob012ar1n02x5 _35166_ (.a(_09609_),
    .b(net147),
    .c(net946),
    .out0(_00507_));
 b15nanb02ar1n02x5 _35167_ (.a(net129),
    .b(\text_in_r[115] ),
    .out0(_09610_));
 b15aob012ar1n02x5 _35168_ (.a(_09610_),
    .b(net148),
    .c(net129),
    .out0(_00508_));
 b15nand02ar1n02x5 _35169_ (.a(net946),
    .b(net149),
    .o1(_09612_));
 b15oai012ar1n02x5 _35170_ (.a(_09612_),
    .b(_09380_),
    .c(net946),
    .o1(_00509_));
 b15nand02ar1n02x5 _35171_ (.a(net945),
    .b(net150),
    .o1(_09613_));
 b15oai012ar1n02x5 _35172_ (.a(_09613_),
    .b(_09389_),
    .c(net945),
    .o1(_00510_));
 b15nand02ar1n02x5 _35173_ (.a(net129),
    .b(net151),
    .o1(_09614_));
 b15oai012ar1n02x5 _35174_ (.a(_09614_),
    .b(_09391_),
    .c(net948),
    .o1(_00511_));
 b15nanb02ar1n02x5 _35175_ (.a(net947),
    .b(\text_in_r[119] ),
    .out0(_09615_));
 b15aob012ar1n02x5 _35176_ (.a(_09615_),
    .b(net152),
    .c(net947),
    .out0(_00512_));
 b15nandp2al1n02x5 _35177_ (.a(net129),
    .b(net154),
    .o1(_09616_));
 b15oai012ar1n02x5 _35178_ (.a(_09616_),
    .b(_09398_),
    .c(net129),
    .o1(_00513_));
 b15nanb02ar1n02x5 _35179_ (.a(net948),
    .b(\text_in_r[121] ),
    .out0(_09618_));
 b15aob012ar1n02x5 _35180_ (.a(_09618_),
    .b(net155),
    .c(net948),
    .out0(_00514_));
 b15nand02al1n04x5 _35181_ (.a(net129),
    .b(net156),
    .o1(_09619_));
 b15oai012ar1n02x5 _35182_ (.a(_09619_),
    .b(_09409_),
    .c(net129),
    .o1(_00515_));
 b15nand02ar1n02x5 _35183_ (.a(net129),
    .b(net157),
    .o1(_09620_));
 b15oai012ar1n02x5 _35184_ (.a(_09620_),
    .b(_09412_),
    .c(net129),
    .o1(_00516_));
 b15nanb02ar1n02x5 _35185_ (.a(net129),
    .b(\text_in_r[124] ),
    .out0(_09621_));
 b15aob012ar1n02x5 _35186_ (.a(_09621_),
    .b(net158),
    .c(net129),
    .out0(_00517_));
 b15nanb02ar1n02x5 _35187_ (.a(net129),
    .b(\text_in_r[125] ),
    .out0(_09622_));
 b15aob012ar1n02x5 _35188_ (.a(_09622_),
    .b(net159),
    .c(net129),
    .out0(_00518_));
 b15nand02ar1n02x5 _35189_ (.a(net129),
    .b(net160),
    .o1(_09624_));
 b15oai012ar1n02x5 _35190_ (.a(_09624_),
    .b(_09424_),
    .c(net129),
    .o1(_00519_));
 b15nand02ar1n02x5 _35191_ (.a(net948),
    .b(net161),
    .o1(_09625_));
 b15oai012ar1n02x5 _35192_ (.a(_09625_),
    .b(_09430_),
    .c(net948),
    .o1(_00520_));
 b15ztpn00an1n08x5 PHY_1 ();
 b15nand03ah1n04x5 _35194_ (.a(\u0.r0.rcnt[0] ),
    .b(\u0.r0.rcnt[1] ),
    .c(\u0.r0.rcnt[2] ),
    .o1(_09627_));
 b15nanb02ar1n02x5 _35195_ (.a(net945),
    .b(_09627_),
    .out0(_00385_));
 b15nor003ah1n02x5 _35196_ (.a(\u0.r0.rcnt[0] ),
    .b(\u0.r0.rcnt[1] ),
    .c(\u0.r0.rcnt[2] ),
    .o1(_09628_));
 b15ztpn00an1n08x5 PHY_0 ();
 b15norp02an1n02x5 _35198_ (.a(\u0.r0.rcnt[3] ),
    .b(_09627_),
    .o1(_09631_));
 b15oab012al1n02x5 _35199_ (.a(net945),
    .b(_09628_),
    .c(_09631_),
    .out0(_00386_));
 b15xnr002ar1n02x5 _35200_ (.a(\u0.r0.rcnt[0] ),
    .b(\u0.r0.rcnt[3] ),
    .out0(_09632_));
 b15nor004al1n02x5 _35201_ (.a(\u0.r0.rcnt[1] ),
    .b(\u0.r0.rcnt[2] ),
    .c(net945),
    .d(_09632_),
    .o1(_00387_));
 b15xor002ar1n02x5 _35202_ (.a(\u0.r0.rcnt[0] ),
    .b(\u0.r0.rcnt[2] ),
    .out0(_09633_));
 b15nanb02al1n02x5 _35203_ (.a(net942),
    .b(\u0.r0.rcnt[1] ),
    .out0(_09634_));
 b15norp03an1n02x5 _35204_ (.a(\u0.r0.rcnt[3] ),
    .b(_09633_),
    .c(_09634_),
    .o1(_00388_));
 b15nand02ar1n02x5 _35205_ (.a(\u0.r0.rcnt[3] ),
    .b(_09628_),
    .o1(_09635_));
 b15nand02al1n03x5 _35206_ (.a(\u0.r0.rcnt[0] ),
    .b(\u0.r0.rcnt[1] ),
    .o1(_09636_));
 b15oaoi13al1n02x5 _35207_ (.a(net942),
    .b(_09635_),
    .c(_09636_),
    .d(\u0.r0.rcnt[3] ),
    .o1(_00389_));
 b15inv020an1n04x5 _35208_ (.a(\u0.r0.rcnt[2] ),
    .o1(_09638_));
 b15xor002ar1n02x5 _35209_ (.a(_09638_),
    .b(\u0.r0.rcnt[3] ),
    .out0(_09639_));
 b15nor004al1n03x5 _35210_ (.a(\u0.r0.rcnt[0] ),
    .b(\u0.r0.rcnt[1] ),
    .c(net942),
    .d(_09639_),
    .o1(_00390_));
 b15nor004al1n02x5 _35211_ (.a(\u0.r0.rcnt[1] ),
    .b(_09638_),
    .c(\u0.r0.rcnt[3] ),
    .d(net942),
    .o1(_09640_));
 b15and002al1n02x5 _35212_ (.a(\u0.r0.rcnt[0] ),
    .b(_09640_),
    .o(_00391_));
 b15nor004ah1n03x5 _35213_ (.a(\u0.r0.rcnt[0] ),
    .b(_09638_),
    .c(\u0.r0.rcnt[3] ),
    .d(_09634_),
    .o1(_00392_));
 b15oai012ar1n02x5 _35214_ (.a(\dcnt[2] ),
    .b(\dcnt[0] ),
    .c(\dcnt[1] ),
    .o1(_09641_));
 b15nanb02ar1n02x5 _35215_ (.a(\dcnt[2] ),
    .b(\dcnt[3] ),
    .out0(_09642_));
 b15oai013ar1n02x5 _35216_ (.a(_09641_),
    .b(_09642_),
    .c(\dcnt[0] ),
    .d(\dcnt[1] ),
    .o1(_09643_));
 b15nano22ar1n02x5 _35217_ (.a(net130),
    .b(_09643_),
    .c(net947),
    .out0(_00524_));
 b15norp02ar1n02x5 _35218_ (.a(\u0.r0.rcnt[0] ),
    .b(net942),
    .o1(_00525_));
 b15xnr002ar1n02x5 _35219_ (.a(\u0.r0.rcnt[0] ),
    .b(\u0.r0.rcnt[1] ),
    .out0(_09645_));
 b15norp02ar1n02x5 _35220_ (.a(net942),
    .b(_09645_),
    .o1(_00526_));
 b15xor002ar1n02x5 _35221_ (.a(\u0.r0.rcnt[2] ),
    .b(_09636_),
    .out0(_09646_));
 b15norp02ar1n02x5 _35222_ (.a(net946),
    .b(_09646_),
    .o1(_00527_));
 b15and002ar1n02x5 _35223_ (.a(\u0.r0.rcnt[3] ),
    .b(_09627_),
    .o(_09647_));
 b15oab012ar1n02x5 _35224_ (.a(net945),
    .b(_09631_),
    .c(_09647_),
    .out0(_00528_));
 b15norp02ar1n02x5 _35225_ (.a(\dcnt[0] ),
    .b(_12504_),
    .o1(_09648_));
 b15oa0012ar1n02x5 _35226_ (.a(net130),
    .b(_09648_),
    .c(net947),
    .o(_00521_));
 b15aoi012ar1n02x5 _35227_ (.a(net947),
    .b(\dcnt[0] ),
    .c(\dcnt[1] ),
    .o1(_09649_));
 b15norp02ar1n02x5 _35228_ (.a(\dcnt[2] ),
    .b(\dcnt[3] ),
    .o1(_09651_));
 b15oai013ar1n02x5 _35229_ (.a(_09649_),
    .b(_09651_),
    .c(\dcnt[0] ),
    .d(\dcnt[1] ),
    .o1(_09652_));
 b15and002ar1n02x5 _35230_ (.a(net130),
    .b(_09652_),
    .o(_00522_));
 b15oai013ar1n02x5 _35231_ (.a(\dcnt[3] ),
    .b(\dcnt[2] ),
    .c(\dcnt[0] ),
    .d(\dcnt[1] ),
    .o1(_09653_));
 b15nanb02ar1n02x5 _35232_ (.a(net947),
    .b(_09653_),
    .out0(_09654_));
 b15and002ar1n02x5 _35233_ (.a(net130),
    .b(_09654_),
    .o(_00523_));
 b15fpn000hn1n04x5 _35234_ (.clk(clknet_leaf_9_clk),
    .d(_00385_),
    .o(\u0.r0.out[24] ));
 b15fpn000hn1n04x5 _35235_ (.clk(clknet_leaf_8_clk),
    .d(_00386_),
    .o(\u0.r0.out[25] ));
 b15fpn000hn1n04x5 _35236_ (.clk(clknet_leaf_8_clk),
    .d(_00387_),
    .o(\u0.r0.out[26] ));
 b15fpn000hn1n04x5 _35237_ (.clk(clknet_leaf_11_clk),
    .d(_00388_),
    .o(\u0.r0.out[27] ));
 b15fpn000hn1n04x5 _35238_ (.clk(clknet_leaf_8_clk),
    .d(_00389_),
    .o(\u0.r0.out[28] ));
 b15fpn000hn1n04x5 _35239_ (.clk(clknet_leaf_10_clk),
    .d(_00390_),
    .o(\u0.r0.out[29] ));
 b15fpn000hn1n04x5 _35240_ (.clk(clknet_leaf_11_clk),
    .d(_00391_),
    .o(\u0.r0.out[30] ));
 b15fpn000hn1n04x5 _35241_ (.clk(clknet_leaf_11_clk),
    .d(_00392_),
    .o(\u0.r0.out[31] ));
 b15fpn000hn1n04x5 _35242_ (.clk(clknet_leaf_7_clk),
    .d(_00393_),
    .o(\text_in_r[0] ));
 b15fpn000hn1n04x5 _35243_ (.clk(clknet_leaf_4_clk),
    .d(_00394_),
    .o(\text_in_r[1] ));
 b15fpn000hn1n04x5 _35244_ (.clk(clknet_leaf_4_clk),
    .d(_00395_),
    .o(\text_in_r[2] ));
 b15fpn000hn1n04x5 _35245_ (.clk(clknet_leaf_10_clk),
    .d(_00396_),
    .o(\text_in_r[3] ));
 b15fpn000hn1n04x5 _35246_ (.clk(clknet_leaf_3_clk),
    .d(_00397_),
    .o(\text_in_r[4] ));
 b15fpn000hn1n04x5 _35247_ (.clk(clknet_leaf_2_clk),
    .d(_00398_),
    .o(\text_in_r[5] ));
 b15fpn000hn1n04x5 _35248_ (.clk(clknet_leaf_4_clk),
    .d(_00399_),
    .o(\text_in_r[6] ));
 b15fpn000hn1n04x5 _35249_ (.clk(clknet_leaf_4_clk),
    .d(_00400_),
    .o(\text_in_r[7] ));
 b15fpn000hn1n04x5 _35250_ (.clk(clknet_leaf_5_clk),
    .d(_00401_),
    .o(\text_in_r[8] ));
 b15fpn000hn1n04x5 _35251_ (.clk(clknet_leaf_3_clk),
    .d(_00402_),
    .o(\text_in_r[9] ));
 b15fpn000hn1n04x5 _35252_ (.clk(clknet_leaf_2_clk),
    .d(_00403_),
    .o(\text_in_r[10] ));
 b15fpn000hn1n04x5 _35253_ (.clk(clknet_leaf_3_clk),
    .d(_00404_),
    .o(\text_in_r[11] ));
 b15fpn000hn1n04x5 _35254_ (.clk(clknet_leaf_3_clk),
    .d(_00405_),
    .o(\text_in_r[12] ));
 b15fpn000hn1n04x5 _35255_ (.clk(clknet_leaf_3_clk),
    .d(_00406_),
    .o(\text_in_r[13] ));
 b15fpn000hn1n04x5 _35256_ (.clk(clknet_leaf_3_clk),
    .d(_00407_),
    .o(\text_in_r[14] ));
 b15fpn000hn1n04x5 _35257_ (.clk(clknet_leaf_3_clk),
    .d(_00408_),
    .o(\text_in_r[15] ));
 b15fpn000hn1n04x5 _35258_ (.clk(clknet_leaf_2_clk),
    .d(_00409_),
    .o(\text_in_r[16] ));
 b15fpn000hn1n04x5 _35259_ (.clk(clknet_leaf_18_clk),
    .d(_00410_),
    .o(\text_in_r[17] ));
 b15fpn000hn1n04x5 _35260_ (.clk(clknet_leaf_18_clk),
    .d(_00411_),
    .o(\text_in_r[18] ));
 b15fpn000hn1n04x5 _35261_ (.clk(clknet_leaf_18_clk),
    .d(_00412_),
    .o(\text_in_r[19] ));
 b15fpn000hn1n04x5 _35262_ (.clk(clknet_leaf_18_clk),
    .d(_00413_),
    .o(\text_in_r[20] ));
 b15fpn000hn1n04x5 _35263_ (.clk(clknet_leaf_18_clk),
    .d(_00414_),
    .o(\text_in_r[21] ));
 b15fpn000hn1n04x5 _35264_ (.clk(clknet_leaf_18_clk),
    .d(_00415_),
    .o(\text_in_r[22] ));
 b15fpn000hn1n04x5 _35265_ (.clk(clknet_leaf_18_clk),
    .d(_00416_),
    .o(\text_in_r[23] ));
 b15fpn000hn1n04x5 _35266_ (.clk(clknet_leaf_2_clk),
    .d(_00417_),
    .o(\text_in_r[24] ));
 b15fpn000hn1n04x5 _35267_ (.clk(clknet_leaf_3_clk),
    .d(_00418_),
    .o(\text_in_r[25] ));
 b15fpn000hn1n04x5 _35268_ (.clk(clknet_leaf_4_clk),
    .d(_00419_),
    .o(\text_in_r[26] ));
 b15fpn000hn1n04x5 _35269_ (.clk(clknet_leaf_2_clk),
    .d(_00420_),
    .o(\text_in_r[27] ));
 b15fpn000hn1n04x5 _35270_ (.clk(clknet_leaf_3_clk),
    .d(_00421_),
    .o(\text_in_r[28] ));
 b15fpn000hn1n04x5 _35271_ (.clk(clknet_leaf_3_clk),
    .d(_00422_),
    .o(\text_in_r[29] ));
 b15fpn000hn1n04x5 _35272_ (.clk(clknet_leaf_3_clk),
    .d(_00423_),
    .o(\text_in_r[30] ));
 b15fpn000hn1n04x5 _35273_ (.clk(clknet_leaf_3_clk),
    .d(_00424_),
    .o(\text_in_r[31] ));
 b15fpn000hn1n04x5 _35274_ (.clk(clknet_leaf_10_clk),
    .d(_00425_),
    .o(\text_in_r[32] ));
 b15fpn000hn1n04x5 _35275_ (.clk(clknet_leaf_16_clk),
    .d(_00426_),
    .o(\text_in_r[33] ));
 b15fpn000hn1n04x5 _35276_ (.clk(clknet_leaf_16_clk),
    .d(_00427_),
    .o(\text_in_r[34] ));
 b15fpn000hn1n04x5 _35277_ (.clk(clknet_leaf_16_clk),
    .d(_00428_),
    .o(\text_in_r[35] ));
 b15fpn000hn1n04x5 _35278_ (.clk(clknet_leaf_16_clk),
    .d(_00429_),
    .o(\text_in_r[36] ));
 b15fpn000hn1n04x5 _35279_ (.clk(clknet_leaf_18_clk),
    .d(_00430_),
    .o(\text_in_r[37] ));
 b15fpn000hn1n04x5 _35280_ (.clk(clknet_leaf_17_clk),
    .d(_00431_),
    .o(\text_in_r[38] ));
 b15fpn000hn1n04x5 _35281_ (.clk(clknet_leaf_17_clk),
    .d(_00432_),
    .o(\text_in_r[39] ));
 b15fpn000hn1n04x5 _35282_ (.clk(clknet_leaf_14_clk),
    .d(_00433_),
    .o(\text_in_r[40] ));
 b15fpn000hn1n04x5 _35283_ (.clk(clknet_leaf_14_clk),
    .d(_00434_),
    .o(\text_in_r[41] ));
 b15fpn000hn1n04x5 _35284_ (.clk(clknet_leaf_15_clk),
    .d(_00435_),
    .o(\text_in_r[42] ));
 b15fpn000hn1n04x5 _35285_ (.clk(clknet_leaf_14_clk),
    .d(_00436_),
    .o(\text_in_r[43] ));
 b15fpn000hn1n04x5 _35286_ (.clk(clknet_leaf_16_clk),
    .d(_00437_),
    .o(\text_in_r[44] ));
 b15fpn000hn1n04x5 _35287_ (.clk(clknet_leaf_17_clk),
    .d(_00438_),
    .o(\text_in_r[45] ));
 b15fpn000hn1n04x5 _35288_ (.clk(clknet_leaf_16_clk),
    .d(_00439_),
    .o(\text_in_r[46] ));
 b15fpn000hn1n04x5 _35289_ (.clk(clknet_leaf_17_clk),
    .d(_00440_),
    .o(\text_in_r[47] ));
 b15fpn000hn1n04x5 _35290_ (.clk(clknet_leaf_17_clk),
    .d(_00441_),
    .o(\text_in_r[48] ));
 b15fpn000hn1n04x5 _35291_ (.clk(clknet_leaf_16_clk),
    .d(_00442_),
    .o(\text_in_r[49] ));
 b15fpn000hn1n04x5 _35292_ (.clk(clknet_leaf_16_clk),
    .d(_00443_),
    .o(\text_in_r[50] ));
 b15fpn000hn1n04x5 _35293_ (.clk(clknet_leaf_17_clk),
    .d(_00444_),
    .o(\text_in_r[51] ));
 b15fpn000hn1n04x5 _35294_ (.clk(clknet_leaf_18_clk),
    .d(_00445_),
    .o(\text_in_r[52] ));
 b15fpn000hn1n04x5 _35295_ (.clk(clknet_leaf_18_clk),
    .d(_00446_),
    .o(\text_in_r[53] ));
 b15fpn000hn1n04x5 _35296_ (.clk(clknet_leaf_18_clk),
    .d(_00447_),
    .o(\text_in_r[54] ));
 b15fpn000hn1n04x5 _35297_ (.clk(clknet_leaf_17_clk),
    .d(_00448_),
    .o(\text_in_r[55] ));
 b15fpn000hn1n04x5 _35298_ (.clk(clknet_leaf_15_clk),
    .d(_00449_),
    .o(\text_in_r[56] ));
 b15fpn000hn1n04x5 _35299_ (.clk(clknet_leaf_15_clk),
    .d(_00450_),
    .o(\text_in_r[57] ));
 b15fpn000hn1n04x5 _35300_ (.clk(clknet_leaf_16_clk),
    .d(_00451_),
    .o(\text_in_r[58] ));
 b15fpn000hn1n04x5 _35301_ (.clk(clknet_leaf_17_clk),
    .d(_00452_),
    .o(\text_in_r[59] ));
 b15fpn000hn1n04x5 _35302_ (.clk(clknet_leaf_16_clk),
    .d(_00453_),
    .o(\text_in_r[60] ));
 b15fpn000hn1n04x5 _35303_ (.clk(clknet_leaf_18_clk),
    .d(_00454_),
    .o(\text_in_r[61] ));
 b15fpn000hn1n04x5 _35304_ (.clk(clknet_leaf_18_clk),
    .d(_00455_),
    .o(\text_in_r[62] ));
 b15fpn000hn1n04x5 _35305_ (.clk(clknet_leaf_17_clk),
    .d(_00456_),
    .o(\text_in_r[63] ));
 b15fpn000hn1n04x5 _35306_ (.clk(clknet_leaf_15_clk),
    .d(_00457_),
    .o(\text_in_r[64] ));
 b15fpn000hn1n04x5 _35307_ (.clk(clknet_leaf_5_clk),
    .d(_00458_),
    .o(\text_in_r[65] ));
 b15fpn000hn1n04x5 _35308_ (.clk(clknet_leaf_10_clk),
    .d(_00459_),
    .o(\text_in_r[66] ));
 b15fpn000hn1n04x5 _35309_ (.clk(clknet_leaf_15_clk),
    .d(_00460_),
    .o(\text_in_r[67] ));
 b15fpn000hn1n04x5 _35310_ (.clk(clknet_leaf_17_clk),
    .d(_00461_),
    .o(\text_in_r[68] ));
 b15fpn000hn1n04x5 _35311_ (.clk(clknet_leaf_18_clk),
    .d(_00462_),
    .o(\text_in_r[69] ));
 b15fpn000hn1n04x5 _35312_ (.clk(clknet_leaf_18_clk),
    .d(_00463_),
    .o(\text_in_r[70] ));
 b15fpn000hn1n04x5 _35313_ (.clk(clknet_leaf_1_clk),
    .d(_00464_),
    .o(\text_in_r[71] ));
 b15fpn000hn1n04x5 _35314_ (.clk(clknet_leaf_15_clk),
    .d(_00465_),
    .o(\text_in_r[72] ));
 b15fpn000hn1n04x5 _35315_ (.clk(clknet_leaf_9_clk),
    .d(_00466_),
    .o(\text_in_r[73] ));
 b15fpn000hn1n04x5 _35316_ (.clk(clknet_leaf_7_clk),
    .d(_00467_),
    .o(\text_in_r[74] ));
 b15fpn000hn1n04x5 _35317_ (.clk(clknet_leaf_8_clk),
    .d(_00468_),
    .o(\text_in_r[75] ));
 b15fpn000hn1n04x5 _35318_ (.clk(clknet_leaf_1_clk),
    .d(_00469_),
    .o(\text_in_r[76] ));
 b15fpn000hn1n04x5 _35319_ (.clk(clknet_leaf_1_clk),
    .d(_00470_),
    .o(\text_in_r[77] ));
 b15fpn000hn1n04x5 _35320_ (.clk(clknet_leaf_1_clk),
    .d(_00471_),
    .o(\text_in_r[78] ));
 b15fpn000hn1n04x5 _35321_ (.clk(clknet_leaf_0_clk),
    .d(_00472_),
    .o(\text_in_r[79] ));
 b15fpn000hn1n04x5 _35322_ (.clk(clknet_leaf_7_clk),
    .d(_00473_),
    .o(\text_in_r[80] ));
 b15fpn000hn1n04x5 _35323_ (.clk(clknet_leaf_9_clk),
    .d(_00474_),
    .o(\text_in_r[81] ));
 b15fpn000hn1n04x5 _35324_ (.clk(clknet_leaf_7_clk),
    .d(_00475_),
    .o(\text_in_r[82] ));
 b15fpn000hn1n04x5 _35325_ (.clk(clknet_leaf_7_clk),
    .d(_00476_),
    .o(\text_in_r[83] ));
 b15fpn000hn1n04x5 _35326_ (.clk(clknet_leaf_4_clk),
    .d(_00477_),
    .o(\text_in_r[84] ));
 b15fpn000hn1n04x5 _35327_ (.clk(clknet_leaf_0_clk),
    .d(_00478_),
    .o(\text_in_r[85] ));
 b15fpn000hn1n04x5 _35328_ (.clk(clknet_leaf_0_clk),
    .d(_00479_),
    .o(\text_in_r[86] ));
 b15fpn000hn1n04x5 _35329_ (.clk(clknet_leaf_4_clk),
    .d(_00480_),
    .o(\text_in_r[87] ));
 b15fpn000hn1n04x5 _35330_ (.clk(clknet_leaf_4_clk),
    .d(_00481_),
    .o(\text_in_r[88] ));
 b15fpn000hn1n04x5 _35331_ (.clk(clknet_leaf_9_clk),
    .d(_00482_),
    .o(\text_in_r[89] ));
 b15fpn000hn1n04x5 _35332_ (.clk(clknet_leaf_4_clk),
    .d(_00483_),
    .o(\text_in_r[90] ));
 b15fpn000hn1n04x5 _35333_ (.clk(clknet_leaf_10_clk),
    .d(_00484_),
    .o(\text_in_r[91] ));
 b15fpn000hn1n04x5 _35334_ (.clk(clknet_leaf_0_clk),
    .d(_00485_),
    .o(\text_in_r[92] ));
 b15fpn000hn1n04x5 _35335_ (.clk(clknet_leaf_0_clk),
    .d(_00486_),
    .o(\text_in_r[93] ));
 b15fpn000hn1n04x5 _35336_ (.clk(clknet_leaf_0_clk),
    .d(_00487_),
    .o(\text_in_r[94] ));
 b15fpn000hn1n04x5 _35337_ (.clk(clknet_leaf_0_clk),
    .d(_00488_),
    .o(\text_in_r[95] ));
 b15fpn000hn1n04x5 _35338_ (.clk(clknet_leaf_8_clk),
    .d(_00489_),
    .o(\text_in_r[96] ));
 b15fpn000hn1n04x5 _35339_ (.clk(clknet_leaf_7_clk),
    .d(_00490_),
    .o(\text_in_r[97] ));
 b15fpn000hn1n04x5 _35340_ (.clk(clknet_leaf_12_clk),
    .d(_00491_),
    .o(\text_in_r[98] ));
 b15fpn000hn1n04x5 _35341_ (.clk(clknet_leaf_12_clk),
    .d(_00492_),
    .o(\text_in_r[99] ));
 b15fpn000hn1n04x5 _35342_ (.clk(clknet_leaf_12_clk),
    .d(_00493_),
    .o(\text_in_r[100] ));
 b15fpn000hn1n04x5 _35343_ (.clk(clknet_leaf_12_clk),
    .d(_00494_),
    .o(\text_in_r[101] ));
 b15fpn000hn1n04x5 _35344_ (.clk(clknet_leaf_14_clk),
    .d(_00495_),
    .o(\text_in_r[102] ));
 b15fpn000hn1n04x5 _35345_ (.clk(clknet_leaf_12_clk),
    .d(_00496_),
    .o(\text_in_r[103] ));
 b15fpn000hn1n04x5 _35346_ (.clk(clknet_leaf_12_clk),
    .d(_00497_),
    .o(\text_in_r[104] ));
 b15fpn000hn1n04x5 _35347_ (.clk(clknet_leaf_12_clk),
    .d(_00498_),
    .o(\text_in_r[105] ));
 b15fpn000hn1n04x5 _35348_ (.clk(clknet_leaf_14_clk),
    .d(_00499_),
    .o(\text_in_r[106] ));
 b15fpn000hn1n04x5 _35349_ (.clk(clknet_leaf_14_clk),
    .d(_00500_),
    .o(\text_in_r[107] ));
 b15fpn000hn1n04x5 _35350_ (.clk(clknet_leaf_14_clk),
    .d(_00501_),
    .o(\text_in_r[108] ));
 b15fpn000hn1n04x5 _35351_ (.clk(clknet_leaf_14_clk),
    .d(_00502_),
    .o(\text_in_r[109] ));
 b15fpn000hn1n04x5 _35352_ (.clk(clknet_leaf_11_clk),
    .d(_00503_),
    .o(\text_in_r[110] ));
 b15fpn000hn1n04x5 _35353_ (.clk(clknet_leaf_14_clk),
    .d(_00504_),
    .o(\text_in_r[111] ));
 b15fpn000hn1n04x5 _35354_ (.clk(clknet_leaf_7_clk),
    .d(_00505_),
    .o(\text_in_r[112] ));
 b15fpn000hn1n04x5 _35355_ (.clk(clknet_leaf_6_clk),
    .d(_00506_),
    .o(\text_in_r[113] ));
 b15fpn000hn1n04x5 _35356_ (.clk(clknet_leaf_7_clk),
    .d(_00507_),
    .o(\text_in_r[114] ));
 b15fpn000hn1n04x5 _35357_ (.clk(clknet_leaf_7_clk),
    .d(_00508_),
    .o(\text_in_r[115] ));
 b15fpn000hn1n04x5 _35358_ (.clk(clknet_leaf_6_clk),
    .d(_00509_),
    .o(\text_in_r[116] ));
 b15fpn000hn1n04x5 _35359_ (.clk(clknet_leaf_9_clk),
    .d(_00510_),
    .o(\text_in_r[117] ));
 b15fpn000hn1n04x5 _35360_ (.clk(clknet_leaf_8_clk),
    .d(_00511_),
    .o(\text_in_r[118] ));
 b15fpn000hn1n04x5 _35361_ (.clk(clknet_leaf_7_clk),
    .d(_00512_),
    .o(\text_in_r[119] ));
 b15fpn000hn1n04x5 _35362_ (.clk(clknet_leaf_13_clk),
    .d(_00513_),
    .o(\text_in_r[120] ));
 b15fpn000hn1n04x5 _35363_ (.clk(clknet_leaf_12_clk),
    .d(_00514_),
    .o(\text_in_r[121] ));
 b15fpn000hn1n04x5 _35364_ (.clk(clknet_leaf_13_clk),
    .d(_00515_),
    .o(\text_in_r[122] ));
 b15fpn000hn1n04x5 _35365_ (.clk(clknet_leaf_12_clk),
    .d(_00516_),
    .o(\text_in_r[123] ));
 b15fpn000hn1n04x5 _35366_ (.clk(clknet_leaf_12_clk),
    .d(_00517_),
    .o(\text_in_r[124] ));
 b15fpn000hn1n04x5 _35367_ (.clk(clknet_leaf_13_clk),
    .d(_00518_),
    .o(\text_in_r[125] ));
 b15fpn000hn1n04x5 _35368_ (.clk(clknet_leaf_13_clk),
    .d(_00519_),
    .o(\text_in_r[126] ));
 b15fpn000hn1n04x5 _35369_ (.clk(clknet_leaf_12_clk),
    .d(_00520_),
    .o(\text_in_r[127] ));
 b15fpn000hn1n04x5 _35370_ (.clk(clknet_leaf_6_clk),
    .d(_00521_),
    .o(\dcnt[0] ));
 b15fpn000hn1n04x5 _35371_ (.clk(clknet_leaf_6_clk),
    .d(_00522_),
    .o(\dcnt[1] ));
 b15fpn000hn1n04x5 _35372_ (.clk(clknet_leaf_6_clk),
    .d(_00523_),
    .o(\dcnt[3] ));
 b15fpn000hn1n04x5 _35373_ (.clk(clknet_leaf_5_clk),
    .d(_00233_),
    .o(net260));
 b15fpn000hn1n04x5 _35374_ (.clk(clknet_leaf_4_clk),
    .d(_00234_),
    .o(net299));
 b15fpn000hn1n04x5 _35375_ (.clk(clknet_leaf_4_clk),
    .d(_00235_),
    .o(net310));
 b15fpn000hn1n04x5 _35376_ (.clk(clknet_leaf_3_clk),
    .d(_00236_),
    .o(net321));
 b15fpn000hn1n04x5 _35377_ (.clk(clknet_leaf_3_clk),
    .d(_00237_),
    .o(net332));
 b15fpn000hn1n04x5 _35378_ (.clk(clknet_leaf_3_clk),
    .d(_00238_),
    .o(net343));
 b15fpn000hn1n04x5 _35379_ (.clk(clknet_leaf_4_clk),
    .d(_00239_),
    .o(net354));
 b15fpn000hn1n04x5 _35380_ (.clk(clknet_leaf_3_clk),
    .d(_00240_),
    .o(net365));
 b15fpn000hn1n04x5 _35381_ (.clk(clknet_leaf_16_clk),
    .d(_00185_),
    .o(net313));
 b15fpn000hn1n04x5 _35382_ (.clk(clknet_leaf_15_clk),
    .d(_00186_),
    .o(net314));
 b15fpn000hn1n04x5 _35383_ (.clk(clknet_leaf_16_clk),
    .d(_00187_),
    .o(net315));
 b15fpn000hn1n04x5 _35384_ (.clk(clknet_leaf_16_clk),
    .d(_00188_),
    .o(net316));
 b15fpn000hn1n04x5 _35385_ (.clk(clknet_leaf_16_clk),
    .d(_00189_),
    .o(net317));
 b15fpn000hn1n04x5 _35386_ (.clk(clknet_leaf_18_clk),
    .d(_00190_),
    .o(net318));
 b15fpn000hn1n04x5 _35387_ (.clk(clknet_leaf_17_clk),
    .d(_00191_),
    .o(net319));
 b15fpn000hn1n04x5 _35388_ (.clk(clknet_leaf_16_clk),
    .d(_00192_),
    .o(net320));
 b15fpn000hn1n04x5 _35389_ (.clk(clknet_leaf_12_clk),
    .d(_00217_),
    .o(net348));
 b15fpn000hn1n04x5 _35390_ (.clk(clknet_leaf_10_clk),
    .d(_00218_),
    .o(net349));
 b15fpn000hn1n04x5 _35391_ (.clk(clknet_leaf_8_clk),
    .d(_00219_),
    .o(net350));
 b15fpn000hn1n04x5 _35392_ (.clk(clknet_leaf_10_clk),
    .d(_00220_),
    .o(net351));
 b15fpn000hn1n04x5 _35393_ (.clk(clknet_leaf_17_clk),
    .d(_00221_),
    .o(net352));
 b15fpn000hn1n04x5 _35394_ (.clk(clknet_leaf_18_clk),
    .d(_00222_),
    .o(net353));
 b15fpn000hn1n04x5 _35395_ (.clk(clknet_leaf_16_clk),
    .d(_00223_),
    .o(net355));
 b15fpn000hn1n04x5 _35396_ (.clk(clknet_leaf_16_clk),
    .d(_00224_),
    .o(net356));
 b15fpn000hn1n04x5 _35397_ (.clk(clknet_leaf_12_clk),
    .d(_00129_),
    .o(net383));
 b15fpn000hn1n04x5 _35398_ (.clk(clknet_leaf_8_clk),
    .d(_00130_),
    .o(net384));
 b15fpn000hn1n04x5 _35399_ (.clk(clknet_leaf_12_clk),
    .d(_00131_),
    .o(net385));
 b15fpn000hn1n04x5 _35400_ (.clk(clknet_leaf_12_clk),
    .d(_00132_),
    .o(net386));
 b15fpn000hn1n04x5 _35401_ (.clk(clknet_leaf_12_clk),
    .d(_00133_),
    .o(net261));
 b15fpn000hn1n04x5 _35402_ (.clk(clknet_leaf_12_clk),
    .d(_00134_),
    .o(net262));
 b15fpn000hn1n04x5 _35403_ (.clk(clknet_leaf_14_clk),
    .d(_00135_),
    .o(net263));
 b15fpn000hn1n04x5 _35404_ (.clk(clknet_leaf_12_clk),
    .d(_00136_),
    .o(net264));
 b15fpn000hn1n04x5 _35405_ (.clk(clknet_leaf_6_clk),
    .d(_00161_),
    .o(net376));
 b15fpn000hn1n04x5 _35406_ (.clk(clknet_leaf_4_clk),
    .d(_00162_),
    .o(net387));
 b15fpn000hn1n04x5 _35407_ (.clk(clknet_leaf_5_clk),
    .d(_00163_),
    .o(net271));
 b15fpn000hn1n04x5 _35408_ (.clk(clknet_leaf_2_clk),
    .d(_00164_),
    .o(net282));
 b15fpn000hn1n04x5 _35409_ (.clk(clknet_leaf_3_clk),
    .d(_00165_),
    .o(net291));
 b15fpn000hn1n04x5 _35410_ (.clk(clknet_leaf_2_clk),
    .d(_00166_),
    .o(net292));
 b15fpn000hn1n04x5 _35411_ (.clk(clknet_leaf_4_clk),
    .d(_00167_),
    .o(net293));
 b15fpn000hn1n04x5 _35412_ (.clk(clknet_leaf_3_clk),
    .d(_00168_),
    .o(net294));
 b15fpn000hn1n04x5 _35413_ (.clk(clknet_leaf_14_clk),
    .d(_00193_),
    .o(net322));
 b15fpn000hn1n04x5 _35414_ (.clk(clknet_leaf_14_clk),
    .d(_00194_),
    .o(net323));
 b15fpn000hn1n04x5 _35415_ (.clk(clknet_leaf_14_clk),
    .d(_00195_),
    .o(net324));
 b15fpn000hn1n04x5 _35416_ (.clk(clknet_leaf_14_clk),
    .d(_00196_),
    .o(net325));
 b15fpn000hn1n04x5 _35417_ (.clk(clknet_leaf_16_clk),
    .d(_00197_),
    .o(net326));
 b15fpn000hn1n04x5 _35418_ (.clk(clknet_leaf_17_clk),
    .d(_00198_),
    .o(net327));
 b15fpn000hn1n04x5 _35419_ (.clk(clknet_leaf_16_clk),
    .d(_00199_),
    .o(net328));
 b15fpn000hn1n04x5 _35420_ (.clk(clknet_leaf_16_clk),
    .d(_00200_),
    .o(net329));
 b15fpn000hn1n04x5 _35421_ (.clk(clknet_leaf_10_clk),
    .d(_00225_),
    .o(net357));
 b15fpn000hn1n04x5 _35422_ (.clk(clknet_leaf_9_clk),
    .d(_00226_),
    .o(net358));
 b15fpn000hn1n04x5 _35423_ (.clk(clknet_leaf_7_clk),
    .d(_00227_),
    .o(net359));
 b15fpn000hn1n04x5 _35424_ (.clk(clknet_leaf_8_clk),
    .d(_00228_),
    .o(net360));
 b15fpn000hn1n04x5 _35425_ (.clk(clknet_leaf_15_clk),
    .d(_00229_),
    .o(net361));
 b15fpn000hn1n04x5 _35426_ (.clk(clknet_leaf_1_clk),
    .d(_00230_),
    .o(net362));
 b15fpn000hn1n04x5 _35427_ (.clk(clknet_leaf_16_clk),
    .d(_00231_),
    .o(net363));
 b15fpn000hn1n04x5 _35428_ (.clk(clknet_leaf_1_clk),
    .d(_00232_),
    .o(net364));
 b15fpn000hn1n04x5 _35429_ (.clk(clknet_leaf_12_clk),
    .d(_00137_),
    .o(net265));
 b15fpn000hn1n04x5 _35430_ (.clk(clknet_leaf_12_clk),
    .d(_00138_),
    .o(net266));
 b15fpn000hn1n04x5 _35431_ (.clk(clknet_leaf_12_clk),
    .d(_00139_),
    .o(net267));
 b15fpn000hn1n04x5 _35432_ (.clk(clknet_leaf_14_clk),
    .d(_00140_),
    .o(net268));
 b15fpn000hn1n04x5 _35433_ (.clk(clknet_leaf_14_clk),
    .d(_00141_),
    .o(net269));
 b15fpn000hn1n04x5 _35434_ (.clk(clknet_leaf_14_clk),
    .d(_00142_),
    .o(net270));
 b15fpn000hn1n04x5 _35435_ (.clk(clknet_leaf_12_clk),
    .d(_00143_),
    .o(net272));
 b15fpn000hn1n04x5 _35436_ (.clk(clknet_leaf_14_clk),
    .d(_00144_),
    .o(net273));
 b15fpn000hn1n04x5 _35437_ (.clk(clknet_leaf_2_clk),
    .d(_00169_),
    .o(net295));
 b15fpn000hn1n04x5 _35438_ (.clk(clknet_leaf_2_clk),
    .d(_00170_),
    .o(net296));
 b15fpn000hn1n04x5 _35439_ (.clk(clknet_leaf_2_clk),
    .d(_00171_),
    .o(net297));
 b15fpn000hn1n04x5 _35440_ (.clk(clknet_leaf_2_clk),
    .d(_00172_),
    .o(net298));
 b15fpn000hn1n04x5 _35441_ (.clk(clknet_leaf_2_clk),
    .d(_00173_),
    .o(net300));
 b15fpn000hn1n04x5 _35442_ (.clk(clknet_leaf_7_clk),
    .d(_00174_),
    .o(net301));
 b15fpn000hn1n04x5 _35443_ (.clk(clknet_leaf_7_clk),
    .d(_00175_),
    .o(net302));
 b15fpn000hn1n04x5 _35444_ (.clk(clknet_leaf_3_clk),
    .d(_00176_),
    .o(net303));
 b15fpn000hn1n04x5 _35445_ (.clk(clknet_leaf_15_clk),
    .d(_00201_),
    .o(net330));
 b15fpn000hn1n04x5 _35446_ (.clk(clknet_leaf_15_clk),
    .d(_00202_),
    .o(net331));
 b15fpn000hn1n04x5 _35447_ (.clk(clknet_leaf_15_clk),
    .d(_00203_),
    .o(net333));
 b15fpn000hn1n04x5 _35448_ (.clk(clknet_leaf_16_clk),
    .d(_00204_),
    .o(net334));
 b15fpn000hn1n04x5 _35449_ (.clk(clknet_leaf_18_clk),
    .d(_00205_),
    .o(net335));
 b15fpn000hn1n04x5 _35450_ (.clk(clknet_leaf_17_clk),
    .d(_00206_),
    .o(net336));
 b15fpn000hn1n04x5 _35451_ (.clk(clknet_leaf_18_clk),
    .d(_00207_),
    .o(net337));
 b15fpn000hn1n04x5 _35452_ (.clk(clknet_leaf_16_clk),
    .d(_00208_),
    .o(net338));
 b15fpn000hn1n04x5 _35453_ (.clk(clknet_leaf_7_clk),
    .d(_00241_),
    .o(net366));
 b15fpn000hn1n04x5 _35454_ (.clk(clknet_leaf_9_clk),
    .d(_00242_),
    .o(net367));
 b15fpn000hn1n04x5 _35455_ (.clk(clknet_leaf_7_clk),
    .d(_00243_),
    .o(net368));
 b15fpn000hn1n04x5 _35456_ (.clk(clknet_leaf_8_clk),
    .d(_00244_),
    .o(net369));
 b15fpn000hn1n04x5 _35457_ (.clk(clknet_leaf_15_clk),
    .d(_00245_),
    .o(net370));
 b15fpn000hn1n04x5 _35458_ (.clk(clknet_leaf_0_clk),
    .d(_00246_),
    .o(net371));
 b15fpn000hn1n04x5 _35459_ (.clk(clknet_leaf_0_clk),
    .d(_00247_),
    .o(net372));
 b15fpn000hn1n04x5 _35460_ (.clk(clknet_leaf_7_clk),
    .d(_00248_),
    .o(net373));
 b15fpn000hn1n04x5 _35461_ (.clk(clknet_leaf_6_clk),
    .d(_00145_),
    .o(net274));
 b15fpn000hn1n04x5 _35462_ (.clk(clknet_leaf_6_clk),
    .d(_00146_),
    .o(net275));
 b15fpn000hn1n04x5 _35463_ (.clk(clknet_leaf_7_clk),
    .d(_00147_),
    .o(net276));
 b15fpn000hn1n04x5 _35464_ (.clk(clknet_leaf_9_clk),
    .d(_00148_),
    .o(net277));
 b15fpn000hn1n04x5 _35465_ (.clk(clknet_leaf_7_clk),
    .d(_00149_),
    .o(net278));
 b15fpn000hn1n04x5 _35466_ (.clk(clknet_leaf_7_clk),
    .d(_00150_),
    .o(net279));
 b15fpn000hn1n04x5 _35467_ (.clk(clknet_leaf_7_clk),
    .d(_00151_),
    .o(net280));
 b15fpn000hn1n04x5 _35468_ (.clk(clknet_leaf_7_clk),
    .d(_00152_),
    .o(net281));
 b15fpn000hn1n04x5 _35469_ (.clk(clknet_leaf_4_clk),
    .d(_00177_),
    .o(net304));
 b15fpn000hn1n04x5 _35470_ (.clk(clknet_leaf_3_clk),
    .d(_00178_),
    .o(net305));
 b15fpn000hn1n04x5 _35471_ (.clk(clknet_leaf_4_clk),
    .d(_00179_),
    .o(net306));
 b15fpn000hn1n04x5 _35472_ (.clk(clknet_leaf_2_clk),
    .d(_00180_),
    .o(net307));
 b15fpn000hn1n04x5 _35473_ (.clk(clknet_leaf_3_clk),
    .d(_00181_),
    .o(net308));
 b15fpn000hn1n04x5 _35474_ (.clk(clknet_leaf_2_clk),
    .d(_00182_),
    .o(net309));
 b15fpn000hn1n04x5 _35475_ (.clk(clknet_leaf_4_clk),
    .d(_00183_),
    .o(net311));
 b15fpn000hn1n04x5 _35476_ (.clk(clknet_leaf_3_clk),
    .d(_00184_),
    .o(net312));
 b15fpn000hn1n04x5 _35477_ (.clk(clknet_leaf_15_clk),
    .d(_00209_),
    .o(net339));
 b15fpn000hn1n04x5 _35478_ (.clk(clknet_leaf_15_clk),
    .d(_00210_),
    .o(net340));
 b15fpn000hn1n04x5 _35479_ (.clk(clknet_leaf_16_clk),
    .d(_00211_),
    .o(net341));
 b15fpn000hn1n04x5 _35480_ (.clk(clknet_leaf_16_clk),
    .d(_00212_),
    .o(net342));
 b15fpn000hn1n04x5 _35481_ (.clk(clknet_leaf_17_clk),
    .d(_00213_),
    .o(net344));
 b15fpn000hn1n04x5 _35482_ (.clk(clknet_leaf_17_clk),
    .d(_00214_),
    .o(net345));
 b15fpn000hn1n04x5 _35483_ (.clk(clknet_leaf_16_clk),
    .d(_00215_),
    .o(net346));
 b15fpn000hn1n04x5 _35484_ (.clk(clknet_leaf_16_clk),
    .d(_00216_),
    .o(net347));
 b15fpn000hn1n04x5 _35485_ (.clk(clknet_leaf_9_clk),
    .d(_00249_),
    .o(net374));
 b15fpn000hn1n04x5 _35486_ (.clk(clknet_leaf_8_clk),
    .d(_00250_),
    .o(net375));
 b15fpn000hn1n04x5 _35487_ (.clk(clknet_leaf_9_clk),
    .d(_00251_),
    .o(net377));
 b15fpn000hn1n04x5 _35488_ (.clk(clknet_leaf_7_clk),
    .d(_00252_),
    .o(net378));
 b15fpn000hn1n04x5 _35489_ (.clk(clknet_leaf_0_clk),
    .d(_00253_),
    .o(net379));
 b15fpn000hn1n04x5 _35490_ (.clk(clknet_leaf_0_clk),
    .d(_00254_),
    .o(net380));
 b15fpn000hn1n04x5 _35491_ (.clk(clknet_leaf_0_clk),
    .d(_00255_),
    .o(net381));
 b15fpn000hn1n04x5 _35492_ (.clk(clknet_leaf_15_clk),
    .d(_00256_),
    .o(net382));
 b15fpn000hn1n04x5 _35493_ (.clk(clknet_leaf_13_clk),
    .d(_00153_),
    .o(net283));
 b15fpn000hn1n04x5 _35494_ (.clk(clknet_leaf_12_clk),
    .d(_00154_),
    .o(net284));
 b15fpn000hn1n04x5 _35495_ (.clk(clknet_leaf_13_clk),
    .d(_00155_),
    .o(net285));
 b15fpn000hn1n04x5 _35496_ (.clk(clknet_leaf_12_clk),
    .d(_00156_),
    .o(net286));
 b15fpn000hn1n04x5 _35497_ (.clk(clknet_leaf_12_clk),
    .d(_00157_),
    .o(net287));
 b15fpn000hn1n04x5 _35498_ (.clk(clknet_leaf_13_clk),
    .d(_00158_),
    .o(net288));
 b15fpn000hn1n04x5 _35499_ (.clk(clknet_leaf_13_clk),
    .d(_00159_),
    .o(net289));
 b15fpn000hn1n04x5 _35500_ (.clk(clknet_leaf_11_clk),
    .d(_00160_),
    .o(net290));
 b15fpn000hn1n04x5 _35501_ (.clk(clknet_leaf_11_clk),
    .d(_00001_),
    .o(\us00.a[0] ));
 b15fpn000hn1n04x5 _35502_ (.clk(clknet_leaf_11_clk),
    .d(_00002_),
    .o(\us00.a[1] ));
 b15fpn000hn1n04x5 _35503_ (.clk(clknet_leaf_12_clk),
    .d(_00003_),
    .o(\us00.a[2] ));
 b15fpn000hn1n04x5 _35504_ (.clk(clknet_leaf_11_clk),
    .d(_00004_),
    .o(\us00.a[3] ));
 b15fpn000hn1n04x5 _35505_ (.clk(clknet_leaf_11_clk),
    .d(_00005_),
    .o(\us00.a[4] ));
 b15fpn000hn1n04x5 _35506_ (.clk(clknet_leaf_11_clk),
    .d(_00006_),
    .o(\us00.a[5] ));
 b15fpn000hn1n04x5 _35507_ (.clk(clknet_leaf_11_clk),
    .d(_00007_),
    .o(\us00.a[6] ));
 b15fpn000hn1n04x5 _35508_ (.clk(clknet_leaf_11_clk),
    .d(_00008_),
    .o(\us00.a[7] ));
 b15fpn000hn1n04x5 _35509_ (.clk(clknet_leaf_6_clk),
    .d(_00033_),
    .o(\us10.a[0] ));
 b15fpn000hn1n04x5 _35510_ (.clk(clknet_leaf_6_clk),
    .d(_00034_),
    .o(\us10.a[1] ));
 b15fpn000hn1n04x5 _35511_ (.clk(clknet_leaf_10_clk),
    .d(_00035_),
    .o(\us10.a[2] ));
 b15fpn000hn1n04x5 _35512_ (.clk(clknet_leaf_9_clk),
    .d(_00036_),
    .o(\us10.a[3] ));
 b15fpn000hn1n04x5 _35513_ (.clk(clknet_leaf_9_clk),
    .d(_00037_),
    .o(\us10.a[4] ));
 b15fpn000hn1n04x5 _35514_ (.clk(clknet_leaf_5_clk),
    .d(_00038_),
    .o(\us10.a[5] ));
 b15fpn000hn1n04x5 _35515_ (.clk(clknet_leaf_4_clk),
    .d(_00039_),
    .o(\us10.a[6] ));
 b15fpn000hn1n04x5 _35516_ (.clk(clknet_leaf_5_clk),
    .d(_00040_),
    .o(\us10.a[7] ));
 b15fpn000hn1n04x5 _35517_ (.clk(clknet_leaf_11_clk),
    .d(_00065_),
    .o(\us20.a[0] ));
 b15fpn000hn1n04x5 _35518_ (.clk(clknet_leaf_11_clk),
    .d(_00066_),
    .o(\us20.a[1] ));
 b15fpn000hn1n04x5 _35519_ (.clk(clknet_leaf_11_clk),
    .d(_00067_),
    .o(\us20.a[2] ));
 b15fpn000hn1n04x5 _35520_ (.clk(clknet_leaf_14_clk),
    .d(_00068_),
    .o(\us20.a[3] ));
 b15fpn000hn1n04x5 _35521_ (.clk(clknet_leaf_14_clk),
    .d(_00069_),
    .o(\us20.a[4] ));
 b15fpn000hn1n04x5 _35522_ (.clk(clknet_leaf_14_clk),
    .d(_00070_),
    .o(\us20.a[5] ));
 b15fpn000hn1n04x5 _35523_ (.clk(clknet_leaf_15_clk),
    .d(_00071_),
    .o(\us20.a[6] ));
 b15fpn000hn1n04x5 _35524_ (.clk(clknet_leaf_14_clk),
    .d(_00072_),
    .o(\us20.a[7] ));
 b15fpn000hn1n04x5 _35525_ (.clk(clknet_leaf_11_clk),
    .d(_00097_),
    .o(\us30.a[0] ));
 b15fpn000hn1n04x5 _35526_ (.clk(clknet_leaf_11_clk),
    .d(_00098_),
    .o(\us30.a[1] ));
 b15fpn000hn1n04x5 _35527_ (.clk(clknet_leaf_11_clk),
    .d(_00099_),
    .o(\us30.a[2] ));
 b15fpn000hn1n04x5 _35528_ (.clk(clknet_leaf_11_clk),
    .d(_00100_),
    .o(\us30.a[3] ));
 b15fpn000hn1n04x5 _35529_ (.clk(clknet_leaf_10_clk),
    .d(_00101_),
    .o(\us30.a[4] ));
 b15fpn000hn1n04x5 _35530_ (.clk(clknet_leaf_10_clk),
    .d(_00102_),
    .o(\us30.a[5] ));
 b15fpn000hn1n04x5 _35531_ (.clk(clknet_leaf_15_clk),
    .d(_00103_),
    .o(\us30.a[6] ));
 b15fpn000hn1n04x5 _35532_ (.clk(clknet_leaf_10_clk),
    .d(_00104_),
    .o(\us30.a[7] ));
 b15fpn000hn1n04x5 _35533_ (.clk(clknet_leaf_5_clk),
    .d(_00009_),
    .o(\us01.a[0] ));
 b15fpn000hn1n04x5 _35534_ (.clk(clknet_leaf_9_clk),
    .d(_00010_),
    .o(\us01.a[1] ));
 b15fpn000hn1n04x5 _35535_ (.clk(clknet_leaf_5_clk),
    .d(_00011_),
    .o(\us01.a[2] ));
 b15fpn000hn1n04x5 _35536_ (.clk(clknet_leaf_10_clk),
    .d(_00012_),
    .o(\us01.a[3] ));
 b15fpn000hn1n04x5 _35537_ (.clk(clknet_leaf_1_clk),
    .d(_00013_),
    .o(\us01.a[4] ));
 b15fpn000hn1n04x5 _35538_ (.clk(clknet_leaf_0_clk),
    .d(_00014_),
    .o(\us01.a[5] ));
 b15fpn000hn1n04x5 _35539_ (.clk(clknet_leaf_0_clk),
    .d(_00015_),
    .o(\us01.a[6] ));
 b15fpn000hn1n04x5 _35540_ (.clk(clknet_leaf_1_clk),
    .d(_00016_),
    .o(\us01.a[7] ));
 b15fpn000hn1n04x5 _35541_ (.clk(clknet_leaf_6_clk),
    .d(_00041_),
    .o(\us11.a[0] ));
 b15fpn000hn1n04x5 _35542_ (.clk(clknet_leaf_6_clk),
    .d(_00042_),
    .o(\us11.a[1] ));
 b15fpn000hn1n04x5 _35543_ (.clk(clknet_leaf_6_clk),
    .d(_00043_),
    .o(\us11.a[2] ));
 b15fpn000hn1n04x5 _35544_ (.clk(clknet_leaf_6_clk),
    .d(_00044_),
    .o(\us11.a[3] ));
 b15fpn000hn1n04x5 _35545_ (.clk(clknet_leaf_1_clk),
    .d(_00045_),
    .o(\us11.a[4] ));
 b15fpn000hn1n04x5 _35546_ (.clk(clknet_leaf_6_clk),
    .d(net389),
    .o(\us11.a[5] ));
 b15fpn000hn1n04x5 _35547_ (.clk(clknet_leaf_6_clk),
    .d(net388),
    .o(\us11.a[6] ));
 b15fpn000hn1n04x5 _35548_ (.clk(clknet_leaf_6_clk),
    .d(_00048_),
    .o(\us11.a[7] ));
 b15fpn000hn1n04x5 _35549_ (.clk(clknet_leaf_5_clk),
    .d(_00073_),
    .o(\us21.a[0] ));
 b15fpn000hn1n04x5 _35550_ (.clk(clknet_leaf_10_clk),
    .d(_00074_),
    .o(\us21.a[1] ));
 b15fpn000hn1n04x5 _35551_ (.clk(clknet_leaf_10_clk),
    .d(_00075_),
    .o(\us21.a[2] ));
 b15fpn000hn1n04x5 _35552_ (.clk(clknet_leaf_10_clk),
    .d(_00076_),
    .o(\us21.a[3] ));
 b15fpn000hn1n04x5 _35553_ (.clk(clknet_leaf_1_clk),
    .d(_00077_),
    .o(\us21.a[4] ));
 b15fpn000hn1n04x5 _35554_ (.clk(clknet_leaf_1_clk),
    .d(_00078_),
    .o(\us21.a[5] ));
 b15fpn000hn1n04x5 _35555_ (.clk(clknet_leaf_1_clk),
    .d(_00079_),
    .o(\us21.a[6] ));
 b15fpn000hn1n04x5 _35556_ (.clk(clknet_leaf_0_clk),
    .d(_00080_),
    .o(\us21.a[7] ));
 b15fpn000hn1n04x5 _35557_ (.clk(clknet_leaf_1_clk),
    .d(_00105_),
    .o(\us31.a[0] ));
 b15fpn000hn1n04x5 _35558_ (.clk(clknet_leaf_5_clk),
    .d(_00106_),
    .o(\us31.a[1] ));
 b15fpn000hn1n04x5 _35559_ (.clk(clknet_leaf_1_clk),
    .d(_00107_),
    .o(\us31.a[2] ));
 b15fpn000hn1n04x5 _35560_ (.clk(clknet_leaf_1_clk),
    .d(_00108_),
    .o(\us31.a[3] ));
 b15fpn000hn1n04x5 _35561_ (.clk(clknet_leaf_1_clk),
    .d(_00109_),
    .o(\us31.a[4] ));
 b15fpn000hn1n04x5 _35562_ (.clk(clknet_leaf_18_clk),
    .d(_00110_),
    .o(\us31.a[5] ));
 b15fpn000hn1n04x5 _35563_ (.clk(clknet_leaf_18_clk),
    .d(_00111_),
    .o(\us31.a[6] ));
 b15fpn000hn1n04x5 _35564_ (.clk(clknet_leaf_0_clk),
    .d(_00112_),
    .o(\us31.a[7] ));
 b15fpn000hn1n04x5 _35565_ (.clk(clknet_leaf_17_clk),
    .d(_00017_),
    .o(\us02.a[0] ));
 b15fpn000hn1n04x5 _35566_ (.clk(clknet_leaf_18_clk),
    .d(_00018_),
    .o(\us02.a[1] ));
 b15fpn000hn1n04x5 _35567_ (.clk(clknet_leaf_17_clk),
    .d(_00019_),
    .o(\us02.a[2] ));
 b15fpn000hn1n04x5 _35568_ (.clk(clknet_leaf_18_clk),
    .d(_00020_),
    .o(\us02.a[3] ));
 b15fpn000hn1n04x5 _35569_ (.clk(clknet_leaf_17_clk),
    .d(_00021_),
    .o(\us02.a[4] ));
 b15fpn000hn1n04x5 _35570_ (.clk(clknet_leaf_17_clk),
    .d(_00022_),
    .o(\us02.a[5] ));
 b15fpn000hn1n04x5 _35571_ (.clk(clknet_leaf_18_clk),
    .d(_00023_),
    .o(\us02.a[6] ));
 b15fpn000hn1n04x5 _35572_ (.clk(clknet_leaf_17_clk),
    .d(_00024_),
    .o(\us02.a[7] ));
 b15fpn000hn1n04x5 _35573_ (.clk(clknet_leaf_0_clk),
    .d(_00049_),
    .o(\us12.a[0] ));
 b15fpn000hn1n04x5 _35574_ (.clk(clknet_leaf_1_clk),
    .d(_00050_),
    .o(\us12.a[1] ));
 b15fpn000hn1n04x5 _35575_ (.clk(clknet_leaf_1_clk),
    .d(_00051_),
    .o(\us12.a[2] ));
 b15fpn000hn1n04x5 _35576_ (.clk(clknet_leaf_1_clk),
    .d(_00052_),
    .o(\us12.a[3] ));
 b15fpn000hn1n04x5 _35577_ (.clk(clknet_leaf_0_clk),
    .d(_00053_),
    .o(\us12.a[4] ));
 b15fpn000hn1n04x5 _35578_ (.clk(clknet_leaf_0_clk),
    .d(_00054_),
    .o(\us12.a[5] ));
 b15fpn000hn1n04x5 _35579_ (.clk(clknet_leaf_0_clk),
    .d(_00055_),
    .o(\us12.a[6] ));
 b15fpn000hn1n04x5 _35580_ (.clk(clknet_leaf_0_clk),
    .d(_00056_),
    .o(\us12.a[7] ));
 b15fpn000hn1n04x5 _35581_ (.clk(clknet_leaf_14_clk),
    .d(_00081_),
    .o(\us22.a[0] ));
 b15fpn000hn1n04x5 _35582_ (.clk(clknet_leaf_14_clk),
    .d(_00082_),
    .o(\us22.a[1] ));
 b15fpn000hn1n04x5 _35583_ (.clk(clknet_leaf_14_clk),
    .d(_00083_),
    .o(\us22.a[2] ));
 b15fpn000hn1n04x5 _35584_ (.clk(clknet_leaf_14_clk),
    .d(_00084_),
    .o(\us22.a[3] ));
 b15fpn000hn1n04x5 _35585_ (.clk(clknet_leaf_14_clk),
    .d(_00085_),
    .o(\us22.a[4] ));
 b15fpn000hn1n04x5 _35586_ (.clk(clknet_leaf_14_clk),
    .d(_00086_),
    .o(\us22.a[5] ));
 b15fpn000hn1n04x5 _35587_ (.clk(clknet_leaf_14_clk),
    .d(_00087_),
    .o(\us22.a[6] ));
 b15fpn000hn1n04x5 _35588_ (.clk(clknet_leaf_14_clk),
    .d(_00088_),
    .o(\us22.a[7] ));
 b15fpn000hn1n04x5 _35589_ (.clk(clknet_leaf_2_clk),
    .d(_00113_),
    .o(\us32.a[0] ));
 b15fpn000hn1n04x5 _35590_ (.clk(clknet_leaf_2_clk),
    .d(_00114_),
    .o(\us32.a[1] ));
 b15fpn000hn1n04x5 _35591_ (.clk(clknet_leaf_2_clk),
    .d(_00115_),
    .o(\us32.a[2] ));
 b15fpn000hn1n04x5 _35592_ (.clk(clknet_leaf_2_clk),
    .d(_00116_),
    .o(\us32.a[3] ));
 b15fpn000hn1n04x5 _35593_ (.clk(clknet_leaf_2_clk),
    .d(_00117_),
    .o(\us32.a[4] ));
 b15fpn000hn1n04x5 _35594_ (.clk(clknet_leaf_2_clk),
    .d(_00118_),
    .o(\us32.a[5] ));
 b15fpn000hn1n04x5 _35595_ (.clk(clknet_leaf_2_clk),
    .d(net390),
    .o(\us32.a[6] ));
 b15fpn000hn1n04x5 _35596_ (.clk(clknet_leaf_2_clk),
    .d(_00120_),
    .o(\us32.a[7] ));
 b15fpn000hn1n04x5 _35597_ (.clk(clknet_leaf_3_clk),
    .d(_00025_),
    .o(\us03.a[0] ));
 b15fpn000hn1n04x5 _35598_ (.clk(clknet_leaf_3_clk),
    .d(_00026_),
    .o(\us03.a[1] ));
 b15fpn000hn1n04x5 _35599_ (.clk(clknet_leaf_3_clk),
    .d(_00027_),
    .o(\us03.a[2] ));
 b15fpn000hn1n04x5 _35600_ (.clk(clknet_leaf_3_clk),
    .d(_00028_),
    .o(\us03.a[3] ));
 b15fpn000hn1n04x5 _35601_ (.clk(clknet_leaf_3_clk),
    .d(_00029_),
    .o(\us03.a[4] ));
 b15fpn000hn1n04x5 _35602_ (.clk(clknet_leaf_3_clk),
    .d(_00030_),
    .o(\us03.a[5] ));
 b15fpn000hn1n04x5 _35603_ (.clk(clknet_leaf_3_clk),
    .d(_00031_),
    .o(\us03.a[6] ));
 b15fpn000hn1n04x5 _35604_ (.clk(clknet_leaf_3_clk),
    .d(_00032_),
    .o(\us03.a[7] ));
 b15fpn000hn1n04x5 _35605_ (.clk(clknet_leaf_0_clk),
    .d(_00057_),
    .o(\us13.a[0] ));
 b15fpn000hn1n04x5 _35606_ (.clk(clknet_leaf_0_clk),
    .d(_00058_),
    .o(\us13.a[1] ));
 b15fpn000hn1n04x5 _35607_ (.clk(clknet_leaf_0_clk),
    .d(_00059_),
    .o(\us13.a[2] ));
 b15fpn000hn1n04x5 _35608_ (.clk(clknet_leaf_0_clk),
    .d(_00060_),
    .o(\us13.a[3] ));
 b15fpn000hn1n04x5 _35609_ (.clk(clknet_leaf_18_clk),
    .d(_00061_),
    .o(\us13.a[4] ));
 b15fpn000hn1n04x5 _35610_ (.clk(clknet_leaf_0_clk),
    .d(_00062_),
    .o(\us13.a[5] ));
 b15fpn000hn1n04x5 _35611_ (.clk(clknet_leaf_18_clk),
    .d(_00063_),
    .o(\us13.a[6] ));
 b15fpn000hn1n04x5 _35612_ (.clk(clknet_leaf_0_clk),
    .d(_00064_),
    .o(\us13.a[7] ));
 b15fpn000hn1n04x5 _35613_ (.clk(clknet_leaf_2_clk),
    .d(_00089_),
    .o(\us23.a[0] ));
 b15fpn000hn1n04x5 _35614_ (.clk(clknet_leaf_2_clk),
    .d(_00090_),
    .o(\us23.a[1] ));
 b15fpn000hn1n04x5 _35615_ (.clk(clknet_leaf_2_clk),
    .d(_00091_),
    .o(\us23.a[2] ));
 b15fpn000hn1n04x5 _35616_ (.clk(clknet_leaf_2_clk),
    .d(_00092_),
    .o(\us23.a[3] ));
 b15fpn000hn1n04x5 _35617_ (.clk(clknet_leaf_2_clk),
    .d(_00093_),
    .o(\us23.a[4] ));
 b15fpn000hn1n04x5 _35618_ (.clk(clknet_leaf_2_clk),
    .d(_00094_),
    .o(\us23.a[5] ));
 b15fpn000hn1n04x5 _35619_ (.clk(clknet_leaf_2_clk),
    .d(_00095_),
    .o(\us23.a[6] ));
 b15fpn000hn1n04x5 _35620_ (.clk(clknet_leaf_2_clk),
    .d(_00096_),
    .o(\us23.a[7] ));
 b15fpn000hn1n04x5 _35621_ (.clk(clknet_leaf_6_clk),
    .d(_00121_),
    .o(\us33.a[0] ));
 b15fpn000hn1n04x5 _35622_ (.clk(clknet_leaf_6_clk),
    .d(_00122_),
    .o(\us33.a[1] ));
 b15fpn000hn1n04x5 _35623_ (.clk(clknet_leaf_6_clk),
    .d(_00123_),
    .o(\us33.a[2] ));
 b15fpn000hn1n04x5 _35624_ (.clk(clknet_leaf_9_clk),
    .d(_00124_),
    .o(\us33.a[3] ));
 b15fpn000hn1n04x5 _35625_ (.clk(clknet_leaf_6_clk),
    .d(_00125_),
    .o(\us33.a[4] ));
 b15fpn000hn1n04x5 _35626_ (.clk(clknet_leaf_6_clk),
    .d(_00126_),
    .o(\us33.a[5] ));
 b15fpn000hn1n04x5 _35627_ (.clk(clknet_leaf_6_clk),
    .d(_00127_),
    .o(\us33.a[6] ));
 b15fpn000hn1n04x5 _35628_ (.clk(clknet_leaf_6_clk),
    .d(_00128_),
    .o(\us33.a[7] ));
 b15fpn000hn1n04x5 _35629_ (.clk(clknet_leaf_1_clk),
    .d(net940),
    .o(ld_r));
 b15fpn000hn1n04x5 _35630_ (.clk(clknet_leaf_6_clk),
    .d(_00000_),
    .o(net259));
 b15fpn000hn1n04x5 _35631_ (.clk(clknet_leaf_6_clk),
    .d(_00524_),
    .o(\dcnt[2] ));
 b15fpn000hn1n04x5 _35632_ (.clk(clknet_leaf_8_clk),
    .d(_00525_),
    .o(\u0.r0.rcnt[0] ));
 b15fpn000hn1n04x5 _35633_ (.clk(clknet_leaf_8_clk),
    .d(_00526_),
    .o(\u0.r0.rcnt[1] ));
 b15fpn000hn1n04x5 _35634_ (.clk(clknet_leaf_8_clk),
    .d(_00527_),
    .o(\u0.r0.rcnt[2] ));
 b15fpn000hn1n04x5 _35635_ (.clk(clknet_leaf_9_clk),
    .d(_00528_),
    .o(\u0.r0.rcnt[3] ));
 b15fpn000hn1n04x5 _35636_ (.clk(clknet_leaf_12_clk),
    .d(_00257_),
    .o(\u0.w[0][0] ));
 b15fpn000hn1n04x5 _35637_ (.clk(clknet_leaf_5_clk),
    .d(_00268_),
    .o(\u0.w[0][1] ));
 b15fpn000hn1n04x5 _35638_ (.clk(clknet_leaf_11_clk),
    .d(_00279_),
    .o(\u0.w[0][2] ));
 b15fpn000hn1n04x5 _35639_ (.clk(clknet_leaf_8_clk),
    .d(_00282_),
    .o(\u0.w[0][3] ));
 b15fpn000hn1n04x5 _35640_ (.clk(clknet_leaf_10_clk),
    .d(_00283_),
    .o(\u0.w[0][4] ));
 b15fpn000hn1n04x5 _35641_ (.clk(clknet_leaf_10_clk),
    .d(_00284_),
    .o(\u0.w[0][5] ));
 b15fpn000hn1n04x5 _35642_ (.clk(clknet_leaf_15_clk),
    .d(_00285_),
    .o(\u0.w[0][6] ));
 b15fpn000hn1n04x5 _35643_ (.clk(clknet_leaf_1_clk),
    .d(_00286_),
    .o(\u0.w[0][7] ));
 b15fpn000hn1n04x5 _35644_ (.clk(clknet_leaf_8_clk),
    .d(_00287_),
    .o(\u0.w[0][8] ));
 b15fpn000hn1n04x5 _35645_ (.clk(clknet_leaf_9_clk),
    .d(_00288_),
    .o(\u0.w[0][9] ));
 b15fpn000hn1n04x5 _35646_ (.clk(clknet_leaf_8_clk),
    .d(_00258_),
    .o(\u0.w[0][10] ));
 b15fpn000hn1n04x5 _35647_ (.clk(clknet_leaf_10_clk),
    .d(_00259_),
    .o(\u0.w[0][11] ));
 b15fpn000hn1n04x5 _35648_ (.clk(clknet_leaf_10_clk),
    .d(_00260_),
    .o(\u0.w[0][12] ));
 b15fpn000hn1n04x5 _35649_ (.clk(clknet_leaf_15_clk),
    .d(_00261_),
    .o(\u0.w[0][13] ));
 b15fpn000hn1n04x5 _35650_ (.clk(clknet_leaf_11_clk),
    .d(_00262_),
    .o(\u0.w[0][14] ));
 b15fpn000hn1n04x5 _35651_ (.clk(clknet_leaf_11_clk),
    .d(_00263_),
    .o(\u0.w[0][15] ));
 b15fpn000hn1n04x5 _35652_ (.clk(clknet_leaf_6_clk),
    .d(_00264_),
    .o(\u0.w[0][16] ));
 b15fpn000hn1n04x5 _35653_ (.clk(clknet_leaf_6_clk),
    .d(_00265_),
    .o(\u0.w[0][17] ));
 b15fpn000hn1n04x5 _35654_ (.clk(clknet_leaf_6_clk),
    .d(_00266_),
    .o(\u0.w[0][18] ));
 b15fpn000hn1n04x5 _35655_ (.clk(clknet_leaf_9_clk),
    .d(_00267_),
    .o(\u0.w[0][19] ));
 b15fpn000hn1n04x5 _35656_ (.clk(clknet_leaf_10_clk),
    .d(_00269_),
    .o(\u0.w[0][20] ));
 b15fpn000hn1n04x5 _35657_ (.clk(clknet_leaf_9_clk),
    .d(_00270_),
    .o(\u0.w[0][21] ));
 b15fpn000hn1n04x5 _35658_ (.clk(clknet_leaf_9_clk),
    .d(_00271_),
    .o(\u0.w[0][22] ));
 b15fpn000hn1n04x5 _35659_ (.clk(clknet_leaf_9_clk),
    .d(_00272_),
    .o(\u0.w[0][23] ));
 b15fpn000hn1n04x5 _35660_ (.clk(clknet_leaf_9_clk),
    .d(_00273_),
    .o(\u0.w[0][24] ));
 b15fpn000hn1n04x5 _35661_ (.clk(clknet_leaf_8_clk),
    .d(_00274_),
    .o(\u0.w[0][25] ));
 b15fpn000hn1n04x5 _35662_ (.clk(clknet_leaf_8_clk),
    .d(_00275_),
    .o(\u0.w[0][26] ));
 b15fpn000hn1n04x5 _35663_ (.clk(clknet_leaf_11_clk),
    .d(_00276_),
    .o(\u0.w[0][27] ));
 b15fpn000hn1n04x5 _35664_ (.clk(clknet_leaf_11_clk),
    .d(_00277_),
    .o(\u0.w[0][28] ));
 b15fpn000hn1n04x5 _35665_ (.clk(clknet_leaf_11_clk),
    .d(_00278_),
    .o(\u0.w[0][29] ));
 b15fpn000hn1n04x5 _35666_ (.clk(clknet_leaf_11_clk),
    .d(_00280_),
    .o(\u0.w[0][30] ));
 b15fpn000hn1n04x5 _35667_ (.clk(clknet_leaf_11_clk),
    .d(_00281_),
    .o(\u0.w[0][31] ));
 b15fpn000hn1n04x5 _35668_ (.clk(clknet_leaf_12_clk),
    .d(_00289_),
    .o(\u0.w[1][0] ));
 b15fpn000hn1n04x5 _35669_ (.clk(clknet_leaf_4_clk),
    .d(_00300_),
    .o(\u0.w[1][1] ));
 b15fpn000hn1n04x5 _35670_ (.clk(clknet_leaf_10_clk),
    .d(_00311_),
    .o(\u0.w[1][2] ));
 b15fpn000hn1n04x5 _35671_ (.clk(clknet_leaf_8_clk),
    .d(_00314_),
    .o(\u0.w[1][3] ));
 b15fpn000hn1n04x5 _35672_ (.clk(clknet_leaf_1_clk),
    .d(_00315_),
    .o(\u0.w[1][4] ));
 b15fpn000hn1n04x5 _35673_ (.clk(clknet_leaf_18_clk),
    .d(_00316_),
    .o(\u0.w[1][5] ));
 b15fpn000hn1n04x5 _35674_ (.clk(clknet_leaf_15_clk),
    .d(_00317_),
    .o(\u0.w[1][6] ));
 b15fpn000hn1n04x5 _35675_ (.clk(clknet_leaf_1_clk),
    .d(_00318_),
    .o(\u0.w[1][7] ));
 b15fpn000hn1n04x5 _35676_ (.clk(clknet_leaf_8_clk),
    .d(_00319_),
    .o(\u0.w[1][8] ));
 b15fpn000hn1n04x5 _35677_ (.clk(clknet_leaf_9_clk),
    .d(_00320_),
    .o(\u0.w[1][9] ));
 b15fpn000hn1n04x5 _35678_ (.clk(clknet_leaf_10_clk),
    .d(_00290_),
    .o(\u0.w[1][10] ));
 b15fpn000hn1n04x5 _35679_ (.clk(clknet_leaf_10_clk),
    .d(_00291_),
    .o(\u0.w[1][11] ));
 b15fpn000hn1n04x5 _35680_ (.clk(clknet_leaf_1_clk),
    .d(_00292_),
    .o(\u0.w[1][12] ));
 b15fpn000hn1n04x5 _35681_ (.clk(clknet_leaf_1_clk),
    .d(_00293_),
    .o(\u0.w[1][13] ));
 b15fpn000hn1n04x5 _35682_ (.clk(clknet_leaf_15_clk),
    .d(_00294_),
    .o(\u0.w[1][14] ));
 b15fpn000hn1n04x5 _35683_ (.clk(clknet_leaf_1_clk),
    .d(_00295_),
    .o(\u0.w[1][15] ));
 b15fpn000hn1n04x5 _35684_ (.clk(clknet_leaf_7_clk),
    .d(_00296_),
    .o(\u0.w[1][16] ));
 b15fpn000hn1n04x5 _35685_ (.clk(clknet_leaf_9_clk),
    .d(_00297_),
    .o(\u0.w[1][17] ));
 b15fpn000hn1n04x5 _35686_ (.clk(clknet_leaf_7_clk),
    .d(_00298_),
    .o(\u0.w[1][18] ));
 b15fpn000hn1n04x5 _35687_ (.clk(clknet_leaf_8_clk),
    .d(_00299_),
    .o(\u0.w[1][19] ));
 b15fpn000hn1n04x5 _35688_ (.clk(clknet_leaf_1_clk),
    .d(_00301_),
    .o(\u0.w[1][20] ));
 b15fpn000hn1n04x5 _35689_ (.clk(clknet_leaf_0_clk),
    .d(_00302_),
    .o(\u0.w[1][21] ));
 b15fpn000hn1n04x5 _35690_ (.clk(clknet_leaf_0_clk),
    .d(_00303_),
    .o(\u0.w[1][22] ));
 b15fpn000hn1n04x5 _35691_ (.clk(clknet_leaf_9_clk),
    .d(_00304_),
    .o(\u0.w[1][23] ));
 b15fpn000hn1n04x5 _35692_ (.clk(clknet_leaf_9_clk),
    .d(_00305_),
    .o(\u0.w[1][24] ));
 b15fpn000hn1n04x5 _35693_ (.clk(clknet_leaf_8_clk),
    .d(_00306_),
    .o(\u0.w[1][25] ));
 b15fpn000hn1n04x5 _35694_ (.clk(clknet_leaf_9_clk),
    .d(_00307_),
    .o(\u0.w[1][26] ));
 b15fpn000hn1n04x5 _35695_ (.clk(clknet_leaf_11_clk),
    .d(_00308_),
    .o(\u0.w[1][27] ));
 b15fpn000hn1n04x5 _35696_ (.clk(clknet_leaf_11_clk),
    .d(_00309_),
    .o(\u0.w[1][28] ));
 b15fpn000hn1n04x5 _35697_ (.clk(clknet_leaf_1_clk),
    .d(_00310_),
    .o(\u0.w[1][29] ));
 b15fpn000hn1n04x5 _35698_ (.clk(clknet_leaf_15_clk),
    .d(_00312_),
    .o(\u0.w[1][30] ));
 b15fpn000hn1n04x5 _35699_ (.clk(clknet_leaf_15_clk),
    .d(_00313_),
    .o(\u0.w[1][31] ));
 b15fpn000hn1n04x5 _35700_ (.clk(clknet_leaf_12_clk),
    .d(_00321_),
    .o(\u0.w[2][0] ));
 b15fpn000hn1n04x5 _35701_ (.clk(clknet_leaf_4_clk),
    .d(_00332_),
    .o(\u0.w[2][1] ));
 b15fpn000hn1n04x5 _35702_ (.clk(clknet_leaf_1_clk),
    .d(_00343_),
    .o(\u0.w[2][2] ));
 b15fpn000hn1n04x5 _35703_ (.clk(clknet_leaf_8_clk),
    .d(_00346_),
    .o(\u0.w[2][3] ));
 b15fpn000hn1n04x5 _35704_ (.clk(clknet_leaf_1_clk),
    .d(_00347_),
    .o(\u0.w[2][4] ));
 b15fpn000hn1n04x5 _35705_ (.clk(clknet_leaf_18_clk),
    .d(_00348_),
    .o(\u0.w[2][5] ));
 b15fpn000hn1n04x5 _35706_ (.clk(clknet_leaf_17_clk),
    .d(_00349_),
    .o(\u0.w[2][6] ));
 b15fpn000hn1n04x5 _35707_ (.clk(clknet_leaf_17_clk),
    .d(_00350_),
    .o(\u0.w[2][7] ));
 b15fpn000hn1n04x5 _35708_ (.clk(clknet_leaf_8_clk),
    .d(_00351_),
    .o(\u0.w[2][8] ));
 b15fpn000hn1n04x5 _35709_ (.clk(clknet_leaf_10_clk),
    .d(_00352_),
    .o(\u0.w[2][9] ));
 b15fpn000hn1n04x5 _35710_ (.clk(clknet_leaf_10_clk),
    .d(_00322_),
    .o(\u0.w[2][10] ));
 b15fpn000hn1n04x5 _35711_ (.clk(clknet_leaf_10_clk),
    .d(_00323_),
    .o(\u0.w[2][11] ));
 b15fpn000hn1n04x5 _35712_ (.clk(clknet_leaf_15_clk),
    .d(_00324_),
    .o(\u0.w[2][12] ));
 b15fpn000hn1n04x5 _35713_ (.clk(clknet_leaf_15_clk),
    .d(_00325_),
    .o(\u0.w[2][13] ));
 b15fpn000hn1n04x5 _35714_ (.clk(clknet_leaf_17_clk),
    .d(_00326_),
    .o(\u0.w[2][14] ));
 b15fpn000hn1n04x5 _35715_ (.clk(clknet_leaf_15_clk),
    .d(_00327_),
    .o(\u0.w[2][15] ));
 b15fpn000hn1n04x5 _35716_ (.clk(clknet_leaf_7_clk),
    .d(_00328_),
    .o(\u0.w[2][16] ));
 b15fpn000hn1n04x5 _35717_ (.clk(clknet_leaf_8_clk),
    .d(_00329_),
    .o(\u0.w[2][17] ));
 b15fpn000hn1n04x5 _35718_ (.clk(clknet_leaf_7_clk),
    .d(_00330_),
    .o(\u0.w[2][18] ));
 b15fpn000hn1n04x5 _35719_ (.clk(clknet_leaf_8_clk),
    .d(_00331_),
    .o(\u0.w[2][19] ));
 b15fpn000hn1n04x5 _35720_ (.clk(clknet_leaf_17_clk),
    .d(_00333_),
    .o(\u0.w[2][20] ));
 b15fpn000hn1n04x5 _35721_ (.clk(clknet_leaf_18_clk),
    .d(_00334_),
    .o(\u0.w[2][21] ));
 b15fpn000hn1n04x5 _35722_ (.clk(clknet_leaf_17_clk),
    .d(_00335_),
    .o(\u0.w[2][22] ));
 b15fpn000hn1n04x5 _35723_ (.clk(clknet_leaf_15_clk),
    .d(_00336_),
    .o(\u0.w[2][23] ));
 b15fpn000hn1n04x5 _35724_ (.clk(clknet_leaf_9_clk),
    .d(_00337_),
    .o(\u0.w[2][24] ));
 b15fpn000hn1n04x5 _35725_ (.clk(clknet_leaf_8_clk),
    .d(_00338_),
    .o(\u0.w[2][25] ));
 b15fpn000hn1n04x5 _35726_ (.clk(clknet_leaf_9_clk),
    .d(_00339_),
    .o(\u0.w[2][26] ));
 b15fpn000hn1n04x5 _35727_ (.clk(clknet_leaf_11_clk),
    .d(_00340_),
    .o(\u0.w[2][27] ));
 b15fpn000hn1n04x5 _35728_ (.clk(clknet_leaf_10_clk),
    .d(_00341_),
    .o(\u0.w[2][28] ));
 b15fpn000hn1n04x5 _35729_ (.clk(clknet_leaf_15_clk),
    .d(_00342_),
    .o(\u0.w[2][29] ));
 b15fpn000hn1n04x5 _35730_ (.clk(clknet_leaf_16_clk),
    .d(_00344_),
    .o(\u0.w[2][30] ));
 b15fpn000hn1n04x5 _35731_ (.clk(clknet_leaf_17_clk),
    .d(_00345_),
    .o(\u0.w[2][31] ));
 b15fpn000hn1n04x5 _35732_ (.clk(clknet_leaf_12_clk),
    .d(_00353_),
    .o(\u0.tmp_w[0] ));
 b15fpn000hn1n04x5 _35733_ (.clk(clknet_leaf_4_clk),
    .d(_00364_),
    .o(\u0.tmp_w[1] ));
 b15fpn000hn1n04x5 _35734_ (.clk(clknet_leaf_4_clk),
    .d(_00375_),
    .o(\u0.tmp_w[2] ));
 b15fpn000hn1n04x5 _35735_ (.clk(clknet_leaf_7_clk),
    .d(_00378_),
    .o(\u0.tmp_w[3] ));
 b15fpn000hn1n04x5 _35736_ (.clk(clknet_leaf_4_clk),
    .d(_00379_),
    .o(\u0.tmp_w[4] ));
 b15fpn000hn1n04x5 _35737_ (.clk(clknet_leaf_17_clk),
    .d(_00380_),
    .o(\u0.tmp_w[5] ));
 b15fpn000hn1n04x5 _35738_ (.clk(clknet_leaf_17_clk),
    .d(_00381_),
    .o(\u0.tmp_w[6] ));
 b15fpn000hn1n04x5 _35739_ (.clk(clknet_leaf_16_clk),
    .d(_00382_),
    .o(\u0.tmp_w[7] ));
 b15fpn000hn1n04x5 _35740_ (.clk(clknet_leaf_7_clk),
    .d(_00383_),
    .o(\u0.tmp_w[8] ));
 b15fpn000hn1n04x5 _35741_ (.clk(clknet_leaf_5_clk),
    .d(_00384_),
    .o(\u0.tmp_w[9] ));
 b15fpn000hn1n04x5 _35742_ (.clk(clknet_leaf_5_clk),
    .d(_00354_),
    .o(\u0.tmp_w[10] ));
 b15fpn000hn1n04x5 _35743_ (.clk(clknet_leaf_10_clk),
    .d(_00355_),
    .o(\u0.tmp_w[11] ));
 b15fpn000hn1n04x5 _35744_ (.clk(clknet_leaf_4_clk),
    .d(_00356_),
    .o(\u0.tmp_w[12] ));
 b15fpn000hn1n04x5 _35745_ (.clk(clknet_leaf_4_clk),
    .d(_00357_),
    .o(\u0.tmp_w[13] ));
 b15fpn000hn1n04x5 _35746_ (.clk(clknet_leaf_4_clk),
    .d(_00358_),
    .o(\u0.tmp_w[14] ));
 b15fpn000hn1n04x5 _35747_ (.clk(clknet_leaf_4_clk),
    .d(_00359_),
    .o(\u0.tmp_w[15] ));
 b15fpn000hn1n04x5 _35748_ (.clk(clknet_leaf_7_clk),
    .d(_00360_),
    .o(\u0.tmp_w[16] ));
 b15fpn000hn1n04x5 _35749_ (.clk(clknet_leaf_8_clk),
    .d(_00361_),
    .o(\u0.tmp_w[17] ));
 b15fpn000hn1n04x5 _35750_ (.clk(clknet_leaf_7_clk),
    .d(_00362_),
    .o(\u0.tmp_w[18] ));
 b15fpn000hn1n04x5 _35751_ (.clk(clknet_leaf_8_clk),
    .d(_00363_),
    .o(\u0.tmp_w[19] ));
 b15fpn000hn1n04x5 _35752_ (.clk(clknet_leaf_15_clk),
    .d(_00365_),
    .o(\u0.tmp_w[20] ));
 b15fpn000hn1n04x5 _35753_ (.clk(clknet_leaf_0_clk),
    .d(_00366_),
    .o(\u0.tmp_w[21] ));
 b15fpn000hn1n04x5 _35754_ (.clk(clknet_leaf_17_clk),
    .d(_00367_),
    .o(\u0.tmp_w[22] ));
 b15fpn000hn1n04x5 _35755_ (.clk(clknet_leaf_15_clk),
    .d(_00368_),
    .o(\u0.tmp_w[23] ));
 b15fpn000hn1n04x5 _35756_ (.clk(clknet_leaf_9_clk),
    .d(_00369_),
    .o(\u0.tmp_w[24] ));
 b15fpn000hn1n04x5 _35757_ (.clk(clknet_leaf_9_clk),
    .d(_00370_),
    .o(\u0.tmp_w[25] ));
 b15fpn000hn1n04x5 _35758_ (.clk(clknet_leaf_6_clk),
    .d(_00371_),
    .o(\u0.tmp_w[26] ));
 b15fpn000hn1n04x5 _35759_ (.clk(clknet_leaf_10_clk),
    .d(_00372_),
    .o(\u0.tmp_w[27] ));
 b15fpn000hn1n04x5 _35760_ (.clk(clknet_leaf_4_clk),
    .d(_00373_),
    .o(\u0.tmp_w[28] ));
 b15fpn000hn1n04x5 _35761_ (.clk(clknet_leaf_4_clk),
    .d(_00374_),
    .o(\u0.tmp_w[29] ));
 b15fpn000hn1n04x5 _35762_ (.clk(clknet_leaf_16_clk),
    .d(_00376_),
    .o(\u0.tmp_w[30] ));
 b15fpn000hn1n04x5 _35763_ (.clk(clknet_leaf_4_clk),
    .d(_00377_),
    .o(\u0.tmp_w[31] ));
 b15zdnd11an1n64x5 FILLER_1_1688 ();
 b15zdnd11an1n64x5 FILLER_1_1752 ();
 b15zdnd11an1n64x5 FILLER_1_1816 ();
 b15zdnd11an1n64x5 FILLER_1_1880 ();
 b15zdnd11an1n64x5 FILLER_1_1944 ();
 b15zdnd11an1n64x5 FILLER_1_2008 ();
 b15zdnd11an1n64x5 FILLER_1_2072 ();
 b15zdnd11an1n64x5 FILLER_1_2136 ();
 b15zdnd11an1n64x5 FILLER_1_2200 ();
 b15zdnd11an1n16x5 FILLER_1_2264 ();
 b15zdnd11an1n04x5 FILLER_1_2280 ();
 b15zdnd11an1n64x5 FILLER_2_8 ();
 b15zdnd11an1n64x5 FILLER_2_72 ();
 b15zdnd11an1n64x5 FILLER_2_136 ();
 b15zdnd11an1n64x5 FILLER_2_200 ();
 b15zdnd11an1n64x5 FILLER_2_264 ();
 b15zdnd11an1n64x5 FILLER_2_328 ();
 b15zdnd11an1n16x5 FILLER_2_392 ();
 b15zdnd11an1n08x5 FILLER_2_408 ();
 b15zdnd11an1n04x5 FILLER_2_416 ();
 b15zdnd11an1n64x5 FILLER_2_427 ();
 b15zdnd11an1n16x5 FILLER_2_491 ();
 b15zdnd11an1n08x5 FILLER_2_507 ();
 b15zdnd00an1n02x5 FILLER_2_515 ();
 b15zdnd11an1n04x5 FILLER_2_522 ();
 b15zdnd11an1n04x5 FILLER_2_542 ();
 b15zdnd11an1n16x5 FILLER_2_551 ();
 b15zdnd11an1n08x5 FILLER_2_567 ();
 b15zdnd00an1n01x5 FILLER_2_575 ();
 b15zdnd11an1n04x5 FILLER_2_584 ();
 b15zdnd11an1n08x5 FILLER_2_600 ();
 b15zdnd00an1n02x5 FILLER_2_608 ();
 b15zdnd00an1n01x5 FILLER_2_610 ();
 b15zdnd11an1n16x5 FILLER_2_626 ();
 b15zdnd11an1n04x5 FILLER_2_642 ();
 b15zdnd00an1n02x5 FILLER_2_646 ();
 b15zdnd00an1n01x5 FILLER_2_648 ();
 b15zdnd11an1n32x5 FILLER_2_653 ();
 b15zdnd11an1n16x5 FILLER_2_685 ();
 b15zdnd00an1n02x5 FILLER_2_701 ();
 b15zdnd11an1n08x5 FILLER_2_707 ();
 b15zdnd00an1n02x5 FILLER_2_715 ();
 b15zdnd00an1n01x5 FILLER_2_717 ();
 b15zdnd11an1n16x5 FILLER_2_726 ();
 b15zdnd00an1n01x5 FILLER_2_742 ();
 b15zdnd11an1n16x5 FILLER_2_759 ();
 b15zdnd11an1n32x5 FILLER_2_782 ();
 b15zdnd11an1n16x5 FILLER_2_814 ();
 b15zdnd00an1n01x5 FILLER_2_830 ();
 b15zdnd11an1n64x5 FILLER_2_836 ();
 b15zdnd11an1n16x5 FILLER_2_900 ();
 b15zdnd11an1n08x5 FILLER_2_916 ();
 b15zdnd00an1n02x5 FILLER_2_924 ();
 b15zdnd00an1n01x5 FILLER_2_926 ();
 b15zdnd11an1n32x5 FILLER_2_931 ();
 b15zdnd11an1n16x5 FILLER_2_963 ();
 b15zdnd11an1n04x5 FILLER_2_979 ();
 b15zdnd00an1n02x5 FILLER_2_983 ();
 b15zdnd00an1n01x5 FILLER_2_985 ();
 b15zdnd11an1n04x5 FILLER_2_990 ();
 b15zdnd11an1n08x5 FILLER_2_997 ();
 b15zdnd00an1n02x5 FILLER_2_1005 ();
 b15zdnd00an1n01x5 FILLER_2_1007 ();
 b15zdnd11an1n04x5 FILLER_2_1012 ();
 b15zdnd11an1n04x5 FILLER_2_1022 ();
 b15zdnd11an1n04x5 FILLER_2_1030 ();
 b15zdnd11an1n04x5 FILLER_2_1038 ();
 b15zdnd11an1n04x5 FILLER_2_1046 ();
 b15zdnd11an1n04x5 FILLER_2_1055 ();
 b15zdnd11an1n08x5 FILLER_2_1063 ();
 b15zdnd11an1n08x5 FILLER_2_1075 ();
 b15zdnd11an1n04x5 FILLER_2_1083 ();
 b15zdnd00an1n02x5 FILLER_2_1087 ();
 b15zdnd00an1n01x5 FILLER_2_1089 ();
 b15zdnd11an1n04x5 FILLER_2_1094 ();
 b15zdnd11an1n04x5 FILLER_2_1102 ();
 b15zdnd00an1n02x5 FILLER_2_1106 ();
 b15zdnd11an1n04x5 FILLER_2_1112 ();
 b15zdnd11an1n08x5 FILLER_2_1121 ();
 b15zdnd00an1n02x5 FILLER_2_1129 ();
 b15zdnd11an1n08x5 FILLER_2_1135 ();
 b15zdnd11an1n04x5 FILLER_2_1143 ();
 b15zdnd11an1n04x5 FILLER_2_1153 ();
 b15zdnd11an1n04x5 FILLER_2_1161 ();
 b15zdnd11an1n04x5 FILLER_2_1170 ();
 b15zdnd00an1n02x5 FILLER_2_1174 ();
 b15zdnd11an1n08x5 FILLER_2_1180 ();
 b15zdnd00an1n02x5 FILLER_2_1188 ();
 b15zdnd11an1n16x5 FILLER_2_1210 ();
 b15zdnd00an1n02x5 FILLER_2_1226 ();
 b15zdnd00an1n01x5 FILLER_2_1228 ();
 b15zdnd11an1n04x5 FILLER_2_1233 ();
 b15zdnd11an1n04x5 FILLER_2_1241 ();
 b15zdnd00an1n01x5 FILLER_2_1245 ();
 b15zdnd11an1n04x5 FILLER_2_1251 ();
 b15zdnd00an1n02x5 FILLER_2_1255 ();
 b15zdnd00an1n01x5 FILLER_2_1257 ();
 b15zdnd11an1n16x5 FILLER_2_1262 ();
 b15zdnd11an1n04x5 FILLER_2_1278 ();
 b15zdnd11an1n08x5 FILLER_2_1288 ();
 b15zdnd11an1n04x5 FILLER_2_1296 ();
 b15zdnd11an1n04x5 FILLER_2_1304 ();
 b15zdnd00an1n02x5 FILLER_2_1308 ();
 b15zdnd11an1n08x5 FILLER_2_1314 ();
 b15zdnd11an1n04x5 FILLER_2_1322 ();
 b15zdnd00an1n02x5 FILLER_2_1326 ();
 b15zdnd11an1n64x5 FILLER_2_1348 ();
 b15zdnd11an1n04x5 FILLER_2_1412 ();
 b15zdnd00an1n02x5 FILLER_2_1416 ();
 b15zdnd00an1n01x5 FILLER_2_1418 ();
 b15zdnd11an1n08x5 FILLER_2_1423 ();
 b15zdnd11an1n04x5 FILLER_2_1431 ();
 b15zdnd11an1n08x5 FILLER_2_1441 ();
 b15zdnd11an1n04x5 FILLER_2_1449 ();
 b15zdnd11an1n32x5 FILLER_2_1457 ();
 b15zdnd00an1n01x5 FILLER_2_1489 ();
 b15zdnd11an1n64x5 FILLER_2_1495 ();
 b15zdnd11an1n16x5 FILLER_2_1559 ();
 b15zdnd11an1n08x5 FILLER_2_1575 ();
 b15zdnd11an1n64x5 FILLER_2_1589 ();
 b15zdnd00an1n02x5 FILLER_2_1653 ();
 b15zdnd11an1n32x5 FILLER_2_1675 ();
 b15zdnd11an1n04x5 FILLER_2_1707 ();
 b15zdnd00an1n02x5 FILLER_2_1711 ();
 b15zdnd11an1n04x5 FILLER_2_1725 ();
 b15zdnd11an1n16x5 FILLER_2_1741 ();
 b15zdnd11an1n64x5 FILLER_2_1773 ();
 b15zdnd11an1n16x5 FILLER_2_1837 ();
 b15zdnd11an1n32x5 FILLER_2_1866 ();
 b15zdnd11an1n16x5 FILLER_2_1898 ();
 b15zdnd11an1n08x5 FILLER_2_1914 ();
 b15zdnd00an1n02x5 FILLER_2_1922 ();
 b15zdnd11an1n16x5 FILLER_2_1931 ();
 b15zdnd11an1n08x5 FILLER_2_1947 ();
 b15zdnd11an1n04x5 FILLER_2_1955 ();
 b15zdnd00an1n02x5 FILLER_2_1959 ();
 b15zdnd11an1n64x5 FILLER_2_1967 ();
 b15zdnd00an1n02x5 FILLER_2_2031 ();
 b15zdnd00an1n01x5 FILLER_2_2033 ();
 b15zdnd11an1n32x5 FILLER_2_2043 ();
 b15zdnd11an1n04x5 FILLER_2_2075 ();
 b15zdnd00an1n02x5 FILLER_2_2079 ();
 b15zdnd00an1n01x5 FILLER_2_2081 ();
 b15zdnd11an1n16x5 FILLER_2_2094 ();
 b15zdnd11an1n08x5 FILLER_2_2110 ();
 b15zdnd00an1n02x5 FILLER_2_2118 ();
 b15zdnd11an1n16x5 FILLER_2_2132 ();
 b15zdnd11an1n04x5 FILLER_2_2148 ();
 b15zdnd00an1n02x5 FILLER_2_2152 ();
 b15zdnd11an1n64x5 FILLER_2_2162 ();
 b15zdnd11an1n32x5 FILLER_2_2226 ();
 b15zdnd11an1n16x5 FILLER_2_2258 ();
 b15zdnd00an1n02x5 FILLER_2_2274 ();
 b15zdnd11an1n64x5 FILLER_3_0 ();
 b15zdnd11an1n64x5 FILLER_3_64 ();
 b15zdnd11an1n64x5 FILLER_3_128 ();
 b15zdnd11an1n64x5 FILLER_3_192 ();
 b15zdnd11an1n64x5 FILLER_3_256 ();
 b15zdnd11an1n64x5 FILLER_3_320 ();
 b15zdnd11an1n08x5 FILLER_3_384 ();
 b15zdnd00an1n01x5 FILLER_3_392 ();
 b15zdnd11an1n04x5 FILLER_3_411 ();
 b15zdnd11an1n04x5 FILLER_3_422 ();
 b15zdnd11an1n04x5 FILLER_3_433 ();
 b15zdnd11an1n08x5 FILLER_3_455 ();
 b15zdnd11an1n04x5 FILLER_3_463 ();
 b15zdnd00an1n02x5 FILLER_3_467 ();
 b15zdnd00an1n01x5 FILLER_3_469 ();
 b15zdnd11an1n08x5 FILLER_3_476 ();
 b15zdnd00an1n01x5 FILLER_3_484 ();
 b15zdnd11an1n04x5 FILLER_3_503 ();
 b15zdnd11an1n04x5 FILLER_3_513 ();
 b15zdnd00an1n02x5 FILLER_3_517 ();
 b15zdnd11an1n08x5 FILLER_3_527 ();
 b15zdnd11an1n04x5 FILLER_3_535 ();
 b15zdnd00an1n01x5 FILLER_3_539 ();
 b15zdnd11an1n16x5 FILLER_3_551 ();
 b15zdnd11an1n08x5 FILLER_3_567 ();
 b15zdnd11an1n04x5 FILLER_3_575 ();
 b15zdnd11an1n04x5 FILLER_3_597 ();
 b15zdnd11an1n04x5 FILLER_3_632 ();
 b15zdnd11an1n04x5 FILLER_3_640 ();
 b15zdnd11an1n04x5 FILLER_3_653 ();
 b15zdnd11an1n04x5 FILLER_3_665 ();
 b15zdnd00an1n01x5 FILLER_3_669 ();
 b15zdnd11an1n04x5 FILLER_3_678 ();
 b15zdnd00an1n01x5 FILLER_3_682 ();
 b15zdnd11an1n08x5 FILLER_3_690 ();
 b15zdnd11an1n16x5 FILLER_3_712 ();
 b15zdnd00an1n01x5 FILLER_3_728 ();
 b15zdnd11an1n16x5 FILLER_3_746 ();
 b15zdnd00an1n01x5 FILLER_3_762 ();
 b15zdnd11an1n04x5 FILLER_3_771 ();
 b15zdnd11an1n16x5 FILLER_3_791 ();
 b15zdnd11an1n04x5 FILLER_3_807 ();
 b15zdnd00an1n02x5 FILLER_3_811 ();
 b15zdnd11an1n04x5 FILLER_3_829 ();
 b15zdnd11an1n04x5 FILLER_3_853 ();
 b15zdnd11an1n64x5 FILLER_3_875 ();
 b15zdnd11an1n08x5 FILLER_3_939 ();
 b15zdnd11an1n04x5 FILLER_3_947 ();
 b15zdnd00an1n01x5 FILLER_3_951 ();
 b15zdnd11an1n16x5 FILLER_3_958 ();
 b15zdnd11an1n08x5 FILLER_3_974 ();
 b15zdnd11an1n04x5 FILLER_3_982 ();
 b15zdnd11an1n04x5 FILLER_3_1006 ();
 b15zdnd11an1n16x5 FILLER_3_1030 ();
 b15zdnd11an1n08x5 FILLER_3_1046 ();
 b15zdnd00an1n01x5 FILLER_3_1054 ();
 b15zdnd11an1n16x5 FILLER_3_1060 ();
 b15zdnd11an1n04x5 FILLER_3_1076 ();
 b15zdnd00an1n01x5 FILLER_3_1080 ();
 b15zdnd11an1n08x5 FILLER_3_1101 ();
 b15zdnd11an1n04x5 FILLER_3_1109 ();
 b15zdnd11an1n04x5 FILLER_3_1117 ();
 b15zdnd00an1n01x5 FILLER_3_1121 ();
 b15zdnd11an1n08x5 FILLER_3_1142 ();
 b15zdnd11an1n04x5 FILLER_3_1150 ();
 b15zdnd11an1n04x5 FILLER_3_1159 ();
 b15zdnd00an1n02x5 FILLER_3_1163 ();
 b15zdnd00an1n01x5 FILLER_3_1165 ();
 b15zdnd11an1n04x5 FILLER_3_1170 ();
 b15zdnd00an1n02x5 FILLER_3_1174 ();
 b15zdnd11an1n04x5 FILLER_3_1180 ();
 b15zdnd00an1n02x5 FILLER_3_1184 ();
 b15zdnd11an1n08x5 FILLER_3_1190 ();
 b15zdnd11an1n04x5 FILLER_3_1202 ();
 b15zdnd00an1n02x5 FILLER_3_1206 ();
 b15zdnd11an1n08x5 FILLER_3_1212 ();
 b15zdnd11an1n04x5 FILLER_3_1223 ();
 b15zdnd11an1n08x5 FILLER_3_1231 ();
 b15zdnd11an1n08x5 FILLER_3_1245 ();
 b15zdnd00an1n01x5 FILLER_3_1253 ();
 b15zdnd11an1n16x5 FILLER_3_1260 ();
 b15zdnd11an1n04x5 FILLER_3_1276 ();
 b15zdnd00an1n01x5 FILLER_3_1280 ();
 b15zdnd11an1n08x5 FILLER_3_1286 ();
 b15zdnd11an1n04x5 FILLER_3_1294 ();
 b15zdnd00an1n02x5 FILLER_3_1298 ();
 b15zdnd00an1n01x5 FILLER_3_1300 ();
 b15zdnd11an1n04x5 FILLER_3_1321 ();
 b15zdnd00an1n01x5 FILLER_3_1325 ();
 b15zdnd11an1n16x5 FILLER_3_1331 ();
 b15zdnd11an1n08x5 FILLER_3_1347 ();
 b15zdnd11an1n32x5 FILLER_3_1375 ();
 b15zdnd11an1n16x5 FILLER_3_1411 ();
 b15zdnd00an1n02x5 FILLER_3_1427 ();
 b15zdnd11an1n16x5 FILLER_3_1449 ();
 b15zdnd11an1n16x5 FILLER_3_1469 ();
 b15zdnd00an1n02x5 FILLER_3_1485 ();
 b15zdnd00an1n01x5 FILLER_3_1487 ();
 b15zdnd11an1n64x5 FILLER_3_1508 ();
 b15zdnd11an1n16x5 FILLER_3_1572 ();
 b15zdnd00an1n01x5 FILLER_3_1588 ();
 b15zdnd11an1n64x5 FILLER_3_1594 ();
 b15zdnd11an1n32x5 FILLER_3_1658 ();
 b15zdnd11an1n16x5 FILLER_3_1690 ();
 b15zdnd11an1n08x5 FILLER_3_1706 ();
 b15zdnd11an1n04x5 FILLER_3_1714 ();
 b15zdnd11an1n16x5 FILLER_3_1739 ();
 b15zdnd11an1n08x5 FILLER_3_1755 ();
 b15zdnd11an1n04x5 FILLER_3_1763 ();
 b15zdnd11an1n04x5 FILLER_3_1788 ();
 b15zdnd11an1n04x5 FILLER_3_1800 ();
 b15zdnd11an1n04x5 FILLER_3_1813 ();
 b15zdnd11an1n04x5 FILLER_3_1833 ();
 b15zdnd11an1n16x5 FILLER_3_1845 ();
 b15zdnd00an1n02x5 FILLER_3_1861 ();
 b15zdnd11an1n04x5 FILLER_3_1877 ();
 b15zdnd11an1n16x5 FILLER_3_1894 ();
 b15zdnd00an1n01x5 FILLER_3_1910 ();
 b15zdnd11an1n08x5 FILLER_3_1927 ();
 b15zdnd11an1n04x5 FILLER_3_1935 ();
 b15zdnd00an1n01x5 FILLER_3_1939 ();
 b15zdnd11an1n04x5 FILLER_3_1946 ();
 b15zdnd11an1n04x5 FILLER_3_1957 ();
 b15zdnd00an1n02x5 FILLER_3_1961 ();
 b15zdnd11an1n04x5 FILLER_3_1970 ();
 b15zdnd11an1n04x5 FILLER_3_1980 ();
 b15zdnd11an1n04x5 FILLER_3_1993 ();
 b15zdnd00an1n01x5 FILLER_3_1997 ();
 b15zdnd11an1n04x5 FILLER_3_2002 ();
 b15zdnd11an1n04x5 FILLER_3_2020 ();
 b15zdnd11an1n08x5 FILLER_3_2030 ();
 b15zdnd11an1n04x5 FILLER_3_2038 ();
 b15zdnd00an1n01x5 FILLER_3_2042 ();
 b15zdnd11an1n04x5 FILLER_3_2055 ();
 b15zdnd11an1n08x5 FILLER_3_2063 ();
 b15zdnd11an1n08x5 FILLER_3_2075 ();
 b15zdnd00an1n02x5 FILLER_3_2083 ();
 b15zdnd11an1n16x5 FILLER_3_2092 ();
 b15zdnd11an1n04x5 FILLER_3_2108 ();
 b15zdnd00an1n01x5 FILLER_3_2112 ();
 b15zdnd11an1n64x5 FILLER_3_2130 ();
 b15zdnd11an1n64x5 FILLER_3_2194 ();
 b15zdnd11an1n16x5 FILLER_3_2258 ();
 b15zdnd11an1n08x5 FILLER_3_2274 ();
 b15zdnd00an1n02x5 FILLER_3_2282 ();
 b15zdnd11an1n64x5 FILLER_4_8 ();
 b15zdnd11an1n64x5 FILLER_4_72 ();
 b15zdnd11an1n64x5 FILLER_4_136 ();
 b15zdnd11an1n64x5 FILLER_4_200 ();
 b15zdnd11an1n64x5 FILLER_4_264 ();
 b15zdnd11an1n64x5 FILLER_4_328 ();
 b15zdnd11an1n16x5 FILLER_4_392 ();
 b15zdnd11an1n04x5 FILLER_4_408 ();
 b15zdnd00an1n01x5 FILLER_4_412 ();
 b15zdnd11an1n16x5 FILLER_4_434 ();
 b15zdnd11an1n04x5 FILLER_4_450 ();
 b15zdnd00an1n02x5 FILLER_4_454 ();
 b15zdnd11an1n04x5 FILLER_4_464 ();
 b15zdnd11an1n08x5 FILLER_4_480 ();
 b15zdnd11an1n04x5 FILLER_4_488 ();
 b15zdnd00an1n02x5 FILLER_4_492 ();
 b15zdnd11an1n04x5 FILLER_4_500 ();
 b15zdnd11an1n64x5 FILLER_4_514 ();
 b15zdnd11an1n16x5 FILLER_4_578 ();
 b15zdnd11an1n08x5 FILLER_4_594 ();
 b15zdnd00an1n02x5 FILLER_4_602 ();
 b15zdnd00an1n01x5 FILLER_4_604 ();
 b15zdnd11an1n08x5 FILLER_4_621 ();
 b15zdnd00an1n02x5 FILLER_4_629 ();
 b15zdnd00an1n01x5 FILLER_4_631 ();
 b15zdnd11an1n08x5 FILLER_4_658 ();
 b15zdnd11an1n04x5 FILLER_4_666 ();
 b15zdnd00an1n01x5 FILLER_4_670 ();
 b15zdnd11an1n32x5 FILLER_4_676 ();
 b15zdnd11an1n08x5 FILLER_4_708 ();
 b15zdnd00an1n02x5 FILLER_4_716 ();
 b15zdnd11an1n04x5 FILLER_4_726 ();
 b15zdnd11an1n04x5 FILLER_4_746 ();
 b15zdnd11an1n16x5 FILLER_4_772 ();
 b15zdnd11an1n08x5 FILLER_4_788 ();
 b15zdnd00an1n01x5 FILLER_4_796 ();
 b15zdnd11an1n16x5 FILLER_4_813 ();
 b15zdnd11an1n08x5 FILLER_4_829 ();
 b15zdnd11an1n04x5 FILLER_4_842 ();
 b15zdnd11an1n64x5 FILLER_4_862 ();
 b15zdnd11an1n16x5 FILLER_4_926 ();
 b15zdnd00an1n02x5 FILLER_4_942 ();
 b15zdnd00an1n01x5 FILLER_4_944 ();
 b15zdnd11an1n16x5 FILLER_4_965 ();
 b15zdnd11an1n08x5 FILLER_4_981 ();
 b15zdnd11an1n04x5 FILLER_4_989 ();
 b15zdnd00an1n01x5 FILLER_4_993 ();
 b15zdnd11an1n16x5 FILLER_4_998 ();
 b15zdnd00an1n02x5 FILLER_4_1014 ();
 b15zdnd00an1n01x5 FILLER_4_1016 ();
 b15zdnd11an1n16x5 FILLER_4_1022 ();
 b15zdnd11an1n04x5 FILLER_4_1038 ();
 b15zdnd00an1n02x5 FILLER_4_1042 ();
 b15zdnd00an1n01x5 FILLER_4_1044 ();
 b15zdnd11an1n32x5 FILLER_4_1065 ();
 b15zdnd11an1n16x5 FILLER_4_1097 ();
 b15zdnd11an1n32x5 FILLER_4_1119 ();
 b15zdnd11an1n16x5 FILLER_4_1151 ();
 b15zdnd11an1n08x5 FILLER_4_1167 ();
 b15zdnd00an1n02x5 FILLER_4_1175 ();
 b15zdnd11an1n16x5 FILLER_4_1181 ();
 b15zdnd11an1n08x5 FILLER_4_1197 ();
 b15zdnd00an1n02x5 FILLER_4_1205 ();
 b15zdnd00an1n01x5 FILLER_4_1207 ();
 b15zdnd11an1n08x5 FILLER_4_1212 ();
 b15zdnd00an1n02x5 FILLER_4_1220 ();
 b15zdnd00an1n01x5 FILLER_4_1222 ();
 b15zdnd11an1n16x5 FILLER_4_1243 ();
 b15zdnd11an1n08x5 FILLER_4_1259 ();
 b15zdnd11an1n04x5 FILLER_4_1267 ();
 b15zdnd11an1n04x5 FILLER_4_1291 ();
 b15zdnd00an1n02x5 FILLER_4_1295 ();
 b15zdnd11an1n64x5 FILLER_4_1317 ();
 b15zdnd11an1n32x5 FILLER_4_1381 ();
 b15zdnd11an1n16x5 FILLER_4_1413 ();
 b15zdnd11an1n08x5 FILLER_4_1429 ();
 b15zdnd00an1n02x5 FILLER_4_1437 ();
 b15zdnd11an1n16x5 FILLER_4_1444 ();
 b15zdnd11an1n04x5 FILLER_4_1460 ();
 b15zdnd00an1n02x5 FILLER_4_1464 ();
 b15zdnd11an1n16x5 FILLER_4_1471 ();
 b15zdnd11an1n08x5 FILLER_4_1487 ();
 b15zdnd11an1n04x5 FILLER_4_1495 ();
 b15zdnd11an1n64x5 FILLER_4_1502 ();
 b15zdnd11an1n16x5 FILLER_4_1566 ();
 b15zdnd11an1n08x5 FILLER_4_1582 ();
 b15zdnd00an1n02x5 FILLER_4_1590 ();
 b15zdnd11an1n64x5 FILLER_4_1612 ();
 b15zdnd11an1n32x5 FILLER_4_1676 ();
 b15zdnd11an1n08x5 FILLER_4_1708 ();
 b15zdnd00an1n02x5 FILLER_4_1716 ();
 b15zdnd00an1n01x5 FILLER_4_1718 ();
 b15zdnd11an1n32x5 FILLER_4_1725 ();
 b15zdnd11an1n16x5 FILLER_4_1757 ();
 b15zdnd11an1n08x5 FILLER_4_1773 ();
 b15zdnd11an1n04x5 FILLER_4_1781 ();
 b15zdnd00an1n01x5 FILLER_4_1785 ();
 b15zdnd11an1n16x5 FILLER_4_1803 ();
 b15zdnd11an1n04x5 FILLER_4_1819 ();
 b15zdnd00an1n01x5 FILLER_4_1823 ();
 b15zdnd11an1n64x5 FILLER_4_1828 ();
 b15zdnd11an1n16x5 FILLER_4_1892 ();
 b15zdnd11an1n08x5 FILLER_4_1908 ();
 b15zdnd00an1n01x5 FILLER_4_1916 ();
 b15zdnd11an1n04x5 FILLER_4_1933 ();
 b15zdnd00an1n01x5 FILLER_4_1937 ();
 b15zdnd11an1n08x5 FILLER_4_1944 ();
 b15zdnd11an1n04x5 FILLER_4_1952 ();
 b15zdnd00an1n01x5 FILLER_4_1956 ();
 b15zdnd11an1n64x5 FILLER_4_1971 ();
 b15zdnd00an1n01x5 FILLER_4_2035 ();
 b15zdnd11an1n04x5 FILLER_4_2041 ();
 b15zdnd11an1n04x5 FILLER_4_2057 ();
 b15zdnd00an1n01x5 FILLER_4_2061 ();
 b15zdnd11an1n04x5 FILLER_4_2072 ();
 b15zdnd00an1n02x5 FILLER_4_2076 ();
 b15zdnd00an1n01x5 FILLER_4_2078 ();
 b15zdnd11an1n04x5 FILLER_4_2094 ();
 b15zdnd11an1n08x5 FILLER_4_2116 ();
 b15zdnd11an1n04x5 FILLER_4_2124 ();
 b15zdnd00an1n02x5 FILLER_4_2128 ();
 b15zdnd00an1n01x5 FILLER_4_2130 ();
 b15zdnd11an1n08x5 FILLER_4_2141 ();
 b15zdnd11an1n04x5 FILLER_4_2149 ();
 b15zdnd00an1n01x5 FILLER_4_2153 ();
 b15zdnd11an1n16x5 FILLER_4_2162 ();
 b15zdnd11an1n04x5 FILLER_4_2178 ();
 b15zdnd11an1n04x5 FILLER_4_2205 ();
 b15zdnd11an1n32x5 FILLER_4_2227 ();
 b15zdnd11an1n16x5 FILLER_4_2259 ();
 b15zdnd00an1n01x5 FILLER_4_2275 ();
 b15zdnd11an1n64x5 FILLER_5_0 ();
 b15zdnd11an1n64x5 FILLER_5_64 ();
 b15zdnd11an1n64x5 FILLER_5_128 ();
 b15zdnd11an1n64x5 FILLER_5_192 ();
 b15zdnd11an1n64x5 FILLER_5_256 ();
 b15zdnd11an1n64x5 FILLER_5_320 ();
 b15zdnd11an1n64x5 FILLER_5_384 ();
 b15zdnd11an1n32x5 FILLER_5_448 ();
 b15zdnd11an1n16x5 FILLER_5_480 ();
 b15zdnd11an1n04x5 FILLER_5_496 ();
 b15zdnd00an1n01x5 FILLER_5_500 ();
 b15zdnd11an1n64x5 FILLER_5_507 ();
 b15zdnd11an1n32x5 FILLER_5_571 ();
 b15zdnd11an1n08x5 FILLER_5_603 ();
 b15zdnd11an1n04x5 FILLER_5_611 ();
 b15zdnd00an1n02x5 FILLER_5_615 ();
 b15zdnd11an1n16x5 FILLER_5_622 ();
 b15zdnd11an1n04x5 FILLER_5_638 ();
 b15zdnd00an1n02x5 FILLER_5_642 ();
 b15zdnd11an1n04x5 FILLER_5_667 ();
 b15zdnd11an1n08x5 FILLER_5_678 ();
 b15zdnd00an1n01x5 FILLER_5_686 ();
 b15zdnd11an1n64x5 FILLER_5_703 ();
 b15zdnd11an1n64x5 FILLER_5_767 ();
 b15zdnd11an1n04x5 FILLER_5_831 ();
 b15zdnd00an1n01x5 FILLER_5_835 ();
 b15zdnd11an1n08x5 FILLER_5_868 ();
 b15zdnd00an1n02x5 FILLER_5_876 ();
 b15zdnd11an1n04x5 FILLER_5_909 ();
 b15zdnd11an1n16x5 FILLER_5_933 ();
 b15zdnd11an1n04x5 FILLER_5_949 ();
 b15zdnd00an1n02x5 FILLER_5_953 ();
 b15zdnd11an1n64x5 FILLER_5_960 ();
 b15zdnd11an1n32x5 FILLER_5_1024 ();
 b15zdnd00an1n01x5 FILLER_5_1056 ();
 b15zdnd11an1n32x5 FILLER_5_1061 ();
 b15zdnd11an1n08x5 FILLER_5_1093 ();
 b15zdnd11an1n04x5 FILLER_5_1101 ();
 b15zdnd00an1n01x5 FILLER_5_1105 ();
 b15zdnd11an1n64x5 FILLER_5_1126 ();
 b15zdnd11an1n16x5 FILLER_5_1210 ();
 b15zdnd11an1n08x5 FILLER_5_1226 ();
 b15zdnd00an1n02x5 FILLER_5_1234 ();
 b15zdnd11an1n64x5 FILLER_5_1241 ();
 b15zdnd11an1n64x5 FILLER_5_1305 ();
 b15zdnd11an1n04x5 FILLER_5_1369 ();
 b15zdnd00an1n02x5 FILLER_5_1373 ();
 b15zdnd11an1n04x5 FILLER_5_1395 ();
 b15zdnd11an1n32x5 FILLER_5_1404 ();
 b15zdnd11an1n16x5 FILLER_5_1436 ();
 b15zdnd11an1n08x5 FILLER_5_1452 ();
 b15zdnd11an1n04x5 FILLER_5_1460 ();
 b15zdnd00an1n01x5 FILLER_5_1464 ();
 b15zdnd11an1n16x5 FILLER_5_1485 ();
 b15zdnd11an1n04x5 FILLER_5_1501 ();
 b15zdnd00an1n02x5 FILLER_5_1505 ();
 b15zdnd11an1n64x5 FILLER_5_1511 ();
 b15zdnd11an1n64x5 FILLER_5_1575 ();
 b15zdnd11an1n32x5 FILLER_5_1639 ();
 b15zdnd11an1n04x5 FILLER_5_1671 ();
 b15zdnd11an1n32x5 FILLER_5_1695 ();
 b15zdnd11an1n08x5 FILLER_5_1727 ();
 b15zdnd11an1n04x5 FILLER_5_1735 ();
 b15zdnd00an1n02x5 FILLER_5_1739 ();
 b15zdnd00an1n01x5 FILLER_5_1741 ();
 b15zdnd11an1n08x5 FILLER_5_1768 ();
 b15zdnd11an1n04x5 FILLER_5_1776 ();
 b15zdnd11an1n08x5 FILLER_5_1803 ();
 b15zdnd11an1n04x5 FILLER_5_1824 ();
 b15zdnd11an1n32x5 FILLER_5_1836 ();
 b15zdnd11an1n08x5 FILLER_5_1868 ();
 b15zdnd00an1n02x5 FILLER_5_1876 ();
 b15zdnd00an1n01x5 FILLER_5_1878 ();
 b15zdnd11an1n08x5 FILLER_5_1897 ();
 b15zdnd11an1n04x5 FILLER_5_1905 ();
 b15zdnd00an1n02x5 FILLER_5_1909 ();
 b15zdnd00an1n01x5 FILLER_5_1911 ();
 b15zdnd11an1n04x5 FILLER_5_1930 ();
 b15zdnd00an1n02x5 FILLER_5_1934 ();
 b15zdnd11an1n08x5 FILLER_5_1950 ();
 b15zdnd11an1n04x5 FILLER_5_1958 ();
 b15zdnd00an1n01x5 FILLER_5_1962 ();
 b15zdnd11an1n32x5 FILLER_5_1969 ();
 b15zdnd11an1n04x5 FILLER_5_2001 ();
 b15zdnd00an1n02x5 FILLER_5_2005 ();
 b15zdnd11an1n32x5 FILLER_5_2013 ();
 b15zdnd00an1n01x5 FILLER_5_2045 ();
 b15zdnd11an1n08x5 FILLER_5_2050 ();
 b15zdnd11an1n04x5 FILLER_5_2058 ();
 b15zdnd00an1n02x5 FILLER_5_2062 ();
 b15zdnd00an1n01x5 FILLER_5_2064 ();
 b15zdnd11an1n32x5 FILLER_5_2089 ();
 b15zdnd11an1n04x5 FILLER_5_2121 ();
 b15zdnd11an1n04x5 FILLER_5_2131 ();
 b15zdnd11an1n64x5 FILLER_5_2156 ();
 b15zdnd11an1n64x5 FILLER_5_2220 ();
 b15zdnd11an1n64x5 FILLER_6_8 ();
 b15zdnd11an1n64x5 FILLER_6_72 ();
 b15zdnd11an1n64x5 FILLER_6_136 ();
 b15zdnd11an1n64x5 FILLER_6_200 ();
 b15zdnd11an1n64x5 FILLER_6_264 ();
 b15zdnd11an1n64x5 FILLER_6_328 ();
 b15zdnd11an1n64x5 FILLER_6_392 ();
 b15zdnd11an1n64x5 FILLER_6_456 ();
 b15zdnd11an1n08x5 FILLER_6_520 ();
 b15zdnd00an1n02x5 FILLER_6_528 ();
 b15zdnd11an1n04x5 FILLER_6_539 ();
 b15zdnd00an1n01x5 FILLER_6_543 ();
 b15zdnd11an1n16x5 FILLER_6_548 ();
 b15zdnd00an1n02x5 FILLER_6_564 ();
 b15zdnd11an1n04x5 FILLER_6_575 ();
 b15zdnd11an1n16x5 FILLER_6_585 ();
 b15zdnd11an1n04x5 FILLER_6_601 ();
 b15zdnd00an1n02x5 FILLER_6_605 ();
 b15zdnd11an1n04x5 FILLER_6_612 ();
 b15zdnd11an1n32x5 FILLER_6_626 ();
 b15zdnd11an1n16x5 FILLER_6_658 ();
 b15zdnd11an1n04x5 FILLER_6_674 ();
 b15zdnd00an1n02x5 FILLER_6_678 ();
 b15zdnd11an1n16x5 FILLER_6_692 ();
 b15zdnd11an1n08x5 FILLER_6_708 ();
 b15zdnd00an1n02x5 FILLER_6_716 ();
 b15zdnd00an1n02x5 FILLER_6_726 ();
 b15zdnd00an1n01x5 FILLER_6_728 ();
 b15zdnd11an1n04x5 FILLER_6_734 ();
 b15zdnd11an1n32x5 FILLER_6_744 ();
 b15zdnd11an1n08x5 FILLER_6_776 ();
 b15zdnd11an1n04x5 FILLER_6_784 ();
 b15zdnd00an1n02x5 FILLER_6_788 ();
 b15zdnd00an1n01x5 FILLER_6_790 ();
 b15zdnd11an1n08x5 FILLER_6_803 ();
 b15zdnd11an1n04x5 FILLER_6_811 ();
 b15zdnd11an1n64x5 FILLER_6_820 ();
 b15zdnd11an1n32x5 FILLER_6_884 ();
 b15zdnd00an1n02x5 FILLER_6_916 ();
 b15zdnd00an1n01x5 FILLER_6_918 ();
 b15zdnd11an1n04x5 FILLER_6_924 ();
 b15zdnd11an1n64x5 FILLER_6_932 ();
 b15zdnd11an1n64x5 FILLER_6_996 ();
 b15zdnd11an1n16x5 FILLER_6_1060 ();
 b15zdnd11an1n08x5 FILLER_6_1076 ();
 b15zdnd00an1n02x5 FILLER_6_1084 ();
 b15zdnd11an1n08x5 FILLER_6_1106 ();
 b15zdnd00an1n01x5 FILLER_6_1114 ();
 b15zdnd11an1n16x5 FILLER_6_1120 ();
 b15zdnd11an1n08x5 FILLER_6_1136 ();
 b15zdnd00an1n01x5 FILLER_6_1144 ();
 b15zdnd11an1n64x5 FILLER_6_1165 ();
 b15zdnd11an1n64x5 FILLER_6_1229 ();
 b15zdnd11an1n08x5 FILLER_6_1293 ();
 b15zdnd11an1n04x5 FILLER_6_1301 ();
 b15zdnd00an1n01x5 FILLER_6_1305 ();
 b15zdnd11an1n64x5 FILLER_6_1326 ();
 b15zdnd00an1n02x5 FILLER_6_1390 ();
 b15zdnd11an1n64x5 FILLER_6_1412 ();
 b15zdnd11an1n04x5 FILLER_6_1476 ();
 b15zdnd11an1n16x5 FILLER_6_1483 ();
 b15zdnd11an1n04x5 FILLER_6_1499 ();
 b15zdnd00an1n02x5 FILLER_6_1503 ();
 b15zdnd11an1n08x5 FILLER_6_1510 ();
 b15zdnd11an1n16x5 FILLER_6_1521 ();
 b15zdnd11an1n04x5 FILLER_6_1537 ();
 b15zdnd00an1n02x5 FILLER_6_1541 ();
 b15zdnd00an1n01x5 FILLER_6_1543 ();
 b15zdnd11an1n04x5 FILLER_6_1564 ();
 b15zdnd11an1n64x5 FILLER_6_1588 ();
 b15zdnd11an1n64x5 FILLER_6_1652 ();
 b15zdnd11an1n32x5 FILLER_6_1716 ();
 b15zdnd11an1n16x5 FILLER_6_1748 ();
 b15zdnd11an1n04x5 FILLER_6_1764 ();
 b15zdnd11an1n16x5 FILLER_6_1778 ();
 b15zdnd00an1n02x5 FILLER_6_1794 ();
 b15zdnd00an1n01x5 FILLER_6_1796 ();
 b15zdnd11an1n08x5 FILLER_6_1810 ();
 b15zdnd00an1n02x5 FILLER_6_1818 ();
 b15zdnd00an1n01x5 FILLER_6_1820 ();
 b15zdnd11an1n16x5 FILLER_6_1828 ();
 b15zdnd11an1n04x5 FILLER_6_1844 ();
 b15zdnd00an1n01x5 FILLER_6_1848 ();
 b15zdnd11an1n04x5 FILLER_6_1853 ();
 b15zdnd11an1n64x5 FILLER_6_1873 ();
 b15zdnd11an1n64x5 FILLER_6_1937 ();
 b15zdnd11an1n08x5 FILLER_6_2001 ();
 b15zdnd11an1n64x5 FILLER_6_2014 ();
 b15zdnd11an1n32x5 FILLER_6_2078 ();
 b15zdnd11an1n08x5 FILLER_6_2110 ();
 b15zdnd00an1n01x5 FILLER_6_2118 ();
 b15zdnd11an1n16x5 FILLER_6_2133 ();
 b15zdnd11an1n04x5 FILLER_6_2149 ();
 b15zdnd00an1n01x5 FILLER_6_2153 ();
 b15zdnd11an1n64x5 FILLER_6_2162 ();
 b15zdnd11an1n32x5 FILLER_6_2226 ();
 b15zdnd11an1n16x5 FILLER_6_2258 ();
 b15zdnd00an1n02x5 FILLER_6_2274 ();
 b15zdnd11an1n64x5 FILLER_7_0 ();
 b15zdnd11an1n64x5 FILLER_7_64 ();
 b15zdnd11an1n64x5 FILLER_7_128 ();
 b15zdnd11an1n64x5 FILLER_7_192 ();
 b15zdnd11an1n64x5 FILLER_7_256 ();
 b15zdnd11an1n64x5 FILLER_7_320 ();
 b15zdnd11an1n08x5 FILLER_7_384 ();
 b15zdnd11an1n04x5 FILLER_7_392 ();
 b15zdnd00an1n02x5 FILLER_7_396 ();
 b15zdnd00an1n01x5 FILLER_7_398 ();
 b15zdnd11an1n32x5 FILLER_7_408 ();
 b15zdnd11an1n16x5 FILLER_7_440 ();
 b15zdnd11an1n04x5 FILLER_7_456 ();
 b15zdnd00an1n01x5 FILLER_7_460 ();
 b15zdnd11an1n08x5 FILLER_7_477 ();
 b15zdnd11an1n04x5 FILLER_7_485 ();
 b15zdnd11an1n16x5 FILLER_7_494 ();
 b15zdnd11an1n08x5 FILLER_7_510 ();
 b15zdnd00an1n02x5 FILLER_7_518 ();
 b15zdnd11an1n04x5 FILLER_7_526 ();
 b15zdnd11an1n32x5 FILLER_7_536 ();
 b15zdnd11an1n08x5 FILLER_7_568 ();
 b15zdnd00an1n01x5 FILLER_7_576 ();
 b15zdnd11an1n04x5 FILLER_7_589 ();
 b15zdnd11an1n32x5 FILLER_7_598 ();
 b15zdnd11an1n08x5 FILLER_7_630 ();
 b15zdnd00an1n02x5 FILLER_7_638 ();
 b15zdnd11an1n64x5 FILLER_7_666 ();
 b15zdnd11an1n32x5 FILLER_7_730 ();
 b15zdnd11an1n08x5 FILLER_7_762 ();
 b15zdnd11an1n32x5 FILLER_7_778 ();
 b15zdnd11an1n04x5 FILLER_7_810 ();
 b15zdnd00an1n02x5 FILLER_7_814 ();
 b15zdnd00an1n01x5 FILLER_7_816 ();
 b15zdnd11an1n08x5 FILLER_7_824 ();
 b15zdnd00an1n01x5 FILLER_7_832 ();
 b15zdnd11an1n04x5 FILLER_7_864 ();
 b15zdnd11an1n64x5 FILLER_7_891 ();
 b15zdnd11an1n16x5 FILLER_7_955 ();
 b15zdnd11an1n08x5 FILLER_7_971 ();
 b15zdnd11an1n04x5 FILLER_7_979 ();
 b15zdnd00an1n02x5 FILLER_7_983 ();
 b15zdnd11an1n64x5 FILLER_7_990 ();
 b15zdnd11an1n64x5 FILLER_7_1054 ();
 b15zdnd11an1n32x5 FILLER_7_1118 ();
 b15zdnd00an1n02x5 FILLER_7_1150 ();
 b15zdnd11an1n64x5 FILLER_7_1172 ();
 b15zdnd11an1n32x5 FILLER_7_1236 ();
 b15zdnd11an1n16x5 FILLER_7_1268 ();
 b15zdnd11an1n08x5 FILLER_7_1284 ();
 b15zdnd11an1n04x5 FILLER_7_1292 ();
 b15zdnd00an1n02x5 FILLER_7_1296 ();
 b15zdnd00an1n01x5 FILLER_7_1298 ();
 b15zdnd11an1n64x5 FILLER_7_1319 ();
 b15zdnd11an1n16x5 FILLER_7_1383 ();
 b15zdnd11an1n04x5 FILLER_7_1399 ();
 b15zdnd11an1n64x5 FILLER_7_1409 ();
 b15zdnd11an1n16x5 FILLER_7_1473 ();
 b15zdnd11an1n08x5 FILLER_7_1489 ();
 b15zdnd11an1n04x5 FILLER_7_1497 ();
 b15zdnd11an1n64x5 FILLER_7_1521 ();
 b15zdnd11an1n64x5 FILLER_7_1585 ();
 b15zdnd11an1n64x5 FILLER_7_1649 ();
 b15zdnd11an1n32x5 FILLER_7_1713 ();
 b15zdnd11an1n16x5 FILLER_7_1745 ();
 b15zdnd11an1n04x5 FILLER_7_1761 ();
 b15zdnd00an1n02x5 FILLER_7_1765 ();
 b15zdnd00an1n01x5 FILLER_7_1767 ();
 b15zdnd11an1n16x5 FILLER_7_1789 ();
 b15zdnd11an1n08x5 FILLER_7_1805 ();
 b15zdnd11an1n04x5 FILLER_7_1813 ();
 b15zdnd00an1n02x5 FILLER_7_1817 ();
 b15zdnd11an1n64x5 FILLER_7_1827 ();
 b15zdnd00an1n01x5 FILLER_7_1891 ();
 b15zdnd11an1n64x5 FILLER_7_1898 ();
 b15zdnd11an1n64x5 FILLER_7_1962 ();
 b15zdnd11an1n08x5 FILLER_7_2026 ();
 b15zdnd00an1n01x5 FILLER_7_2034 ();
 b15zdnd11an1n64x5 FILLER_7_2053 ();
 b15zdnd11an1n16x5 FILLER_7_2117 ();
 b15zdnd11an1n04x5 FILLER_7_2133 ();
 b15zdnd11an1n64x5 FILLER_7_2160 ();
 b15zdnd11an1n32x5 FILLER_7_2224 ();
 b15zdnd11an1n16x5 FILLER_7_2256 ();
 b15zdnd11an1n08x5 FILLER_7_2272 ();
 b15zdnd11an1n04x5 FILLER_7_2280 ();
 b15zdnd11an1n64x5 FILLER_8_8 ();
 b15zdnd11an1n64x5 FILLER_8_72 ();
 b15zdnd11an1n64x5 FILLER_8_136 ();
 b15zdnd11an1n64x5 FILLER_8_200 ();
 b15zdnd11an1n64x5 FILLER_8_264 ();
 b15zdnd11an1n64x5 FILLER_8_328 ();
 b15zdnd11an1n08x5 FILLER_8_392 ();
 b15zdnd00an1n02x5 FILLER_8_400 ();
 b15zdnd00an1n01x5 FILLER_8_402 ();
 b15zdnd11an1n04x5 FILLER_8_409 ();
 b15zdnd00an1n01x5 FILLER_8_413 ();
 b15zdnd11an1n64x5 FILLER_8_435 ();
 b15zdnd11an1n16x5 FILLER_8_499 ();
 b15zdnd11an1n04x5 FILLER_8_515 ();
 b15zdnd00an1n02x5 FILLER_8_519 ();
 b15zdnd00an1n01x5 FILLER_8_521 ();
 b15zdnd11an1n32x5 FILLER_8_529 ();
 b15zdnd11an1n32x5 FILLER_8_577 ();
 b15zdnd11an1n04x5 FILLER_8_609 ();
 b15zdnd00an1n02x5 FILLER_8_613 ();
 b15zdnd00an1n01x5 FILLER_8_615 ();
 b15zdnd11an1n32x5 FILLER_8_622 ();
 b15zdnd11an1n08x5 FILLER_8_654 ();
 b15zdnd11an1n04x5 FILLER_8_662 ();
 b15zdnd00an1n02x5 FILLER_8_666 ();
 b15zdnd00an1n01x5 FILLER_8_668 ();
 b15zdnd11an1n32x5 FILLER_8_675 ();
 b15zdnd11an1n08x5 FILLER_8_707 ();
 b15zdnd00an1n02x5 FILLER_8_715 ();
 b15zdnd00an1n01x5 FILLER_8_717 ();
 b15zdnd11an1n32x5 FILLER_8_726 ();
 b15zdnd11an1n08x5 FILLER_8_758 ();
 b15zdnd11an1n32x5 FILLER_8_773 ();
 b15zdnd11an1n08x5 FILLER_8_805 ();
 b15zdnd00an1n01x5 FILLER_8_813 ();
 b15zdnd11an1n08x5 FILLER_8_827 ();
 b15zdnd11an1n04x5 FILLER_8_835 ();
 b15zdnd00an1n01x5 FILLER_8_839 ();
 b15zdnd11an1n64x5 FILLER_8_852 ();
 b15zdnd11an1n32x5 FILLER_8_916 ();
 b15zdnd11an1n16x5 FILLER_8_948 ();
 b15zdnd11an1n08x5 FILLER_8_964 ();
 b15zdnd11an1n04x5 FILLER_8_972 ();
 b15zdnd11an1n16x5 FILLER_8_996 ();
 b15zdnd11an1n08x5 FILLER_8_1012 ();
 b15zdnd00an1n02x5 FILLER_8_1020 ();
 b15zdnd11an1n64x5 FILLER_8_1042 ();
 b15zdnd11an1n64x5 FILLER_8_1106 ();
 b15zdnd11an1n64x5 FILLER_8_1170 ();
 b15zdnd11an1n32x5 FILLER_8_1234 ();
 b15zdnd11an1n08x5 FILLER_8_1266 ();
 b15zdnd11an1n04x5 FILLER_8_1274 ();
 b15zdnd11an1n16x5 FILLER_8_1282 ();
 b15zdnd11an1n08x5 FILLER_8_1298 ();
 b15zdnd00an1n02x5 FILLER_8_1306 ();
 b15zdnd11an1n64x5 FILLER_8_1328 ();
 b15zdnd11an1n64x5 FILLER_8_1392 ();
 b15zdnd11an1n64x5 FILLER_8_1456 ();
 b15zdnd11an1n64x5 FILLER_8_1520 ();
 b15zdnd11an1n64x5 FILLER_8_1584 ();
 b15zdnd11an1n64x5 FILLER_8_1648 ();
 b15zdnd11an1n32x5 FILLER_8_1712 ();
 b15zdnd11an1n16x5 FILLER_8_1744 ();
 b15zdnd11an1n08x5 FILLER_8_1760 ();
 b15zdnd11an1n16x5 FILLER_8_1780 ();
 b15zdnd00an1n02x5 FILLER_8_1796 ();
 b15zdnd11an1n04x5 FILLER_8_1812 ();
 b15zdnd11an1n08x5 FILLER_8_1826 ();
 b15zdnd11an1n04x5 FILLER_8_1834 ();
 b15zdnd00an1n01x5 FILLER_8_1838 ();
 b15zdnd11an1n64x5 FILLER_8_1843 ();
 b15zdnd11an1n08x5 FILLER_8_1907 ();
 b15zdnd11an1n04x5 FILLER_8_1915 ();
 b15zdnd00an1n02x5 FILLER_8_1919 ();
 b15zdnd00an1n01x5 FILLER_8_1921 ();
 b15zdnd11an1n04x5 FILLER_8_1929 ();
 b15zdnd11an1n64x5 FILLER_8_1947 ();
 b15zdnd11an1n64x5 FILLER_8_2011 ();
 b15zdnd11an1n16x5 FILLER_8_2075 ();
 b15zdnd11an1n04x5 FILLER_8_2091 ();
 b15zdnd00an1n02x5 FILLER_8_2095 ();
 b15zdnd00an1n01x5 FILLER_8_2097 ();
 b15zdnd11an1n08x5 FILLER_8_2115 ();
 b15zdnd11an1n04x5 FILLER_8_2123 ();
 b15zdnd00an1n02x5 FILLER_8_2127 ();
 b15zdnd00an1n01x5 FILLER_8_2129 ();
 b15zdnd11an1n08x5 FILLER_8_2146 ();
 b15zdnd11an1n16x5 FILLER_8_2162 ();
 b15zdnd11an1n08x5 FILLER_8_2178 ();
 b15zdnd00an1n01x5 FILLER_8_2186 ();
 b15zdnd11an1n04x5 FILLER_8_2203 ();
 b15zdnd11an1n32x5 FILLER_8_2225 ();
 b15zdnd11an1n16x5 FILLER_8_2257 ();
 b15zdnd00an1n02x5 FILLER_8_2273 ();
 b15zdnd00an1n01x5 FILLER_8_2275 ();
 b15zdnd11an1n64x5 FILLER_9_0 ();
 b15zdnd11an1n64x5 FILLER_9_64 ();
 b15zdnd11an1n64x5 FILLER_9_128 ();
 b15zdnd11an1n64x5 FILLER_9_192 ();
 b15zdnd11an1n64x5 FILLER_9_256 ();
 b15zdnd11an1n64x5 FILLER_9_320 ();
 b15zdnd11an1n16x5 FILLER_9_384 ();
 b15zdnd00an1n02x5 FILLER_9_400 ();
 b15zdnd00an1n01x5 FILLER_9_402 ();
 b15zdnd11an1n08x5 FILLER_9_417 ();
 b15zdnd11an1n04x5 FILLER_9_425 ();
 b15zdnd11an1n32x5 FILLER_9_433 ();
 b15zdnd00an1n02x5 FILLER_9_465 ();
 b15zdnd00an1n01x5 FILLER_9_467 ();
 b15zdnd11an1n16x5 FILLER_9_478 ();
 b15zdnd00an1n02x5 FILLER_9_494 ();
 b15zdnd11an1n16x5 FILLER_9_506 ();
 b15zdnd00an1n02x5 FILLER_9_522 ();
 b15zdnd11an1n64x5 FILLER_9_533 ();
 b15zdnd11an1n16x5 FILLER_9_597 ();
 b15zdnd11an1n04x5 FILLER_9_613 ();
 b15zdnd00an1n02x5 FILLER_9_617 ();
 b15zdnd11an1n04x5 FILLER_9_625 ();
 b15zdnd00an1n01x5 FILLER_9_629 ();
 b15zdnd11an1n64x5 FILLER_9_646 ();
 b15zdnd11an1n32x5 FILLER_9_710 ();
 b15zdnd11an1n16x5 FILLER_9_742 ();
 b15zdnd11an1n04x5 FILLER_9_758 ();
 b15zdnd00an1n02x5 FILLER_9_762 ();
 b15zdnd11an1n08x5 FILLER_9_774 ();
 b15zdnd11an1n04x5 FILLER_9_782 ();
 b15zdnd11an1n16x5 FILLER_9_794 ();
 b15zdnd00an1n02x5 FILLER_9_810 ();
 b15zdnd00an1n01x5 FILLER_9_812 ();
 b15zdnd11an1n32x5 FILLER_9_817 ();
 b15zdnd11an1n16x5 FILLER_9_849 ();
 b15zdnd11an1n08x5 FILLER_9_865 ();
 b15zdnd11an1n04x5 FILLER_9_873 ();
 b15zdnd11an1n04x5 FILLER_9_895 ();
 b15zdnd11an1n32x5 FILLER_9_915 ();
 b15zdnd11an1n04x5 FILLER_9_947 ();
 b15zdnd11an1n32x5 FILLER_9_955 ();
 b15zdnd00an1n02x5 FILLER_9_987 ();
 b15zdnd00an1n01x5 FILLER_9_989 ();
 b15zdnd11an1n32x5 FILLER_9_995 ();
 b15zdnd11an1n16x5 FILLER_9_1027 ();
 b15zdnd11an1n08x5 FILLER_9_1043 ();
 b15zdnd11an1n04x5 FILLER_9_1051 ();
 b15zdnd00an1n01x5 FILLER_9_1055 ();
 b15zdnd11an1n64x5 FILLER_9_1060 ();
 b15zdnd11an1n16x5 FILLER_9_1124 ();
 b15zdnd11an1n08x5 FILLER_9_1140 ();
 b15zdnd11an1n64x5 FILLER_9_1152 ();
 b15zdnd11an1n04x5 FILLER_9_1216 ();
 b15zdnd00an1n01x5 FILLER_9_1220 ();
 b15zdnd11an1n64x5 FILLER_9_1232 ();
 b15zdnd11an1n64x5 FILLER_9_1296 ();
 b15zdnd11an1n64x5 FILLER_9_1360 ();
 b15zdnd11an1n16x5 FILLER_9_1424 ();
 b15zdnd00an1n02x5 FILLER_9_1440 ();
 b15zdnd00an1n01x5 FILLER_9_1442 ();
 b15zdnd11an1n64x5 FILLER_9_1463 ();
 b15zdnd11an1n32x5 FILLER_9_1527 ();
 b15zdnd11an1n16x5 FILLER_9_1559 ();
 b15zdnd11an1n08x5 FILLER_9_1575 ();
 b15zdnd11an1n04x5 FILLER_9_1583 ();
 b15zdnd00an1n02x5 FILLER_9_1587 ();
 b15zdnd11an1n64x5 FILLER_9_1609 ();
 b15zdnd11an1n16x5 FILLER_9_1673 ();
 b15zdnd11an1n04x5 FILLER_9_1689 ();
 b15zdnd11an1n32x5 FILLER_9_1713 ();
 b15zdnd11an1n04x5 FILLER_9_1745 ();
 b15zdnd11an1n04x5 FILLER_9_1765 ();
 b15zdnd11an1n08x5 FILLER_9_1778 ();
 b15zdnd11an1n08x5 FILLER_9_1806 ();
 b15zdnd00an1n02x5 FILLER_9_1814 ();
 b15zdnd00an1n01x5 FILLER_9_1816 ();
 b15zdnd11an1n04x5 FILLER_9_1835 ();
 b15zdnd00an1n01x5 FILLER_9_1839 ();
 b15zdnd11an1n64x5 FILLER_9_1852 ();
 b15zdnd11an1n32x5 FILLER_9_1916 ();
 b15zdnd11an1n04x5 FILLER_9_1948 ();
 b15zdnd11an1n04x5 FILLER_9_1958 ();
 b15zdnd11an1n04x5 FILLER_9_1968 ();
 b15zdnd11an1n16x5 FILLER_9_1982 ();
 b15zdnd11an1n08x5 FILLER_9_1998 ();
 b15zdnd11an1n04x5 FILLER_9_2006 ();
 b15zdnd00an1n02x5 FILLER_9_2010 ();
 b15zdnd11an1n16x5 FILLER_9_2019 ();
 b15zdnd11an1n08x5 FILLER_9_2035 ();
 b15zdnd11an1n64x5 FILLER_9_2049 ();
 b15zdnd11an1n16x5 FILLER_9_2113 ();
 b15zdnd11an1n64x5 FILLER_9_2138 ();
 b15zdnd11an1n64x5 FILLER_9_2202 ();
 b15zdnd11an1n16x5 FILLER_9_2266 ();
 b15zdnd00an1n02x5 FILLER_9_2282 ();
 b15zdnd11an1n64x5 FILLER_10_8 ();
 b15zdnd11an1n64x5 FILLER_10_72 ();
 b15zdnd11an1n64x5 FILLER_10_136 ();
 b15zdnd11an1n64x5 FILLER_10_200 ();
 b15zdnd11an1n64x5 FILLER_10_264 ();
 b15zdnd11an1n64x5 FILLER_10_328 ();
 b15zdnd11an1n08x5 FILLER_10_392 ();
 b15zdnd00an1n02x5 FILLER_10_400 ();
 b15zdnd11an1n04x5 FILLER_10_411 ();
 b15zdnd00an1n02x5 FILLER_10_415 ();
 b15zdnd00an1n01x5 FILLER_10_417 ();
 b15zdnd11an1n16x5 FILLER_10_438 ();
 b15zdnd11an1n08x5 FILLER_10_454 ();
 b15zdnd00an1n02x5 FILLER_10_462 ();
 b15zdnd11an1n64x5 FILLER_10_485 ();
 b15zdnd11an1n32x5 FILLER_10_549 ();
 b15zdnd11an1n16x5 FILLER_10_581 ();
 b15zdnd00an1n02x5 FILLER_10_597 ();
 b15zdnd11an1n32x5 FILLER_10_605 ();
 b15zdnd11an1n16x5 FILLER_10_637 ();
 b15zdnd11an1n08x5 FILLER_10_653 ();
 b15zdnd11an1n16x5 FILLER_10_668 ();
 b15zdnd11an1n08x5 FILLER_10_684 ();
 b15zdnd11an1n04x5 FILLER_10_692 ();
 b15zdnd00an1n01x5 FILLER_10_696 ();
 b15zdnd11an1n04x5 FILLER_10_713 ();
 b15zdnd00an1n01x5 FILLER_10_717 ();
 b15zdnd11an1n08x5 FILLER_10_726 ();
 b15zdnd11an1n04x5 FILLER_10_734 ();
 b15zdnd11an1n16x5 FILLER_10_748 ();
 b15zdnd11an1n08x5 FILLER_10_764 ();
 b15zdnd00an1n01x5 FILLER_10_772 ();
 b15zdnd11an1n08x5 FILLER_10_779 ();
 b15zdnd00an1n02x5 FILLER_10_787 ();
 b15zdnd00an1n01x5 FILLER_10_789 ();
 b15zdnd11an1n32x5 FILLER_10_806 ();
 b15zdnd00an1n02x5 FILLER_10_838 ();
 b15zdnd00an1n01x5 FILLER_10_840 ();
 b15zdnd11an1n64x5 FILLER_10_872 ();
 b15zdnd11an1n08x5 FILLER_10_936 ();
 b15zdnd00an1n02x5 FILLER_10_944 ();
 b15zdnd11an1n64x5 FILLER_10_951 ();
 b15zdnd11an1n32x5 FILLER_10_1015 ();
 b15zdnd11an1n04x5 FILLER_10_1047 ();
 b15zdnd11an1n64x5 FILLER_10_1056 ();
 b15zdnd11an1n64x5 FILLER_10_1120 ();
 b15zdnd11an1n04x5 FILLER_10_1184 ();
 b15zdnd00an1n01x5 FILLER_10_1188 ();
 b15zdnd11an1n16x5 FILLER_10_1195 ();
 b15zdnd11an1n08x5 FILLER_10_1211 ();
 b15zdnd11an1n04x5 FILLER_10_1219 ();
 b15zdnd00an1n02x5 FILLER_10_1223 ();
 b15zdnd11an1n16x5 FILLER_10_1245 ();
 b15zdnd11an1n08x5 FILLER_10_1261 ();
 b15zdnd11an1n04x5 FILLER_10_1269 ();
 b15zdnd11an1n64x5 FILLER_10_1278 ();
 b15zdnd11an1n64x5 FILLER_10_1342 ();
 b15zdnd11an1n16x5 FILLER_10_1406 ();
 b15zdnd11an1n08x5 FILLER_10_1422 ();
 b15zdnd11an1n04x5 FILLER_10_1430 ();
 b15zdnd00an1n02x5 FILLER_10_1434 ();
 b15zdnd00an1n01x5 FILLER_10_1436 ();
 b15zdnd11an1n32x5 FILLER_10_1449 ();
 b15zdnd11an1n16x5 FILLER_10_1481 ();
 b15zdnd11an1n04x5 FILLER_10_1497 ();
 b15zdnd11an1n04x5 FILLER_10_1514 ();
 b15zdnd11an1n08x5 FILLER_10_1527 ();
 b15zdnd00an1n02x5 FILLER_10_1535 ();
 b15zdnd00an1n01x5 FILLER_10_1537 ();
 b15zdnd11an1n16x5 FILLER_10_1549 ();
 b15zdnd11an1n04x5 FILLER_10_1565 ();
 b15zdnd00an1n02x5 FILLER_10_1569 ();
 b15zdnd11an1n16x5 FILLER_10_1580 ();
 b15zdnd00an1n01x5 FILLER_10_1596 ();
 b15zdnd11an1n16x5 FILLER_10_1615 ();
 b15zdnd11an1n08x5 FILLER_10_1631 ();
 b15zdnd11an1n04x5 FILLER_10_1639 ();
 b15zdnd11an1n08x5 FILLER_10_1652 ();
 b15zdnd00an1n01x5 FILLER_10_1660 ();
 b15zdnd11an1n16x5 FILLER_10_1681 ();
 b15zdnd11an1n04x5 FILLER_10_1697 ();
 b15zdnd00an1n02x5 FILLER_10_1701 ();
 b15zdnd11an1n08x5 FILLER_10_1723 ();
 b15zdnd00an1n01x5 FILLER_10_1731 ();
 b15zdnd11an1n04x5 FILLER_10_1758 ();
 b15zdnd00an1n02x5 FILLER_10_1762 ();
 b15zdnd00an1n01x5 FILLER_10_1764 ();
 b15zdnd11an1n16x5 FILLER_10_1788 ();
 b15zdnd11an1n08x5 FILLER_10_1804 ();
 b15zdnd11an1n04x5 FILLER_10_1812 ();
 b15zdnd00an1n02x5 FILLER_10_1816 ();
 b15zdnd00an1n01x5 FILLER_10_1818 ();
 b15zdnd11an1n08x5 FILLER_10_1845 ();
 b15zdnd11an1n04x5 FILLER_10_1853 ();
 b15zdnd00an1n02x5 FILLER_10_1857 ();
 b15zdnd11an1n32x5 FILLER_10_1868 ();
 b15zdnd11an1n08x5 FILLER_10_1906 ();
 b15zdnd11an1n04x5 FILLER_10_1914 ();
 b15zdnd00an1n02x5 FILLER_10_1918 ();
 b15zdnd00an1n01x5 FILLER_10_1920 ();
 b15zdnd11an1n08x5 FILLER_10_1930 ();
 b15zdnd00an1n02x5 FILLER_10_1938 ();
 b15zdnd11an1n04x5 FILLER_10_1950 ();
 b15zdnd00an1n02x5 FILLER_10_1954 ();
 b15zdnd11an1n04x5 FILLER_10_1963 ();
 b15zdnd11an1n08x5 FILLER_10_1980 ();
 b15zdnd00an1n02x5 FILLER_10_1988 ();
 b15zdnd00an1n01x5 FILLER_10_1990 ();
 b15zdnd11an1n04x5 FILLER_10_2014 ();
 b15zdnd11an1n08x5 FILLER_10_2034 ();
 b15zdnd11an1n04x5 FILLER_10_2042 ();
 b15zdnd00an1n02x5 FILLER_10_2046 ();
 b15zdnd00an1n01x5 FILLER_10_2048 ();
 b15zdnd11an1n04x5 FILLER_10_2054 ();
 b15zdnd11an1n16x5 FILLER_10_2065 ();
 b15zdnd00an1n01x5 FILLER_10_2081 ();
 b15zdnd11an1n64x5 FILLER_10_2089 ();
 b15zdnd00an1n01x5 FILLER_10_2153 ();
 b15zdnd00an1n02x5 FILLER_10_2162 ();
 b15zdnd11an1n04x5 FILLER_10_2184 ();
 b15zdnd11an1n04x5 FILLER_10_2201 ();
 b15zdnd11an1n32x5 FILLER_10_2223 ();
 b15zdnd11an1n16x5 FILLER_10_2255 ();
 b15zdnd11an1n04x5 FILLER_10_2271 ();
 b15zdnd00an1n01x5 FILLER_10_2275 ();
 b15zdnd11an1n64x5 FILLER_11_0 ();
 b15zdnd11an1n64x5 FILLER_11_64 ();
 b15zdnd11an1n64x5 FILLER_11_128 ();
 b15zdnd11an1n64x5 FILLER_11_192 ();
 b15zdnd11an1n64x5 FILLER_11_256 ();
 b15zdnd11an1n64x5 FILLER_11_320 ();
 b15zdnd11an1n64x5 FILLER_11_384 ();
 b15zdnd11an1n64x5 FILLER_11_448 ();
 b15zdnd11an1n16x5 FILLER_11_512 ();
 b15zdnd11an1n04x5 FILLER_11_528 ();
 b15zdnd11an1n16x5 FILLER_11_537 ();
 b15zdnd11an1n04x5 FILLER_11_553 ();
 b15zdnd00an1n02x5 FILLER_11_557 ();
 b15zdnd11an1n04x5 FILLER_11_571 ();
 b15zdnd00an1n02x5 FILLER_11_575 ();
 b15zdnd11an1n64x5 FILLER_11_584 ();
 b15zdnd11an1n04x5 FILLER_11_648 ();
 b15zdnd00an1n02x5 FILLER_11_652 ();
 b15zdnd00an1n01x5 FILLER_11_654 ();
 b15zdnd11an1n04x5 FILLER_11_660 ();
 b15zdnd11an1n16x5 FILLER_11_671 ();
 b15zdnd11an1n08x5 FILLER_11_687 ();
 b15zdnd11an1n04x5 FILLER_11_695 ();
 b15zdnd11an1n04x5 FILLER_11_704 ();
 b15zdnd11an1n08x5 FILLER_11_712 ();
 b15zdnd00an1n01x5 FILLER_11_720 ();
 b15zdnd11an1n08x5 FILLER_11_733 ();
 b15zdnd00an1n02x5 FILLER_11_741 ();
 b15zdnd11an1n08x5 FILLER_11_749 ();
 b15zdnd11an1n04x5 FILLER_11_757 ();
 b15zdnd11an1n64x5 FILLER_11_777 ();
 b15zdnd11an1n16x5 FILLER_11_841 ();
 b15zdnd11an1n08x5 FILLER_11_857 ();
 b15zdnd11an1n04x5 FILLER_11_865 ();
 b15zdnd00an1n02x5 FILLER_11_869 ();
 b15zdnd00an1n01x5 FILLER_11_871 ();
 b15zdnd11an1n04x5 FILLER_11_904 ();
 b15zdnd11an1n08x5 FILLER_11_928 ();
 b15zdnd00an1n02x5 FILLER_11_936 ();
 b15zdnd11an1n32x5 FILLER_11_958 ();
 b15zdnd11an1n16x5 FILLER_11_990 ();
 b15zdnd11an1n16x5 FILLER_11_1015 ();
 b15zdnd11an1n08x5 FILLER_11_1031 ();
 b15zdnd11an1n04x5 FILLER_11_1039 ();
 b15zdnd00an1n02x5 FILLER_11_1043 ();
 b15zdnd11an1n08x5 FILLER_11_1065 ();
 b15zdnd00an1n02x5 FILLER_11_1073 ();
 b15zdnd00an1n01x5 FILLER_11_1075 ();
 b15zdnd11an1n16x5 FILLER_11_1096 ();
 b15zdnd11an1n08x5 FILLER_11_1112 ();
 b15zdnd00an1n01x5 FILLER_11_1120 ();
 b15zdnd11an1n32x5 FILLER_11_1126 ();
 b15zdnd11an1n16x5 FILLER_11_1158 ();
 b15zdnd11an1n08x5 FILLER_11_1174 ();
 b15zdnd00an1n01x5 FILLER_11_1182 ();
 b15zdnd11an1n08x5 FILLER_11_1203 ();
 b15zdnd00an1n02x5 FILLER_11_1211 ();
 b15zdnd00an1n01x5 FILLER_11_1213 ();
 b15zdnd11an1n32x5 FILLER_11_1234 ();
 b15zdnd00an1n02x5 FILLER_11_1266 ();
 b15zdnd11an1n64x5 FILLER_11_1273 ();
 b15zdnd11an1n08x5 FILLER_11_1337 ();
 b15zdnd11an1n04x5 FILLER_11_1345 ();
 b15zdnd00an1n02x5 FILLER_11_1349 ();
 b15zdnd11an1n64x5 FILLER_11_1355 ();
 b15zdnd11an1n32x5 FILLER_11_1419 ();
 b15zdnd11an1n04x5 FILLER_11_1451 ();
 b15zdnd00an1n02x5 FILLER_11_1455 ();
 b15zdnd00an1n01x5 FILLER_11_1457 ();
 b15zdnd11an1n64x5 FILLER_11_1478 ();
 b15zdnd11an1n16x5 FILLER_11_1542 ();
 b15zdnd11an1n08x5 FILLER_11_1558 ();
 b15zdnd00an1n01x5 FILLER_11_1566 ();
 b15zdnd11an1n64x5 FILLER_11_1576 ();
 b15zdnd11an1n64x5 FILLER_11_1640 ();
 b15zdnd11an1n32x5 FILLER_11_1704 ();
 b15zdnd11an1n08x5 FILLER_11_1736 ();
 b15zdnd11an1n04x5 FILLER_11_1744 ();
 b15zdnd11an1n04x5 FILLER_11_1764 ();
 b15zdnd11an1n16x5 FILLER_11_1788 ();
 b15zdnd11an1n08x5 FILLER_11_1804 ();
 b15zdnd00an1n02x5 FILLER_11_1812 ();
 b15zdnd00an1n01x5 FILLER_11_1814 ();
 b15zdnd11an1n16x5 FILLER_11_1825 ();
 b15zdnd00an1n02x5 FILLER_11_1841 ();
 b15zdnd00an1n01x5 FILLER_11_1843 ();
 b15zdnd11an1n32x5 FILLER_11_1854 ();
 b15zdnd11an1n16x5 FILLER_11_1886 ();
 b15zdnd11an1n08x5 FILLER_11_1902 ();
 b15zdnd11an1n04x5 FILLER_11_1910 ();
 b15zdnd00an1n02x5 FILLER_11_1914 ();
 b15zdnd11an1n64x5 FILLER_11_1925 ();
 b15zdnd11an1n16x5 FILLER_11_1989 ();
 b15zdnd11an1n08x5 FILLER_11_2005 ();
 b15zdnd11an1n04x5 FILLER_11_2013 ();
 b15zdnd00an1n02x5 FILLER_11_2017 ();
 b15zdnd00an1n01x5 FILLER_11_2019 ();
 b15zdnd11an1n16x5 FILLER_11_2027 ();
 b15zdnd11an1n08x5 FILLER_11_2043 ();
 b15zdnd11an1n08x5 FILLER_11_2066 ();
 b15zdnd11an1n04x5 FILLER_11_2074 ();
 b15zdnd00an1n02x5 FILLER_11_2078 ();
 b15zdnd11an1n04x5 FILLER_11_2100 ();
 b15zdnd11an1n04x5 FILLER_11_2127 ();
 b15zdnd11an1n16x5 FILLER_11_2141 ();
 b15zdnd00an1n01x5 FILLER_11_2157 ();
 b15zdnd11an1n04x5 FILLER_11_2190 ();
 b15zdnd11an1n64x5 FILLER_11_2218 ();
 b15zdnd00an1n02x5 FILLER_11_2282 ();
 b15zdnd11an1n64x5 FILLER_12_8 ();
 b15zdnd11an1n64x5 FILLER_12_72 ();
 b15zdnd11an1n16x5 FILLER_12_136 ();
 b15zdnd00an1n02x5 FILLER_12_152 ();
 b15zdnd11an1n64x5 FILLER_12_159 ();
 b15zdnd11an1n64x5 FILLER_12_223 ();
 b15zdnd11an1n64x5 FILLER_12_287 ();
 b15zdnd11an1n64x5 FILLER_12_351 ();
 b15zdnd11an1n04x5 FILLER_12_415 ();
 b15zdnd00an1n01x5 FILLER_12_419 ();
 b15zdnd11an1n04x5 FILLER_12_434 ();
 b15zdnd11an1n16x5 FILLER_12_453 ();
 b15zdnd00an1n01x5 FILLER_12_469 ();
 b15zdnd11an1n08x5 FILLER_12_477 ();
 b15zdnd11an1n04x5 FILLER_12_485 ();
 b15zdnd00an1n02x5 FILLER_12_489 ();
 b15zdnd00an1n01x5 FILLER_12_491 ();
 b15zdnd11an1n04x5 FILLER_12_513 ();
 b15zdnd11an1n04x5 FILLER_12_527 ();
 b15zdnd11an1n16x5 FILLER_12_547 ();
 b15zdnd11an1n08x5 FILLER_12_563 ();
 b15zdnd00an1n01x5 FILLER_12_571 ();
 b15zdnd11an1n32x5 FILLER_12_585 ();
 b15zdnd11an1n16x5 FILLER_12_617 ();
 b15zdnd11an1n08x5 FILLER_12_633 ();
 b15zdnd11an1n04x5 FILLER_12_641 ();
 b15zdnd00an1n01x5 FILLER_12_645 ();
 b15zdnd11an1n32x5 FILLER_12_652 ();
 b15zdnd11an1n04x5 FILLER_12_700 ();
 b15zdnd11an1n08x5 FILLER_12_710 ();
 b15zdnd11an1n32x5 FILLER_12_726 ();
 b15zdnd11an1n04x5 FILLER_12_758 ();
 b15zdnd00an1n02x5 FILLER_12_762 ();
 b15zdnd00an1n01x5 FILLER_12_764 ();
 b15zdnd11an1n64x5 FILLER_12_778 ();
 b15zdnd11an1n32x5 FILLER_12_842 ();
 b15zdnd11an1n16x5 FILLER_12_874 ();
 b15zdnd00an1n02x5 FILLER_12_890 ();
 b15zdnd00an1n01x5 FILLER_12_892 ();
 b15zdnd11an1n04x5 FILLER_12_911 ();
 b15zdnd11an1n08x5 FILLER_12_941 ();
 b15zdnd00an1n02x5 FILLER_12_949 ();
 b15zdnd11an1n64x5 FILLER_12_955 ();
 b15zdnd11an1n32x5 FILLER_12_1019 ();
 b15zdnd11an1n08x5 FILLER_12_1051 ();
 b15zdnd11an1n16x5 FILLER_12_1063 ();
 b15zdnd11an1n08x5 FILLER_12_1079 ();
 b15zdnd11an1n04x5 FILLER_12_1087 ();
 b15zdnd11an1n04x5 FILLER_12_1111 ();
 b15zdnd11an1n04x5 FILLER_12_1135 ();
 b15zdnd11an1n16x5 FILLER_12_1148 ();
 b15zdnd00an1n02x5 FILLER_12_1164 ();
 b15zdnd11an1n04x5 FILLER_12_1186 ();
 b15zdnd11an1n16x5 FILLER_12_1195 ();
 b15zdnd11an1n08x5 FILLER_12_1211 ();
 b15zdnd11an1n04x5 FILLER_12_1219 ();
 b15zdnd11an1n32x5 FILLER_12_1232 ();
 b15zdnd11an1n04x5 FILLER_12_1264 ();
 b15zdnd00an1n01x5 FILLER_12_1268 ();
 b15zdnd11an1n64x5 FILLER_12_1289 ();
 b15zdnd11an1n16x5 FILLER_12_1353 ();
 b15zdnd11an1n04x5 FILLER_12_1369 ();
 b15zdnd11an1n04x5 FILLER_12_1393 ();
 b15zdnd00an1n02x5 FILLER_12_1397 ();
 b15zdnd00an1n01x5 FILLER_12_1399 ();
 b15zdnd11an1n32x5 FILLER_12_1420 ();
 b15zdnd11an1n16x5 FILLER_12_1452 ();
 b15zdnd11an1n04x5 FILLER_12_1468 ();
 b15zdnd00an1n02x5 FILLER_12_1472 ();
 b15zdnd11an1n64x5 FILLER_12_1496 ();
 b15zdnd11an1n64x5 FILLER_12_1560 ();
 b15zdnd11an1n32x5 FILLER_12_1624 ();
 b15zdnd11an1n04x5 FILLER_12_1656 ();
 b15zdnd00an1n02x5 FILLER_12_1660 ();
 b15zdnd00an1n01x5 FILLER_12_1662 ();
 b15zdnd11an1n04x5 FILLER_12_1672 ();
 b15zdnd00an1n02x5 FILLER_12_1676 ();
 b15zdnd00an1n01x5 FILLER_12_1678 ();
 b15zdnd11an1n64x5 FILLER_12_1699 ();
 b15zdnd11an1n16x5 FILLER_12_1763 ();
 b15zdnd11an1n08x5 FILLER_12_1779 ();
 b15zdnd11an1n04x5 FILLER_12_1792 ();
 b15zdnd11an1n32x5 FILLER_12_1804 ();
 b15zdnd11an1n04x5 FILLER_12_1836 ();
 b15zdnd00an1n02x5 FILLER_12_1840 ();
 b15zdnd00an1n01x5 FILLER_12_1842 ();
 b15zdnd11an1n32x5 FILLER_12_1856 ();
 b15zdnd11an1n08x5 FILLER_12_1888 ();
 b15zdnd11an1n04x5 FILLER_12_1896 ();
 b15zdnd00an1n02x5 FILLER_12_1900 ();
 b15zdnd11an1n04x5 FILLER_12_1909 ();
 b15zdnd11an1n16x5 FILLER_12_1919 ();
 b15zdnd11an1n64x5 FILLER_12_1949 ();
 b15zdnd11an1n32x5 FILLER_12_2013 ();
 b15zdnd11an1n16x5 FILLER_12_2045 ();
 b15zdnd00an1n02x5 FILLER_12_2061 ();
 b15zdnd11an1n32x5 FILLER_12_2067 ();
 b15zdnd11an1n16x5 FILLER_12_2099 ();
 b15zdnd11an1n08x5 FILLER_12_2115 ();
 b15zdnd11an1n04x5 FILLER_12_2123 ();
 b15zdnd00an1n02x5 FILLER_12_2151 ();
 b15zdnd00an1n01x5 FILLER_12_2153 ();
 b15zdnd11an1n32x5 FILLER_12_2162 ();
 b15zdnd11an1n04x5 FILLER_12_2194 ();
 b15zdnd11an1n32x5 FILLER_12_2216 ();
 b15zdnd11an1n16x5 FILLER_12_2248 ();
 b15zdnd11an1n08x5 FILLER_12_2264 ();
 b15zdnd11an1n04x5 FILLER_12_2272 ();
 b15zdnd11an1n64x5 FILLER_13_0 ();
 b15zdnd11an1n32x5 FILLER_13_64 ();
 b15zdnd11an1n16x5 FILLER_13_96 ();
 b15zdnd11an1n04x5 FILLER_13_112 ();
 b15zdnd00an1n01x5 FILLER_13_116 ();
 b15zdnd11an1n04x5 FILLER_13_126 ();
 b15zdnd00an1n02x5 FILLER_13_130 ();
 b15zdnd11an1n04x5 FILLER_13_137 ();
 b15zdnd00an1n01x5 FILLER_13_141 ();
 b15zdnd11an1n04x5 FILLER_13_148 ();
 b15zdnd00an1n02x5 FILLER_13_152 ();
 b15zdnd11an1n64x5 FILLER_13_169 ();
 b15zdnd11an1n64x5 FILLER_13_233 ();
 b15zdnd11an1n64x5 FILLER_13_297 ();
 b15zdnd11an1n64x5 FILLER_13_361 ();
 b15zdnd00an1n01x5 FILLER_13_425 ();
 b15zdnd11an1n32x5 FILLER_13_446 ();
 b15zdnd11an1n16x5 FILLER_13_478 ();
 b15zdnd00an1n02x5 FILLER_13_494 ();
 b15zdnd00an1n01x5 FILLER_13_496 ();
 b15zdnd11an1n32x5 FILLER_13_521 ();
 b15zdnd11an1n16x5 FILLER_13_553 ();
 b15zdnd11an1n08x5 FILLER_13_569 ();
 b15zdnd11an1n04x5 FILLER_13_577 ();
 b15zdnd00an1n02x5 FILLER_13_581 ();
 b15zdnd00an1n01x5 FILLER_13_583 ();
 b15zdnd11an1n16x5 FILLER_13_592 ();
 b15zdnd11an1n08x5 FILLER_13_608 ();
 b15zdnd11an1n04x5 FILLER_13_616 ();
 b15zdnd11an1n04x5 FILLER_13_627 ();
 b15zdnd11an1n04x5 FILLER_13_635 ();
 b15zdnd11an1n04x5 FILLER_13_651 ();
 b15zdnd11an1n32x5 FILLER_13_681 ();
 b15zdnd11an1n08x5 FILLER_13_713 ();
 b15zdnd11an1n04x5 FILLER_13_721 ();
 b15zdnd11an1n64x5 FILLER_13_731 ();
 b15zdnd00an1n02x5 FILLER_13_795 ();
 b15zdnd11an1n16x5 FILLER_13_801 ();
 b15zdnd11an1n08x5 FILLER_13_817 ();
 b15zdnd11an1n04x5 FILLER_13_825 ();
 b15zdnd00an1n02x5 FILLER_13_829 ();
 b15zdnd11an1n08x5 FILLER_13_840 ();
 b15zdnd00an1n02x5 FILLER_13_848 ();
 b15zdnd00an1n01x5 FILLER_13_850 ();
 b15zdnd11an1n16x5 FILLER_13_871 ();
 b15zdnd00an1n02x5 FILLER_13_887 ();
 b15zdnd11an1n64x5 FILLER_13_905 ();
 b15zdnd11an1n08x5 FILLER_13_969 ();
 b15zdnd11an1n04x5 FILLER_13_977 ();
 b15zdnd00an1n02x5 FILLER_13_981 ();
 b15zdnd00an1n01x5 FILLER_13_983 ();
 b15zdnd11an1n04x5 FILLER_13_1004 ();
 b15zdnd11an1n64x5 FILLER_13_1020 ();
 b15zdnd11an1n32x5 FILLER_13_1084 ();
 b15zdnd11an1n08x5 FILLER_13_1116 ();
 b15zdnd00an1n02x5 FILLER_13_1124 ();
 b15zdnd11an1n32x5 FILLER_13_1130 ();
 b15zdnd11an1n16x5 FILLER_13_1162 ();
 b15zdnd11an1n04x5 FILLER_13_1178 ();
 b15zdnd00an1n02x5 FILLER_13_1182 ();
 b15zdnd00an1n01x5 FILLER_13_1184 ();
 b15zdnd11an1n64x5 FILLER_13_1193 ();
 b15zdnd11an1n32x5 FILLER_13_1257 ();
 b15zdnd11an1n08x5 FILLER_13_1289 ();
 b15zdnd00an1n02x5 FILLER_13_1297 ();
 b15zdnd00an1n01x5 FILLER_13_1299 ();
 b15zdnd11an1n32x5 FILLER_13_1306 ();
 b15zdnd11an1n64x5 FILLER_13_1343 ();
 b15zdnd11an1n32x5 FILLER_13_1407 ();
 b15zdnd00an1n02x5 FILLER_13_1439 ();
 b15zdnd00an1n01x5 FILLER_13_1441 ();
 b15zdnd11an1n04x5 FILLER_13_1453 ();
 b15zdnd11an1n64x5 FILLER_13_1466 ();
 b15zdnd11an1n64x5 FILLER_13_1530 ();
 b15zdnd11an1n64x5 FILLER_13_1594 ();
 b15zdnd11an1n64x5 FILLER_13_1658 ();
 b15zdnd11an1n16x5 FILLER_13_1722 ();
 b15zdnd11an1n04x5 FILLER_13_1738 ();
 b15zdnd11an1n08x5 FILLER_13_1755 ();
 b15zdnd11an1n04x5 FILLER_13_1763 ();
 b15zdnd00an1n02x5 FILLER_13_1767 ();
 b15zdnd11an1n08x5 FILLER_13_1779 ();
 b15zdnd11an1n04x5 FILLER_13_1787 ();
 b15zdnd00an1n01x5 FILLER_13_1791 ();
 b15zdnd11an1n08x5 FILLER_13_1797 ();
 b15zdnd11an1n04x5 FILLER_13_1805 ();
 b15zdnd00an1n01x5 FILLER_13_1809 ();
 b15zdnd11an1n04x5 FILLER_13_1816 ();
 b15zdnd11an1n16x5 FILLER_13_1826 ();
 b15zdnd11an1n04x5 FILLER_13_1842 ();
 b15zdnd11an1n32x5 FILLER_13_1852 ();
 b15zdnd11an1n16x5 FILLER_13_1884 ();
 b15zdnd11an1n04x5 FILLER_13_1905 ();
 b15zdnd00an1n02x5 FILLER_13_1909 ();
 b15zdnd00an1n01x5 FILLER_13_1911 ();
 b15zdnd11an1n08x5 FILLER_13_1922 ();
 b15zdnd11an1n04x5 FILLER_13_1930 ();
 b15zdnd00an1n02x5 FILLER_13_1934 ();
 b15zdnd11an1n32x5 FILLER_13_1942 ();
 b15zdnd11an1n04x5 FILLER_13_1974 ();
 b15zdnd00an1n02x5 FILLER_13_1978 ();
 b15zdnd11an1n16x5 FILLER_13_1985 ();
 b15zdnd11an1n08x5 FILLER_13_2001 ();
 b15zdnd11an1n04x5 FILLER_13_2009 ();
 b15zdnd00an1n02x5 FILLER_13_2013 ();
 b15zdnd11an1n64x5 FILLER_13_2021 ();
 b15zdnd11an1n32x5 FILLER_13_2085 ();
 b15zdnd11an1n08x5 FILLER_13_2117 ();
 b15zdnd00an1n02x5 FILLER_13_2125 ();
 b15zdnd11an1n16x5 FILLER_13_2142 ();
 b15zdnd11an1n08x5 FILLER_13_2158 ();
 b15zdnd11an1n64x5 FILLER_13_2198 ();
 b15zdnd11an1n16x5 FILLER_13_2262 ();
 b15zdnd11an1n04x5 FILLER_13_2278 ();
 b15zdnd00an1n02x5 FILLER_13_2282 ();
 b15zdnd11an1n64x5 FILLER_14_8 ();
 b15zdnd11an1n32x5 FILLER_14_72 ();
 b15zdnd11an1n16x5 FILLER_14_104 ();
 b15zdnd00an1n02x5 FILLER_14_120 ();
 b15zdnd11an1n08x5 FILLER_14_140 ();
 b15zdnd00an1n02x5 FILLER_14_148 ();
 b15zdnd00an1n01x5 FILLER_14_150 ();
 b15zdnd11an1n16x5 FILLER_14_158 ();
 b15zdnd11an1n08x5 FILLER_14_174 ();
 b15zdnd11an1n04x5 FILLER_14_182 ();
 b15zdnd00an1n02x5 FILLER_14_186 ();
 b15zdnd00an1n01x5 FILLER_14_188 ();
 b15zdnd11an1n04x5 FILLER_14_198 ();
 b15zdnd11an1n08x5 FILLER_14_208 ();
 b15zdnd11an1n04x5 FILLER_14_216 ();
 b15zdnd00an1n02x5 FILLER_14_220 ();
 b15zdnd11an1n64x5 FILLER_14_234 ();
 b15zdnd11an1n64x5 FILLER_14_298 ();
 b15zdnd11an1n32x5 FILLER_14_362 ();
 b15zdnd11an1n08x5 FILLER_14_394 ();
 b15zdnd11an1n04x5 FILLER_14_402 ();
 b15zdnd00an1n02x5 FILLER_14_406 ();
 b15zdnd11an1n32x5 FILLER_14_426 ();
 b15zdnd11an1n16x5 FILLER_14_458 ();
 b15zdnd00an1n02x5 FILLER_14_474 ();
 b15zdnd00an1n01x5 FILLER_14_476 ();
 b15zdnd11an1n64x5 FILLER_14_491 ();
 b15zdnd11an1n32x5 FILLER_14_555 ();
 b15zdnd00an1n02x5 FILLER_14_587 ();
 b15zdnd00an1n01x5 FILLER_14_589 ();
 b15zdnd11an1n08x5 FILLER_14_597 ();
 b15zdnd11an1n04x5 FILLER_14_611 ();
 b15zdnd11an1n32x5 FILLER_14_625 ();
 b15zdnd11an1n08x5 FILLER_14_657 ();
 b15zdnd11an1n04x5 FILLER_14_665 ();
 b15zdnd00an1n02x5 FILLER_14_669 ();
 b15zdnd11an1n32x5 FILLER_14_677 ();
 b15zdnd11an1n08x5 FILLER_14_709 ();
 b15zdnd00an1n01x5 FILLER_14_717 ();
 b15zdnd11an1n04x5 FILLER_14_726 ();
 b15zdnd00an1n01x5 FILLER_14_730 ();
 b15zdnd11an1n08x5 FILLER_14_739 ();
 b15zdnd11an1n32x5 FILLER_14_752 ();
 b15zdnd11an1n16x5 FILLER_14_784 ();
 b15zdnd11an1n08x5 FILLER_14_800 ();
 b15zdnd00an1n02x5 FILLER_14_808 ();
 b15zdnd00an1n01x5 FILLER_14_810 ();
 b15zdnd11an1n16x5 FILLER_14_815 ();
 b15zdnd11an1n08x5 FILLER_14_831 ();
 b15zdnd11an1n64x5 FILLER_14_854 ();
 b15zdnd11an1n64x5 FILLER_14_918 ();
 b15zdnd11an1n32x5 FILLER_14_982 ();
 b15zdnd11an1n16x5 FILLER_14_1014 ();
 b15zdnd11an1n08x5 FILLER_14_1030 ();
 b15zdnd11an1n04x5 FILLER_14_1038 ();
 b15zdnd11an1n64x5 FILLER_14_1046 ();
 b15zdnd11an1n64x5 FILLER_14_1110 ();
 b15zdnd11an1n32x5 FILLER_14_1174 ();
 b15zdnd11an1n16x5 FILLER_14_1206 ();
 b15zdnd00an1n02x5 FILLER_14_1222 ();
 b15zdnd11an1n32x5 FILLER_14_1234 ();
 b15zdnd11an1n16x5 FILLER_14_1266 ();
 b15zdnd11an1n08x5 FILLER_14_1282 ();
 b15zdnd11an1n04x5 FILLER_14_1290 ();
 b15zdnd00an1n02x5 FILLER_14_1294 ();
 b15zdnd00an1n01x5 FILLER_14_1296 ();
 b15zdnd11an1n08x5 FILLER_14_1317 ();
 b15zdnd11an1n04x5 FILLER_14_1325 ();
 b15zdnd00an1n02x5 FILLER_14_1329 ();
 b15zdnd11an1n64x5 FILLER_14_1351 ();
 b15zdnd11an1n64x5 FILLER_14_1415 ();
 b15zdnd11an1n32x5 FILLER_14_1479 ();
 b15zdnd11an1n16x5 FILLER_14_1511 ();
 b15zdnd11an1n08x5 FILLER_14_1527 ();
 b15zdnd00an1n01x5 FILLER_14_1535 ();
 b15zdnd11an1n32x5 FILLER_14_1544 ();
 b15zdnd11an1n08x5 FILLER_14_1576 ();
 b15zdnd11an1n04x5 FILLER_14_1584 ();
 b15zdnd00an1n01x5 FILLER_14_1588 ();
 b15zdnd11an1n08x5 FILLER_14_1596 ();
 b15zdnd11an1n04x5 FILLER_14_1604 ();
 b15zdnd11an1n64x5 FILLER_14_1614 ();
 b15zdnd11an1n64x5 FILLER_14_1678 ();
 b15zdnd11an1n08x5 FILLER_14_1742 ();
 b15zdnd11an1n08x5 FILLER_14_1776 ();
 b15zdnd11an1n04x5 FILLER_14_1784 ();
 b15zdnd00an1n02x5 FILLER_14_1788 ();
 b15zdnd11an1n16x5 FILLER_14_1797 ();
 b15zdnd00an1n02x5 FILLER_14_1813 ();
 b15zdnd11an1n64x5 FILLER_14_1822 ();
 b15zdnd11an1n32x5 FILLER_14_1886 ();
 b15zdnd11an1n16x5 FILLER_14_1918 ();
 b15zdnd11an1n04x5 FILLER_14_1934 ();
 b15zdnd00an1n02x5 FILLER_14_1938 ();
 b15zdnd11an1n16x5 FILLER_14_1952 ();
 b15zdnd11an1n08x5 FILLER_14_1968 ();
 b15zdnd11an1n04x5 FILLER_14_1976 ();
 b15zdnd00an1n02x5 FILLER_14_1980 ();
 b15zdnd00an1n01x5 FILLER_14_1982 ();
 b15zdnd11an1n16x5 FILLER_14_1989 ();
 b15zdnd11an1n08x5 FILLER_14_2005 ();
 b15zdnd11an1n16x5 FILLER_14_2022 ();
 b15zdnd11an1n04x5 FILLER_14_2038 ();
 b15zdnd00an1n02x5 FILLER_14_2042 ();
 b15zdnd00an1n01x5 FILLER_14_2044 ();
 b15zdnd11an1n04x5 FILLER_14_2051 ();
 b15zdnd00an1n02x5 FILLER_14_2055 ();
 b15zdnd00an1n01x5 FILLER_14_2057 ();
 b15zdnd11an1n16x5 FILLER_14_2067 ();
 b15zdnd11an1n08x5 FILLER_14_2083 ();
 b15zdnd11an1n04x5 FILLER_14_2091 ();
 b15zdnd00an1n01x5 FILLER_14_2095 ();
 b15zdnd11an1n32x5 FILLER_14_2111 ();
 b15zdnd11an1n08x5 FILLER_14_2143 ();
 b15zdnd00an1n02x5 FILLER_14_2151 ();
 b15zdnd00an1n01x5 FILLER_14_2153 ();
 b15zdnd11an1n04x5 FILLER_14_2162 ();
 b15zdnd00an1n01x5 FILLER_14_2166 ();
 b15zdnd11an1n64x5 FILLER_14_2182 ();
 b15zdnd11an1n16x5 FILLER_14_2246 ();
 b15zdnd11an1n08x5 FILLER_14_2262 ();
 b15zdnd11an1n04x5 FILLER_14_2270 ();
 b15zdnd00an1n02x5 FILLER_14_2274 ();
 b15zdnd11an1n64x5 FILLER_15_0 ();
 b15zdnd11an1n16x5 FILLER_15_64 ();
 b15zdnd11an1n08x5 FILLER_15_80 ();
 b15zdnd11an1n04x5 FILLER_15_88 ();
 b15zdnd11an1n16x5 FILLER_15_108 ();
 b15zdnd11an1n04x5 FILLER_15_124 ();
 b15zdnd11an1n08x5 FILLER_15_148 ();
 b15zdnd11an1n04x5 FILLER_15_156 ();
 b15zdnd00an1n01x5 FILLER_15_160 ();
 b15zdnd11an1n04x5 FILLER_15_166 ();
 b15zdnd11an1n04x5 FILLER_15_176 ();
 b15zdnd11an1n08x5 FILLER_15_197 ();
 b15zdnd11an1n04x5 FILLER_15_205 ();
 b15zdnd00an1n01x5 FILLER_15_209 ();
 b15zdnd11an1n16x5 FILLER_15_217 ();
 b15zdnd11an1n04x5 FILLER_15_233 ();
 b15zdnd00an1n01x5 FILLER_15_237 ();
 b15zdnd11an1n32x5 FILLER_15_242 ();
 b15zdnd11an1n16x5 FILLER_15_274 ();
 b15zdnd11an1n64x5 FILLER_15_302 ();
 b15zdnd11an1n32x5 FILLER_15_366 ();
 b15zdnd11an1n08x5 FILLER_15_398 ();
 b15zdnd11an1n04x5 FILLER_15_406 ();
 b15zdnd00an1n02x5 FILLER_15_410 ();
 b15zdnd00an1n01x5 FILLER_15_412 ();
 b15zdnd11an1n04x5 FILLER_15_429 ();
 b15zdnd11an1n16x5 FILLER_15_464 ();
 b15zdnd11an1n08x5 FILLER_15_480 ();
 b15zdnd00an1n02x5 FILLER_15_488 ();
 b15zdnd11an1n04x5 FILLER_15_497 ();
 b15zdnd11an1n04x5 FILLER_15_515 ();
 b15zdnd11an1n64x5 FILLER_15_524 ();
 b15zdnd00an1n02x5 FILLER_15_588 ();
 b15zdnd11an1n64x5 FILLER_15_597 ();
 b15zdnd11an1n04x5 FILLER_15_661 ();
 b15zdnd00an1n02x5 FILLER_15_665 ();
 b15zdnd11an1n16x5 FILLER_15_674 ();
 b15zdnd11an1n08x5 FILLER_15_690 ();
 b15zdnd11an1n32x5 FILLER_15_703 ();
 b15zdnd11an1n04x5 FILLER_15_735 ();
 b15zdnd11an1n16x5 FILLER_15_751 ();
 b15zdnd11an1n08x5 FILLER_15_767 ();
 b15zdnd11an1n04x5 FILLER_15_775 ();
 b15zdnd00an1n02x5 FILLER_15_779 ();
 b15zdnd00an1n01x5 FILLER_15_781 ();
 b15zdnd11an1n04x5 FILLER_15_814 ();
 b15zdnd11an1n16x5 FILLER_15_823 ();
 b15zdnd11an1n04x5 FILLER_15_839 ();
 b15zdnd00an1n01x5 FILLER_15_843 ();
 b15zdnd11an1n16x5 FILLER_15_850 ();
 b15zdnd11an1n04x5 FILLER_15_866 ();
 b15zdnd11an1n64x5 FILLER_15_888 ();
 b15zdnd11an1n64x5 FILLER_15_952 ();
 b15zdnd11an1n64x5 FILLER_15_1016 ();
 b15zdnd11an1n64x5 FILLER_15_1080 ();
 b15zdnd11an1n64x5 FILLER_15_1144 ();
 b15zdnd11an1n16x5 FILLER_15_1208 ();
 b15zdnd11an1n04x5 FILLER_15_1224 ();
 b15zdnd11an1n16x5 FILLER_15_1249 ();
 b15zdnd11an1n08x5 FILLER_15_1265 ();
 b15zdnd11an1n04x5 FILLER_15_1273 ();
 b15zdnd11an1n16x5 FILLER_15_1281 ();
 b15zdnd11an1n04x5 FILLER_15_1297 ();
 b15zdnd00an1n01x5 FILLER_15_1301 ();
 b15zdnd11an1n32x5 FILLER_15_1307 ();
 b15zdnd00an1n02x5 FILLER_15_1339 ();
 b15zdnd11an1n64x5 FILLER_15_1344 ();
 b15zdnd11an1n64x5 FILLER_15_1408 ();
 b15zdnd11an1n32x5 FILLER_15_1472 ();
 b15zdnd11an1n04x5 FILLER_15_1504 ();
 b15zdnd00an1n01x5 FILLER_15_1508 ();
 b15zdnd11an1n16x5 FILLER_15_1514 ();
 b15zdnd11an1n08x5 FILLER_15_1530 ();
 b15zdnd00an1n02x5 FILLER_15_1538 ();
 b15zdnd11an1n04x5 FILLER_15_1558 ();
 b15zdnd11an1n08x5 FILLER_15_1574 ();
 b15zdnd11an1n04x5 FILLER_15_1582 ();
 b15zdnd00an1n02x5 FILLER_15_1586 ();
 b15zdnd11an1n04x5 FILLER_15_1597 ();
 b15zdnd11an1n16x5 FILLER_15_1608 ();
 b15zdnd00an1n01x5 FILLER_15_1624 ();
 b15zdnd11an1n04x5 FILLER_15_1637 ();
 b15zdnd00an1n01x5 FILLER_15_1641 ();
 b15zdnd11an1n64x5 FILLER_15_1652 ();
 b15zdnd11an1n16x5 FILLER_15_1716 ();
 b15zdnd11an1n08x5 FILLER_15_1732 ();
 b15zdnd00an1n01x5 FILLER_15_1740 ();
 b15zdnd11an1n08x5 FILLER_15_1747 ();
 b15zdnd11an1n04x5 FILLER_15_1755 ();
 b15zdnd00an1n01x5 FILLER_15_1759 ();
 b15zdnd11an1n08x5 FILLER_15_1772 ();
 b15zdnd00an1n02x5 FILLER_15_1780 ();
 b15zdnd11an1n08x5 FILLER_15_1791 ();
 b15zdnd00an1n01x5 FILLER_15_1799 ();
 b15zdnd11an1n04x5 FILLER_15_1806 ();
 b15zdnd11an1n32x5 FILLER_15_1822 ();
 b15zdnd11an1n04x5 FILLER_15_1854 ();
 b15zdnd11an1n16x5 FILLER_15_1878 ();
 b15zdnd11an1n08x5 FILLER_15_1894 ();
 b15zdnd11an1n04x5 FILLER_15_1902 ();
 b15zdnd00an1n01x5 FILLER_15_1906 ();
 b15zdnd11an1n16x5 FILLER_15_1913 ();
 b15zdnd11an1n08x5 FILLER_15_1929 ();
 b15zdnd00an1n02x5 FILLER_15_1937 ();
 b15zdnd00an1n01x5 FILLER_15_1939 ();
 b15zdnd11an1n16x5 FILLER_15_1951 ();
 b15zdnd11an1n08x5 FILLER_15_1967 ();
 b15zdnd11an1n04x5 FILLER_15_1975 ();
 b15zdnd00an1n01x5 FILLER_15_1979 ();
 b15zdnd11an1n32x5 FILLER_15_1984 ();
 b15zdnd11an1n16x5 FILLER_15_2016 ();
 b15zdnd11an1n08x5 FILLER_15_2032 ();
 b15zdnd00an1n01x5 FILLER_15_2040 ();
 b15zdnd11an1n16x5 FILLER_15_2047 ();
 b15zdnd11an1n16x5 FILLER_15_2070 ();
 b15zdnd00an1n01x5 FILLER_15_2086 ();
 b15zdnd11an1n64x5 FILLER_15_2092 ();
 b15zdnd11an1n04x5 FILLER_15_2156 ();
 b15zdnd00an1n01x5 FILLER_15_2160 ();
 b15zdnd11an1n32x5 FILLER_15_2175 ();
 b15zdnd00an1n01x5 FILLER_15_2207 ();
 b15zdnd11an1n04x5 FILLER_15_2213 ();
 b15zdnd11an1n32x5 FILLER_15_2226 ();
 b15zdnd11an1n16x5 FILLER_15_2258 ();
 b15zdnd11an1n08x5 FILLER_15_2274 ();
 b15zdnd00an1n02x5 FILLER_15_2282 ();
 b15zdnd11an1n16x5 FILLER_16_8 ();
 b15zdnd11an1n08x5 FILLER_16_24 ();
 b15zdnd11an1n04x5 FILLER_16_32 ();
 b15zdnd00an1n02x5 FILLER_16_36 ();
 b15zdnd00an1n01x5 FILLER_16_38 ();
 b15zdnd11an1n04x5 FILLER_16_62 ();
 b15zdnd11an1n08x5 FILLER_16_91 ();
 b15zdnd11an1n64x5 FILLER_16_122 ();
 b15zdnd11an1n32x5 FILLER_16_186 ();
 b15zdnd11an1n16x5 FILLER_16_218 ();
 b15zdnd11an1n04x5 FILLER_16_234 ();
 b15zdnd00an1n01x5 FILLER_16_238 ();
 b15zdnd11an1n04x5 FILLER_16_249 ();
 b15zdnd11an1n08x5 FILLER_16_277 ();
 b15zdnd00an1n02x5 FILLER_16_285 ();
 b15zdnd11an1n04x5 FILLER_16_294 ();
 b15zdnd11an1n04x5 FILLER_16_310 ();
 b15zdnd00an1n01x5 FILLER_16_314 ();
 b15zdnd11an1n16x5 FILLER_16_320 ();
 b15zdnd11an1n08x5 FILLER_16_336 ();
 b15zdnd11an1n04x5 FILLER_16_344 ();
 b15zdnd00an1n02x5 FILLER_16_348 ();
 b15zdnd11an1n32x5 FILLER_16_381 ();
 b15zdnd00an1n02x5 FILLER_16_413 ();
 b15zdnd11an1n32x5 FILLER_16_429 ();
 b15zdnd11an1n08x5 FILLER_16_471 ();
 b15zdnd11an1n04x5 FILLER_16_479 ();
 b15zdnd00an1n01x5 FILLER_16_483 ();
 b15zdnd11an1n04x5 FILLER_16_490 ();
 b15zdnd11an1n32x5 FILLER_16_499 ();
 b15zdnd00an1n02x5 FILLER_16_531 ();
 b15zdnd00an1n01x5 FILLER_16_533 ();
 b15zdnd11an1n04x5 FILLER_16_539 ();
 b15zdnd11an1n32x5 FILLER_16_551 ();
 b15zdnd11an1n16x5 FILLER_16_583 ();
 b15zdnd11an1n04x5 FILLER_16_599 ();
 b15zdnd00an1n01x5 FILLER_16_603 ();
 b15zdnd11an1n08x5 FILLER_16_609 ();
 b15zdnd11an1n04x5 FILLER_16_617 ();
 b15zdnd00an1n02x5 FILLER_16_621 ();
 b15zdnd11an1n04x5 FILLER_16_637 ();
 b15zdnd11an1n08x5 FILLER_16_653 ();
 b15zdnd11an1n04x5 FILLER_16_661 ();
 b15zdnd00an1n02x5 FILLER_16_665 ();
 b15zdnd00an1n01x5 FILLER_16_667 ();
 b15zdnd11an1n08x5 FILLER_16_684 ();
 b15zdnd00an1n02x5 FILLER_16_716 ();
 b15zdnd11an1n16x5 FILLER_16_726 ();
 b15zdnd11an1n08x5 FILLER_16_742 ();
 b15zdnd11an1n04x5 FILLER_16_750 ();
 b15zdnd00an1n02x5 FILLER_16_754 ();
 b15zdnd11an1n04x5 FILLER_16_765 ();
 b15zdnd11an1n04x5 FILLER_16_775 ();
 b15zdnd11an1n16x5 FILLER_16_788 ();
 b15zdnd11an1n04x5 FILLER_16_804 ();
 b15zdnd00an1n01x5 FILLER_16_808 ();
 b15zdnd11an1n04x5 FILLER_16_815 ();
 b15zdnd11an1n16x5 FILLER_16_824 ();
 b15zdnd00an1n02x5 FILLER_16_840 ();
 b15zdnd00an1n01x5 FILLER_16_842 ();
 b15zdnd11an1n04x5 FILLER_16_850 ();
 b15zdnd00an1n02x5 FILLER_16_854 ();
 b15zdnd00an1n01x5 FILLER_16_856 ();
 b15zdnd11an1n16x5 FILLER_16_867 ();
 b15zdnd00an1n02x5 FILLER_16_883 ();
 b15zdnd11an1n64x5 FILLER_16_911 ();
 b15zdnd11an1n04x5 FILLER_16_975 ();
 b15zdnd00an1n02x5 FILLER_16_979 ();
 b15zdnd00an1n01x5 FILLER_16_981 ();
 b15zdnd11an1n32x5 FILLER_16_986 ();
 b15zdnd11an1n04x5 FILLER_16_1018 ();
 b15zdnd00an1n01x5 FILLER_16_1022 ();
 b15zdnd11an1n64x5 FILLER_16_1028 ();
 b15zdnd11an1n64x5 FILLER_16_1092 ();
 b15zdnd11an1n08x5 FILLER_16_1156 ();
 b15zdnd11an1n32x5 FILLER_16_1184 ();
 b15zdnd11an1n16x5 FILLER_16_1216 ();
 b15zdnd11an1n08x5 FILLER_16_1232 ();
 b15zdnd11an1n04x5 FILLER_16_1240 ();
 b15zdnd00an1n02x5 FILLER_16_1244 ();
 b15zdnd11an1n04x5 FILLER_16_1267 ();
 b15zdnd00an1n01x5 FILLER_16_1271 ();
 b15zdnd11an1n64x5 FILLER_16_1277 ();
 b15zdnd11an1n32x5 FILLER_16_1341 ();
 b15zdnd11an1n16x5 FILLER_16_1373 ();
 b15zdnd11an1n04x5 FILLER_16_1389 ();
 b15zdnd00an1n01x5 FILLER_16_1393 ();
 b15zdnd11an1n04x5 FILLER_16_1400 ();
 b15zdnd11an1n32x5 FILLER_16_1414 ();
 b15zdnd00an1n02x5 FILLER_16_1446 ();
 b15zdnd11an1n32x5 FILLER_16_1452 ();
 b15zdnd11an1n04x5 FILLER_16_1484 ();
 b15zdnd11an1n04x5 FILLER_16_1497 ();
 b15zdnd00an1n01x5 FILLER_16_1501 ();
 b15zdnd11an1n16x5 FILLER_16_1512 ();
 b15zdnd00an1n02x5 FILLER_16_1528 ();
 b15zdnd11an1n04x5 FILLER_16_1546 ();
 b15zdnd00an1n01x5 FILLER_16_1550 ();
 b15zdnd11an1n32x5 FILLER_16_1556 ();
 b15zdnd11an1n08x5 FILLER_16_1588 ();
 b15zdnd11an1n04x5 FILLER_16_1596 ();
 b15zdnd11an1n04x5 FILLER_16_1608 ();
 b15zdnd11an1n08x5 FILLER_16_1619 ();
 b15zdnd00an1n02x5 FILLER_16_1627 ();
 b15zdnd11an1n04x5 FILLER_16_1636 ();
 b15zdnd00an1n02x5 FILLER_16_1640 ();
 b15zdnd00an1n01x5 FILLER_16_1642 ();
 b15zdnd11an1n08x5 FILLER_16_1650 ();
 b15zdnd11an1n32x5 FILLER_16_1676 ();
 b15zdnd11an1n16x5 FILLER_16_1708 ();
 b15zdnd11an1n04x5 FILLER_16_1724 ();
 b15zdnd00an1n02x5 FILLER_16_1728 ();
 b15zdnd11an1n04x5 FILLER_16_1737 ();
 b15zdnd00an1n01x5 FILLER_16_1741 ();
 b15zdnd11an1n04x5 FILLER_16_1755 ();
 b15zdnd11an1n16x5 FILLER_16_1766 ();
 b15zdnd11an1n04x5 FILLER_16_1782 ();
 b15zdnd00an1n02x5 FILLER_16_1786 ();
 b15zdnd11an1n32x5 FILLER_16_1814 ();
 b15zdnd11an1n08x5 FILLER_16_1846 ();
 b15zdnd00an1n01x5 FILLER_16_1854 ();
 b15zdnd11an1n16x5 FILLER_16_1861 ();
 b15zdnd11an1n04x5 FILLER_16_1877 ();
 b15zdnd11an1n16x5 FILLER_16_1886 ();
 b15zdnd11an1n04x5 FILLER_16_1902 ();
 b15zdnd00an1n02x5 FILLER_16_1906 ();
 b15zdnd11an1n32x5 FILLER_16_1916 ();
 b15zdnd00an1n02x5 FILLER_16_1948 ();
 b15zdnd11an1n04x5 FILLER_16_1955 ();
 b15zdnd11an1n08x5 FILLER_16_1979 ();
 b15zdnd11an1n04x5 FILLER_16_1987 ();
 b15zdnd00an1n01x5 FILLER_16_1991 ();
 b15zdnd11an1n04x5 FILLER_16_2001 ();
 b15zdnd11an1n08x5 FILLER_16_2009 ();
 b15zdnd11an1n16x5 FILLER_16_2022 ();
 b15zdnd11an1n08x5 FILLER_16_2038 ();
 b15zdnd00an1n01x5 FILLER_16_2046 ();
 b15zdnd11an1n16x5 FILLER_16_2063 ();
 b15zdnd11an1n08x5 FILLER_16_2079 ();
 b15zdnd11an1n08x5 FILLER_16_2095 ();
 b15zdnd11an1n16x5 FILLER_16_2107 ();
 b15zdnd11an1n04x5 FILLER_16_2123 ();
 b15zdnd11an1n08x5 FILLER_16_2143 ();
 b15zdnd00an1n02x5 FILLER_16_2151 ();
 b15zdnd00an1n01x5 FILLER_16_2153 ();
 b15zdnd11an1n32x5 FILLER_16_2162 ();
 b15zdnd11an1n04x5 FILLER_16_2206 ();
 b15zdnd11an1n32x5 FILLER_16_2226 ();
 b15zdnd11an1n16x5 FILLER_16_2258 ();
 b15zdnd00an1n02x5 FILLER_16_2274 ();
 b15zdnd11an1n64x5 FILLER_17_0 ();
 b15zdnd11an1n32x5 FILLER_17_64 ();
 b15zdnd00an1n01x5 FILLER_17_96 ();
 b15zdnd11an1n64x5 FILLER_17_129 ();
 b15zdnd11an1n16x5 FILLER_17_193 ();
 b15zdnd11an1n04x5 FILLER_17_214 ();
 b15zdnd11an1n08x5 FILLER_17_223 ();
 b15zdnd11an1n04x5 FILLER_17_231 ();
 b15zdnd00an1n01x5 FILLER_17_235 ();
 b15zdnd11an1n08x5 FILLER_17_257 ();
 b15zdnd11an1n04x5 FILLER_17_265 ();
 b15zdnd00an1n02x5 FILLER_17_269 ();
 b15zdnd00an1n01x5 FILLER_17_271 ();
 b15zdnd11an1n16x5 FILLER_17_284 ();
 b15zdnd11an1n08x5 FILLER_17_300 ();
 b15zdnd11an1n16x5 FILLER_17_312 ();
 b15zdnd11an1n04x5 FILLER_17_328 ();
 b15zdnd11an1n64x5 FILLER_17_336 ();
 b15zdnd11an1n32x5 FILLER_17_400 ();
 b15zdnd11an1n04x5 FILLER_17_432 ();
 b15zdnd00an1n01x5 FILLER_17_436 ();
 b15zdnd11an1n32x5 FILLER_17_441 ();
 b15zdnd11an1n04x5 FILLER_17_473 ();
 b15zdnd11an1n04x5 FILLER_17_492 ();
 b15zdnd00an1n02x5 FILLER_17_496 ();
 b15zdnd11an1n64x5 FILLER_17_504 ();
 b15zdnd00an1n02x5 FILLER_17_568 ();
 b15zdnd00an1n01x5 FILLER_17_570 ();
 b15zdnd11an1n32x5 FILLER_17_576 ();
 b15zdnd11an1n16x5 FILLER_17_608 ();
 b15zdnd00an1n02x5 FILLER_17_624 ();
 b15zdnd00an1n01x5 FILLER_17_626 ();
 b15zdnd11an1n32x5 FILLER_17_634 ();
 b15zdnd00an1n02x5 FILLER_17_666 ();
 b15zdnd00an1n01x5 FILLER_17_668 ();
 b15zdnd11an1n64x5 FILLER_17_674 ();
 b15zdnd11an1n64x5 FILLER_17_738 ();
 b15zdnd11an1n32x5 FILLER_17_802 ();
 b15zdnd11an1n16x5 FILLER_17_834 ();
 b15zdnd11an1n08x5 FILLER_17_850 ();
 b15zdnd11an1n04x5 FILLER_17_858 ();
 b15zdnd00an1n01x5 FILLER_17_862 ();
 b15zdnd11an1n64x5 FILLER_17_873 ();
 b15zdnd11an1n08x5 FILLER_17_937 ();
 b15zdnd00an1n01x5 FILLER_17_945 ();
 b15zdnd11an1n04x5 FILLER_17_966 ();
 b15zdnd11an1n32x5 FILLER_17_975 ();
 b15zdnd11an1n08x5 FILLER_17_1007 ();
 b15zdnd00an1n02x5 FILLER_17_1015 ();
 b15zdnd00an1n01x5 FILLER_17_1017 ();
 b15zdnd11an1n32x5 FILLER_17_1038 ();
 b15zdnd11an1n08x5 FILLER_17_1070 ();
 b15zdnd00an1n02x5 FILLER_17_1078 ();
 b15zdnd11an1n08x5 FILLER_17_1100 ();
 b15zdnd00an1n02x5 FILLER_17_1108 ();
 b15zdnd11an1n16x5 FILLER_17_1116 ();
 b15zdnd11an1n04x5 FILLER_17_1132 ();
 b15zdnd00an1n02x5 FILLER_17_1136 ();
 b15zdnd00an1n01x5 FILLER_17_1138 ();
 b15zdnd11an1n64x5 FILLER_17_1152 ();
 b15zdnd11an1n32x5 FILLER_17_1216 ();
 b15zdnd11an1n16x5 FILLER_17_1248 ();
 b15zdnd11an1n08x5 FILLER_17_1264 ();
 b15zdnd11an1n64x5 FILLER_17_1292 ();
 b15zdnd11an1n32x5 FILLER_17_1356 ();
 b15zdnd11an1n08x5 FILLER_17_1388 ();
 b15zdnd00an1n02x5 FILLER_17_1396 ();
 b15zdnd00an1n01x5 FILLER_17_1398 ();
 b15zdnd11an1n04x5 FILLER_17_1404 ();
 b15zdnd00an1n02x5 FILLER_17_1408 ();
 b15zdnd11an1n08x5 FILLER_17_1434 ();
 b15zdnd11an1n08x5 FILLER_17_1450 ();
 b15zdnd11an1n04x5 FILLER_17_1458 ();
 b15zdnd00an1n02x5 FILLER_17_1462 ();
 b15zdnd00an1n01x5 FILLER_17_1464 ();
 b15zdnd11an1n32x5 FILLER_17_1472 ();
 b15zdnd11an1n16x5 FILLER_17_1504 ();
 b15zdnd11an1n08x5 FILLER_17_1520 ();
 b15zdnd00an1n02x5 FILLER_17_1528 ();
 b15zdnd11an1n08x5 FILLER_17_1542 ();
 b15zdnd11an1n04x5 FILLER_17_1550 ();
 b15zdnd11an1n32x5 FILLER_17_1567 ();
 b15zdnd11an1n08x5 FILLER_17_1599 ();
 b15zdnd00an1n01x5 FILLER_17_1607 ();
 b15zdnd11an1n32x5 FILLER_17_1621 ();
 b15zdnd11an1n08x5 FILLER_17_1653 ();
 b15zdnd00an1n02x5 FILLER_17_1661 ();
 b15zdnd00an1n01x5 FILLER_17_1663 ();
 b15zdnd11an1n64x5 FILLER_17_1682 ();
 b15zdnd11an1n64x5 FILLER_17_1746 ();
 b15zdnd11an1n32x5 FILLER_17_1810 ();
 b15zdnd11an1n08x5 FILLER_17_1842 ();
 b15zdnd00an1n01x5 FILLER_17_1850 ();
 b15zdnd11an1n16x5 FILLER_17_1856 ();
 b15zdnd11an1n04x5 FILLER_17_1872 ();
 b15zdnd00an1n02x5 FILLER_17_1876 ();
 b15zdnd00an1n01x5 FILLER_17_1878 ();
 b15zdnd11an1n64x5 FILLER_17_1893 ();
 b15zdnd11an1n64x5 FILLER_17_1957 ();
 b15zdnd11an1n08x5 FILLER_17_2021 ();
 b15zdnd00an1n01x5 FILLER_17_2029 ();
 b15zdnd11an1n32x5 FILLER_17_2051 ();
 b15zdnd11an1n16x5 FILLER_17_2083 ();
 b15zdnd11an1n08x5 FILLER_17_2099 ();
 b15zdnd11an1n32x5 FILLER_17_2112 ();
 b15zdnd11an1n16x5 FILLER_17_2144 ();
 b15zdnd11an1n08x5 FILLER_17_2160 ();
 b15zdnd11an1n04x5 FILLER_17_2168 ();
 b15zdnd00an1n02x5 FILLER_17_2172 ();
 b15zdnd11an1n32x5 FILLER_17_2178 ();
 b15zdnd11an1n64x5 FILLER_17_2215 ();
 b15zdnd11an1n04x5 FILLER_17_2279 ();
 b15zdnd00an1n01x5 FILLER_17_2283 ();
 b15zdnd11an1n32x5 FILLER_18_8 ();
 b15zdnd11an1n16x5 FILLER_18_40 ();
 b15zdnd00an1n01x5 FILLER_18_56 ();
 b15zdnd11an1n04x5 FILLER_18_73 ();
 b15zdnd11an1n16x5 FILLER_18_109 ();
 b15zdnd00an1n01x5 FILLER_18_125 ();
 b15zdnd11an1n04x5 FILLER_18_131 ();
 b15zdnd11an1n64x5 FILLER_18_150 ();
 b15zdnd11an1n32x5 FILLER_18_214 ();
 b15zdnd11an1n16x5 FILLER_18_246 ();
 b15zdnd11an1n08x5 FILLER_18_262 ();
 b15zdnd11an1n04x5 FILLER_18_270 ();
 b15zdnd00an1n02x5 FILLER_18_274 ();
 b15zdnd11an1n64x5 FILLER_18_286 ();
 b15zdnd11an1n64x5 FILLER_18_350 ();
 b15zdnd11an1n16x5 FILLER_18_414 ();
 b15zdnd00an1n02x5 FILLER_18_430 ();
 b15zdnd00an1n01x5 FILLER_18_432 ();
 b15zdnd11an1n64x5 FILLER_18_446 ();
 b15zdnd11an1n16x5 FILLER_18_510 ();
 b15zdnd11an1n08x5 FILLER_18_526 ();
 b15zdnd11an1n16x5 FILLER_18_554 ();
 b15zdnd00an1n01x5 FILLER_18_570 ();
 b15zdnd11an1n16x5 FILLER_18_577 ();
 b15zdnd00an1n01x5 FILLER_18_593 ();
 b15zdnd11an1n64x5 FILLER_18_600 ();
 b15zdnd11an1n08x5 FILLER_18_664 ();
 b15zdnd00an1n01x5 FILLER_18_672 ();
 b15zdnd11an1n32x5 FILLER_18_679 ();
 b15zdnd11an1n04x5 FILLER_18_711 ();
 b15zdnd00an1n02x5 FILLER_18_715 ();
 b15zdnd00an1n01x5 FILLER_18_717 ();
 b15zdnd11an1n08x5 FILLER_18_726 ();
 b15zdnd00an1n01x5 FILLER_18_734 ();
 b15zdnd11an1n64x5 FILLER_18_749 ();
 b15zdnd11an1n04x5 FILLER_18_813 ();
 b15zdnd00an1n02x5 FILLER_18_817 ();
 b15zdnd11an1n16x5 FILLER_18_839 ();
 b15zdnd11an1n08x5 FILLER_18_855 ();
 b15zdnd11an1n04x5 FILLER_18_863 ();
 b15zdnd11an1n64x5 FILLER_18_880 ();
 b15zdnd11an1n04x5 FILLER_18_944 ();
 b15zdnd11an1n16x5 FILLER_18_968 ();
 b15zdnd11an1n04x5 FILLER_18_984 ();
 b15zdnd11an1n16x5 FILLER_18_1008 ();
 b15zdnd11an1n08x5 FILLER_18_1024 ();
 b15zdnd00an1n01x5 FILLER_18_1032 ();
 b15zdnd11an1n64x5 FILLER_18_1036 ();
 b15zdnd11an1n04x5 FILLER_18_1100 ();
 b15zdnd00an1n02x5 FILLER_18_1104 ();
 b15zdnd11an1n08x5 FILLER_18_1126 ();
 b15zdnd11an1n04x5 FILLER_18_1134 ();
 b15zdnd00an1n02x5 FILLER_18_1138 ();
 b15zdnd00an1n01x5 FILLER_18_1140 ();
 b15zdnd11an1n32x5 FILLER_18_1159 ();
 b15zdnd11an1n04x5 FILLER_18_1191 ();
 b15zdnd00an1n02x5 FILLER_18_1195 ();
 b15zdnd11an1n64x5 FILLER_18_1203 ();
 b15zdnd11an1n16x5 FILLER_18_1267 ();
 b15zdnd00an1n02x5 FILLER_18_1283 ();
 b15zdnd11an1n16x5 FILLER_18_1311 ();
 b15zdnd11an1n08x5 FILLER_18_1327 ();
 b15zdnd11an1n64x5 FILLER_18_1353 ();
 b15zdnd11an1n08x5 FILLER_18_1417 ();
 b15zdnd11an1n04x5 FILLER_18_1425 ();
 b15zdnd00an1n01x5 FILLER_18_1429 ();
 b15zdnd11an1n32x5 FILLER_18_1440 ();
 b15zdnd11an1n16x5 FILLER_18_1472 ();
 b15zdnd11an1n08x5 FILLER_18_1488 ();
 b15zdnd11an1n04x5 FILLER_18_1496 ();
 b15zdnd00an1n02x5 FILLER_18_1500 ();
 b15zdnd11an1n64x5 FILLER_18_1506 ();
 b15zdnd11an1n16x5 FILLER_18_1570 ();
 b15zdnd11an1n04x5 FILLER_18_1586 ();
 b15zdnd11an1n64x5 FILLER_18_1601 ();
 b15zdnd11an1n64x5 FILLER_18_1665 ();
 b15zdnd11an1n32x5 FILLER_18_1729 ();
 b15zdnd11an1n16x5 FILLER_18_1761 ();
 b15zdnd11an1n08x5 FILLER_18_1777 ();
 b15zdnd11an1n04x5 FILLER_18_1785 ();
 b15zdnd11an1n16x5 FILLER_18_1802 ();
 b15zdnd11an1n08x5 FILLER_18_1818 ();
 b15zdnd00an1n02x5 FILLER_18_1826 ();
 b15zdnd11an1n16x5 FILLER_18_1843 ();
 b15zdnd00an1n02x5 FILLER_18_1859 ();
 b15zdnd00an1n01x5 FILLER_18_1861 ();
 b15zdnd11an1n16x5 FILLER_18_1871 ();
 b15zdnd11an1n08x5 FILLER_18_1887 ();
 b15zdnd11an1n04x5 FILLER_18_1895 ();
 b15zdnd00an1n01x5 FILLER_18_1899 ();
 b15zdnd11an1n64x5 FILLER_18_1906 ();
 b15zdnd11an1n64x5 FILLER_18_1970 ();
 b15zdnd11an1n08x5 FILLER_18_2034 ();
 b15zdnd00an1n01x5 FILLER_18_2042 ();
 b15zdnd11an1n04x5 FILLER_18_2053 ();
 b15zdnd11an1n16x5 FILLER_18_2062 ();
 b15zdnd11an1n04x5 FILLER_18_2078 ();
 b15zdnd00an1n01x5 FILLER_18_2082 ();
 b15zdnd11an1n04x5 FILLER_18_2099 ();
 b15zdnd00an1n02x5 FILLER_18_2103 ();
 b15zdnd00an1n01x5 FILLER_18_2105 ();
 b15zdnd11an1n16x5 FILLER_18_2112 ();
 b15zdnd11an1n04x5 FILLER_18_2128 ();
 b15zdnd00an1n02x5 FILLER_18_2132 ();
 b15zdnd00an1n02x5 FILLER_18_2152 ();
 b15zdnd11an1n08x5 FILLER_18_2162 ();
 b15zdnd11an1n04x5 FILLER_18_2174 ();
 b15zdnd11an1n64x5 FILLER_18_2191 ();
 b15zdnd11an1n16x5 FILLER_18_2255 ();
 b15zdnd11an1n04x5 FILLER_18_2271 ();
 b15zdnd00an1n01x5 FILLER_18_2275 ();
 b15zdnd11an1n32x5 FILLER_19_0 ();
 b15zdnd11an1n16x5 FILLER_19_32 ();
 b15zdnd11an1n16x5 FILLER_19_60 ();
 b15zdnd00an1n02x5 FILLER_19_76 ();
 b15zdnd00an1n01x5 FILLER_19_78 ();
 b15zdnd11an1n16x5 FILLER_19_111 ();
 b15zdnd11an1n08x5 FILLER_19_127 ();
 b15zdnd00an1n02x5 FILLER_19_135 ();
 b15zdnd11an1n32x5 FILLER_19_153 ();
 b15zdnd11an1n08x5 FILLER_19_185 ();
 b15zdnd00an1n01x5 FILLER_19_193 ();
 b15zdnd11an1n32x5 FILLER_19_200 ();
 b15zdnd00an1n02x5 FILLER_19_232 ();
 b15zdnd11an1n32x5 FILLER_19_238 ();
 b15zdnd11an1n08x5 FILLER_19_270 ();
 b15zdnd00an1n02x5 FILLER_19_278 ();
 b15zdnd11an1n32x5 FILLER_19_285 ();
 b15zdnd11an1n08x5 FILLER_19_317 ();
 b15zdnd11an1n04x5 FILLER_19_330 ();
 b15zdnd11an1n32x5 FILLER_19_350 ();
 b15zdnd11an1n16x5 FILLER_19_382 ();
 b15zdnd11an1n08x5 FILLER_19_398 ();
 b15zdnd11an1n04x5 FILLER_19_406 ();
 b15zdnd00an1n02x5 FILLER_19_410 ();
 b15zdnd00an1n01x5 FILLER_19_412 ();
 b15zdnd11an1n04x5 FILLER_19_429 ();
 b15zdnd00an1n01x5 FILLER_19_433 ();
 b15zdnd11an1n32x5 FILLER_19_447 ();
 b15zdnd11an1n08x5 FILLER_19_479 ();
 b15zdnd00an1n02x5 FILLER_19_487 ();
 b15zdnd00an1n01x5 FILLER_19_489 ();
 b15zdnd11an1n08x5 FILLER_19_500 ();
 b15zdnd11an1n04x5 FILLER_19_508 ();
 b15zdnd00an1n02x5 FILLER_19_512 ();
 b15zdnd11an1n08x5 FILLER_19_527 ();
 b15zdnd11an1n04x5 FILLER_19_535 ();
 b15zdnd00an1n02x5 FILLER_19_539 ();
 b15zdnd11an1n16x5 FILLER_19_553 ();
 b15zdnd11an1n08x5 FILLER_19_569 ();
 b15zdnd00an1n01x5 FILLER_19_577 ();
 b15zdnd11an1n64x5 FILLER_19_590 ();
 b15zdnd00an1n02x5 FILLER_19_654 ();
 b15zdnd11an1n32x5 FILLER_19_661 ();
 b15zdnd11an1n04x5 FILLER_19_693 ();
 b15zdnd00an1n02x5 FILLER_19_697 ();
 b15zdnd11an1n16x5 FILLER_19_714 ();
 b15zdnd11an1n08x5 FILLER_19_730 ();
 b15zdnd11an1n32x5 FILLER_19_743 ();
 b15zdnd11an1n16x5 FILLER_19_775 ();
 b15zdnd11an1n08x5 FILLER_19_791 ();
 b15zdnd11an1n04x5 FILLER_19_799 ();
 b15zdnd00an1n01x5 FILLER_19_803 ();
 b15zdnd11an1n64x5 FILLER_19_808 ();
 b15zdnd11an1n64x5 FILLER_19_872 ();
 b15zdnd11an1n16x5 FILLER_19_936 ();
 b15zdnd11an1n08x5 FILLER_19_952 ();
 b15zdnd11an1n04x5 FILLER_19_960 ();
 b15zdnd11an1n64x5 FILLER_19_967 ();
 b15zdnd11an1n32x5 FILLER_19_1031 ();
 b15zdnd11an1n04x5 FILLER_19_1063 ();
 b15zdnd00an1n02x5 FILLER_19_1067 ();
 b15zdnd00an1n01x5 FILLER_19_1069 ();
 b15zdnd11an1n16x5 FILLER_19_1074 ();
 b15zdnd11an1n04x5 FILLER_19_1110 ();
 b15zdnd11an1n64x5 FILLER_19_1119 ();
 b15zdnd11an1n08x5 FILLER_19_1183 ();
 b15zdnd11an1n64x5 FILLER_19_1211 ();
 b15zdnd11an1n64x5 FILLER_19_1275 ();
 b15zdnd11an1n08x5 FILLER_19_1339 ();
 b15zdnd00an1n01x5 FILLER_19_1347 ();
 b15zdnd11an1n08x5 FILLER_19_1360 ();
 b15zdnd00an1n01x5 FILLER_19_1368 ();
 b15zdnd11an1n32x5 FILLER_19_1377 ();
 b15zdnd11an1n08x5 FILLER_19_1409 ();
 b15zdnd11an1n16x5 FILLER_19_1433 ();
 b15zdnd11an1n08x5 FILLER_19_1449 ();
 b15zdnd11an1n04x5 FILLER_19_1457 ();
 b15zdnd00an1n01x5 FILLER_19_1461 ();
 b15zdnd11an1n04x5 FILLER_19_1467 ();
 b15zdnd11an1n16x5 FILLER_19_1478 ();
 b15zdnd11an1n08x5 FILLER_19_1494 ();
 b15zdnd00an1n02x5 FILLER_19_1502 ();
 b15zdnd11an1n04x5 FILLER_19_1519 ();
 b15zdnd11an1n32x5 FILLER_19_1529 ();
 b15zdnd11an1n04x5 FILLER_19_1561 ();
 b15zdnd00an1n02x5 FILLER_19_1565 ();
 b15zdnd11an1n04x5 FILLER_19_1582 ();
 b15zdnd11an1n64x5 FILLER_19_1594 ();
 b15zdnd11an1n04x5 FILLER_19_1658 ();
 b15zdnd00an1n02x5 FILLER_19_1662 ();
 b15zdnd11an1n64x5 FILLER_19_1687 ();
 b15zdnd00an1n02x5 FILLER_19_1751 ();
 b15zdnd11an1n08x5 FILLER_19_1761 ();
 b15zdnd00an1n02x5 FILLER_19_1769 ();
 b15zdnd00an1n01x5 FILLER_19_1771 ();
 b15zdnd11an1n04x5 FILLER_19_1776 ();
 b15zdnd11an1n08x5 FILLER_19_1786 ();
 b15zdnd00an1n02x5 FILLER_19_1794 ();
 b15zdnd00an1n01x5 FILLER_19_1796 ();
 b15zdnd11an1n16x5 FILLER_19_1803 ();
 b15zdnd11an1n08x5 FILLER_19_1819 ();
 b15zdnd11an1n04x5 FILLER_19_1827 ();
 b15zdnd00an1n01x5 FILLER_19_1831 ();
 b15zdnd11an1n16x5 FILLER_19_1838 ();
 b15zdnd11an1n08x5 FILLER_19_1854 ();
 b15zdnd11an1n04x5 FILLER_19_1862 ();
 b15zdnd11an1n16x5 FILLER_19_1871 ();
 b15zdnd11an1n08x5 FILLER_19_1887 ();
 b15zdnd11an1n04x5 FILLER_19_1895 ();
 b15zdnd00an1n02x5 FILLER_19_1899 ();
 b15zdnd11an1n16x5 FILLER_19_1909 ();
 b15zdnd11an1n08x5 FILLER_19_1925 ();
 b15zdnd11an1n04x5 FILLER_19_1933 ();
 b15zdnd00an1n01x5 FILLER_19_1937 ();
 b15zdnd11an1n16x5 FILLER_19_1942 ();
 b15zdnd11an1n04x5 FILLER_19_1958 ();
 b15zdnd00an1n02x5 FILLER_19_1962 ();
 b15zdnd00an1n01x5 FILLER_19_1964 ();
 b15zdnd11an1n64x5 FILLER_19_1972 ();
 b15zdnd11an1n32x5 FILLER_19_2036 ();
 b15zdnd11an1n08x5 FILLER_19_2068 ();
 b15zdnd00an1n02x5 FILLER_19_2076 ();
 b15zdnd11an1n32x5 FILLER_19_2088 ();
 b15zdnd11an1n08x5 FILLER_19_2120 ();
 b15zdnd11an1n04x5 FILLER_19_2128 ();
 b15zdnd11an1n32x5 FILLER_19_2150 ();
 b15zdnd11an1n16x5 FILLER_19_2182 ();
 b15zdnd11an1n04x5 FILLER_19_2198 ();
 b15zdnd00an1n01x5 FILLER_19_2202 ();
 b15zdnd11an1n04x5 FILLER_19_2208 ();
 b15zdnd11an1n32x5 FILLER_19_2227 ();
 b15zdnd11an1n16x5 FILLER_19_2259 ();
 b15zdnd11an1n08x5 FILLER_19_2275 ();
 b15zdnd00an1n01x5 FILLER_19_2283 ();
 b15zdnd11an1n16x5 FILLER_20_8 ();
 b15zdnd11an1n08x5 FILLER_20_24 ();
 b15zdnd11an1n04x5 FILLER_20_32 ();
 b15zdnd00an1n01x5 FILLER_20_36 ();
 b15zdnd11an1n32x5 FILLER_20_60 ();
 b15zdnd11an1n16x5 FILLER_20_92 ();
 b15zdnd11an1n04x5 FILLER_20_108 ();
 b15zdnd00an1n02x5 FILLER_20_112 ();
 b15zdnd00an1n01x5 FILLER_20_114 ();
 b15zdnd11an1n32x5 FILLER_20_133 ();
 b15zdnd00an1n01x5 FILLER_20_165 ();
 b15zdnd11an1n32x5 FILLER_20_171 ();
 b15zdnd11an1n16x5 FILLER_20_203 ();
 b15zdnd11an1n08x5 FILLER_20_219 ();
 b15zdnd11an1n04x5 FILLER_20_227 ();
 b15zdnd00an1n02x5 FILLER_20_231 ();
 b15zdnd00an1n01x5 FILLER_20_233 ();
 b15zdnd11an1n64x5 FILLER_20_243 ();
 b15zdnd11an1n64x5 FILLER_20_307 ();
 b15zdnd11an1n08x5 FILLER_20_371 ();
 b15zdnd00an1n02x5 FILLER_20_379 ();
 b15zdnd11an1n08x5 FILLER_20_397 ();
 b15zdnd11an1n04x5 FILLER_20_405 ();
 b15zdnd00an1n01x5 FILLER_20_409 ();
 b15zdnd11an1n04x5 FILLER_20_414 ();
 b15zdnd11an1n16x5 FILLER_20_432 ();
 b15zdnd11an1n08x5 FILLER_20_448 ();
 b15zdnd11an1n04x5 FILLER_20_456 ();
 b15zdnd11an1n64x5 FILLER_20_468 ();
 b15zdnd11an1n32x5 FILLER_20_532 ();
 b15zdnd11an1n16x5 FILLER_20_564 ();
 b15zdnd00an1n02x5 FILLER_20_580 ();
 b15zdnd00an1n01x5 FILLER_20_582 ();
 b15zdnd11an1n08x5 FILLER_20_589 ();
 b15zdnd00an1n02x5 FILLER_20_597 ();
 b15zdnd11an1n32x5 FILLER_20_603 ();
 b15zdnd11an1n16x5 FILLER_20_635 ();
 b15zdnd11an1n32x5 FILLER_20_655 ();
 b15zdnd11an1n16x5 FILLER_20_687 ();
 b15zdnd11an1n08x5 FILLER_20_703 ();
 b15zdnd11an1n04x5 FILLER_20_711 ();
 b15zdnd00an1n02x5 FILLER_20_715 ();
 b15zdnd00an1n01x5 FILLER_20_717 ();
 b15zdnd11an1n32x5 FILLER_20_726 ();
 b15zdnd11an1n04x5 FILLER_20_758 ();
 b15zdnd00an1n01x5 FILLER_20_762 ();
 b15zdnd11an1n08x5 FILLER_20_769 ();
 b15zdnd11an1n04x5 FILLER_20_777 ();
 b15zdnd00an1n02x5 FILLER_20_781 ();
 b15zdnd00an1n01x5 FILLER_20_783 ();
 b15zdnd11an1n64x5 FILLER_20_795 ();
 b15zdnd00an1n01x5 FILLER_20_859 ();
 b15zdnd11an1n04x5 FILLER_20_867 ();
 b15zdnd00an1n02x5 FILLER_20_871 ();
 b15zdnd00an1n01x5 FILLER_20_873 ();
 b15zdnd11an1n04x5 FILLER_20_878 ();
 b15zdnd00an1n02x5 FILLER_20_882 ();
 b15zdnd11an1n04x5 FILLER_20_910 ();
 b15zdnd11an1n64x5 FILLER_20_940 ();
 b15zdnd11an1n16x5 FILLER_20_1004 ();
 b15zdnd11an1n08x5 FILLER_20_1020 ();
 b15zdnd00an1n01x5 FILLER_20_1028 ();
 b15zdnd11an1n64x5 FILLER_20_1033 ();
 b15zdnd11an1n64x5 FILLER_20_1097 ();
 b15zdnd11an1n32x5 FILLER_20_1161 ();
 b15zdnd11an1n04x5 FILLER_20_1193 ();
 b15zdnd00an1n01x5 FILLER_20_1197 ();
 b15zdnd11an1n32x5 FILLER_20_1203 ();
 b15zdnd11an1n16x5 FILLER_20_1235 ();
 b15zdnd11an1n08x5 FILLER_20_1251 ();
 b15zdnd11an1n64x5 FILLER_20_1263 ();
 b15zdnd11an1n08x5 FILLER_20_1358 ();
 b15zdnd11an1n64x5 FILLER_20_1382 ();
 b15zdnd11an1n08x5 FILLER_20_1452 ();
 b15zdnd11an1n04x5 FILLER_20_1471 ();
 b15zdnd11an1n32x5 FILLER_20_1479 ();
 b15zdnd11an1n04x5 FILLER_20_1511 ();
 b15zdnd00an1n02x5 FILLER_20_1515 ();
 b15zdnd00an1n01x5 FILLER_20_1517 ();
 b15zdnd11an1n16x5 FILLER_20_1534 ();
 b15zdnd11an1n04x5 FILLER_20_1550 ();
 b15zdnd00an1n02x5 FILLER_20_1554 ();
 b15zdnd00an1n01x5 FILLER_20_1556 ();
 b15zdnd11an1n64x5 FILLER_20_1573 ();
 b15zdnd00an1n01x5 FILLER_20_1637 ();
 b15zdnd11an1n64x5 FILLER_20_1652 ();
 b15zdnd11an1n16x5 FILLER_20_1716 ();
 b15zdnd00an1n02x5 FILLER_20_1732 ();
 b15zdnd00an1n01x5 FILLER_20_1734 ();
 b15zdnd11an1n04x5 FILLER_20_1761 ();
 b15zdnd11an1n32x5 FILLER_20_1791 ();
 b15zdnd11an1n08x5 FILLER_20_1823 ();
 b15zdnd00an1n01x5 FILLER_20_1831 ();
 b15zdnd11an1n16x5 FILLER_20_1838 ();
 b15zdnd11an1n04x5 FILLER_20_1854 ();
 b15zdnd11an1n16x5 FILLER_20_1872 ();
 b15zdnd00an1n02x5 FILLER_20_1888 ();
 b15zdnd11an1n08x5 FILLER_20_1896 ();
 b15zdnd11an1n04x5 FILLER_20_1904 ();
 b15zdnd00an1n02x5 FILLER_20_1908 ();
 b15zdnd11an1n08x5 FILLER_20_1924 ();
 b15zdnd00an1n02x5 FILLER_20_1932 ();
 b15zdnd00an1n01x5 FILLER_20_1934 ();
 b15zdnd11an1n16x5 FILLER_20_1951 ();
 b15zdnd00an1n02x5 FILLER_20_1967 ();
 b15zdnd00an1n01x5 FILLER_20_1969 ();
 b15zdnd11an1n08x5 FILLER_20_1982 ();
 b15zdnd11an1n04x5 FILLER_20_1990 ();
 b15zdnd11an1n04x5 FILLER_20_2001 ();
 b15zdnd00an1n02x5 FILLER_20_2005 ();
 b15zdnd00an1n01x5 FILLER_20_2007 ();
 b15zdnd11an1n32x5 FILLER_20_2015 ();
 b15zdnd00an1n01x5 FILLER_20_2047 ();
 b15zdnd11an1n16x5 FILLER_20_2052 ();
 b15zdnd11an1n08x5 FILLER_20_2068 ();
 b15zdnd00an1n02x5 FILLER_20_2076 ();
 b15zdnd11an1n04x5 FILLER_20_2092 ();
 b15zdnd11an1n32x5 FILLER_20_2101 ();
 b15zdnd11an1n16x5 FILLER_20_2133 ();
 b15zdnd11an1n04x5 FILLER_20_2149 ();
 b15zdnd00an1n01x5 FILLER_20_2153 ();
 b15zdnd11an1n16x5 FILLER_20_2162 ();
 b15zdnd11an1n04x5 FILLER_20_2178 ();
 b15zdnd11an1n16x5 FILLER_20_2189 ();
 b15zdnd11an1n08x5 FILLER_20_2205 ();
 b15zdnd00an1n02x5 FILLER_20_2213 ();
 b15zdnd11an1n32x5 FILLER_20_2231 ();
 b15zdnd11an1n08x5 FILLER_20_2263 ();
 b15zdnd11an1n04x5 FILLER_20_2271 ();
 b15zdnd00an1n01x5 FILLER_20_2275 ();
 b15zdnd11an1n64x5 FILLER_21_0 ();
 b15zdnd11an1n64x5 FILLER_21_64 ();
 b15zdnd00an1n01x5 FILLER_21_128 ();
 b15zdnd11an1n16x5 FILLER_21_143 ();
 b15zdnd11an1n04x5 FILLER_21_159 ();
 b15zdnd00an1n02x5 FILLER_21_163 ();
 b15zdnd11an1n04x5 FILLER_21_175 ();
 b15zdnd00an1n01x5 FILLER_21_179 ();
 b15zdnd11an1n04x5 FILLER_21_200 ();
 b15zdnd11an1n08x5 FILLER_21_214 ();
 b15zdnd11an1n04x5 FILLER_21_222 ();
 b15zdnd00an1n02x5 FILLER_21_226 ();
 b15zdnd00an1n01x5 FILLER_21_228 ();
 b15zdnd11an1n08x5 FILLER_21_234 ();
 b15zdnd00an1n02x5 FILLER_21_242 ();
 b15zdnd11an1n16x5 FILLER_21_258 ();
 b15zdnd11an1n08x5 FILLER_21_274 ();
 b15zdnd00an1n01x5 FILLER_21_282 ();
 b15zdnd11an1n04x5 FILLER_21_295 ();
 b15zdnd11an1n08x5 FILLER_21_314 ();
 b15zdnd11an1n08x5 FILLER_21_330 ();
 b15zdnd11an1n04x5 FILLER_21_338 ();
 b15zdnd00an1n01x5 FILLER_21_342 ();
 b15zdnd11an1n32x5 FILLER_21_357 ();
 b15zdnd11an1n08x5 FILLER_21_389 ();
 b15zdnd11an1n04x5 FILLER_21_397 ();
 b15zdnd00an1n02x5 FILLER_21_401 ();
 b15zdnd00an1n01x5 FILLER_21_403 ();
 b15zdnd11an1n32x5 FILLER_21_418 ();
 b15zdnd00an1n02x5 FILLER_21_450 ();
 b15zdnd11an1n04x5 FILLER_21_458 ();
 b15zdnd11an1n08x5 FILLER_21_468 ();
 b15zdnd11an1n04x5 FILLER_21_476 ();
 b15zdnd00an1n02x5 FILLER_21_480 ();
 b15zdnd00an1n01x5 FILLER_21_482 ();
 b15zdnd11an1n32x5 FILLER_21_490 ();
 b15zdnd00an1n01x5 FILLER_21_522 ();
 b15zdnd11an1n16x5 FILLER_21_529 ();
 b15zdnd11an1n08x5 FILLER_21_545 ();
 b15zdnd11an1n04x5 FILLER_21_553 ();
 b15zdnd00an1n02x5 FILLER_21_557 ();
 b15zdnd11an1n04x5 FILLER_21_563 ();
 b15zdnd11an1n16x5 FILLER_21_583 ();
 b15zdnd11an1n04x5 FILLER_21_605 ();
 b15zdnd11an1n16x5 FILLER_21_619 ();
 b15zdnd11an1n08x5 FILLER_21_635 ();
 b15zdnd00an1n02x5 FILLER_21_643 ();
 b15zdnd11an1n08x5 FILLER_21_666 ();
 b15zdnd11an1n04x5 FILLER_21_674 ();
 b15zdnd00an1n02x5 FILLER_21_678 ();
 b15zdnd11an1n08x5 FILLER_21_696 ();
 b15zdnd11an1n04x5 FILLER_21_704 ();
 b15zdnd00an1n01x5 FILLER_21_708 ();
 b15zdnd11an1n16x5 FILLER_21_715 ();
 b15zdnd11an1n08x5 FILLER_21_731 ();
 b15zdnd11an1n04x5 FILLER_21_739 ();
 b15zdnd00an1n02x5 FILLER_21_743 ();
 b15zdnd11an1n04x5 FILLER_21_752 ();
 b15zdnd11an1n04x5 FILLER_21_773 ();
 b15zdnd11an1n32x5 FILLER_21_789 ();
 b15zdnd00an1n02x5 FILLER_21_821 ();
 b15zdnd11an1n08x5 FILLER_21_829 ();
 b15zdnd00an1n01x5 FILLER_21_837 ();
 b15zdnd11an1n04x5 FILLER_21_844 ();
 b15zdnd11an1n04x5 FILLER_21_854 ();
 b15zdnd11an1n08x5 FILLER_21_884 ();
 b15zdnd00an1n02x5 FILLER_21_892 ();
 b15zdnd11an1n64x5 FILLER_21_899 ();
 b15zdnd11an1n64x5 FILLER_21_963 ();
 b15zdnd11an1n64x5 FILLER_21_1027 ();
 b15zdnd11an1n64x5 FILLER_21_1091 ();
 b15zdnd11an1n64x5 FILLER_21_1155 ();
 b15zdnd11an1n64x5 FILLER_21_1219 ();
 b15zdnd11an1n32x5 FILLER_21_1283 ();
 b15zdnd11an1n04x5 FILLER_21_1315 ();
 b15zdnd00an1n01x5 FILLER_21_1319 ();
 b15zdnd11an1n32x5 FILLER_21_1330 ();
 b15zdnd11an1n04x5 FILLER_21_1362 ();
 b15zdnd00an1n02x5 FILLER_21_1366 ();
 b15zdnd11an1n32x5 FILLER_21_1378 ();
 b15zdnd11an1n08x5 FILLER_21_1410 ();
 b15zdnd11an1n04x5 FILLER_21_1418 ();
 b15zdnd00an1n01x5 FILLER_21_1422 ();
 b15zdnd11an1n04x5 FILLER_21_1444 ();
 b15zdnd11an1n64x5 FILLER_21_1454 ();
 b15zdnd11an1n32x5 FILLER_21_1518 ();
 b15zdnd11an1n04x5 FILLER_21_1550 ();
 b15zdnd00an1n02x5 FILLER_21_1554 ();
 b15zdnd11an1n32x5 FILLER_21_1562 ();
 b15zdnd00an1n02x5 FILLER_21_1594 ();
 b15zdnd00an1n01x5 FILLER_21_1596 ();
 b15zdnd11an1n04x5 FILLER_21_1605 ();
 b15zdnd11an1n04x5 FILLER_21_1625 ();
 b15zdnd11an1n04x5 FILLER_21_1647 ();
 b15zdnd11an1n32x5 FILLER_21_1658 ();
 b15zdnd11an1n16x5 FILLER_21_1690 ();
 b15zdnd11an1n08x5 FILLER_21_1706 ();
 b15zdnd00an1n02x5 FILLER_21_1714 ();
 b15zdnd11an1n08x5 FILLER_21_1742 ();
 b15zdnd11an1n04x5 FILLER_21_1750 ();
 b15zdnd00an1n01x5 FILLER_21_1754 ();
 b15zdnd11an1n08x5 FILLER_21_1760 ();
 b15zdnd11an1n04x5 FILLER_21_1768 ();
 b15zdnd00an1n02x5 FILLER_21_1772 ();
 b15zdnd11an1n32x5 FILLER_21_1780 ();
 b15zdnd11an1n16x5 FILLER_21_1812 ();
 b15zdnd00an1n01x5 FILLER_21_1828 ();
 b15zdnd11an1n04x5 FILLER_21_1843 ();
 b15zdnd00an1n01x5 FILLER_21_1847 ();
 b15zdnd11an1n32x5 FILLER_21_1855 ();
 b15zdnd11an1n04x5 FILLER_21_1887 ();
 b15zdnd00an1n02x5 FILLER_21_1891 ();
 b15zdnd11an1n64x5 FILLER_21_1905 ();
 b15zdnd11an1n08x5 FILLER_21_1969 ();
 b15zdnd00an1n02x5 FILLER_21_1977 ();
 b15zdnd00an1n01x5 FILLER_21_1979 ();
 b15zdnd11an1n04x5 FILLER_21_1995 ();
 b15zdnd00an1n02x5 FILLER_21_1999 ();
 b15zdnd00an1n01x5 FILLER_21_2001 ();
 b15zdnd11an1n64x5 FILLER_21_2012 ();
 b15zdnd11an1n08x5 FILLER_21_2076 ();
 b15zdnd00an1n02x5 FILLER_21_2084 ();
 b15zdnd00an1n01x5 FILLER_21_2086 ();
 b15zdnd11an1n04x5 FILLER_21_2097 ();
 b15zdnd00an1n01x5 FILLER_21_2101 ();
 b15zdnd11an1n32x5 FILLER_21_2128 ();
 b15zdnd11an1n04x5 FILLER_21_2160 ();
 b15zdnd00an1n02x5 FILLER_21_2164 ();
 b15zdnd00an1n01x5 FILLER_21_2166 ();
 b15zdnd11an1n64x5 FILLER_21_2198 ();
 b15zdnd11an1n16x5 FILLER_21_2262 ();
 b15zdnd11an1n04x5 FILLER_21_2278 ();
 b15zdnd00an1n02x5 FILLER_21_2282 ();
 b15zdnd11an1n32x5 FILLER_22_8 ();
 b15zdnd00an1n02x5 FILLER_22_40 ();
 b15zdnd11an1n16x5 FILLER_22_58 ();
 b15zdnd11an1n08x5 FILLER_22_74 ();
 b15zdnd11an1n04x5 FILLER_22_82 ();
 b15zdnd00an1n02x5 FILLER_22_86 ();
 b15zdnd00an1n01x5 FILLER_22_88 ();
 b15zdnd11an1n16x5 FILLER_22_95 ();
 b15zdnd00an1n01x5 FILLER_22_111 ();
 b15zdnd11an1n64x5 FILLER_22_118 ();
 b15zdnd11an1n16x5 FILLER_22_182 ();
 b15zdnd00an1n02x5 FILLER_22_198 ();
 b15zdnd00an1n01x5 FILLER_22_200 ();
 b15zdnd11an1n16x5 FILLER_22_206 ();
 b15zdnd11an1n04x5 FILLER_22_222 ();
 b15zdnd00an1n02x5 FILLER_22_226 ();
 b15zdnd11an1n16x5 FILLER_22_235 ();
 b15zdnd11an1n08x5 FILLER_22_251 ();
 b15zdnd00an1n02x5 FILLER_22_259 ();
 b15zdnd00an1n01x5 FILLER_22_261 ();
 b15zdnd11an1n64x5 FILLER_22_270 ();
 b15zdnd11an1n64x5 FILLER_22_334 ();
 b15zdnd11an1n08x5 FILLER_22_398 ();
 b15zdnd11an1n04x5 FILLER_22_406 ();
 b15zdnd00an1n01x5 FILLER_22_410 ();
 b15zdnd11an1n16x5 FILLER_22_416 ();
 b15zdnd11an1n08x5 FILLER_22_432 ();
 b15zdnd00an1n02x5 FILLER_22_440 ();
 b15zdnd00an1n01x5 FILLER_22_442 ();
 b15zdnd11an1n32x5 FILLER_22_447 ();
 b15zdnd11an1n04x5 FILLER_22_479 ();
 b15zdnd11an1n04x5 FILLER_22_489 ();
 b15zdnd00an1n02x5 FILLER_22_493 ();
 b15zdnd11an1n08x5 FILLER_22_510 ();
 b15zdnd11an1n04x5 FILLER_22_518 ();
 b15zdnd11an1n16x5 FILLER_22_536 ();
 b15zdnd11an1n08x5 FILLER_22_552 ();
 b15zdnd11an1n04x5 FILLER_22_560 ();
 b15zdnd11an1n08x5 FILLER_22_581 ();
 b15zdnd11an1n04x5 FILLER_22_589 ();
 b15zdnd11an1n64x5 FILLER_22_602 ();
 b15zdnd11an1n08x5 FILLER_22_666 ();
 b15zdnd11an1n04x5 FILLER_22_674 ();
 b15zdnd00an1n02x5 FILLER_22_678 ();
 b15zdnd00an1n01x5 FILLER_22_680 ();
 b15zdnd11an1n32x5 FILLER_22_685 ();
 b15zdnd00an1n01x5 FILLER_22_717 ();
 b15zdnd11an1n04x5 FILLER_22_726 ();
 b15zdnd00an1n02x5 FILLER_22_730 ();
 b15zdnd00an1n01x5 FILLER_22_732 ();
 b15zdnd11an1n32x5 FILLER_22_742 ();
 b15zdnd11an1n16x5 FILLER_22_774 ();
 b15zdnd11an1n08x5 FILLER_22_790 ();
 b15zdnd11an1n04x5 FILLER_22_798 ();
 b15zdnd00an1n01x5 FILLER_22_802 ();
 b15zdnd11an1n08x5 FILLER_22_811 ();
 b15zdnd11an1n04x5 FILLER_22_819 ();
 b15zdnd11an1n64x5 FILLER_22_830 ();
 b15zdnd00an1n02x5 FILLER_22_894 ();
 b15zdnd00an1n01x5 FILLER_22_896 ();
 b15zdnd11an1n16x5 FILLER_22_904 ();
 b15zdnd11an1n04x5 FILLER_22_920 ();
 b15zdnd00an1n02x5 FILLER_22_924 ();
 b15zdnd00an1n01x5 FILLER_22_926 ();
 b15zdnd11an1n64x5 FILLER_22_947 ();
 b15zdnd11an1n16x5 FILLER_22_1011 ();
 b15zdnd00an1n01x5 FILLER_22_1027 ();
 b15zdnd11an1n08x5 FILLER_22_1033 ();
 b15zdnd00an1n02x5 FILLER_22_1041 ();
 b15zdnd00an1n01x5 FILLER_22_1043 ();
 b15zdnd11an1n16x5 FILLER_22_1047 ();
 b15zdnd11an1n04x5 FILLER_22_1063 ();
 b15zdnd11an1n16x5 FILLER_22_1072 ();
 b15zdnd11an1n08x5 FILLER_22_1088 ();
 b15zdnd11an1n04x5 FILLER_22_1096 ();
 b15zdnd00an1n02x5 FILLER_22_1100 ();
 b15zdnd00an1n01x5 FILLER_22_1102 ();
 b15zdnd11an1n32x5 FILLER_22_1107 ();
 b15zdnd00an1n02x5 FILLER_22_1139 ();
 b15zdnd00an1n01x5 FILLER_22_1141 ();
 b15zdnd11an1n64x5 FILLER_22_1146 ();
 b15zdnd11an1n32x5 FILLER_22_1210 ();
 b15zdnd11an1n16x5 FILLER_22_1242 ();
 b15zdnd11an1n08x5 FILLER_22_1258 ();
 b15zdnd00an1n02x5 FILLER_22_1266 ();
 b15zdnd11an1n16x5 FILLER_22_1288 ();
 b15zdnd11an1n08x5 FILLER_22_1304 ();
 b15zdnd00an1n02x5 FILLER_22_1312 ();
 b15zdnd11an1n32x5 FILLER_22_1332 ();
 b15zdnd11an1n04x5 FILLER_22_1364 ();
 b15zdnd11an1n16x5 FILLER_22_1386 ();
 b15zdnd11an1n04x5 FILLER_22_1402 ();
 b15zdnd11an1n32x5 FILLER_22_1410 ();
 b15zdnd11an1n04x5 FILLER_22_1442 ();
 b15zdnd00an1n02x5 FILLER_22_1446 ();
 b15zdnd00an1n01x5 FILLER_22_1448 ();
 b15zdnd11an1n04x5 FILLER_22_1461 ();
 b15zdnd11an1n64x5 FILLER_22_1472 ();
 b15zdnd11an1n16x5 FILLER_22_1536 ();
 b15zdnd11an1n04x5 FILLER_22_1552 ();
 b15zdnd00an1n01x5 FILLER_22_1556 ();
 b15zdnd11an1n16x5 FILLER_22_1570 ();
 b15zdnd11an1n04x5 FILLER_22_1586 ();
 b15zdnd00an1n02x5 FILLER_22_1590 ();
 b15zdnd11an1n04x5 FILLER_22_1602 ();
 b15zdnd00an1n02x5 FILLER_22_1606 ();
 b15zdnd11an1n04x5 FILLER_22_1618 ();
 b15zdnd00an1n01x5 FILLER_22_1622 ();
 b15zdnd11an1n04x5 FILLER_22_1630 ();
 b15zdnd11an1n08x5 FILLER_22_1654 ();
 b15zdnd00an1n02x5 FILLER_22_1662 ();
 b15zdnd00an1n01x5 FILLER_22_1664 ();
 b15zdnd11an1n64x5 FILLER_22_1681 ();
 b15zdnd11an1n16x5 FILLER_22_1758 ();
 b15zdnd11an1n04x5 FILLER_22_1774 ();
 b15zdnd00an1n01x5 FILLER_22_1778 ();
 b15zdnd11an1n04x5 FILLER_22_1784 ();
 b15zdnd11an1n64x5 FILLER_22_1800 ();
 b15zdnd11an1n64x5 FILLER_22_1864 ();
 b15zdnd11an1n64x5 FILLER_22_1928 ();
 b15zdnd11an1n16x5 FILLER_22_1992 ();
 b15zdnd11an1n04x5 FILLER_22_2008 ();
 b15zdnd00an1n02x5 FILLER_22_2012 ();
 b15zdnd00an1n01x5 FILLER_22_2014 ();
 b15zdnd11an1n04x5 FILLER_22_2041 ();
 b15zdnd11an1n64x5 FILLER_22_2051 ();
 b15zdnd11an1n08x5 FILLER_22_2115 ();
 b15zdnd11an1n04x5 FILLER_22_2123 ();
 b15zdnd00an1n02x5 FILLER_22_2127 ();
 b15zdnd00an1n01x5 FILLER_22_2129 ();
 b15zdnd11an1n08x5 FILLER_22_2139 ();
 b15zdnd11an1n04x5 FILLER_22_2147 ();
 b15zdnd00an1n02x5 FILLER_22_2151 ();
 b15zdnd00an1n01x5 FILLER_22_2153 ();
 b15zdnd11an1n16x5 FILLER_22_2162 ();
 b15zdnd11an1n08x5 FILLER_22_2178 ();
 b15zdnd00an1n02x5 FILLER_22_2186 ();
 b15zdnd00an1n01x5 FILLER_22_2188 ();
 b15zdnd11an1n64x5 FILLER_22_2203 ();
 b15zdnd11an1n08x5 FILLER_22_2267 ();
 b15zdnd00an1n01x5 FILLER_22_2275 ();
 b15zdnd11an1n32x5 FILLER_23_0 ();
 b15zdnd11an1n08x5 FILLER_23_32 ();
 b15zdnd11an1n04x5 FILLER_23_40 ();
 b15zdnd00an1n01x5 FILLER_23_44 ();
 b15zdnd11an1n08x5 FILLER_23_77 ();
 b15zdnd00an1n02x5 FILLER_23_85 ();
 b15zdnd00an1n01x5 FILLER_23_87 ();
 b15zdnd11an1n04x5 FILLER_23_92 ();
 b15zdnd11an1n08x5 FILLER_23_107 ();
 b15zdnd11an1n04x5 FILLER_23_120 ();
 b15zdnd11an1n08x5 FILLER_23_140 ();
 b15zdnd11an1n04x5 FILLER_23_148 ();
 b15zdnd00an1n02x5 FILLER_23_152 ();
 b15zdnd11an1n04x5 FILLER_23_166 ();
 b15zdnd11an1n16x5 FILLER_23_176 ();
 b15zdnd11an1n08x5 FILLER_23_192 ();
 b15zdnd00an1n02x5 FILLER_23_200 ();
 b15zdnd00an1n01x5 FILLER_23_202 ();
 b15zdnd11an1n64x5 FILLER_23_210 ();
 b15zdnd11an1n32x5 FILLER_23_274 ();
 b15zdnd11an1n08x5 FILLER_23_306 ();
 b15zdnd11an1n04x5 FILLER_23_314 ();
 b15zdnd11an1n64x5 FILLER_23_338 ();
 b15zdnd11an1n64x5 FILLER_23_402 ();
 b15zdnd11an1n16x5 FILLER_23_466 ();
 b15zdnd11an1n04x5 FILLER_23_482 ();
 b15zdnd11an1n16x5 FILLER_23_495 ();
 b15zdnd11an1n04x5 FILLER_23_511 ();
 b15zdnd00an1n02x5 FILLER_23_515 ();
 b15zdnd11an1n32x5 FILLER_23_533 ();
 b15zdnd00an1n02x5 FILLER_23_565 ();
 b15zdnd00an1n01x5 FILLER_23_567 ();
 b15zdnd11an1n64x5 FILLER_23_575 ();
 b15zdnd11an1n08x5 FILLER_23_639 ();
 b15zdnd11an1n04x5 FILLER_23_647 ();
 b15zdnd11an1n08x5 FILLER_23_663 ();
 b15zdnd11an1n04x5 FILLER_23_671 ();
 b15zdnd00an1n01x5 FILLER_23_675 ();
 b15zdnd11an1n04x5 FILLER_23_683 ();
 b15zdnd00an1n02x5 FILLER_23_687 ();
 b15zdnd11an1n32x5 FILLER_23_694 ();
 b15zdnd11an1n04x5 FILLER_23_726 ();
 b15zdnd00an1n01x5 FILLER_23_730 ();
 b15zdnd11an1n04x5 FILLER_23_737 ();
 b15zdnd11an1n32x5 FILLER_23_745 ();
 b15zdnd00an1n01x5 FILLER_23_777 ();
 b15zdnd11an1n32x5 FILLER_23_798 ();
 b15zdnd11an1n16x5 FILLER_23_830 ();
 b15zdnd00an1n02x5 FILLER_23_846 ();
 b15zdnd00an1n01x5 FILLER_23_848 ();
 b15zdnd11an1n64x5 FILLER_23_863 ();
 b15zdnd11an1n32x5 FILLER_23_927 ();
 b15zdnd11an1n16x5 FILLER_23_959 ();
 b15zdnd11an1n08x5 FILLER_23_975 ();
 b15zdnd11an1n08x5 FILLER_23_987 ();
 b15zdnd11an1n16x5 FILLER_23_1006 ();
 b15zdnd11an1n04x5 FILLER_23_1022 ();
 b15zdnd00an1n02x5 FILLER_23_1026 ();
 b15zdnd00an1n01x5 FILLER_23_1028 ();
 b15zdnd11an1n16x5 FILLER_23_1049 ();
 b15zdnd11an1n04x5 FILLER_23_1065 ();
 b15zdnd11an1n08x5 FILLER_23_1089 ();
 b15zdnd00an1n02x5 FILLER_23_1097 ();
 b15zdnd11an1n32x5 FILLER_23_1104 ();
 b15zdnd00an1n02x5 FILLER_23_1136 ();
 b15zdnd11an1n16x5 FILLER_23_1143 ();
 b15zdnd11an1n04x5 FILLER_23_1159 ();
 b15zdnd11an1n04x5 FILLER_23_1183 ();
 b15zdnd00an1n02x5 FILLER_23_1187 ();
 b15zdnd00an1n01x5 FILLER_23_1189 ();
 b15zdnd11an1n16x5 FILLER_23_1194 ();
 b15zdnd11an1n08x5 FILLER_23_1210 ();
 b15zdnd00an1n02x5 FILLER_23_1218 ();
 b15zdnd00an1n01x5 FILLER_23_1220 ();
 b15zdnd11an1n04x5 FILLER_23_1241 ();
 b15zdnd00an1n02x5 FILLER_23_1245 ();
 b15zdnd11an1n32x5 FILLER_23_1252 ();
 b15zdnd11an1n08x5 FILLER_23_1284 ();
 b15zdnd11an1n16x5 FILLER_23_1315 ();
 b15zdnd11an1n04x5 FILLER_23_1331 ();
 b15zdnd11an1n16x5 FILLER_23_1339 ();
 b15zdnd11an1n04x5 FILLER_23_1355 ();
 b15zdnd11an1n32x5 FILLER_23_1364 ();
 b15zdnd00an1n02x5 FILLER_23_1396 ();
 b15zdnd11an1n32x5 FILLER_23_1412 ();
 b15zdnd11an1n16x5 FILLER_23_1444 ();
 b15zdnd11an1n08x5 FILLER_23_1460 ();
 b15zdnd11an1n32x5 FILLER_23_1474 ();
 b15zdnd11an1n04x5 FILLER_23_1506 ();
 b15zdnd00an1n01x5 FILLER_23_1510 ();
 b15zdnd11an1n04x5 FILLER_23_1523 ();
 b15zdnd11an1n16x5 FILLER_23_1533 ();
 b15zdnd11an1n08x5 FILLER_23_1549 ();
 b15zdnd00an1n02x5 FILLER_23_1557 ();
 b15zdnd00an1n01x5 FILLER_23_1559 ();
 b15zdnd11an1n16x5 FILLER_23_1570 ();
 b15zdnd11an1n08x5 FILLER_23_1586 ();
 b15zdnd11an1n32x5 FILLER_23_1606 ();
 b15zdnd00an1n02x5 FILLER_23_1638 ();
 b15zdnd00an1n01x5 FILLER_23_1640 ();
 b15zdnd11an1n08x5 FILLER_23_1665 ();
 b15zdnd11an1n16x5 FILLER_23_1693 ();
 b15zdnd11an1n08x5 FILLER_23_1709 ();
 b15zdnd00an1n02x5 FILLER_23_1717 ();
 b15zdnd11an1n16x5 FILLER_23_1745 ();
 b15zdnd00an1n01x5 FILLER_23_1761 ();
 b15zdnd11an1n08x5 FILLER_23_1773 ();
 b15zdnd11an1n04x5 FILLER_23_1781 ();
 b15zdnd00an1n01x5 FILLER_23_1785 ();
 b15zdnd11an1n04x5 FILLER_23_1805 ();
 b15zdnd11an1n16x5 FILLER_23_1819 ();
 b15zdnd11an1n04x5 FILLER_23_1835 ();
 b15zdnd00an1n02x5 FILLER_23_1839 ();
 b15zdnd00an1n01x5 FILLER_23_1841 ();
 b15zdnd11an1n32x5 FILLER_23_1852 ();
 b15zdnd11an1n16x5 FILLER_23_1884 ();
 b15zdnd11an1n08x5 FILLER_23_1900 ();
 b15zdnd00an1n02x5 FILLER_23_1908 ();
 b15zdnd11an1n04x5 FILLER_23_1928 ();
 b15zdnd11an1n08x5 FILLER_23_1958 ();
 b15zdnd11an1n04x5 FILLER_23_1966 ();
 b15zdnd11an1n32x5 FILLER_23_1978 ();
 b15zdnd11an1n16x5 FILLER_23_2010 ();
 b15zdnd11an1n04x5 FILLER_23_2026 ();
 b15zdnd11an1n08x5 FILLER_23_2035 ();
 b15zdnd00an1n02x5 FILLER_23_2043 ();
 b15zdnd11an1n32x5 FILLER_23_2057 ();
 b15zdnd11an1n04x5 FILLER_23_2089 ();
 b15zdnd00an1n02x5 FILLER_23_2093 ();
 b15zdnd11an1n64x5 FILLER_23_2110 ();
 b15zdnd11an1n64x5 FILLER_23_2174 ();
 b15zdnd11an1n32x5 FILLER_23_2238 ();
 b15zdnd11an1n08x5 FILLER_23_2270 ();
 b15zdnd11an1n04x5 FILLER_23_2278 ();
 b15zdnd00an1n02x5 FILLER_23_2282 ();
 b15zdnd11an1n32x5 FILLER_24_8 ();
 b15zdnd11an1n04x5 FILLER_24_40 ();
 b15zdnd00an1n02x5 FILLER_24_44 ();
 b15zdnd00an1n01x5 FILLER_24_46 ();
 b15zdnd11an1n16x5 FILLER_24_63 ();
 b15zdnd11an1n04x5 FILLER_24_79 ();
 b15zdnd00an1n01x5 FILLER_24_83 ();
 b15zdnd11an1n32x5 FILLER_24_92 ();
 b15zdnd00an1n01x5 FILLER_24_124 ();
 b15zdnd11an1n32x5 FILLER_24_134 ();
 b15zdnd00an1n02x5 FILLER_24_166 ();
 b15zdnd00an1n01x5 FILLER_24_168 ();
 b15zdnd11an1n64x5 FILLER_24_174 ();
 b15zdnd11an1n32x5 FILLER_24_238 ();
 b15zdnd11an1n04x5 FILLER_24_270 ();
 b15zdnd11an1n64x5 FILLER_24_279 ();
 b15zdnd11an1n64x5 FILLER_24_343 ();
 b15zdnd11an1n64x5 FILLER_24_407 ();
 b15zdnd11an1n32x5 FILLER_24_471 ();
 b15zdnd11an1n16x5 FILLER_24_503 ();
 b15zdnd11an1n04x5 FILLER_24_519 ();
 b15zdnd00an1n01x5 FILLER_24_523 ();
 b15zdnd11an1n08x5 FILLER_24_532 ();
 b15zdnd11an1n04x5 FILLER_24_540 ();
 b15zdnd00an1n02x5 FILLER_24_544 ();
 b15zdnd00an1n01x5 FILLER_24_546 ();
 b15zdnd11an1n08x5 FILLER_24_559 ();
 b15zdnd00an1n01x5 FILLER_24_567 ();
 b15zdnd11an1n32x5 FILLER_24_580 ();
 b15zdnd11an1n16x5 FILLER_24_612 ();
 b15zdnd11an1n08x5 FILLER_24_628 ();
 b15zdnd00an1n02x5 FILLER_24_636 ();
 b15zdnd11an1n32x5 FILLER_24_656 ();
 b15zdnd11an1n04x5 FILLER_24_688 ();
 b15zdnd00an1n02x5 FILLER_24_692 ();
 b15zdnd11an1n04x5 FILLER_24_701 ();
 b15zdnd00an1n02x5 FILLER_24_716 ();
 b15zdnd11an1n16x5 FILLER_24_726 ();
 b15zdnd00an1n02x5 FILLER_24_742 ();
 b15zdnd11an1n16x5 FILLER_24_757 ();
 b15zdnd11an1n08x5 FILLER_24_773 ();
 b15zdnd11an1n04x5 FILLER_24_781 ();
 b15zdnd11an1n64x5 FILLER_24_794 ();
 b15zdnd11an1n08x5 FILLER_24_863 ();
 b15zdnd00an1n01x5 FILLER_24_871 ();
 b15zdnd11an1n04x5 FILLER_24_882 ();
 b15zdnd11an1n64x5 FILLER_24_897 ();
 b15zdnd11an1n16x5 FILLER_24_961 ();
 b15zdnd11an1n04x5 FILLER_24_977 ();
 b15zdnd11an1n08x5 FILLER_24_986 ();
 b15zdnd11an1n04x5 FILLER_24_994 ();
 b15zdnd11an1n64x5 FILLER_24_1018 ();
 b15zdnd11an1n16x5 FILLER_24_1082 ();
 b15zdnd00an1n02x5 FILLER_24_1098 ();
 b15zdnd00an1n01x5 FILLER_24_1100 ();
 b15zdnd11an1n08x5 FILLER_24_1121 ();
 b15zdnd11an1n04x5 FILLER_24_1129 ();
 b15zdnd00an1n01x5 FILLER_24_1133 ();
 b15zdnd11an1n32x5 FILLER_24_1154 ();
 b15zdnd11an1n16x5 FILLER_24_1186 ();
 b15zdnd11an1n08x5 FILLER_24_1202 ();
 b15zdnd11an1n04x5 FILLER_24_1210 ();
 b15zdnd00an1n02x5 FILLER_24_1214 ();
 b15zdnd00an1n01x5 FILLER_24_1216 ();
 b15zdnd11an1n04x5 FILLER_24_1237 ();
 b15zdnd11an1n32x5 FILLER_24_1245 ();
 b15zdnd11an1n16x5 FILLER_24_1277 ();
 b15zdnd11an1n08x5 FILLER_24_1293 ();
 b15zdnd11an1n08x5 FILLER_24_1321 ();
 b15zdnd11an1n04x5 FILLER_24_1329 ();
 b15zdnd11an1n04x5 FILLER_24_1345 ();
 b15zdnd00an1n02x5 FILLER_24_1349 ();
 b15zdnd00an1n01x5 FILLER_24_1351 ();
 b15zdnd11an1n16x5 FILLER_24_1364 ();
 b15zdnd00an1n02x5 FILLER_24_1380 ();
 b15zdnd00an1n01x5 FILLER_24_1382 ();
 b15zdnd11an1n08x5 FILLER_24_1406 ();
 b15zdnd11an1n04x5 FILLER_24_1414 ();
 b15zdnd11an1n32x5 FILLER_24_1426 ();
 b15zdnd11an1n16x5 FILLER_24_1458 ();
 b15zdnd11an1n04x5 FILLER_24_1474 ();
 b15zdnd00an1n02x5 FILLER_24_1478 ();
 b15zdnd11an1n16x5 FILLER_24_1491 ();
 b15zdnd11an1n08x5 FILLER_24_1507 ();
 b15zdnd11an1n04x5 FILLER_24_1515 ();
 b15zdnd00an1n02x5 FILLER_24_1519 ();
 b15zdnd11an1n64x5 FILLER_24_1527 ();
 b15zdnd11an1n64x5 FILLER_24_1591 ();
 b15zdnd11an1n64x5 FILLER_24_1655 ();
 b15zdnd11an1n16x5 FILLER_24_1719 ();
 b15zdnd11an1n08x5 FILLER_24_1735 ();
 b15zdnd11an1n04x5 FILLER_24_1743 ();
 b15zdnd00an1n02x5 FILLER_24_1747 ();
 b15zdnd11an1n04x5 FILLER_24_1754 ();
 b15zdnd00an1n02x5 FILLER_24_1758 ();
 b15zdnd11an1n32x5 FILLER_24_1769 ();
 b15zdnd11an1n08x5 FILLER_24_1808 ();
 b15zdnd00an1n02x5 FILLER_24_1816 ();
 b15zdnd11an1n16x5 FILLER_24_1824 ();
 b15zdnd11an1n04x5 FILLER_24_1840 ();
 b15zdnd00an1n02x5 FILLER_24_1844 ();
 b15zdnd00an1n01x5 FILLER_24_1846 ();
 b15zdnd11an1n16x5 FILLER_24_1858 ();
 b15zdnd11an1n08x5 FILLER_24_1889 ();
 b15zdnd00an1n02x5 FILLER_24_1897 ();
 b15zdnd11an1n08x5 FILLER_24_1913 ();
 b15zdnd11an1n04x5 FILLER_24_1935 ();
 b15zdnd00an1n02x5 FILLER_24_1939 ();
 b15zdnd00an1n01x5 FILLER_24_1941 ();
 b15zdnd11an1n04x5 FILLER_24_1947 ();
 b15zdnd11an1n16x5 FILLER_24_1958 ();
 b15zdnd11an1n08x5 FILLER_24_1974 ();
 b15zdnd11an1n04x5 FILLER_24_1982 ();
 b15zdnd11an1n32x5 FILLER_24_2000 ();
 b15zdnd11an1n04x5 FILLER_24_2032 ();
 b15zdnd00an1n02x5 FILLER_24_2036 ();
 b15zdnd00an1n01x5 FILLER_24_2038 ();
 b15zdnd11an1n04x5 FILLER_24_2044 ();
 b15zdnd00an1n02x5 FILLER_24_2048 ();
 b15zdnd11an1n32x5 FILLER_24_2057 ();
 b15zdnd11an1n16x5 FILLER_24_2089 ();
 b15zdnd11an1n08x5 FILLER_24_2105 ();
 b15zdnd00an1n02x5 FILLER_24_2113 ();
 b15zdnd11an1n04x5 FILLER_24_2129 ();
 b15zdnd11an1n16x5 FILLER_24_2137 ();
 b15zdnd00an1n01x5 FILLER_24_2153 ();
 b15zdnd11an1n32x5 FILLER_24_2162 ();
 b15zdnd00an1n02x5 FILLER_24_2194 ();
 b15zdnd00an1n01x5 FILLER_24_2196 ();
 b15zdnd11an1n64x5 FILLER_24_2205 ();
 b15zdnd11an1n04x5 FILLER_24_2269 ();
 b15zdnd00an1n02x5 FILLER_24_2273 ();
 b15zdnd00an1n01x5 FILLER_24_2275 ();
 b15zdnd11an1n32x5 FILLER_25_0 ();
 b15zdnd11an1n08x5 FILLER_25_32 ();
 b15zdnd11an1n04x5 FILLER_25_40 ();
 b15zdnd00an1n02x5 FILLER_25_44 ();
 b15zdnd00an1n01x5 FILLER_25_46 ();
 b15zdnd11an1n04x5 FILLER_25_65 ();
 b15zdnd11an1n64x5 FILLER_25_87 ();
 b15zdnd11an1n04x5 FILLER_25_151 ();
 b15zdnd11an1n16x5 FILLER_25_170 ();
 b15zdnd11an1n08x5 FILLER_25_186 ();
 b15zdnd00an1n02x5 FILLER_25_194 ();
 b15zdnd11an1n32x5 FILLER_25_202 ();
 b15zdnd11an1n08x5 FILLER_25_234 ();
 b15zdnd11an1n04x5 FILLER_25_242 ();
 b15zdnd11an1n04x5 FILLER_25_252 ();
 b15zdnd11an1n04x5 FILLER_25_264 ();
 b15zdnd11an1n32x5 FILLER_25_275 ();
 b15zdnd11an1n16x5 FILLER_25_307 ();
 b15zdnd11an1n04x5 FILLER_25_323 ();
 b15zdnd00an1n01x5 FILLER_25_327 ();
 b15zdnd11an1n04x5 FILLER_25_333 ();
 b15zdnd11an1n04x5 FILLER_25_351 ();
 b15zdnd11an1n32x5 FILLER_25_386 ();
 b15zdnd11an1n04x5 FILLER_25_418 ();
 b15zdnd00an1n01x5 FILLER_25_422 ();
 b15zdnd11an1n16x5 FILLER_25_432 ();
 b15zdnd11an1n08x5 FILLER_25_448 ();
 b15zdnd00an1n02x5 FILLER_25_456 ();
 b15zdnd00an1n01x5 FILLER_25_458 ();
 b15zdnd11an1n64x5 FILLER_25_471 ();
 b15zdnd11an1n04x5 FILLER_25_535 ();
 b15zdnd11an1n04x5 FILLER_25_563 ();
 b15zdnd11an1n16x5 FILLER_25_573 ();
 b15zdnd11an1n08x5 FILLER_25_589 ();
 b15zdnd11an1n04x5 FILLER_25_597 ();
 b15zdnd00an1n02x5 FILLER_25_601 ();
 b15zdnd00an1n01x5 FILLER_25_603 ();
 b15zdnd11an1n16x5 FILLER_25_610 ();
 b15zdnd11an1n08x5 FILLER_25_626 ();
 b15zdnd11an1n04x5 FILLER_25_634 ();
 b15zdnd11an1n32x5 FILLER_25_655 ();
 b15zdnd11an1n08x5 FILLER_25_687 ();
 b15zdnd11an1n32x5 FILLER_25_706 ();
 b15zdnd11an1n08x5 FILLER_25_738 ();
 b15zdnd00an1n02x5 FILLER_25_746 ();
 b15zdnd00an1n01x5 FILLER_25_748 ();
 b15zdnd11an1n16x5 FILLER_25_764 ();
 b15zdnd00an1n02x5 FILLER_25_780 ();
 b15zdnd11an1n04x5 FILLER_25_787 ();
 b15zdnd11an1n32x5 FILLER_25_807 ();
 b15zdnd11an1n04x5 FILLER_25_839 ();
 b15zdnd11an1n04x5 FILLER_25_847 ();
 b15zdnd00an1n01x5 FILLER_25_851 ();
 b15zdnd11an1n16x5 FILLER_25_861 ();
 b15zdnd11an1n08x5 FILLER_25_877 ();
 b15zdnd00an1n02x5 FILLER_25_885 ();
 b15zdnd00an1n01x5 FILLER_25_887 ();
 b15zdnd11an1n04x5 FILLER_25_894 ();
 b15zdnd11an1n64x5 FILLER_25_902 ();
 b15zdnd11an1n04x5 FILLER_25_966 ();
 b15zdnd00an1n01x5 FILLER_25_970 ();
 b15zdnd11an1n04x5 FILLER_25_991 ();
 b15zdnd11an1n64x5 FILLER_25_1004 ();
 b15zdnd11an1n16x5 FILLER_25_1068 ();
 b15zdnd11an1n08x5 FILLER_25_1084 ();
 b15zdnd11an1n04x5 FILLER_25_1092 ();
 b15zdnd00an1n02x5 FILLER_25_1096 ();
 b15zdnd11an1n16x5 FILLER_25_1107 ();
 b15zdnd11an1n08x5 FILLER_25_1123 ();
 b15zdnd11an1n04x5 FILLER_25_1131 ();
 b15zdnd00an1n02x5 FILLER_25_1135 ();
 b15zdnd00an1n01x5 FILLER_25_1137 ();
 b15zdnd11an1n64x5 FILLER_25_1141 ();
 b15zdnd11an1n64x5 FILLER_25_1205 ();
 b15zdnd11an1n64x5 FILLER_25_1269 ();
 b15zdnd11an1n16x5 FILLER_25_1333 ();
 b15zdnd11an1n64x5 FILLER_25_1354 ();
 b15zdnd11an1n32x5 FILLER_25_1418 ();
 b15zdnd11an1n04x5 FILLER_25_1450 ();
 b15zdnd00an1n02x5 FILLER_25_1454 ();
 b15zdnd11an1n32x5 FILLER_25_1473 ();
 b15zdnd11an1n08x5 FILLER_25_1505 ();
 b15zdnd11an1n04x5 FILLER_25_1513 ();
 b15zdnd00an1n01x5 FILLER_25_1517 ();
 b15zdnd11an1n16x5 FILLER_25_1533 ();
 b15zdnd11an1n08x5 FILLER_25_1549 ();
 b15zdnd11an1n04x5 FILLER_25_1557 ();
 b15zdnd11an1n64x5 FILLER_25_1573 ();
 b15zdnd11an1n64x5 FILLER_25_1637 ();
 b15zdnd11an1n32x5 FILLER_25_1701 ();
 b15zdnd11an1n08x5 FILLER_25_1733 ();
 b15zdnd00an1n01x5 FILLER_25_1741 ();
 b15zdnd11an1n04x5 FILLER_25_1749 ();
 b15zdnd00an1n01x5 FILLER_25_1753 ();
 b15zdnd11an1n64x5 FILLER_25_1763 ();
 b15zdnd11an1n64x5 FILLER_25_1827 ();
 b15zdnd11an1n32x5 FILLER_25_1891 ();
 b15zdnd11an1n08x5 FILLER_25_1923 ();
 b15zdnd11an1n32x5 FILLER_25_1935 ();
 b15zdnd11an1n04x5 FILLER_25_1967 ();
 b15zdnd00an1n01x5 FILLER_25_1971 ();
 b15zdnd11an1n32x5 FILLER_25_1980 ();
 b15zdnd11an1n04x5 FILLER_25_2022 ();
 b15zdnd11an1n08x5 FILLER_25_2039 ();
 b15zdnd11an1n04x5 FILLER_25_2047 ();
 b15zdnd00an1n01x5 FILLER_25_2051 ();
 b15zdnd11an1n32x5 FILLER_25_2072 ();
 b15zdnd11an1n04x5 FILLER_25_2120 ();
 b15zdnd11an1n32x5 FILLER_25_2129 ();
 b15zdnd11an1n04x5 FILLER_25_2161 ();
 b15zdnd00an1n02x5 FILLER_25_2165 ();
 b15zdnd11an1n16x5 FILLER_25_2171 ();
 b15zdnd00an1n01x5 FILLER_25_2187 ();
 b15zdnd11an1n04x5 FILLER_25_2192 ();
 b15zdnd00an1n01x5 FILLER_25_2196 ();
 b15zdnd11an1n04x5 FILLER_25_2207 ();
 b15zdnd11an1n64x5 FILLER_25_2215 ();
 b15zdnd11an1n04x5 FILLER_25_2279 ();
 b15zdnd00an1n01x5 FILLER_25_2283 ();
 b15zdnd11an1n64x5 FILLER_26_8 ();
 b15zdnd11an1n32x5 FILLER_26_72 ();
 b15zdnd11an1n16x5 FILLER_26_104 ();
 b15zdnd11an1n04x5 FILLER_26_120 ();
 b15zdnd00an1n01x5 FILLER_26_124 ();
 b15zdnd11an1n04x5 FILLER_26_129 ();
 b15zdnd11an1n04x5 FILLER_26_139 ();
 b15zdnd11an1n32x5 FILLER_26_157 ();
 b15zdnd00an1n02x5 FILLER_26_189 ();
 b15zdnd11an1n04x5 FILLER_26_196 ();
 b15zdnd11an1n04x5 FILLER_26_205 ();
 b15zdnd11an1n32x5 FILLER_26_217 ();
 b15zdnd11an1n16x5 FILLER_26_249 ();
 b15zdnd11an1n04x5 FILLER_26_265 ();
 b15zdnd00an1n02x5 FILLER_26_269 ();
 b15zdnd00an1n01x5 FILLER_26_271 ();
 b15zdnd11an1n16x5 FILLER_26_286 ();
 b15zdnd00an1n02x5 FILLER_26_302 ();
 b15zdnd00an1n01x5 FILLER_26_304 ();
 b15zdnd11an1n04x5 FILLER_26_326 ();
 b15zdnd11an1n64x5 FILLER_26_336 ();
 b15zdnd11an1n16x5 FILLER_26_400 ();
 b15zdnd11an1n08x5 FILLER_26_416 ();
 b15zdnd00an1n02x5 FILLER_26_424 ();
 b15zdnd11an1n04x5 FILLER_26_456 ();
 b15zdnd11an1n04x5 FILLER_26_472 ();
 b15zdnd11an1n32x5 FILLER_26_483 ();
 b15zdnd11an1n16x5 FILLER_26_515 ();
 b15zdnd11an1n08x5 FILLER_26_531 ();
 b15zdnd00an1n02x5 FILLER_26_539 ();
 b15zdnd00an1n01x5 FILLER_26_541 ();
 b15zdnd11an1n64x5 FILLER_26_554 ();
 b15zdnd11an1n16x5 FILLER_26_618 ();
 b15zdnd11an1n08x5 FILLER_26_634 ();
 b15zdnd00an1n02x5 FILLER_26_642 ();
 b15zdnd00an1n01x5 FILLER_26_644 ();
 b15zdnd11an1n32x5 FILLER_26_657 ();
 b15zdnd11an1n16x5 FILLER_26_689 ();
 b15zdnd00an1n02x5 FILLER_26_705 ();
 b15zdnd00an1n01x5 FILLER_26_707 ();
 b15zdnd00an1n02x5 FILLER_26_716 ();
 b15zdnd11an1n08x5 FILLER_26_726 ();
 b15zdnd11an1n04x5 FILLER_26_734 ();
 b15zdnd00an1n02x5 FILLER_26_738 ();
 b15zdnd11an1n32x5 FILLER_26_748 ();
 b15zdnd11an1n16x5 FILLER_26_780 ();
 b15zdnd00an1n01x5 FILLER_26_796 ();
 b15zdnd11an1n16x5 FILLER_26_807 ();
 b15zdnd11an1n08x5 FILLER_26_823 ();
 b15zdnd11an1n04x5 FILLER_26_831 ();
 b15zdnd00an1n02x5 FILLER_26_835 ();
 b15zdnd00an1n01x5 FILLER_26_837 ();
 b15zdnd11an1n32x5 FILLER_26_849 ();
 b15zdnd11an1n04x5 FILLER_26_881 ();
 b15zdnd00an1n02x5 FILLER_26_885 ();
 b15zdnd00an1n01x5 FILLER_26_887 ();
 b15zdnd11an1n64x5 FILLER_26_892 ();
 b15zdnd11an1n64x5 FILLER_26_956 ();
 b15zdnd11an1n64x5 FILLER_26_1020 ();
 b15zdnd11an1n64x5 FILLER_26_1084 ();
 b15zdnd11an1n32x5 FILLER_26_1148 ();
 b15zdnd11an1n08x5 FILLER_26_1180 ();
 b15zdnd11an1n04x5 FILLER_26_1188 ();
 b15zdnd00an1n02x5 FILLER_26_1192 ();
 b15zdnd11an1n64x5 FILLER_26_1203 ();
 b15zdnd11an1n16x5 FILLER_26_1267 ();
 b15zdnd11an1n04x5 FILLER_26_1283 ();
 b15zdnd00an1n02x5 FILLER_26_1287 ();
 b15zdnd00an1n01x5 FILLER_26_1289 ();
 b15zdnd11an1n16x5 FILLER_26_1302 ();
 b15zdnd11an1n32x5 FILLER_26_1336 ();
 b15zdnd11an1n08x5 FILLER_26_1368 ();
 b15zdnd11an1n04x5 FILLER_26_1376 ();
 b15zdnd00an1n02x5 FILLER_26_1380 ();
 b15zdnd00an1n01x5 FILLER_26_1382 ();
 b15zdnd11an1n04x5 FILLER_26_1387 ();
 b15zdnd11an1n64x5 FILLER_26_1396 ();
 b15zdnd11an1n64x5 FILLER_26_1460 ();
 b15zdnd11an1n32x5 FILLER_26_1524 ();
 b15zdnd11an1n04x5 FILLER_26_1574 ();
 b15zdnd00an1n01x5 FILLER_26_1578 ();
 b15zdnd11an1n32x5 FILLER_26_1583 ();
 b15zdnd11an1n04x5 FILLER_26_1615 ();
 b15zdnd00an1n02x5 FILLER_26_1619 ();
 b15zdnd11an1n04x5 FILLER_26_1627 ();
 b15zdnd11an1n04x5 FILLER_26_1636 ();
 b15zdnd11an1n08x5 FILLER_26_1647 ();
 b15zdnd00an1n02x5 FILLER_26_1655 ();
 b15zdnd11an1n64x5 FILLER_26_1662 ();
 b15zdnd11an1n64x5 FILLER_26_1726 ();
 b15zdnd00an1n02x5 FILLER_26_1790 ();
 b15zdnd11an1n64x5 FILLER_26_1813 ();
 b15zdnd11an1n04x5 FILLER_26_1877 ();
 b15zdnd00an1n02x5 FILLER_26_1881 ();
 b15zdnd00an1n01x5 FILLER_26_1883 ();
 b15zdnd11an1n04x5 FILLER_26_1893 ();
 b15zdnd11an1n16x5 FILLER_26_1903 ();
 b15zdnd11an1n04x5 FILLER_26_1919 ();
 b15zdnd00an1n02x5 FILLER_26_1923 ();
 b15zdnd11an1n32x5 FILLER_26_1930 ();
 b15zdnd11an1n08x5 FILLER_26_1962 ();
 b15zdnd11an1n04x5 FILLER_26_1970 ();
 b15zdnd00an1n02x5 FILLER_26_1974 ();
 b15zdnd11an1n16x5 FILLER_26_1982 ();
 b15zdnd00an1n02x5 FILLER_26_1998 ();
 b15zdnd00an1n01x5 FILLER_26_2000 ();
 b15zdnd11an1n08x5 FILLER_26_2007 ();
 b15zdnd11an1n04x5 FILLER_26_2015 ();
 b15zdnd00an1n02x5 FILLER_26_2019 ();
 b15zdnd00an1n01x5 FILLER_26_2021 ();
 b15zdnd11an1n08x5 FILLER_26_2050 ();
 b15zdnd00an1n01x5 FILLER_26_2058 ();
 b15zdnd11an1n64x5 FILLER_26_2069 ();
 b15zdnd00an1n02x5 FILLER_26_2133 ();
 b15zdnd00an1n01x5 FILLER_26_2135 ();
 b15zdnd00an1n02x5 FILLER_26_2152 ();
 b15zdnd11an1n16x5 FILLER_26_2162 ();
 b15zdnd11an1n04x5 FILLER_26_2178 ();
 b15zdnd00an1n02x5 FILLER_26_2182 ();
 b15zdnd00an1n01x5 FILLER_26_2184 ();
 b15zdnd11an1n04x5 FILLER_26_2192 ();
 b15zdnd11an1n64x5 FILLER_26_2208 ();
 b15zdnd11an1n04x5 FILLER_26_2272 ();
 b15zdnd11an1n32x5 FILLER_27_0 ();
 b15zdnd11an1n08x5 FILLER_27_32 ();
 b15zdnd00an1n02x5 FILLER_27_40 ();
 b15zdnd11an1n08x5 FILLER_27_52 ();
 b15zdnd00an1n02x5 FILLER_27_60 ();
 b15zdnd00an1n01x5 FILLER_27_62 ();
 b15zdnd11an1n04x5 FILLER_27_81 ();
 b15zdnd00an1n02x5 FILLER_27_85 ();
 b15zdnd00an1n01x5 FILLER_27_87 ();
 b15zdnd11an1n04x5 FILLER_27_110 ();
 b15zdnd11an1n32x5 FILLER_27_120 ();
 b15zdnd11an1n08x5 FILLER_27_152 ();
 b15zdnd11an1n04x5 FILLER_27_160 ();
 b15zdnd00an1n02x5 FILLER_27_164 ();
 b15zdnd11an1n16x5 FILLER_27_170 ();
 b15zdnd11an1n04x5 FILLER_27_186 ();
 b15zdnd00an1n02x5 FILLER_27_190 ();
 b15zdnd11an1n16x5 FILLER_27_199 ();
 b15zdnd11an1n08x5 FILLER_27_215 ();
 b15zdnd00an1n02x5 FILLER_27_223 ();
 b15zdnd00an1n01x5 FILLER_27_225 ();
 b15zdnd11an1n32x5 FILLER_27_238 ();
 b15zdnd11an1n08x5 FILLER_27_270 ();
 b15zdnd00an1n02x5 FILLER_27_278 ();
 b15zdnd11an1n16x5 FILLER_27_285 ();
 b15zdnd11an1n08x5 FILLER_27_301 ();
 b15zdnd11an1n08x5 FILLER_27_319 ();
 b15zdnd11an1n04x5 FILLER_27_327 ();
 b15zdnd11an1n64x5 FILLER_27_338 ();
 b15zdnd11an1n64x5 FILLER_27_402 ();
 b15zdnd11an1n16x5 FILLER_27_466 ();
 b15zdnd11an1n08x5 FILLER_27_482 ();
 b15zdnd00an1n01x5 FILLER_27_490 ();
 b15zdnd11an1n04x5 FILLER_27_497 ();
 b15zdnd00an1n01x5 FILLER_27_501 ();
 b15zdnd11an1n64x5 FILLER_27_510 ();
 b15zdnd11an1n04x5 FILLER_27_574 ();
 b15zdnd00an1n02x5 FILLER_27_578 ();
 b15zdnd00an1n01x5 FILLER_27_580 ();
 b15zdnd11an1n04x5 FILLER_27_597 ();
 b15zdnd11an1n16x5 FILLER_27_607 ();
 b15zdnd11an1n04x5 FILLER_27_623 ();
 b15zdnd11an1n04x5 FILLER_27_633 ();
 b15zdnd00an1n02x5 FILLER_27_637 ();
 b15zdnd00an1n01x5 FILLER_27_639 ();
 b15zdnd11an1n16x5 FILLER_27_646 ();
 b15zdnd11an1n08x5 FILLER_27_662 ();
 b15zdnd11an1n04x5 FILLER_27_670 ();
 b15zdnd11an1n08x5 FILLER_27_686 ();
 b15zdnd11an1n04x5 FILLER_27_694 ();
 b15zdnd00an1n02x5 FILLER_27_698 ();
 b15zdnd00an1n01x5 FILLER_27_700 ();
 b15zdnd11an1n32x5 FILLER_27_707 ();
 b15zdnd11an1n04x5 FILLER_27_739 ();
 b15zdnd00an1n01x5 FILLER_27_743 ();
 b15zdnd11an1n32x5 FILLER_27_750 ();
 b15zdnd11an1n08x5 FILLER_27_782 ();
 b15zdnd11an1n04x5 FILLER_27_790 ();
 b15zdnd00an1n02x5 FILLER_27_794 ();
 b15zdnd11an1n16x5 FILLER_27_810 ();
 b15zdnd11an1n08x5 FILLER_27_826 ();
 b15zdnd00an1n01x5 FILLER_27_834 ();
 b15zdnd11an1n04x5 FILLER_27_853 ();
 b15zdnd11an1n64x5 FILLER_27_862 ();
 b15zdnd11an1n32x5 FILLER_27_926 ();
 b15zdnd11an1n16x5 FILLER_27_958 ();
 b15zdnd11an1n08x5 FILLER_27_974 ();
 b15zdnd11an1n64x5 FILLER_27_991 ();
 b15zdnd11an1n16x5 FILLER_27_1055 ();
 b15zdnd11an1n04x5 FILLER_27_1071 ();
 b15zdnd00an1n02x5 FILLER_27_1075 ();
 b15zdnd11an1n64x5 FILLER_27_1087 ();
 b15zdnd11an1n64x5 FILLER_27_1151 ();
 b15zdnd11an1n08x5 FILLER_27_1215 ();
 b15zdnd11an1n04x5 FILLER_27_1223 ();
 b15zdnd11an1n04x5 FILLER_27_1239 ();
 b15zdnd11an1n16x5 FILLER_27_1268 ();
 b15zdnd00an1n01x5 FILLER_27_1284 ();
 b15zdnd11an1n16x5 FILLER_27_1303 ();
 b15zdnd11an1n08x5 FILLER_27_1319 ();
 b15zdnd00an1n02x5 FILLER_27_1327 ();
 b15zdnd11an1n04x5 FILLER_27_1353 ();
 b15zdnd11an1n08x5 FILLER_27_1369 ();
 b15zdnd11an1n04x5 FILLER_27_1377 ();
 b15zdnd11an1n04x5 FILLER_27_1391 ();
 b15zdnd11an1n04x5 FILLER_27_1400 ();
 b15zdnd11an1n04x5 FILLER_27_1411 ();
 b15zdnd11an1n04x5 FILLER_27_1420 ();
 b15zdnd11an1n16x5 FILLER_27_1429 ();
 b15zdnd11an1n04x5 FILLER_27_1445 ();
 b15zdnd11an1n32x5 FILLER_27_1455 ();
 b15zdnd11an1n04x5 FILLER_27_1487 ();
 b15zdnd00an1n02x5 FILLER_27_1491 ();
 b15zdnd00an1n01x5 FILLER_27_1493 ();
 b15zdnd11an1n08x5 FILLER_27_1506 ();
 b15zdnd11an1n04x5 FILLER_27_1514 ();
 b15zdnd00an1n01x5 FILLER_27_1518 ();
 b15zdnd11an1n32x5 FILLER_27_1528 ();
 b15zdnd11an1n16x5 FILLER_27_1560 ();
 b15zdnd11an1n04x5 FILLER_27_1576 ();
 b15zdnd11an1n04x5 FILLER_27_1586 ();
 b15zdnd11an1n16x5 FILLER_27_1600 ();
 b15zdnd11an1n08x5 FILLER_27_1616 ();
 b15zdnd11an1n04x5 FILLER_27_1624 ();
 b15zdnd11an1n04x5 FILLER_27_1642 ();
 b15zdnd11an1n64x5 FILLER_27_1666 ();
 b15zdnd11an1n32x5 FILLER_27_1730 ();
 b15zdnd11an1n16x5 FILLER_27_1762 ();
 b15zdnd00an1n02x5 FILLER_27_1778 ();
 b15zdnd11an1n32x5 FILLER_27_1785 ();
 b15zdnd11an1n16x5 FILLER_27_1817 ();
 b15zdnd11an1n08x5 FILLER_27_1833 ();
 b15zdnd00an1n02x5 FILLER_27_1841 ();
 b15zdnd11an1n32x5 FILLER_27_1851 ();
 b15zdnd11an1n08x5 FILLER_27_1883 ();
 b15zdnd00an1n02x5 FILLER_27_1891 ();
 b15zdnd00an1n01x5 FILLER_27_1893 ();
 b15zdnd11an1n32x5 FILLER_27_1899 ();
 b15zdnd11an1n16x5 FILLER_27_1931 ();
 b15zdnd11an1n08x5 FILLER_27_1947 ();
 b15zdnd11an1n32x5 FILLER_27_1960 ();
 b15zdnd11an1n16x5 FILLER_27_1992 ();
 b15zdnd11an1n04x5 FILLER_27_2008 ();
 b15zdnd00an1n02x5 FILLER_27_2012 ();
 b15zdnd00an1n01x5 FILLER_27_2014 ();
 b15zdnd11an1n32x5 FILLER_27_2035 ();
 b15zdnd11an1n04x5 FILLER_27_2067 ();
 b15zdnd00an1n01x5 FILLER_27_2071 ();
 b15zdnd11an1n04x5 FILLER_27_2077 ();
 b15zdnd11an1n32x5 FILLER_27_2090 ();
 b15zdnd11an1n16x5 FILLER_27_2122 ();
 b15zdnd11an1n04x5 FILLER_27_2138 ();
 b15zdnd00an1n01x5 FILLER_27_2142 ();
 b15zdnd11an1n04x5 FILLER_27_2149 ();
 b15zdnd11an1n16x5 FILLER_27_2168 ();
 b15zdnd00an1n01x5 FILLER_27_2184 ();
 b15zdnd11an1n08x5 FILLER_27_2195 ();
 b15zdnd00an1n01x5 FILLER_27_2203 ();
 b15zdnd11an1n64x5 FILLER_27_2212 ();
 b15zdnd11an1n08x5 FILLER_27_2276 ();
 b15zdnd11an1n16x5 FILLER_28_8 ();
 b15zdnd11an1n08x5 FILLER_28_24 ();
 b15zdnd11an1n04x5 FILLER_28_32 ();
 b15zdnd00an1n01x5 FILLER_28_36 ();
 b15zdnd11an1n16x5 FILLER_28_45 ();
 b15zdnd11an1n04x5 FILLER_28_61 ();
 b15zdnd11an1n16x5 FILLER_28_72 ();
 b15zdnd11an1n08x5 FILLER_28_88 ();
 b15zdnd00an1n02x5 FILLER_28_96 ();
 b15zdnd11an1n04x5 FILLER_28_104 ();
 b15zdnd11an1n08x5 FILLER_28_114 ();
 b15zdnd11an1n04x5 FILLER_28_122 ();
 b15zdnd00an1n02x5 FILLER_28_126 ();
 b15zdnd00an1n01x5 FILLER_28_128 ();
 b15zdnd11an1n16x5 FILLER_28_135 ();
 b15zdnd11an1n08x5 FILLER_28_151 ();
 b15zdnd11an1n04x5 FILLER_28_159 ();
 b15zdnd00an1n02x5 FILLER_28_163 ();
 b15zdnd00an1n01x5 FILLER_28_165 ();
 b15zdnd11an1n16x5 FILLER_28_171 ();
 b15zdnd11an1n04x5 FILLER_28_187 ();
 b15zdnd00an1n02x5 FILLER_28_191 ();
 b15zdnd00an1n01x5 FILLER_28_193 ();
 b15zdnd11an1n16x5 FILLER_28_199 ();
 b15zdnd11an1n08x5 FILLER_28_215 ();
 b15zdnd11an1n04x5 FILLER_28_223 ();
 b15zdnd00an1n01x5 FILLER_28_227 ();
 b15zdnd11an1n16x5 FILLER_28_237 ();
 b15zdnd11an1n08x5 FILLER_28_253 ();
 b15zdnd11an1n04x5 FILLER_28_261 ();
 b15zdnd00an1n02x5 FILLER_28_265 ();
 b15zdnd00an1n01x5 FILLER_28_267 ();
 b15zdnd11an1n64x5 FILLER_28_274 ();
 b15zdnd11an1n64x5 FILLER_28_338 ();
 b15zdnd11an1n64x5 FILLER_28_402 ();
 b15zdnd11an1n16x5 FILLER_28_466 ();
 b15zdnd11an1n04x5 FILLER_28_491 ();
 b15zdnd11an1n08x5 FILLER_28_502 ();
 b15zdnd11an1n04x5 FILLER_28_510 ();
 b15zdnd00an1n01x5 FILLER_28_514 ();
 b15zdnd11an1n16x5 FILLER_28_527 ();
 b15zdnd11an1n04x5 FILLER_28_543 ();
 b15zdnd11an1n32x5 FILLER_28_553 ();
 b15zdnd11an1n08x5 FILLER_28_585 ();
 b15zdnd11an1n04x5 FILLER_28_593 ();
 b15zdnd00an1n01x5 FILLER_28_597 ();
 b15zdnd11an1n32x5 FILLER_28_610 ();
 b15zdnd11an1n08x5 FILLER_28_642 ();
 b15zdnd11an1n04x5 FILLER_28_650 ();
 b15zdnd00an1n02x5 FILLER_28_654 ();
 b15zdnd00an1n01x5 FILLER_28_656 ();
 b15zdnd11an1n04x5 FILLER_28_665 ();
 b15zdnd00an1n02x5 FILLER_28_669 ();
 b15zdnd11an1n32x5 FILLER_28_686 ();
 b15zdnd11an1n32x5 FILLER_28_726 ();
 b15zdnd00an1n02x5 FILLER_28_758 ();
 b15zdnd00an1n01x5 FILLER_28_760 ();
 b15zdnd11an1n16x5 FILLER_28_773 ();
 b15zdnd00an1n02x5 FILLER_28_789 ();
 b15zdnd11an1n64x5 FILLER_28_797 ();
 b15zdnd11an1n08x5 FILLER_28_861 ();
 b15zdnd11an1n04x5 FILLER_28_878 ();
 b15zdnd11an1n64x5 FILLER_28_900 ();
 b15zdnd11an1n16x5 FILLER_28_964 ();
 b15zdnd11an1n04x5 FILLER_28_980 ();
 b15zdnd00an1n01x5 FILLER_28_984 ();
 b15zdnd11an1n32x5 FILLER_28_996 ();
 b15zdnd00an1n01x5 FILLER_28_1028 ();
 b15zdnd11an1n32x5 FILLER_28_1040 ();
 b15zdnd11an1n32x5 FILLER_28_1089 ();
 b15zdnd00an1n02x5 FILLER_28_1121 ();
 b15zdnd00an1n01x5 FILLER_28_1123 ();
 b15zdnd11an1n32x5 FILLER_28_1137 ();
 b15zdnd11an1n04x5 FILLER_28_1169 ();
 b15zdnd00an1n02x5 FILLER_28_1173 ();
 b15zdnd11an1n16x5 FILLER_28_1185 ();
 b15zdnd00an1n02x5 FILLER_28_1201 ();
 b15zdnd00an1n01x5 FILLER_28_1203 ();
 b15zdnd11an1n64x5 FILLER_28_1208 ();
 b15zdnd11an1n32x5 FILLER_28_1272 ();
 b15zdnd11an1n16x5 FILLER_28_1304 ();
 b15zdnd11an1n08x5 FILLER_28_1320 ();
 b15zdnd11an1n32x5 FILLER_28_1338 ();
 b15zdnd11an1n16x5 FILLER_28_1370 ();
 b15zdnd11an1n04x5 FILLER_28_1386 ();
 b15zdnd00an1n02x5 FILLER_28_1390 ();
 b15zdnd11an1n04x5 FILLER_28_1397 ();
 b15zdnd11an1n08x5 FILLER_28_1411 ();
 b15zdnd00an1n02x5 FILLER_28_1419 ();
 b15zdnd00an1n01x5 FILLER_28_1421 ();
 b15zdnd11an1n08x5 FILLER_28_1438 ();
 b15zdnd11an1n04x5 FILLER_28_1446 ();
 b15zdnd00an1n02x5 FILLER_28_1450 ();
 b15zdnd00an1n01x5 FILLER_28_1452 ();
 b15zdnd11an1n04x5 FILLER_28_1460 ();
 b15zdnd11an1n32x5 FILLER_28_1473 ();
 b15zdnd11an1n16x5 FILLER_28_1505 ();
 b15zdnd11an1n04x5 FILLER_28_1521 ();
 b15zdnd11an1n64x5 FILLER_28_1531 ();
 b15zdnd11an1n64x5 FILLER_28_1595 ();
 b15zdnd11an1n16x5 FILLER_28_1659 ();
 b15zdnd11an1n08x5 FILLER_28_1675 ();
 b15zdnd11an1n32x5 FILLER_28_1703 ();
 b15zdnd11an1n16x5 FILLER_28_1735 ();
 b15zdnd11an1n08x5 FILLER_28_1751 ();
 b15zdnd11an1n04x5 FILLER_28_1759 ();
 b15zdnd00an1n01x5 FILLER_28_1763 ();
 b15zdnd11an1n08x5 FILLER_28_1769 ();
 b15zdnd00an1n02x5 FILLER_28_1777 ();
 b15zdnd00an1n01x5 FILLER_28_1779 ();
 b15zdnd11an1n04x5 FILLER_28_1787 ();
 b15zdnd11an1n16x5 FILLER_28_1795 ();
 b15zdnd11an1n08x5 FILLER_28_1823 ();
 b15zdnd11an1n04x5 FILLER_28_1831 ();
 b15zdnd00an1n01x5 FILLER_28_1835 ();
 b15zdnd11an1n04x5 FILLER_28_1852 ();
 b15zdnd11an1n32x5 FILLER_28_1865 ();
 b15zdnd11an1n04x5 FILLER_28_1897 ();
 b15zdnd00an1n01x5 FILLER_28_1901 ();
 b15zdnd11an1n16x5 FILLER_28_1909 ();
 b15zdnd11an1n04x5 FILLER_28_1925 ();
 b15zdnd00an1n01x5 FILLER_28_1929 ();
 b15zdnd11an1n08x5 FILLER_28_1943 ();
 b15zdnd00an1n02x5 FILLER_28_1951 ();
 b15zdnd00an1n01x5 FILLER_28_1953 ();
 b15zdnd11an1n32x5 FILLER_28_1966 ();
 b15zdnd11an1n16x5 FILLER_28_1998 ();
 b15zdnd11an1n08x5 FILLER_28_2014 ();
 b15zdnd11an1n04x5 FILLER_28_2022 ();
 b15zdnd00an1n02x5 FILLER_28_2026 ();
 b15zdnd11an1n32x5 FILLER_28_2042 ();
 b15zdnd00an1n02x5 FILLER_28_2074 ();
 b15zdnd11an1n04x5 FILLER_28_2096 ();
 b15zdnd11an1n04x5 FILLER_28_2120 ();
 b15zdnd11an1n16x5 FILLER_28_2131 ();
 b15zdnd11an1n04x5 FILLER_28_2147 ();
 b15zdnd00an1n02x5 FILLER_28_2151 ();
 b15zdnd00an1n01x5 FILLER_28_2153 ();
 b15zdnd11an1n16x5 FILLER_28_2162 ();
 b15zdnd11an1n08x5 FILLER_28_2178 ();
 b15zdnd00an1n01x5 FILLER_28_2186 ();
 b15zdnd11an1n64x5 FILLER_28_2192 ();
 b15zdnd11an1n16x5 FILLER_28_2256 ();
 b15zdnd11an1n04x5 FILLER_28_2272 ();
 b15zdnd11an1n64x5 FILLER_29_0 ();
 b15zdnd11an1n04x5 FILLER_29_64 ();
 b15zdnd00an1n02x5 FILLER_29_68 ();
 b15zdnd00an1n01x5 FILLER_29_70 ();
 b15zdnd11an1n16x5 FILLER_29_78 ();
 b15zdnd11an1n04x5 FILLER_29_94 ();
 b15zdnd00an1n01x5 FILLER_29_98 ();
 b15zdnd11an1n32x5 FILLER_29_113 ();
 b15zdnd11an1n08x5 FILLER_29_145 ();
 b15zdnd11an1n04x5 FILLER_29_153 ();
 b15zdnd00an1n02x5 FILLER_29_157 ();
 b15zdnd00an1n01x5 FILLER_29_159 ();
 b15zdnd11an1n64x5 FILLER_29_168 ();
 b15zdnd11an1n08x5 FILLER_29_232 ();
 b15zdnd11an1n16x5 FILLER_29_245 ();
 b15zdnd11an1n64x5 FILLER_29_270 ();
 b15zdnd11an1n64x5 FILLER_29_339 ();
 b15zdnd11an1n32x5 FILLER_29_403 ();
 b15zdnd11an1n16x5 FILLER_29_435 ();
 b15zdnd00an1n02x5 FILLER_29_451 ();
 b15zdnd11an1n32x5 FILLER_29_462 ();
 b15zdnd11an1n04x5 FILLER_29_494 ();
 b15zdnd00an1n02x5 FILLER_29_498 ();
 b15zdnd11an1n04x5 FILLER_29_512 ();
 b15zdnd11an1n32x5 FILLER_29_523 ();
 b15zdnd11an1n16x5 FILLER_29_555 ();
 b15zdnd11an1n04x5 FILLER_29_571 ();
 b15zdnd00an1n01x5 FILLER_29_575 ();
 b15zdnd11an1n04x5 FILLER_29_594 ();
 b15zdnd11an1n32x5 FILLER_29_603 ();
 b15zdnd11an1n08x5 FILLER_29_635 ();
 b15zdnd11an1n04x5 FILLER_29_643 ();
 b15zdnd00an1n02x5 FILLER_29_647 ();
 b15zdnd00an1n01x5 FILLER_29_649 ();
 b15zdnd11an1n08x5 FILLER_29_658 ();
 b15zdnd11an1n04x5 FILLER_29_666 ();
 b15zdnd00an1n02x5 FILLER_29_670 ();
 b15zdnd11an1n16x5 FILLER_29_677 ();
 b15zdnd11an1n04x5 FILLER_29_693 ();
 b15zdnd11an1n32x5 FILLER_29_706 ();
 b15zdnd00an1n01x5 FILLER_29_738 ();
 b15zdnd11an1n08x5 FILLER_29_755 ();
 b15zdnd00an1n01x5 FILLER_29_763 ();
 b15zdnd11an1n08x5 FILLER_29_769 ();
 b15zdnd11an1n04x5 FILLER_29_777 ();
 b15zdnd00an1n01x5 FILLER_29_781 ();
 b15zdnd11an1n64x5 FILLER_29_796 ();
 b15zdnd11an1n08x5 FILLER_29_860 ();
 b15zdnd11an1n04x5 FILLER_29_868 ();
 b15zdnd00an1n02x5 FILLER_29_872 ();
 b15zdnd00an1n01x5 FILLER_29_874 ();
 b15zdnd11an1n32x5 FILLER_29_882 ();
 b15zdnd11an1n08x5 FILLER_29_914 ();
 b15zdnd00an1n02x5 FILLER_29_922 ();
 b15zdnd11an1n16x5 FILLER_29_944 ();
 b15zdnd11an1n08x5 FILLER_29_960 ();
 b15zdnd11an1n04x5 FILLER_29_968 ();
 b15zdnd00an1n01x5 FILLER_29_972 ();
 b15zdnd11an1n16x5 FILLER_29_1004 ();
 b15zdnd11an1n08x5 FILLER_29_1020 ();
 b15zdnd00an1n01x5 FILLER_29_1028 ();
 b15zdnd11an1n64x5 FILLER_29_1044 ();
 b15zdnd11an1n16x5 FILLER_29_1108 ();
 b15zdnd11an1n04x5 FILLER_29_1124 ();
 b15zdnd11an1n16x5 FILLER_29_1153 ();
 b15zdnd11an1n08x5 FILLER_29_1169 ();
 b15zdnd00an1n02x5 FILLER_29_1177 ();
 b15zdnd11an1n64x5 FILLER_29_1204 ();
 b15zdnd11an1n08x5 FILLER_29_1268 ();
 b15zdnd11an1n04x5 FILLER_29_1276 ();
 b15zdnd00an1n02x5 FILLER_29_1280 ();
 b15zdnd00an1n01x5 FILLER_29_1282 ();
 b15zdnd11an1n04x5 FILLER_29_1288 ();
 b15zdnd11an1n16x5 FILLER_29_1310 ();
 b15zdnd11an1n04x5 FILLER_29_1326 ();
 b15zdnd00an1n02x5 FILLER_29_1330 ();
 b15zdnd00an1n01x5 FILLER_29_1332 ();
 b15zdnd11an1n64x5 FILLER_29_1351 ();
 b15zdnd11an1n32x5 FILLER_29_1415 ();
 b15zdnd11an1n04x5 FILLER_29_1447 ();
 b15zdnd00an1n02x5 FILLER_29_1451 ();
 b15zdnd00an1n01x5 FILLER_29_1453 ();
 b15zdnd11an1n32x5 FILLER_29_1460 ();
 b15zdnd11an1n08x5 FILLER_29_1492 ();
 b15zdnd00an1n02x5 FILLER_29_1500 ();
 b15zdnd00an1n01x5 FILLER_29_1502 ();
 b15zdnd11an1n08x5 FILLER_29_1513 ();
 b15zdnd00an1n02x5 FILLER_29_1521 ();
 b15zdnd11an1n16x5 FILLER_29_1529 ();
 b15zdnd11an1n08x5 FILLER_29_1545 ();
 b15zdnd11an1n04x5 FILLER_29_1553 ();
 b15zdnd00an1n01x5 FILLER_29_1557 ();
 b15zdnd11an1n04x5 FILLER_29_1566 ();
 b15zdnd11an1n04x5 FILLER_29_1575 ();
 b15zdnd00an1n01x5 FILLER_29_1579 ();
 b15zdnd11an1n16x5 FILLER_29_1596 ();
 b15zdnd00an1n01x5 FILLER_29_1612 ();
 b15zdnd11an1n16x5 FILLER_29_1622 ();
 b15zdnd11an1n08x5 FILLER_29_1638 ();
 b15zdnd11an1n04x5 FILLER_29_1646 ();
 b15zdnd00an1n01x5 FILLER_29_1650 ();
 b15zdnd11an1n64x5 FILLER_29_1669 ();
 b15zdnd11an1n32x5 FILLER_29_1733 ();
 b15zdnd11an1n16x5 FILLER_29_1765 ();
 b15zdnd00an1n02x5 FILLER_29_1781 ();
 b15zdnd11an1n16x5 FILLER_29_1795 ();
 b15zdnd11an1n04x5 FILLER_29_1811 ();
 b15zdnd00an1n01x5 FILLER_29_1815 ();
 b15zdnd11an1n16x5 FILLER_29_1824 ();
 b15zdnd11an1n08x5 FILLER_29_1840 ();
 b15zdnd00an1n02x5 FILLER_29_1848 ();
 b15zdnd11an1n32x5 FILLER_29_1862 ();
 b15zdnd11an1n08x5 FILLER_29_1894 ();
 b15zdnd00an1n02x5 FILLER_29_1902 ();
 b15zdnd11an1n16x5 FILLER_29_1915 ();
 b15zdnd11an1n08x5 FILLER_29_1931 ();
 b15zdnd00an1n02x5 FILLER_29_1939 ();
 b15zdnd11an1n64x5 FILLER_29_1947 ();
 b15zdnd11an1n16x5 FILLER_29_2011 ();
 b15zdnd00an1n01x5 FILLER_29_2027 ();
 b15zdnd11an1n64x5 FILLER_29_2033 ();
 b15zdnd11an1n32x5 FILLER_29_2097 ();
 b15zdnd00an1n02x5 FILLER_29_2129 ();
 b15zdnd00an1n01x5 FILLER_29_2131 ();
 b15zdnd11an1n32x5 FILLER_29_2143 ();
 b15zdnd11an1n08x5 FILLER_29_2175 ();
 b15zdnd00an1n01x5 FILLER_29_2183 ();
 b15zdnd11an1n64x5 FILLER_29_2198 ();
 b15zdnd11an1n16x5 FILLER_29_2262 ();
 b15zdnd11an1n04x5 FILLER_29_2278 ();
 b15zdnd00an1n02x5 FILLER_29_2282 ();
 b15zdnd11an1n16x5 FILLER_30_8 ();
 b15zdnd11an1n08x5 FILLER_30_24 ();
 b15zdnd00an1n01x5 FILLER_30_32 ();
 b15zdnd11an1n04x5 FILLER_30_64 ();
 b15zdnd11an1n64x5 FILLER_30_86 ();
 b15zdnd11an1n32x5 FILLER_30_150 ();
 b15zdnd11an1n04x5 FILLER_30_182 ();
 b15zdnd00an1n02x5 FILLER_30_186 ();
 b15zdnd00an1n01x5 FILLER_30_188 ();
 b15zdnd11an1n32x5 FILLER_30_194 ();
 b15zdnd11an1n08x5 FILLER_30_226 ();
 b15zdnd00an1n02x5 FILLER_30_234 ();
 b15zdnd00an1n01x5 FILLER_30_236 ();
 b15zdnd11an1n08x5 FILLER_30_244 ();
 b15zdnd11an1n04x5 FILLER_30_252 ();
 b15zdnd00an1n02x5 FILLER_30_256 ();
 b15zdnd11an1n32x5 FILLER_30_264 ();
 b15zdnd00an1n01x5 FILLER_30_296 ();
 b15zdnd11an1n16x5 FILLER_30_309 ();
 b15zdnd11an1n08x5 FILLER_30_325 ();
 b15zdnd11an1n64x5 FILLER_30_337 ();
 b15zdnd00an1n01x5 FILLER_30_401 ();
 b15zdnd11an1n04x5 FILLER_30_421 ();
 b15zdnd11an1n32x5 FILLER_30_440 ();
 b15zdnd00an1n01x5 FILLER_30_472 ();
 b15zdnd11an1n16x5 FILLER_30_498 ();
 b15zdnd00an1n01x5 FILLER_30_514 ();
 b15zdnd11an1n64x5 FILLER_30_526 ();
 b15zdnd11an1n32x5 FILLER_30_590 ();
 b15zdnd11an1n16x5 FILLER_30_622 ();
 b15zdnd11an1n08x5 FILLER_30_638 ();
 b15zdnd11an1n04x5 FILLER_30_646 ();
 b15zdnd00an1n02x5 FILLER_30_650 ();
 b15zdnd11an1n32x5 FILLER_30_658 ();
 b15zdnd11an1n08x5 FILLER_30_690 ();
 b15zdnd00an1n02x5 FILLER_30_698 ();
 b15zdnd00an1n01x5 FILLER_30_700 ();
 b15zdnd11an1n04x5 FILLER_30_713 ();
 b15zdnd00an1n01x5 FILLER_30_717 ();
 b15zdnd11an1n04x5 FILLER_30_726 ();
 b15zdnd11an1n04x5 FILLER_30_739 ();
 b15zdnd11an1n64x5 FILLER_30_764 ();
 b15zdnd11an1n32x5 FILLER_30_828 ();
 b15zdnd11an1n08x5 FILLER_30_860 ();
 b15zdnd11an1n04x5 FILLER_30_868 ();
 b15zdnd00an1n02x5 FILLER_30_872 ();
 b15zdnd00an1n01x5 FILLER_30_874 ();
 b15zdnd11an1n04x5 FILLER_30_880 ();
 b15zdnd00an1n02x5 FILLER_30_884 ();
 b15zdnd11an1n64x5 FILLER_30_896 ();
 b15zdnd11an1n04x5 FILLER_30_960 ();
 b15zdnd00an1n02x5 FILLER_30_964 ();
 b15zdnd11an1n32x5 FILLER_30_983 ();
 b15zdnd11an1n16x5 FILLER_30_1015 ();
 b15zdnd00an1n02x5 FILLER_30_1031 ();
 b15zdnd11an1n32x5 FILLER_30_1043 ();
 b15zdnd11an1n16x5 FILLER_30_1075 ();
 b15zdnd11an1n08x5 FILLER_30_1091 ();
 b15zdnd00an1n02x5 FILLER_30_1099 ();
 b15zdnd00an1n01x5 FILLER_30_1101 ();
 b15zdnd11an1n32x5 FILLER_30_1112 ();
 b15zdnd11an1n16x5 FILLER_30_1144 ();
 b15zdnd00an1n02x5 FILLER_30_1160 ();
 b15zdnd11an1n04x5 FILLER_30_1171 ();
 b15zdnd11an1n64x5 FILLER_30_1179 ();
 b15zdnd11an1n64x5 FILLER_30_1243 ();
 b15zdnd11an1n16x5 FILLER_30_1307 ();
 b15zdnd00an1n02x5 FILLER_30_1323 ();
 b15zdnd11an1n16x5 FILLER_30_1330 ();
 b15zdnd11an1n08x5 FILLER_30_1346 ();
 b15zdnd00an1n02x5 FILLER_30_1354 ();
 b15zdnd11an1n04x5 FILLER_30_1364 ();
 b15zdnd11an1n64x5 FILLER_30_1380 ();
 b15zdnd11an1n64x5 FILLER_30_1444 ();
 b15zdnd11an1n32x5 FILLER_30_1508 ();
 b15zdnd00an1n01x5 FILLER_30_1540 ();
 b15zdnd11an1n08x5 FILLER_30_1556 ();
 b15zdnd11an1n04x5 FILLER_30_1564 ();
 b15zdnd00an1n02x5 FILLER_30_1568 ();
 b15zdnd11an1n16x5 FILLER_30_1582 ();
 b15zdnd11an1n08x5 FILLER_30_1598 ();
 b15zdnd00an1n02x5 FILLER_30_1606 ();
 b15zdnd00an1n01x5 FILLER_30_1608 ();
 b15zdnd11an1n32x5 FILLER_30_1619 ();
 b15zdnd11an1n04x5 FILLER_30_1651 ();
 b15zdnd00an1n02x5 FILLER_30_1655 ();
 b15zdnd11an1n64x5 FILLER_30_1662 ();
 b15zdnd11an1n08x5 FILLER_30_1726 ();
 b15zdnd11an1n04x5 FILLER_30_1734 ();
 b15zdnd00an1n01x5 FILLER_30_1738 ();
 b15zdnd11an1n32x5 FILLER_30_1755 ();
 b15zdnd11an1n16x5 FILLER_30_1787 ();
 b15zdnd11an1n08x5 FILLER_30_1803 ();
 b15zdnd11an1n04x5 FILLER_30_1811 ();
 b15zdnd00an1n01x5 FILLER_30_1815 ();
 b15zdnd11an1n04x5 FILLER_30_1825 ();
 b15zdnd00an1n01x5 FILLER_30_1829 ();
 b15zdnd11an1n32x5 FILLER_30_1836 ();
 b15zdnd11an1n16x5 FILLER_30_1868 ();
 b15zdnd11an1n08x5 FILLER_30_1884 ();
 b15zdnd00an1n01x5 FILLER_30_1892 ();
 b15zdnd11an1n32x5 FILLER_30_1898 ();
 b15zdnd11an1n08x5 FILLER_30_1930 ();
 b15zdnd00an1n02x5 FILLER_30_1938 ();
 b15zdnd00an1n01x5 FILLER_30_1940 ();
 b15zdnd11an1n16x5 FILLER_30_1950 ();
 b15zdnd11an1n04x5 FILLER_30_1966 ();
 b15zdnd00an1n02x5 FILLER_30_1970 ();
 b15zdnd11an1n04x5 FILLER_30_1984 ();
 b15zdnd11an1n08x5 FILLER_30_1994 ();
 b15zdnd00an1n02x5 FILLER_30_2002 ();
 b15zdnd00an1n01x5 FILLER_30_2004 ();
 b15zdnd11an1n64x5 FILLER_30_2013 ();
 b15zdnd11an1n04x5 FILLER_30_2077 ();
 b15zdnd11an1n64x5 FILLER_30_2087 ();
 b15zdnd00an1n02x5 FILLER_30_2151 ();
 b15zdnd00an1n01x5 FILLER_30_2153 ();
 b15zdnd11an1n64x5 FILLER_30_2162 ();
 b15zdnd11an1n32x5 FILLER_30_2226 ();
 b15zdnd11an1n16x5 FILLER_30_2258 ();
 b15zdnd00an1n02x5 FILLER_30_2274 ();
 b15zdnd11an1n32x5 FILLER_31_0 ();
 b15zdnd11an1n08x5 FILLER_31_32 ();
 b15zdnd00an1n01x5 FILLER_31_40 ();
 b15zdnd11an1n16x5 FILLER_31_54 ();
 b15zdnd11an1n04x5 FILLER_31_70 ();
 b15zdnd11an1n32x5 FILLER_31_81 ();
 b15zdnd00an1n02x5 FILLER_31_113 ();
 b15zdnd00an1n01x5 FILLER_31_115 ();
 b15zdnd11an1n64x5 FILLER_31_122 ();
 b15zdnd11an1n32x5 FILLER_31_186 ();
 b15zdnd11an1n16x5 FILLER_31_218 ();
 b15zdnd00an1n02x5 FILLER_31_234 ();
 b15zdnd11an1n32x5 FILLER_31_241 ();
 b15zdnd11an1n04x5 FILLER_31_282 ();
 b15zdnd00an1n02x5 FILLER_31_286 ();
 b15zdnd00an1n01x5 FILLER_31_288 ();
 b15zdnd11an1n04x5 FILLER_31_295 ();
 b15zdnd11an1n16x5 FILLER_31_311 ();
 b15zdnd11an1n04x5 FILLER_31_327 ();
 b15zdnd00an1n01x5 FILLER_31_331 ();
 b15zdnd11an1n04x5 FILLER_31_344 ();
 b15zdnd11an1n32x5 FILLER_31_360 ();
 b15zdnd11an1n16x5 FILLER_31_392 ();
 b15zdnd11an1n04x5 FILLER_31_408 ();
 b15zdnd11an1n04x5 FILLER_31_417 ();
 b15zdnd11an1n16x5 FILLER_31_432 ();
 b15zdnd11an1n08x5 FILLER_31_448 ();
 b15zdnd00an1n01x5 FILLER_31_456 ();
 b15zdnd11an1n64x5 FILLER_31_460 ();
 b15zdnd11an1n16x5 FILLER_31_524 ();
 b15zdnd11an1n08x5 FILLER_31_540 ();
 b15zdnd11an1n16x5 FILLER_31_552 ();
 b15zdnd11an1n08x5 FILLER_31_568 ();
 b15zdnd00an1n01x5 FILLER_31_576 ();
 b15zdnd11an1n16x5 FILLER_31_586 ();
 b15zdnd00an1n02x5 FILLER_31_602 ();
 b15zdnd00an1n01x5 FILLER_31_604 ();
 b15zdnd11an1n64x5 FILLER_31_622 ();
 b15zdnd11an1n64x5 FILLER_31_686 ();
 b15zdnd11an1n32x5 FILLER_31_750 ();
 b15zdnd11an1n08x5 FILLER_31_782 ();
 b15zdnd00an1n02x5 FILLER_31_790 ();
 b15zdnd11an1n04x5 FILLER_31_798 ();
 b15zdnd11an1n32x5 FILLER_31_809 ();
 b15zdnd11an1n08x5 FILLER_31_841 ();
 b15zdnd00an1n02x5 FILLER_31_849 ();
 b15zdnd00an1n01x5 FILLER_31_851 ();
 b15zdnd11an1n32x5 FILLER_31_857 ();
 b15zdnd00an1n01x5 FILLER_31_889 ();
 b15zdnd11an1n64x5 FILLER_31_895 ();
 b15zdnd11an1n64x5 FILLER_31_959 ();
 b15zdnd11an1n32x5 FILLER_31_1023 ();
 b15zdnd11an1n16x5 FILLER_31_1055 ();
 b15zdnd11an1n64x5 FILLER_31_1083 ();
 b15zdnd11an1n08x5 FILLER_31_1147 ();
 b15zdnd11an1n04x5 FILLER_31_1155 ();
 b15zdnd00an1n01x5 FILLER_31_1159 ();
 b15zdnd11an1n64x5 FILLER_31_1164 ();
 b15zdnd11an1n64x5 FILLER_31_1228 ();
 b15zdnd11an1n32x5 FILLER_31_1292 ();
 b15zdnd11an1n04x5 FILLER_31_1324 ();
 b15zdnd00an1n02x5 FILLER_31_1328 ();
 b15zdnd11an1n16x5 FILLER_31_1335 ();
 b15zdnd11an1n04x5 FILLER_31_1351 ();
 b15zdnd00an1n02x5 FILLER_31_1355 ();
 b15zdnd00an1n01x5 FILLER_31_1357 ();
 b15zdnd11an1n32x5 FILLER_31_1363 ();
 b15zdnd11an1n04x5 FILLER_31_1408 ();
 b15zdnd11an1n32x5 FILLER_31_1421 ();
 b15zdnd11an1n16x5 FILLER_31_1453 ();
 b15zdnd11an1n08x5 FILLER_31_1469 ();
 b15zdnd00an1n02x5 FILLER_31_1477 ();
 b15zdnd00an1n01x5 FILLER_31_1479 ();
 b15zdnd11an1n08x5 FILLER_31_1486 ();
 b15zdnd00an1n02x5 FILLER_31_1494 ();
 b15zdnd11an1n08x5 FILLER_31_1520 ();
 b15zdnd00an1n02x5 FILLER_31_1528 ();
 b15zdnd00an1n01x5 FILLER_31_1530 ();
 b15zdnd11an1n64x5 FILLER_31_1539 ();
 b15zdnd11an1n16x5 FILLER_31_1603 ();
 b15zdnd11an1n08x5 FILLER_31_1619 ();
 b15zdnd00an1n02x5 FILLER_31_1627 ();
 b15zdnd00an1n01x5 FILLER_31_1629 ();
 b15zdnd11an1n04x5 FILLER_31_1635 ();
 b15zdnd11an1n04x5 FILLER_31_1652 ();
 b15zdnd11an1n16x5 FILLER_31_1663 ();
 b15zdnd11an1n64x5 FILLER_31_1686 ();
 b15zdnd00an1n01x5 FILLER_31_1750 ();
 b15zdnd11an1n64x5 FILLER_31_1757 ();
 b15zdnd11an1n32x5 FILLER_31_1821 ();
 b15zdnd11an1n08x5 FILLER_31_1853 ();
 b15zdnd11an1n04x5 FILLER_31_1861 ();
 b15zdnd00an1n02x5 FILLER_31_1865 ();
 b15zdnd11an1n16x5 FILLER_31_1871 ();
 b15zdnd00an1n02x5 FILLER_31_1887 ();
 b15zdnd00an1n01x5 FILLER_31_1889 ();
 b15zdnd11an1n32x5 FILLER_31_1901 ();
 b15zdnd11an1n08x5 FILLER_31_1933 ();
 b15zdnd11an1n04x5 FILLER_31_1941 ();
 b15zdnd00an1n01x5 FILLER_31_1945 ();
 b15zdnd11an1n08x5 FILLER_31_1961 ();
 b15zdnd00an1n02x5 FILLER_31_1969 ();
 b15zdnd00an1n01x5 FILLER_31_1971 ();
 b15zdnd11an1n64x5 FILLER_31_1993 ();
 b15zdnd11an1n16x5 FILLER_31_2057 ();
 b15zdnd11an1n08x5 FILLER_31_2073 ();
 b15zdnd11an1n16x5 FILLER_31_2087 ();
 b15zdnd11an1n04x5 FILLER_31_2103 ();
 b15zdnd11an1n04x5 FILLER_31_2112 ();
 b15zdnd11an1n64x5 FILLER_31_2130 ();
 b15zdnd11an1n08x5 FILLER_31_2194 ();
 b15zdnd00an1n02x5 FILLER_31_2202 ();
 b15zdnd00an1n01x5 FILLER_31_2204 ();
 b15zdnd11an1n64x5 FILLER_31_2210 ();
 b15zdnd11an1n08x5 FILLER_31_2274 ();
 b15zdnd00an1n02x5 FILLER_31_2282 ();
 b15zdnd11an1n16x5 FILLER_32_8 ();
 b15zdnd00an1n01x5 FILLER_32_24 ();
 b15zdnd11an1n16x5 FILLER_32_45 ();
 b15zdnd11an1n08x5 FILLER_32_61 ();
 b15zdnd11an1n04x5 FILLER_32_69 ();
 b15zdnd11an1n32x5 FILLER_32_83 ();
 b15zdnd11an1n04x5 FILLER_32_115 ();
 b15zdnd00an1n01x5 FILLER_32_119 ();
 b15zdnd11an1n04x5 FILLER_32_125 ();
 b15zdnd11an1n08x5 FILLER_32_139 ();
 b15zdnd11an1n04x5 FILLER_32_147 ();
 b15zdnd00an1n02x5 FILLER_32_151 ();
 b15zdnd11an1n04x5 FILLER_32_160 ();
 b15zdnd11an1n08x5 FILLER_32_176 ();
 b15zdnd11an1n04x5 FILLER_32_184 ();
 b15zdnd00an1n02x5 FILLER_32_188 ();
 b15zdnd11an1n16x5 FILLER_32_194 ();
 b15zdnd11an1n08x5 FILLER_32_210 ();
 b15zdnd00an1n01x5 FILLER_32_218 ();
 b15zdnd11an1n16x5 FILLER_32_235 ();
 b15zdnd11an1n04x5 FILLER_32_251 ();
 b15zdnd00an1n02x5 FILLER_32_255 ();
 b15zdnd11an1n64x5 FILLER_32_262 ();
 b15zdnd11an1n16x5 FILLER_32_326 ();
 b15zdnd00an1n02x5 FILLER_32_342 ();
 b15zdnd00an1n01x5 FILLER_32_344 ();
 b15zdnd11an1n32x5 FILLER_32_361 ();
 b15zdnd11an1n16x5 FILLER_32_393 ();
 b15zdnd00an1n02x5 FILLER_32_409 ();
 b15zdnd11an1n32x5 FILLER_32_417 ();
 b15zdnd11an1n08x5 FILLER_32_449 ();
 b15zdnd00an1n02x5 FILLER_32_457 ();
 b15zdnd11an1n16x5 FILLER_32_471 ();
 b15zdnd11an1n04x5 FILLER_32_487 ();
 b15zdnd00an1n02x5 FILLER_32_491 ();
 b15zdnd00an1n01x5 FILLER_32_493 ();
 b15zdnd11an1n16x5 FILLER_32_500 ();
 b15zdnd11an1n04x5 FILLER_32_516 ();
 b15zdnd00an1n02x5 FILLER_32_520 ();
 b15zdnd00an1n01x5 FILLER_32_522 ();
 b15zdnd11an1n32x5 FILLER_32_535 ();
 b15zdnd00an1n02x5 FILLER_32_567 ();
 b15zdnd11an1n08x5 FILLER_32_574 ();
 b15zdnd11an1n04x5 FILLER_32_582 ();
 b15zdnd00an1n02x5 FILLER_32_586 ();
 b15zdnd11an1n04x5 FILLER_32_593 ();
 b15zdnd00an1n01x5 FILLER_32_597 ();
 b15zdnd11an1n64x5 FILLER_32_606 ();
 b15zdnd11an1n16x5 FILLER_32_670 ();
 b15zdnd11an1n08x5 FILLER_32_686 ();
 b15zdnd00an1n02x5 FILLER_32_694 ();
 b15zdnd00an1n01x5 FILLER_32_696 ();
 b15zdnd11an1n08x5 FILLER_32_710 ();
 b15zdnd11an1n64x5 FILLER_32_726 ();
 b15zdnd11an1n04x5 FILLER_32_805 ();
 b15zdnd11an1n16x5 FILLER_32_818 ();
 b15zdnd00an1n01x5 FILLER_32_834 ();
 b15zdnd11an1n04x5 FILLER_32_844 ();
 b15zdnd00an1n01x5 FILLER_32_848 ();
 b15zdnd11an1n64x5 FILLER_32_856 ();
 b15zdnd11an1n32x5 FILLER_32_920 ();
 b15zdnd11an1n16x5 FILLER_32_952 ();
 b15zdnd11an1n04x5 FILLER_32_968 ();
 b15zdnd00an1n01x5 FILLER_32_972 ();
 b15zdnd11an1n04x5 FILLER_32_997 ();
 b15zdnd11an1n16x5 FILLER_32_1013 ();
 b15zdnd00an1n02x5 FILLER_32_1029 ();
 b15zdnd00an1n01x5 FILLER_32_1031 ();
 b15zdnd11an1n16x5 FILLER_32_1041 ();
 b15zdnd00an1n02x5 FILLER_32_1057 ();
 b15zdnd11an1n64x5 FILLER_32_1080 ();
 b15zdnd11an1n32x5 FILLER_32_1144 ();
 b15zdnd11an1n16x5 FILLER_32_1176 ();
 b15zdnd00an1n02x5 FILLER_32_1192 ();
 b15zdnd00an1n01x5 FILLER_32_1194 ();
 b15zdnd11an1n16x5 FILLER_32_1200 ();
 b15zdnd11an1n08x5 FILLER_32_1216 ();
 b15zdnd00an1n02x5 FILLER_32_1224 ();
 b15zdnd00an1n01x5 FILLER_32_1226 ();
 b15zdnd11an1n64x5 FILLER_32_1231 ();
 b15zdnd11an1n16x5 FILLER_32_1295 ();
 b15zdnd00an1n02x5 FILLER_32_1311 ();
 b15zdnd11an1n04x5 FILLER_32_1325 ();
 b15zdnd11an1n04x5 FILLER_32_1335 ();
 b15zdnd00an1n01x5 FILLER_32_1339 ();
 b15zdnd11an1n04x5 FILLER_32_1349 ();
 b15zdnd00an1n01x5 FILLER_32_1353 ();
 b15zdnd11an1n32x5 FILLER_32_1358 ();
 b15zdnd11an1n16x5 FILLER_32_1390 ();
 b15zdnd11an1n04x5 FILLER_32_1406 ();
 b15zdnd00an1n02x5 FILLER_32_1410 ();
 b15zdnd11an1n32x5 FILLER_32_1423 ();
 b15zdnd11an1n64x5 FILLER_32_1460 ();
 b15zdnd11an1n32x5 FILLER_32_1524 ();
 b15zdnd11an1n16x5 FILLER_32_1556 ();
 b15zdnd00an1n02x5 FILLER_32_1572 ();
 b15zdnd00an1n01x5 FILLER_32_1574 ();
 b15zdnd11an1n16x5 FILLER_32_1587 ();
 b15zdnd11an1n08x5 FILLER_32_1603 ();
 b15zdnd00an1n01x5 FILLER_32_1611 ();
 b15zdnd11an1n32x5 FILLER_32_1626 ();
 b15zdnd11an1n04x5 FILLER_32_1663 ();
 b15zdnd00an1n02x5 FILLER_32_1667 ();
 b15zdnd11an1n32x5 FILLER_32_1681 ();
 b15zdnd11an1n16x5 FILLER_32_1713 ();
 b15zdnd11an1n08x5 FILLER_32_1729 ();
 b15zdnd11an1n04x5 FILLER_32_1737 ();
 b15zdnd00an1n02x5 FILLER_32_1741 ();
 b15zdnd00an1n01x5 FILLER_32_1743 ();
 b15zdnd11an1n08x5 FILLER_32_1749 ();
 b15zdnd00an1n02x5 FILLER_32_1757 ();
 b15zdnd11an1n04x5 FILLER_32_1772 ();
 b15zdnd11an1n64x5 FILLER_32_1785 ();
 b15zdnd11an1n16x5 FILLER_32_1849 ();
 b15zdnd11an1n04x5 FILLER_32_1865 ();
 b15zdnd11an1n32x5 FILLER_32_1876 ();
 b15zdnd11an1n04x5 FILLER_32_1908 ();
 b15zdnd11an1n16x5 FILLER_32_1924 ();
 b15zdnd11an1n08x5 FILLER_32_1940 ();
 b15zdnd00an1n02x5 FILLER_32_1948 ();
 b15zdnd11an1n32x5 FILLER_32_1964 ();
 b15zdnd11an1n04x5 FILLER_32_1996 ();
 b15zdnd00an1n01x5 FILLER_32_2000 ();
 b15zdnd11an1n04x5 FILLER_32_2012 ();
 b15zdnd00an1n01x5 FILLER_32_2016 ();
 b15zdnd11an1n04x5 FILLER_32_2043 ();
 b15zdnd00an1n02x5 FILLER_32_2047 ();
 b15zdnd11an1n04x5 FILLER_32_2056 ();
 b15zdnd00an1n02x5 FILLER_32_2060 ();
 b15zdnd11an1n04x5 FILLER_32_2076 ();
 b15zdnd00an1n02x5 FILLER_32_2080 ();
 b15zdnd11an1n32x5 FILLER_32_2094 ();
 b15zdnd11an1n16x5 FILLER_32_2126 ();
 b15zdnd11an1n08x5 FILLER_32_2142 ();
 b15zdnd11an1n04x5 FILLER_32_2150 ();
 b15zdnd11an1n08x5 FILLER_32_2162 ();
 b15zdnd00an1n01x5 FILLER_32_2170 ();
 b15zdnd11an1n04x5 FILLER_32_2184 ();
 b15zdnd11an1n08x5 FILLER_32_2197 ();
 b15zdnd11an1n32x5 FILLER_32_2214 ();
 b15zdnd11an1n16x5 FILLER_32_2246 ();
 b15zdnd11an1n08x5 FILLER_32_2262 ();
 b15zdnd11an1n04x5 FILLER_32_2270 ();
 b15zdnd00an1n02x5 FILLER_32_2274 ();
 b15zdnd11an1n64x5 FILLER_33_0 ();
 b15zdnd11an1n08x5 FILLER_33_64 ();
 b15zdnd00an1n02x5 FILLER_33_72 ();
 b15zdnd00an1n01x5 FILLER_33_74 ();
 b15zdnd11an1n04x5 FILLER_33_82 ();
 b15zdnd11an1n16x5 FILLER_33_97 ();
 b15zdnd11an1n08x5 FILLER_33_113 ();
 b15zdnd00an1n01x5 FILLER_33_121 ();
 b15zdnd11an1n16x5 FILLER_33_138 ();
 b15zdnd11an1n08x5 FILLER_33_154 ();
 b15zdnd00an1n02x5 FILLER_33_162 ();
 b15zdnd11an1n32x5 FILLER_33_172 ();
 b15zdnd11an1n08x5 FILLER_33_204 ();
 b15zdnd11an1n04x5 FILLER_33_212 ();
 b15zdnd00an1n02x5 FILLER_33_216 ();
 b15zdnd00an1n01x5 FILLER_33_218 ();
 b15zdnd11an1n64x5 FILLER_33_228 ();
 b15zdnd11an1n04x5 FILLER_33_292 ();
 b15zdnd00an1n02x5 FILLER_33_296 ();
 b15zdnd11an1n04x5 FILLER_33_303 ();
 b15zdnd00an1n01x5 FILLER_33_307 ();
 b15zdnd11an1n64x5 FILLER_33_321 ();
 b15zdnd11an1n64x5 FILLER_33_385 ();
 b15zdnd11an1n08x5 FILLER_33_449 ();
 b15zdnd11an1n04x5 FILLER_33_457 ();
 b15zdnd00an1n02x5 FILLER_33_461 ();
 b15zdnd11an1n16x5 FILLER_33_477 ();
 b15zdnd00an1n01x5 FILLER_33_493 ();
 b15zdnd11an1n16x5 FILLER_33_498 ();
 b15zdnd11an1n08x5 FILLER_33_514 ();
 b15zdnd00an1n02x5 FILLER_33_522 ();
 b15zdnd00an1n01x5 FILLER_33_524 ();
 b15zdnd11an1n08x5 FILLER_33_530 ();
 b15zdnd11an1n08x5 FILLER_33_547 ();
 b15zdnd11an1n04x5 FILLER_33_555 ();
 b15zdnd00an1n01x5 FILLER_33_559 ();
 b15zdnd11an1n64x5 FILLER_33_567 ();
 b15zdnd00an1n02x5 FILLER_33_631 ();
 b15zdnd00an1n01x5 FILLER_33_633 ();
 b15zdnd11an1n08x5 FILLER_33_639 ();
 b15zdnd11an1n04x5 FILLER_33_647 ();
 b15zdnd00an1n01x5 FILLER_33_651 ();
 b15zdnd11an1n08x5 FILLER_33_658 ();
 b15zdnd00an1n02x5 FILLER_33_666 ();
 b15zdnd11an1n04x5 FILLER_33_674 ();
 b15zdnd00an1n02x5 FILLER_33_678 ();
 b15zdnd11an1n32x5 FILLER_33_701 ();
 b15zdnd11an1n16x5 FILLER_33_733 ();
 b15zdnd00an1n02x5 FILLER_33_749 ();
 b15zdnd00an1n01x5 FILLER_33_751 ();
 b15zdnd11an1n32x5 FILLER_33_762 ();
 b15zdnd11an1n16x5 FILLER_33_794 ();
 b15zdnd00an1n02x5 FILLER_33_810 ();
 b15zdnd00an1n01x5 FILLER_33_812 ();
 b15zdnd11an1n04x5 FILLER_33_819 ();
 b15zdnd11an1n04x5 FILLER_33_829 ();
 b15zdnd11an1n64x5 FILLER_33_859 ();
 b15zdnd11an1n32x5 FILLER_33_923 ();
 b15zdnd11an1n16x5 FILLER_33_955 ();
 b15zdnd11an1n04x5 FILLER_33_971 ();
 b15zdnd00an1n02x5 FILLER_33_975 ();
 b15zdnd11an1n04x5 FILLER_33_987 ();
 b15zdnd11an1n08x5 FILLER_33_1003 ();
 b15zdnd11an1n04x5 FILLER_33_1011 ();
 b15zdnd00an1n02x5 FILLER_33_1015 ();
 b15zdnd11an1n64x5 FILLER_33_1042 ();
 b15zdnd11an1n32x5 FILLER_33_1106 ();
 b15zdnd11an1n08x5 FILLER_33_1138 ();
 b15zdnd11an1n04x5 FILLER_33_1146 ();
 b15zdnd00an1n01x5 FILLER_33_1150 ();
 b15zdnd11an1n32x5 FILLER_33_1156 ();
 b15zdnd00an1n02x5 FILLER_33_1188 ();
 b15zdnd00an1n01x5 FILLER_33_1190 ();
 b15zdnd11an1n32x5 FILLER_33_1211 ();
 b15zdnd11an1n16x5 FILLER_33_1243 ();
 b15zdnd00an1n02x5 FILLER_33_1259 ();
 b15zdnd11an1n16x5 FILLER_33_1272 ();
 b15zdnd00an1n01x5 FILLER_33_1288 ();
 b15zdnd11an1n32x5 FILLER_33_1310 ();
 b15zdnd11an1n04x5 FILLER_33_1342 ();
 b15zdnd11an1n32x5 FILLER_33_1358 ();
 b15zdnd11an1n04x5 FILLER_33_1390 ();
 b15zdnd00an1n01x5 FILLER_33_1394 ();
 b15zdnd11an1n08x5 FILLER_33_1398 ();
 b15zdnd11an1n04x5 FILLER_33_1406 ();
 b15zdnd11an1n32x5 FILLER_33_1414 ();
 b15zdnd11an1n08x5 FILLER_33_1446 ();
 b15zdnd00an1n02x5 FILLER_33_1454 ();
 b15zdnd11an1n04x5 FILLER_33_1462 ();
 b15zdnd11an1n32x5 FILLER_33_1471 ();
 b15zdnd11an1n04x5 FILLER_33_1503 ();
 b15zdnd00an1n01x5 FILLER_33_1507 ();
 b15zdnd11an1n16x5 FILLER_33_1517 ();
 b15zdnd11an1n04x5 FILLER_33_1533 ();
 b15zdnd00an1n01x5 FILLER_33_1537 ();
 b15zdnd11an1n32x5 FILLER_33_1543 ();
 b15zdnd00an1n02x5 FILLER_33_1575 ();
 b15zdnd11an1n32x5 FILLER_33_1582 ();
 b15zdnd00an1n01x5 FILLER_33_1614 ();
 b15zdnd11an1n08x5 FILLER_33_1620 ();
 b15zdnd11an1n04x5 FILLER_33_1628 ();
 b15zdnd11an1n16x5 FILLER_33_1641 ();
 b15zdnd11an1n08x5 FILLER_33_1657 ();
 b15zdnd00an1n01x5 FILLER_33_1665 ();
 b15zdnd11an1n64x5 FILLER_33_1671 ();
 b15zdnd11an1n16x5 FILLER_33_1735 ();
 b15zdnd11an1n08x5 FILLER_33_1751 ();
 b15zdnd11an1n04x5 FILLER_33_1759 ();
 b15zdnd00an1n01x5 FILLER_33_1763 ();
 b15zdnd11an1n32x5 FILLER_33_1790 ();
 b15zdnd11an1n04x5 FILLER_33_1822 ();
 b15zdnd00an1n02x5 FILLER_33_1826 ();
 b15zdnd00an1n01x5 FILLER_33_1828 ();
 b15zdnd11an1n08x5 FILLER_33_1835 ();
 b15zdnd11an1n04x5 FILLER_33_1843 ();
 b15zdnd00an1n02x5 FILLER_33_1847 ();
 b15zdnd00an1n01x5 FILLER_33_1849 ();
 b15zdnd11an1n16x5 FILLER_33_1855 ();
 b15zdnd11an1n04x5 FILLER_33_1871 ();
 b15zdnd00an1n02x5 FILLER_33_1875 ();
 b15zdnd00an1n01x5 FILLER_33_1877 ();
 b15zdnd11an1n64x5 FILLER_33_1883 ();
 b15zdnd11an1n64x5 FILLER_33_1947 ();
 b15zdnd11an1n32x5 FILLER_33_2011 ();
 b15zdnd11an1n08x5 FILLER_33_2043 ();
 b15zdnd11an1n04x5 FILLER_33_2064 ();
 b15zdnd11an1n32x5 FILLER_33_2079 ();
 b15zdnd00an1n02x5 FILLER_33_2111 ();
 b15zdnd00an1n01x5 FILLER_33_2113 ();
 b15zdnd11an1n04x5 FILLER_33_2122 ();
 b15zdnd11an1n08x5 FILLER_33_2140 ();
 b15zdnd11an1n04x5 FILLER_33_2148 ();
 b15zdnd00an1n01x5 FILLER_33_2152 ();
 b15zdnd11an1n04x5 FILLER_33_2158 ();
 b15zdnd11an1n04x5 FILLER_33_2169 ();
 b15zdnd00an1n02x5 FILLER_33_2173 ();
 b15zdnd11an1n04x5 FILLER_33_2182 ();
 b15zdnd00an1n02x5 FILLER_33_2186 ();
 b15zdnd11an1n16x5 FILLER_33_2192 ();
 b15zdnd00an1n01x5 FILLER_33_2208 ();
 b15zdnd11an1n64x5 FILLER_33_2213 ();
 b15zdnd11an1n04x5 FILLER_33_2277 ();
 b15zdnd00an1n02x5 FILLER_33_2281 ();
 b15zdnd00an1n01x5 FILLER_33_2283 ();
 b15zdnd11an1n16x5 FILLER_34_8 ();
 b15zdnd11an1n08x5 FILLER_34_24 ();
 b15zdnd11an1n04x5 FILLER_34_32 ();
 b15zdnd11an1n16x5 FILLER_34_48 ();
 b15zdnd11an1n08x5 FILLER_34_64 ();
 b15zdnd11an1n04x5 FILLER_34_72 ();
 b15zdnd00an1n02x5 FILLER_34_76 ();
 b15zdnd11an1n08x5 FILLER_34_82 ();
 b15zdnd11an1n04x5 FILLER_34_90 ();
 b15zdnd00an1n02x5 FILLER_34_94 ();
 b15zdnd11an1n04x5 FILLER_34_119 ();
 b15zdnd11an1n16x5 FILLER_34_130 ();
 b15zdnd11an1n08x5 FILLER_34_146 ();
 b15zdnd11an1n64x5 FILLER_34_160 ();
 b15zdnd11an1n64x5 FILLER_34_224 ();
 b15zdnd11an1n08x5 FILLER_34_288 ();
 b15zdnd00an1n02x5 FILLER_34_296 ();
 b15zdnd00an1n01x5 FILLER_34_298 ();
 b15zdnd11an1n32x5 FILLER_34_311 ();
 b15zdnd11an1n08x5 FILLER_34_343 ();
 b15zdnd11an1n04x5 FILLER_34_351 ();
 b15zdnd11an1n32x5 FILLER_34_369 ();
 b15zdnd11an1n08x5 FILLER_34_401 ();
 b15zdnd11an1n04x5 FILLER_34_409 ();
 b15zdnd11an1n32x5 FILLER_34_423 ();
 b15zdnd11an1n08x5 FILLER_34_455 ();
 b15zdnd00an1n02x5 FILLER_34_463 ();
 b15zdnd00an1n01x5 FILLER_34_465 ();
 b15zdnd11an1n32x5 FILLER_34_471 ();
 b15zdnd11an1n08x5 FILLER_34_503 ();
 b15zdnd11an1n04x5 FILLER_34_511 ();
 b15zdnd11an1n16x5 FILLER_34_521 ();
 b15zdnd00an1n02x5 FILLER_34_537 ();
 b15zdnd11an1n16x5 FILLER_34_543 ();
 b15zdnd11an1n08x5 FILLER_34_563 ();
 b15zdnd11an1n04x5 FILLER_34_571 ();
 b15zdnd00an1n02x5 FILLER_34_575 ();
 b15zdnd00an1n01x5 FILLER_34_577 ();
 b15zdnd11an1n04x5 FILLER_34_590 ();
 b15zdnd11an1n16x5 FILLER_34_601 ();
 b15zdnd11an1n08x5 FILLER_34_617 ();
 b15zdnd00an1n01x5 FILLER_34_625 ();
 b15zdnd11an1n04x5 FILLER_34_632 ();
 b15zdnd00an1n01x5 FILLER_34_636 ();
 b15zdnd11an1n16x5 FILLER_34_643 ();
 b15zdnd11an1n08x5 FILLER_34_659 ();
 b15zdnd11an1n04x5 FILLER_34_667 ();
 b15zdnd00an1n01x5 FILLER_34_671 ();
 b15zdnd11an1n32x5 FILLER_34_685 ();
 b15zdnd00an1n01x5 FILLER_34_717 ();
 b15zdnd11an1n08x5 FILLER_34_726 ();
 b15zdnd00an1n02x5 FILLER_34_734 ();
 b15zdnd00an1n01x5 FILLER_34_736 ();
 b15zdnd11an1n16x5 FILLER_34_743 ();
 b15zdnd11an1n04x5 FILLER_34_759 ();
 b15zdnd00an1n02x5 FILLER_34_763 ();
 b15zdnd00an1n01x5 FILLER_34_765 ();
 b15zdnd11an1n08x5 FILLER_34_773 ();
 b15zdnd11an1n04x5 FILLER_34_781 ();
 b15zdnd00an1n02x5 FILLER_34_785 ();
 b15zdnd11an1n08x5 FILLER_34_799 ();
 b15zdnd11an1n64x5 FILLER_34_816 ();
 b15zdnd00an1n02x5 FILLER_34_880 ();
 b15zdnd00an1n01x5 FILLER_34_882 ();
 b15zdnd11an1n08x5 FILLER_34_887 ();
 b15zdnd11an1n04x5 FILLER_34_895 ();
 b15zdnd00an1n02x5 FILLER_34_899 ();
 b15zdnd00an1n01x5 FILLER_34_901 ();
 b15zdnd11an1n32x5 FILLER_34_911 ();
 b15zdnd11an1n16x5 FILLER_34_943 ();
 b15zdnd11an1n04x5 FILLER_34_959 ();
 b15zdnd00an1n02x5 FILLER_34_963 ();
 b15zdnd11an1n32x5 FILLER_34_996 ();
 b15zdnd00an1n01x5 FILLER_34_1028 ();
 b15zdnd11an1n16x5 FILLER_34_1038 ();
 b15zdnd11an1n04x5 FILLER_34_1054 ();
 b15zdnd00an1n01x5 FILLER_34_1058 ();
 b15zdnd11an1n32x5 FILLER_34_1087 ();
 b15zdnd11an1n16x5 FILLER_34_1119 ();
 b15zdnd00an1n02x5 FILLER_34_1135 ();
 b15zdnd00an1n01x5 FILLER_34_1137 ();
 b15zdnd11an1n16x5 FILLER_34_1158 ();
 b15zdnd00an1n01x5 FILLER_34_1174 ();
 b15zdnd11an1n64x5 FILLER_34_1180 ();
 b15zdnd11an1n32x5 FILLER_34_1244 ();
 b15zdnd11an1n08x5 FILLER_34_1276 ();
 b15zdnd11an1n16x5 FILLER_34_1315 ();
 b15zdnd11an1n08x5 FILLER_34_1331 ();
 b15zdnd00an1n02x5 FILLER_34_1339 ();
 b15zdnd00an1n01x5 FILLER_34_1341 ();
 b15zdnd11an1n04x5 FILLER_34_1356 ();
 b15zdnd11an1n16x5 FILLER_34_1366 ();
 b15zdnd00an1n02x5 FILLER_34_1382 ();
 b15zdnd00an1n01x5 FILLER_34_1384 ();
 b15zdnd11an1n16x5 FILLER_34_1392 ();
 b15zdnd00an1n02x5 FILLER_34_1408 ();
 b15zdnd11an1n32x5 FILLER_34_1421 ();
 b15zdnd11an1n04x5 FILLER_34_1453 ();
 b15zdnd11an1n04x5 FILLER_34_1464 ();
 b15zdnd00an1n02x5 FILLER_34_1468 ();
 b15zdnd00an1n01x5 FILLER_34_1470 ();
 b15zdnd11an1n16x5 FILLER_34_1477 ();
 b15zdnd11an1n08x5 FILLER_34_1493 ();
 b15zdnd00an1n01x5 FILLER_34_1501 ();
 b15zdnd11an1n16x5 FILLER_34_1511 ();
 b15zdnd11an1n08x5 FILLER_34_1527 ();
 b15zdnd11an1n04x5 FILLER_34_1535 ();
 b15zdnd00an1n02x5 FILLER_34_1539 ();
 b15zdnd11an1n08x5 FILLER_34_1547 ();
 b15zdnd11an1n04x5 FILLER_34_1555 ();
 b15zdnd00an1n02x5 FILLER_34_1559 ();
 b15zdnd11an1n04x5 FILLER_34_1569 ();
 b15zdnd11an1n32x5 FILLER_34_1585 ();
 b15zdnd11an1n16x5 FILLER_34_1617 ();
 b15zdnd11an1n04x5 FILLER_34_1633 ();
 b15zdnd00an1n02x5 FILLER_34_1637 ();
 b15zdnd00an1n01x5 FILLER_34_1639 ();
 b15zdnd11an1n64x5 FILLER_34_1651 ();
 b15zdnd11an1n32x5 FILLER_34_1715 ();
 b15zdnd11an1n08x5 FILLER_34_1747 ();
 b15zdnd00an1n02x5 FILLER_34_1755 ();
 b15zdnd00an1n01x5 FILLER_34_1757 ();
 b15zdnd11an1n04x5 FILLER_34_1767 ();
 b15zdnd11an1n04x5 FILLER_34_1791 ();
 b15zdnd11an1n16x5 FILLER_34_1799 ();
 b15zdnd11an1n08x5 FILLER_34_1815 ();
 b15zdnd00an1n02x5 FILLER_34_1823 ();
 b15zdnd11an1n04x5 FILLER_34_1831 ();
 b15zdnd11an1n04x5 FILLER_34_1841 ();
 b15zdnd11an1n16x5 FILLER_34_1850 ();
 b15zdnd00an1n02x5 FILLER_34_1866 ();
 b15zdnd00an1n01x5 FILLER_34_1868 ();
 b15zdnd11an1n04x5 FILLER_34_1885 ();
 b15zdnd11an1n16x5 FILLER_34_1905 ();
 b15zdnd11an1n08x5 FILLER_34_1921 ();
 b15zdnd11an1n32x5 FILLER_34_1953 ();
 b15zdnd11an1n08x5 FILLER_34_1991 ();
 b15zdnd00an1n02x5 FILLER_34_1999 ();
 b15zdnd11an1n04x5 FILLER_34_2006 ();
 b15zdnd00an1n02x5 FILLER_34_2010 ();
 b15zdnd11an1n16x5 FILLER_34_2024 ();
 b15zdnd11an1n32x5 FILLER_34_2061 ();
 b15zdnd11an1n08x5 FILLER_34_2093 ();
 b15zdnd00an1n01x5 FILLER_34_2101 ();
 b15zdnd11an1n04x5 FILLER_34_2108 ();
 b15zdnd11an1n16x5 FILLER_34_2126 ();
 b15zdnd11an1n08x5 FILLER_34_2142 ();
 b15zdnd11an1n04x5 FILLER_34_2150 ();
 b15zdnd00an1n02x5 FILLER_34_2162 ();
 b15zdnd11an1n64x5 FILLER_34_2169 ();
 b15zdnd11an1n32x5 FILLER_34_2233 ();
 b15zdnd11an1n08x5 FILLER_34_2265 ();
 b15zdnd00an1n02x5 FILLER_34_2273 ();
 b15zdnd00an1n01x5 FILLER_34_2275 ();
 b15zdnd11an1n32x5 FILLER_35_0 ();
 b15zdnd11an1n08x5 FILLER_35_32 ();
 b15zdnd11an1n08x5 FILLER_35_54 ();
 b15zdnd00an1n01x5 FILLER_35_62 ();
 b15zdnd11an1n32x5 FILLER_35_75 ();
 b15zdnd11an1n08x5 FILLER_35_107 ();
 b15zdnd00an1n02x5 FILLER_35_115 ();
 b15zdnd11an1n04x5 FILLER_35_122 ();
 b15zdnd11an1n32x5 FILLER_35_131 ();
 b15zdnd11an1n16x5 FILLER_35_163 ();
 b15zdnd11an1n04x5 FILLER_35_179 ();
 b15zdnd00an1n02x5 FILLER_35_183 ();
 b15zdnd00an1n01x5 FILLER_35_185 ();
 b15zdnd11an1n04x5 FILLER_35_191 ();
 b15zdnd11an1n08x5 FILLER_35_201 ();
 b15zdnd11an1n04x5 FILLER_35_209 ();
 b15zdnd00an1n02x5 FILLER_35_213 ();
 b15zdnd00an1n01x5 FILLER_35_215 ();
 b15zdnd11an1n04x5 FILLER_35_225 ();
 b15zdnd11an1n04x5 FILLER_35_234 ();
 b15zdnd11an1n64x5 FILLER_35_245 ();
 b15zdnd11an1n64x5 FILLER_35_309 ();
 b15zdnd11an1n64x5 FILLER_35_373 ();
 b15zdnd11an1n16x5 FILLER_35_437 ();
 b15zdnd11an1n08x5 FILLER_35_453 ();
 b15zdnd00an1n02x5 FILLER_35_461 ();
 b15zdnd00an1n01x5 FILLER_35_463 ();
 b15zdnd11an1n16x5 FILLER_35_478 ();
 b15zdnd11an1n04x5 FILLER_35_494 ();
 b15zdnd00an1n01x5 FILLER_35_498 ();
 b15zdnd11an1n64x5 FILLER_35_511 ();
 b15zdnd11an1n16x5 FILLER_35_575 ();
 b15zdnd00an1n01x5 FILLER_35_591 ();
 b15zdnd11an1n32x5 FILLER_35_599 ();
 b15zdnd11an1n08x5 FILLER_35_631 ();
 b15zdnd11an1n08x5 FILLER_35_643 ();
 b15zdnd11an1n32x5 FILLER_35_679 ();
 b15zdnd11an1n08x5 FILLER_35_711 ();
 b15zdnd00an1n01x5 FILLER_35_719 ();
 b15zdnd11an1n08x5 FILLER_35_730 ();
 b15zdnd00an1n01x5 FILLER_35_738 ();
 b15zdnd11an1n08x5 FILLER_35_750 ();
 b15zdnd11an1n04x5 FILLER_35_758 ();
 b15zdnd00an1n02x5 FILLER_35_762 ();
 b15zdnd11an1n64x5 FILLER_35_780 ();
 b15zdnd11an1n16x5 FILLER_35_844 ();
 b15zdnd11an1n04x5 FILLER_35_865 ();
 b15zdnd11an1n04x5 FILLER_35_878 ();
 b15zdnd00an1n02x5 FILLER_35_882 ();
 b15zdnd11an1n64x5 FILLER_35_892 ();
 b15zdnd11an1n64x5 FILLER_35_956 ();
 b15zdnd11an1n32x5 FILLER_35_1020 ();
 b15zdnd11an1n08x5 FILLER_35_1052 ();
 b15zdnd11an1n08x5 FILLER_35_1069 ();
 b15zdnd11an1n04x5 FILLER_35_1077 ();
 b15zdnd00an1n02x5 FILLER_35_1081 ();
 b15zdnd11an1n04x5 FILLER_35_1114 ();
 b15zdnd00an1n01x5 FILLER_35_1118 ();
 b15zdnd11an1n08x5 FILLER_35_1139 ();
 b15zdnd00an1n02x5 FILLER_35_1147 ();
 b15zdnd00an1n01x5 FILLER_35_1149 ();
 b15zdnd11an1n16x5 FILLER_35_1154 ();
 b15zdnd11an1n64x5 FILLER_35_1190 ();
 b15zdnd11an1n64x5 FILLER_35_1254 ();
 b15zdnd11an1n32x5 FILLER_35_1318 ();
 b15zdnd11an1n16x5 FILLER_35_1350 ();
 b15zdnd11an1n08x5 FILLER_35_1366 ();
 b15zdnd11an1n04x5 FILLER_35_1374 ();
 b15zdnd11an1n08x5 FILLER_35_1385 ();
 b15zdnd11an1n04x5 FILLER_35_1393 ();
 b15zdnd00an1n02x5 FILLER_35_1397 ();
 b15zdnd00an1n01x5 FILLER_35_1399 ();
 b15zdnd11an1n32x5 FILLER_35_1406 ();
 b15zdnd11an1n16x5 FILLER_35_1438 ();
 b15zdnd11an1n08x5 FILLER_35_1454 ();
 b15zdnd11an1n04x5 FILLER_35_1462 ();
 b15zdnd00an1n02x5 FILLER_35_1466 ();
 b15zdnd00an1n01x5 FILLER_35_1468 ();
 b15zdnd11an1n16x5 FILLER_35_1475 ();
 b15zdnd11an1n08x5 FILLER_35_1491 ();
 b15zdnd11an1n04x5 FILLER_35_1499 ();
 b15zdnd00an1n01x5 FILLER_35_1503 ();
 b15zdnd11an1n16x5 FILLER_35_1522 ();
 b15zdnd00an1n02x5 FILLER_35_1538 ();
 b15zdnd00an1n01x5 FILLER_35_1540 ();
 b15zdnd11an1n64x5 FILLER_35_1546 ();
 b15zdnd11an1n64x5 FILLER_35_1610 ();
 b15zdnd11an1n16x5 FILLER_35_1674 ();
 b15zdnd00an1n02x5 FILLER_35_1690 ();
 b15zdnd00an1n01x5 FILLER_35_1692 ();
 b15zdnd11an1n16x5 FILLER_35_1713 ();
 b15zdnd11an1n04x5 FILLER_35_1729 ();
 b15zdnd11an1n08x5 FILLER_35_1759 ();
 b15zdnd11an1n04x5 FILLER_35_1779 ();
 b15zdnd11an1n32x5 FILLER_35_1797 ();
 b15zdnd11an1n16x5 FILLER_35_1829 ();
 b15zdnd11an1n04x5 FILLER_35_1851 ();
 b15zdnd11an1n16x5 FILLER_35_1864 ();
 b15zdnd11an1n08x5 FILLER_35_1880 ();
 b15zdnd11an1n04x5 FILLER_35_1888 ();
 b15zdnd00an1n01x5 FILLER_35_1892 ();
 b15zdnd11an1n08x5 FILLER_35_1905 ();
 b15zdnd00an1n02x5 FILLER_35_1913 ();
 b15zdnd11an1n08x5 FILLER_35_1925 ();
 b15zdnd00an1n01x5 FILLER_35_1933 ();
 b15zdnd11an1n16x5 FILLER_35_1953 ();
 b15zdnd11an1n08x5 FILLER_35_1969 ();
 b15zdnd00an1n01x5 FILLER_35_1977 ();
 b15zdnd11an1n32x5 FILLER_35_1985 ();
 b15zdnd00an1n02x5 FILLER_35_2017 ();
 b15zdnd11an1n64x5 FILLER_35_2024 ();
 b15zdnd11an1n08x5 FILLER_35_2088 ();
 b15zdnd11an1n04x5 FILLER_35_2096 ();
 b15zdnd11an1n04x5 FILLER_35_2114 ();
 b15zdnd11an1n64x5 FILLER_35_2124 ();
 b15zdnd11an1n08x5 FILLER_35_2188 ();
 b15zdnd11an1n64x5 FILLER_35_2211 ();
 b15zdnd11an1n08x5 FILLER_35_2275 ();
 b15zdnd00an1n01x5 FILLER_35_2283 ();
 b15zdnd11an1n16x5 FILLER_36_8 ();
 b15zdnd11an1n08x5 FILLER_36_24 ();
 b15zdnd00an1n02x5 FILLER_36_32 ();
 b15zdnd00an1n01x5 FILLER_36_34 ();
 b15zdnd11an1n64x5 FILLER_36_51 ();
 b15zdnd11an1n32x5 FILLER_36_115 ();
 b15zdnd11an1n16x5 FILLER_36_147 ();
 b15zdnd11an1n08x5 FILLER_36_163 ();
 b15zdnd11an1n08x5 FILLER_36_176 ();
 b15zdnd11an1n04x5 FILLER_36_184 ();
 b15zdnd11an1n32x5 FILLER_36_194 ();
 b15zdnd11an1n16x5 FILLER_36_226 ();
 b15zdnd11an1n08x5 FILLER_36_242 ();
 b15zdnd00an1n02x5 FILLER_36_250 ();
 b15zdnd11an1n04x5 FILLER_36_259 ();
 b15zdnd00an1n02x5 FILLER_36_263 ();
 b15zdnd11an1n16x5 FILLER_36_277 ();
 b15zdnd00an1n01x5 FILLER_36_293 ();
 b15zdnd11an1n04x5 FILLER_36_302 ();
 b15zdnd11an1n64x5 FILLER_36_312 ();
 b15zdnd11an1n32x5 FILLER_36_376 ();
 b15zdnd11an1n08x5 FILLER_36_408 ();
 b15zdnd00an1n01x5 FILLER_36_416 ();
 b15zdnd11an1n04x5 FILLER_36_423 ();
 b15zdnd11an1n32x5 FILLER_36_439 ();
 b15zdnd11an1n16x5 FILLER_36_471 ();
 b15zdnd11an1n08x5 FILLER_36_487 ();
 b15zdnd11an1n04x5 FILLER_36_495 ();
 b15zdnd11an1n04x5 FILLER_36_505 ();
 b15zdnd11an1n16x5 FILLER_36_521 ();
 b15zdnd11an1n04x5 FILLER_36_537 ();
 b15zdnd00an1n02x5 FILLER_36_541 ();
 b15zdnd11an1n64x5 FILLER_36_548 ();
 b15zdnd11an1n32x5 FILLER_36_612 ();
 b15zdnd11an1n08x5 FILLER_36_644 ();
 b15zdnd00an1n02x5 FILLER_36_652 ();
 b15zdnd11an1n32x5 FILLER_36_658 ();
 b15zdnd11an1n16x5 FILLER_36_690 ();
 b15zdnd11an1n08x5 FILLER_36_706 ();
 b15zdnd11an1n04x5 FILLER_36_714 ();
 b15zdnd11an1n08x5 FILLER_36_726 ();
 b15zdnd11an1n04x5 FILLER_36_734 ();
 b15zdnd00an1n01x5 FILLER_36_738 ();
 b15zdnd11an1n04x5 FILLER_36_744 ();
 b15zdnd11an1n16x5 FILLER_36_768 ();
 b15zdnd00an1n02x5 FILLER_36_784 ();
 b15zdnd11an1n32x5 FILLER_36_791 ();
 b15zdnd11an1n16x5 FILLER_36_823 ();
 b15zdnd11an1n08x5 FILLER_36_839 ();
 b15zdnd00an1n01x5 FILLER_36_847 ();
 b15zdnd11an1n04x5 FILLER_36_868 ();
 b15zdnd11an1n04x5 FILLER_36_888 ();
 b15zdnd11an1n04x5 FILLER_36_902 ();
 b15zdnd11an1n32x5 FILLER_36_926 ();
 b15zdnd11an1n04x5 FILLER_36_963 ();
 b15zdnd00an1n02x5 FILLER_36_967 ();
 b15zdnd11an1n64x5 FILLER_36_973 ();
 b15zdnd11an1n16x5 FILLER_36_1037 ();
 b15zdnd11an1n08x5 FILLER_36_1053 ();
 b15zdnd00an1n02x5 FILLER_36_1061 ();
 b15zdnd00an1n01x5 FILLER_36_1063 ();
 b15zdnd11an1n64x5 FILLER_36_1085 ();
 b15zdnd11an1n32x5 FILLER_36_1149 ();
 b15zdnd00an1n02x5 FILLER_36_1181 ();
 b15zdnd11an1n16x5 FILLER_36_1186 ();
 b15zdnd11an1n08x5 FILLER_36_1202 ();
 b15zdnd11an1n04x5 FILLER_36_1210 ();
 b15zdnd00an1n02x5 FILLER_36_1214 ();
 b15zdnd11an1n64x5 FILLER_36_1221 ();
 b15zdnd11an1n32x5 FILLER_36_1285 ();
 b15zdnd11an1n04x5 FILLER_36_1317 ();
 b15zdnd11an1n32x5 FILLER_36_1326 ();
 b15zdnd11an1n16x5 FILLER_36_1358 ();
 b15zdnd11an1n04x5 FILLER_36_1374 ();
 b15zdnd00an1n01x5 FILLER_36_1378 ();
 b15zdnd11an1n16x5 FILLER_36_1389 ();
 b15zdnd11an1n04x5 FILLER_36_1419 ();
 b15zdnd00an1n01x5 FILLER_36_1423 ();
 b15zdnd11an1n32x5 FILLER_36_1434 ();
 b15zdnd11an1n04x5 FILLER_36_1466 ();
 b15zdnd00an1n02x5 FILLER_36_1470 ();
 b15zdnd11an1n04x5 FILLER_36_1487 ();
 b15zdnd11an1n04x5 FILLER_36_1496 ();
 b15zdnd11an1n32x5 FILLER_36_1505 ();
 b15zdnd11an1n08x5 FILLER_36_1537 ();
 b15zdnd00an1n01x5 FILLER_36_1545 ();
 b15zdnd11an1n32x5 FILLER_36_1552 ();
 b15zdnd11an1n08x5 FILLER_36_1584 ();
 b15zdnd00an1n01x5 FILLER_36_1592 ();
 b15zdnd11an1n16x5 FILLER_36_1597 ();
 b15zdnd11an1n08x5 FILLER_36_1613 ();
 b15zdnd11an1n04x5 FILLER_36_1621 ();
 b15zdnd00an1n01x5 FILLER_36_1625 ();
 b15zdnd11an1n16x5 FILLER_36_1632 ();
 b15zdnd11an1n08x5 FILLER_36_1648 ();
 b15zdnd00an1n02x5 FILLER_36_1656 ();
 b15zdnd00an1n01x5 FILLER_36_1658 ();
 b15zdnd11an1n64x5 FILLER_36_1666 ();
 b15zdnd11an1n64x5 FILLER_36_1730 ();
 b15zdnd11an1n08x5 FILLER_36_1794 ();
 b15zdnd11an1n04x5 FILLER_36_1802 ();
 b15zdnd00an1n02x5 FILLER_36_1806 ();
 b15zdnd11an1n64x5 FILLER_36_1814 ();
 b15zdnd11an1n32x5 FILLER_36_1878 ();
 b15zdnd11an1n04x5 FILLER_36_1910 ();
 b15zdnd11an1n04x5 FILLER_36_1926 ();
 b15zdnd11an1n32x5 FILLER_36_1945 ();
 b15zdnd00an1n02x5 FILLER_36_1977 ();
 b15zdnd11an1n16x5 FILLER_36_1986 ();
 b15zdnd11an1n08x5 FILLER_36_2002 ();
 b15zdnd00an1n01x5 FILLER_36_2010 ();
 b15zdnd11an1n16x5 FILLER_36_2015 ();
 b15zdnd11an1n08x5 FILLER_36_2031 ();
 b15zdnd11an1n04x5 FILLER_36_2039 ();
 b15zdnd00an1n02x5 FILLER_36_2043 ();
 b15zdnd11an1n64x5 FILLER_36_2049 ();
 b15zdnd11an1n08x5 FILLER_36_2113 ();
 b15zdnd00an1n01x5 FILLER_36_2121 ();
 b15zdnd11an1n16x5 FILLER_36_2135 ();
 b15zdnd00an1n02x5 FILLER_36_2151 ();
 b15zdnd00an1n01x5 FILLER_36_2153 ();
 b15zdnd11an1n32x5 FILLER_36_2162 ();
 b15zdnd11an1n08x5 FILLER_36_2194 ();
 b15zdnd11an1n32x5 FILLER_36_2218 ();
 b15zdnd11an1n16x5 FILLER_36_2250 ();
 b15zdnd11an1n08x5 FILLER_36_2266 ();
 b15zdnd00an1n02x5 FILLER_36_2274 ();
 b15zdnd11an1n64x5 FILLER_37_0 ();
 b15zdnd11an1n04x5 FILLER_37_64 ();
 b15zdnd11an1n32x5 FILLER_37_80 ();
 b15zdnd11an1n16x5 FILLER_37_112 ();
 b15zdnd11an1n08x5 FILLER_37_128 ();
 b15zdnd00an1n01x5 FILLER_37_136 ();
 b15zdnd11an1n32x5 FILLER_37_149 ();
 b15zdnd11an1n16x5 FILLER_37_181 ();
 b15zdnd11an1n08x5 FILLER_37_197 ();
 b15zdnd00an1n02x5 FILLER_37_205 ();
 b15zdnd00an1n01x5 FILLER_37_207 ();
 b15zdnd11an1n16x5 FILLER_37_218 ();
 b15zdnd11an1n08x5 FILLER_37_234 ();
 b15zdnd11an1n04x5 FILLER_37_272 ();
 b15zdnd11an1n04x5 FILLER_37_290 ();
 b15zdnd11an1n08x5 FILLER_37_305 ();
 b15zdnd00an1n02x5 FILLER_37_313 ();
 b15zdnd11an1n64x5 FILLER_37_320 ();
 b15zdnd11an1n32x5 FILLER_37_384 ();
 b15zdnd00an1n02x5 FILLER_37_416 ();
 b15zdnd11an1n04x5 FILLER_37_424 ();
 b15zdnd11an1n32x5 FILLER_37_434 ();
 b15zdnd11an1n16x5 FILLER_37_466 ();
 b15zdnd11an1n08x5 FILLER_37_482 ();
 b15zdnd11an1n04x5 FILLER_37_490 ();
 b15zdnd00an1n01x5 FILLER_37_494 ();
 b15zdnd11an1n16x5 FILLER_37_509 ();
 b15zdnd11an1n08x5 FILLER_37_525 ();
 b15zdnd00an1n02x5 FILLER_37_533 ();
 b15zdnd00an1n01x5 FILLER_37_535 ();
 b15zdnd11an1n32x5 FILLER_37_546 ();
 b15zdnd11an1n04x5 FILLER_37_578 ();
 b15zdnd11an1n32x5 FILLER_37_588 ();
 b15zdnd11an1n08x5 FILLER_37_620 ();
 b15zdnd11an1n04x5 FILLER_37_628 ();
 b15zdnd00an1n02x5 FILLER_37_632 ();
 b15zdnd00an1n01x5 FILLER_37_634 ();
 b15zdnd11an1n32x5 FILLER_37_641 ();
 b15zdnd00an1n02x5 FILLER_37_673 ();
 b15zdnd00an1n01x5 FILLER_37_675 ();
 b15zdnd11an1n04x5 FILLER_37_684 ();
 b15zdnd11an1n16x5 FILLER_37_699 ();
 b15zdnd11an1n04x5 FILLER_37_715 ();
 b15zdnd11an1n64x5 FILLER_37_733 ();
 b15zdnd11an1n08x5 FILLER_37_797 ();
 b15zdnd11an1n04x5 FILLER_37_805 ();
 b15zdnd00an1n02x5 FILLER_37_809 ();
 b15zdnd11an1n04x5 FILLER_37_818 ();
 b15zdnd11an1n64x5 FILLER_37_834 ();
 b15zdnd11an1n32x5 FILLER_37_898 ();
 b15zdnd11an1n16x5 FILLER_37_930 ();
 b15zdnd11an1n08x5 FILLER_37_946 ();
 b15zdnd11an1n04x5 FILLER_37_954 ();
 b15zdnd00an1n01x5 FILLER_37_958 ();
 b15zdnd11an1n32x5 FILLER_37_979 ();
 b15zdnd11an1n08x5 FILLER_37_1036 ();
 b15zdnd11an1n04x5 FILLER_37_1044 ();
 b15zdnd00an1n02x5 FILLER_37_1048 ();
 b15zdnd00an1n01x5 FILLER_37_1050 ();
 b15zdnd11an1n32x5 FILLER_37_1061 ();
 b15zdnd11an1n16x5 FILLER_37_1093 ();
 b15zdnd11an1n04x5 FILLER_37_1109 ();
 b15zdnd00an1n01x5 FILLER_37_1113 ();
 b15zdnd11an1n32x5 FILLER_37_1123 ();
 b15zdnd00an1n02x5 FILLER_37_1155 ();
 b15zdnd00an1n01x5 FILLER_37_1157 ();
 b15zdnd11an1n32x5 FILLER_37_1168 ();
 b15zdnd11an1n08x5 FILLER_37_1200 ();
 b15zdnd00an1n02x5 FILLER_37_1208 ();
 b15zdnd11an1n64x5 FILLER_37_1219 ();
 b15zdnd11an1n32x5 FILLER_37_1283 ();
 b15zdnd00an1n02x5 FILLER_37_1315 ();
 b15zdnd00an1n01x5 FILLER_37_1317 ();
 b15zdnd11an1n04x5 FILLER_37_1322 ();
 b15zdnd00an1n01x5 FILLER_37_1326 ();
 b15zdnd11an1n64x5 FILLER_37_1332 ();
 b15zdnd11an1n08x5 FILLER_37_1396 ();
 b15zdnd11an1n04x5 FILLER_37_1404 ();
 b15zdnd00an1n01x5 FILLER_37_1408 ();
 b15zdnd11an1n08x5 FILLER_37_1415 ();
 b15zdnd00an1n02x5 FILLER_37_1423 ();
 b15zdnd00an1n01x5 FILLER_37_1425 ();
 b15zdnd11an1n32x5 FILLER_37_1444 ();
 b15zdnd11an1n16x5 FILLER_37_1476 ();
 b15zdnd00an1n01x5 FILLER_37_1492 ();
 b15zdnd11an1n08x5 FILLER_37_1503 ();
 b15zdnd00an1n01x5 FILLER_37_1511 ();
 b15zdnd11an1n04x5 FILLER_37_1517 ();
 b15zdnd11an1n04x5 FILLER_37_1542 ();
 b15zdnd11an1n04x5 FILLER_37_1556 ();
 b15zdnd00an1n01x5 FILLER_37_1560 ();
 b15zdnd11an1n32x5 FILLER_37_1566 ();
 b15zdnd11an1n08x5 FILLER_37_1598 ();
 b15zdnd00an1n02x5 FILLER_37_1606 ();
 b15zdnd00an1n01x5 FILLER_37_1608 ();
 b15zdnd11an1n04x5 FILLER_37_1624 ();
 b15zdnd11an1n08x5 FILLER_37_1633 ();
 b15zdnd11an1n04x5 FILLER_37_1641 ();
 b15zdnd00an1n01x5 FILLER_37_1645 ();
 b15zdnd11an1n08x5 FILLER_37_1653 ();
 b15zdnd11an1n64x5 FILLER_37_1674 ();
 b15zdnd11an1n08x5 FILLER_37_1738 ();
 b15zdnd11an1n04x5 FILLER_37_1746 ();
 b15zdnd00an1n02x5 FILLER_37_1750 ();
 b15zdnd11an1n04x5 FILLER_37_1759 ();
 b15zdnd11an1n16x5 FILLER_37_1769 ();
 b15zdnd11an1n08x5 FILLER_37_1785 ();
 b15zdnd11an1n04x5 FILLER_37_1793 ();
 b15zdnd00an1n01x5 FILLER_37_1797 ();
 b15zdnd11an1n32x5 FILLER_37_1809 ();
 b15zdnd11an1n16x5 FILLER_37_1841 ();
 b15zdnd11an1n08x5 FILLER_37_1857 ();
 b15zdnd11an1n04x5 FILLER_37_1865 ();
 b15zdnd11an1n32x5 FILLER_37_1884 ();
 b15zdnd00an1n02x5 FILLER_37_1916 ();
 b15zdnd11an1n16x5 FILLER_37_1938 ();
 b15zdnd00an1n01x5 FILLER_37_1954 ();
 b15zdnd11an1n16x5 FILLER_37_1960 ();
 b15zdnd00an1n01x5 FILLER_37_1976 ();
 b15zdnd11an1n64x5 FILLER_37_1989 ();
 b15zdnd11an1n32x5 FILLER_37_2053 ();
 b15zdnd00an1n02x5 FILLER_37_2085 ();
 b15zdnd00an1n01x5 FILLER_37_2087 ();
 b15zdnd11an1n32x5 FILLER_37_2096 ();
 b15zdnd11an1n08x5 FILLER_37_2128 ();
 b15zdnd11an1n04x5 FILLER_37_2136 ();
 b15zdnd00an1n01x5 FILLER_37_2140 ();
 b15zdnd11an1n32x5 FILLER_37_2159 ();
 b15zdnd00an1n02x5 FILLER_37_2191 ();
 b15zdnd11an1n04x5 FILLER_37_2199 ();
 b15zdnd11an1n64x5 FILLER_37_2215 ();
 b15zdnd11an1n04x5 FILLER_37_2279 ();
 b15zdnd00an1n01x5 FILLER_37_2283 ();
 b15zdnd11an1n16x5 FILLER_38_8 ();
 b15zdnd11an1n08x5 FILLER_38_24 ();
 b15zdnd11an1n04x5 FILLER_38_48 ();
 b15zdnd11an1n08x5 FILLER_38_56 ();
 b15zdnd00an1n02x5 FILLER_38_64 ();
 b15zdnd00an1n01x5 FILLER_38_66 ();
 b15zdnd11an1n64x5 FILLER_38_73 ();
 b15zdnd11an1n16x5 FILLER_38_137 ();
 b15zdnd00an1n02x5 FILLER_38_153 ();
 b15zdnd11an1n08x5 FILLER_38_159 ();
 b15zdnd00an1n01x5 FILLER_38_167 ();
 b15zdnd11an1n08x5 FILLER_38_175 ();
 b15zdnd11an1n04x5 FILLER_38_183 ();
 b15zdnd00an1n02x5 FILLER_38_187 ();
 b15zdnd00an1n01x5 FILLER_38_189 ();
 b15zdnd11an1n64x5 FILLER_38_203 ();
 b15zdnd11an1n64x5 FILLER_38_267 ();
 b15zdnd00an1n01x5 FILLER_38_331 ();
 b15zdnd11an1n04x5 FILLER_38_343 ();
 b15zdnd11an1n04x5 FILLER_38_352 ();
 b15zdnd00an1n01x5 FILLER_38_356 ();
 b15zdnd11an1n64x5 FILLER_38_366 ();
 b15zdnd11an1n16x5 FILLER_38_430 ();
 b15zdnd11an1n04x5 FILLER_38_446 ();
 b15zdnd00an1n02x5 FILLER_38_450 ();
 b15zdnd11an1n16x5 FILLER_38_458 ();
 b15zdnd11an1n08x5 FILLER_38_474 ();
 b15zdnd11an1n32x5 FILLER_38_486 ();
 b15zdnd11an1n64x5 FILLER_38_532 ();
 b15zdnd11an1n04x5 FILLER_38_596 ();
 b15zdnd00an1n02x5 FILLER_38_600 ();
 b15zdnd11an1n64x5 FILLER_38_606 ();
 b15zdnd11an1n16x5 FILLER_38_670 ();
 b15zdnd11an1n08x5 FILLER_38_686 ();
 b15zdnd00an1n02x5 FILLER_38_694 ();
 b15zdnd00an1n01x5 FILLER_38_696 ();
 b15zdnd11an1n08x5 FILLER_38_707 ();
 b15zdnd00an1n02x5 FILLER_38_715 ();
 b15zdnd00an1n01x5 FILLER_38_717 ();
 b15zdnd11an1n64x5 FILLER_38_726 ();
 b15zdnd11an1n04x5 FILLER_38_790 ();
 b15zdnd00an1n02x5 FILLER_38_794 ();
 b15zdnd00an1n01x5 FILLER_38_796 ();
 b15zdnd11an1n32x5 FILLER_38_801 ();
 b15zdnd11an1n08x5 FILLER_38_833 ();
 b15zdnd00an1n01x5 FILLER_38_841 ();
 b15zdnd11an1n64x5 FILLER_38_854 ();
 b15zdnd00an1n02x5 FILLER_38_918 ();
 b15zdnd11an1n64x5 FILLER_38_941 ();
 b15zdnd11an1n32x5 FILLER_38_1005 ();
 b15zdnd11an1n16x5 FILLER_38_1037 ();
 b15zdnd00an1n02x5 FILLER_38_1053 ();
 b15zdnd00an1n01x5 FILLER_38_1055 ();
 b15zdnd11an1n64x5 FILLER_38_1066 ();
 b15zdnd11an1n16x5 FILLER_38_1130 ();
 b15zdnd11an1n04x5 FILLER_38_1146 ();
 b15zdnd11an1n32x5 FILLER_38_1154 ();
 b15zdnd11an1n16x5 FILLER_38_1186 ();
 b15zdnd11an1n08x5 FILLER_38_1202 ();
 b15zdnd11an1n04x5 FILLER_38_1210 ();
 b15zdnd00an1n02x5 FILLER_38_1214 ();
 b15zdnd00an1n01x5 FILLER_38_1216 ();
 b15zdnd11an1n32x5 FILLER_38_1237 ();
 b15zdnd11an1n16x5 FILLER_38_1269 ();
 b15zdnd11an1n04x5 FILLER_38_1285 ();
 b15zdnd00an1n02x5 FILLER_38_1289 ();
 b15zdnd00an1n01x5 FILLER_38_1291 ();
 b15zdnd11an1n16x5 FILLER_38_1297 ();
 b15zdnd11an1n04x5 FILLER_38_1313 ();
 b15zdnd00an1n02x5 FILLER_38_1317 ();
 b15zdnd00an1n01x5 FILLER_38_1319 ();
 b15zdnd11an1n16x5 FILLER_38_1325 ();
 b15zdnd00an1n02x5 FILLER_38_1341 ();
 b15zdnd11an1n64x5 FILLER_38_1358 ();
 b15zdnd11an1n16x5 FILLER_38_1422 ();
 b15zdnd11an1n08x5 FILLER_38_1438 ();
 b15zdnd11an1n04x5 FILLER_38_1446 ();
 b15zdnd00an1n02x5 FILLER_38_1450 ();
 b15zdnd00an1n01x5 FILLER_38_1452 ();
 b15zdnd11an1n64x5 FILLER_38_1458 ();
 b15zdnd11an1n32x5 FILLER_38_1522 ();
 b15zdnd11an1n16x5 FILLER_38_1554 ();
 b15zdnd11an1n08x5 FILLER_38_1570 ();
 b15zdnd00an1n02x5 FILLER_38_1578 ();
 b15zdnd00an1n01x5 FILLER_38_1580 ();
 b15zdnd11an1n04x5 FILLER_38_1586 ();
 b15zdnd00an1n02x5 FILLER_38_1590 ();
 b15zdnd11an1n08x5 FILLER_38_1599 ();
 b15zdnd00an1n01x5 FILLER_38_1607 ();
 b15zdnd11an1n04x5 FILLER_38_1617 ();
 b15zdnd00an1n02x5 FILLER_38_1621 ();
 b15zdnd11an1n04x5 FILLER_38_1636 ();
 b15zdnd00an1n02x5 FILLER_38_1640 ();
 b15zdnd11an1n16x5 FILLER_38_1653 ();
 b15zdnd11an1n04x5 FILLER_38_1669 ();
 b15zdnd00an1n02x5 FILLER_38_1673 ();
 b15zdnd11an1n64x5 FILLER_38_1681 ();
 b15zdnd11an1n16x5 FILLER_38_1745 ();
 b15zdnd00an1n01x5 FILLER_38_1761 ();
 b15zdnd11an1n16x5 FILLER_38_1771 ();
 b15zdnd11an1n04x5 FILLER_38_1787 ();
 b15zdnd00an1n02x5 FILLER_38_1791 ();
 b15zdnd00an1n01x5 FILLER_38_1793 ();
 b15zdnd11an1n32x5 FILLER_38_1801 ();
 b15zdnd00an1n02x5 FILLER_38_1833 ();
 b15zdnd00an1n01x5 FILLER_38_1835 ();
 b15zdnd11an1n64x5 FILLER_38_1846 ();
 b15zdnd11an1n64x5 FILLER_38_1910 ();
 b15zdnd11an1n64x5 FILLER_38_1974 ();
 b15zdnd11an1n08x5 FILLER_38_2038 ();
 b15zdnd11an1n04x5 FILLER_38_2046 ();
 b15zdnd00an1n01x5 FILLER_38_2050 ();
 b15zdnd11an1n64x5 FILLER_38_2059 ();
 b15zdnd11an1n08x5 FILLER_38_2123 ();
 b15zdnd00an1n01x5 FILLER_38_2131 ();
 b15zdnd11an1n08x5 FILLER_38_2142 ();
 b15zdnd11an1n04x5 FILLER_38_2150 ();
 b15zdnd11an1n04x5 FILLER_38_2162 ();
 b15zdnd00an1n01x5 FILLER_38_2166 ();
 b15zdnd11an1n04x5 FILLER_38_2175 ();
 b15zdnd11an1n64x5 FILLER_38_2190 ();
 b15zdnd11an1n16x5 FILLER_38_2254 ();
 b15zdnd11an1n04x5 FILLER_38_2270 ();
 b15zdnd00an1n02x5 FILLER_38_2274 ();
 b15zdnd11an1n32x5 FILLER_39_0 ();
 b15zdnd11an1n08x5 FILLER_39_32 ();
 b15zdnd00an1n02x5 FILLER_39_40 ();
 b15zdnd11an1n16x5 FILLER_39_49 ();
 b15zdnd11an1n04x5 FILLER_39_65 ();
 b15zdnd00an1n01x5 FILLER_39_69 ();
 b15zdnd11an1n08x5 FILLER_39_84 ();
 b15zdnd00an1n01x5 FILLER_39_92 ();
 b15zdnd11an1n04x5 FILLER_39_98 ();
 b15zdnd00an1n02x5 FILLER_39_102 ();
 b15zdnd00an1n01x5 FILLER_39_104 ();
 b15zdnd11an1n08x5 FILLER_39_110 ();
 b15zdnd11an1n04x5 FILLER_39_118 ();
 b15zdnd00an1n01x5 FILLER_39_122 ();
 b15zdnd11an1n16x5 FILLER_39_134 ();
 b15zdnd00an1n01x5 FILLER_39_150 ();
 b15zdnd11an1n04x5 FILLER_39_163 ();
 b15zdnd11an1n04x5 FILLER_39_171 ();
 b15zdnd00an1n01x5 FILLER_39_175 ();
 b15zdnd11an1n04x5 FILLER_39_189 ();
 b15zdnd11an1n08x5 FILLER_39_213 ();
 b15zdnd00an1n02x5 FILLER_39_221 ();
 b15zdnd00an1n01x5 FILLER_39_223 ();
 b15zdnd11an1n08x5 FILLER_39_228 ();
 b15zdnd11an1n04x5 FILLER_39_236 ();
 b15zdnd11an1n32x5 FILLER_39_250 ();
 b15zdnd11an1n16x5 FILLER_39_282 ();
 b15zdnd00an1n01x5 FILLER_39_298 ();
 b15zdnd11an1n32x5 FILLER_39_307 ();
 b15zdnd11an1n04x5 FILLER_39_339 ();
 b15zdnd11an1n64x5 FILLER_39_350 ();
 b15zdnd11an1n16x5 FILLER_39_414 ();
 b15zdnd11an1n04x5 FILLER_39_430 ();
 b15zdnd11an1n16x5 FILLER_39_446 ();
 b15zdnd11an1n04x5 FILLER_39_462 ();
 b15zdnd00an1n01x5 FILLER_39_466 ();
 b15zdnd11an1n04x5 FILLER_39_483 ();
 b15zdnd11an1n16x5 FILLER_39_499 ();
 b15zdnd11an1n04x5 FILLER_39_515 ();
 b15zdnd00an1n01x5 FILLER_39_519 ();
 b15zdnd11an1n32x5 FILLER_39_533 ();
 b15zdnd11an1n16x5 FILLER_39_565 ();
 b15zdnd11an1n08x5 FILLER_39_581 ();
 b15zdnd00an1n02x5 FILLER_39_589 ();
 b15zdnd11an1n64x5 FILLER_39_603 ();
 b15zdnd11an1n08x5 FILLER_39_667 ();
 b15zdnd00an1n02x5 FILLER_39_675 ();
 b15zdnd00an1n01x5 FILLER_39_677 ();
 b15zdnd11an1n16x5 FILLER_39_685 ();
 b15zdnd11an1n08x5 FILLER_39_701 ();
 b15zdnd11an1n04x5 FILLER_39_709 ();
 b15zdnd11an1n32x5 FILLER_39_731 ();
 b15zdnd00an1n02x5 FILLER_39_763 ();
 b15zdnd11an1n16x5 FILLER_39_771 ();
 b15zdnd11an1n64x5 FILLER_39_796 ();
 b15zdnd11an1n64x5 FILLER_39_860 ();
 b15zdnd11an1n32x5 FILLER_39_924 ();
 b15zdnd11an1n16x5 FILLER_39_956 ();
 b15zdnd00an1n02x5 FILLER_39_972 ();
 b15zdnd11an1n04x5 FILLER_39_983 ();
 b15zdnd00an1n02x5 FILLER_39_987 ();
 b15zdnd11an1n16x5 FILLER_39_999 ();
 b15zdnd11an1n08x5 FILLER_39_1015 ();
 b15zdnd11an1n04x5 FILLER_39_1023 ();
 b15zdnd00an1n02x5 FILLER_39_1027 ();
 b15zdnd11an1n08x5 FILLER_39_1041 ();
 b15zdnd00an1n02x5 FILLER_39_1049 ();
 b15zdnd11an1n04x5 FILLER_39_1069 ();
 b15zdnd11an1n64x5 FILLER_39_1084 ();
 b15zdnd11an1n04x5 FILLER_39_1148 ();
 b15zdnd11an1n08x5 FILLER_39_1173 ();
 b15zdnd00an1n02x5 FILLER_39_1181 ();
 b15zdnd00an1n01x5 FILLER_39_1183 ();
 b15zdnd11an1n32x5 FILLER_39_1212 ();
 b15zdnd11an1n16x5 FILLER_39_1244 ();
 b15zdnd11an1n04x5 FILLER_39_1260 ();
 b15zdnd11an1n08x5 FILLER_39_1290 ();
 b15zdnd11an1n64x5 FILLER_39_1307 ();
 b15zdnd11an1n64x5 FILLER_39_1377 ();
 b15zdnd11an1n64x5 FILLER_39_1441 ();
 b15zdnd11an1n64x5 FILLER_39_1505 ();
 b15zdnd11an1n04x5 FILLER_39_1569 ();
 b15zdnd00an1n02x5 FILLER_39_1573 ();
 b15zdnd00an1n01x5 FILLER_39_1575 ();
 b15zdnd11an1n64x5 FILLER_39_1585 ();
 b15zdnd11an1n64x5 FILLER_39_1649 ();
 b15zdnd11an1n64x5 FILLER_39_1713 ();
 b15zdnd00an1n02x5 FILLER_39_1777 ();
 b15zdnd11an1n32x5 FILLER_39_1788 ();
 b15zdnd00an1n01x5 FILLER_39_1820 ();
 b15zdnd11an1n16x5 FILLER_39_1825 ();
 b15zdnd11an1n04x5 FILLER_39_1846 ();
 b15zdnd11an1n04x5 FILLER_39_1860 ();
 b15zdnd11an1n04x5 FILLER_39_1876 ();
 b15zdnd11an1n08x5 FILLER_39_1889 ();
 b15zdnd00an1n01x5 FILLER_39_1897 ();
 b15zdnd11an1n64x5 FILLER_39_1906 ();
 b15zdnd11an1n32x5 FILLER_39_1970 ();
 b15zdnd11an1n08x5 FILLER_39_2012 ();
 b15zdnd00an1n02x5 FILLER_39_2020 ();
 b15zdnd00an1n01x5 FILLER_39_2022 ();
 b15zdnd11an1n16x5 FILLER_39_2028 ();
 b15zdnd11an1n08x5 FILLER_39_2044 ();
 b15zdnd00an1n02x5 FILLER_39_2052 ();
 b15zdnd11an1n04x5 FILLER_39_2061 ();
 b15zdnd11an1n04x5 FILLER_39_2081 ();
 b15zdnd11an1n32x5 FILLER_39_2099 ();
 b15zdnd11an1n08x5 FILLER_39_2131 ();
 b15zdnd11an1n32x5 FILLER_39_2145 ();
 b15zdnd11an1n08x5 FILLER_39_2177 ();
 b15zdnd00an1n02x5 FILLER_39_2185 ();
 b15zdnd11an1n64x5 FILLER_39_2193 ();
 b15zdnd11an1n16x5 FILLER_39_2257 ();
 b15zdnd11an1n08x5 FILLER_39_2273 ();
 b15zdnd00an1n02x5 FILLER_39_2281 ();
 b15zdnd00an1n01x5 FILLER_39_2283 ();
 b15zdnd11an1n32x5 FILLER_40_8 ();
 b15zdnd00an1n02x5 FILLER_40_40 ();
 b15zdnd11an1n32x5 FILLER_40_46 ();
 b15zdnd11an1n04x5 FILLER_40_78 ();
 b15zdnd00an1n02x5 FILLER_40_82 ();
 b15zdnd00an1n01x5 FILLER_40_84 ();
 b15zdnd11an1n04x5 FILLER_40_96 ();
 b15zdnd11an1n04x5 FILLER_40_112 ();
 b15zdnd11an1n04x5 FILLER_40_137 ();
 b15zdnd11an1n32x5 FILLER_40_151 ();
 b15zdnd11an1n16x5 FILLER_40_183 ();
 b15zdnd11an1n04x5 FILLER_40_199 ();
 b15zdnd11an1n04x5 FILLER_40_213 ();
 b15zdnd11an1n16x5 FILLER_40_227 ();
 b15zdnd11an1n08x5 FILLER_40_243 ();
 b15zdnd11an1n04x5 FILLER_40_251 ();
 b15zdnd00an1n02x5 FILLER_40_255 ();
 b15zdnd00an1n01x5 FILLER_40_257 ();
 b15zdnd11an1n04x5 FILLER_40_270 ();
 b15zdnd11an1n04x5 FILLER_40_280 ();
 b15zdnd00an1n02x5 FILLER_40_284 ();
 b15zdnd11an1n04x5 FILLER_40_290 ();
 b15zdnd11an1n04x5 FILLER_40_301 ();
 b15zdnd11an1n16x5 FILLER_40_309 ();
 b15zdnd11an1n08x5 FILLER_40_325 ();
 b15zdnd11an1n04x5 FILLER_40_333 ();
 b15zdnd11an1n64x5 FILLER_40_343 ();
 b15zdnd11an1n08x5 FILLER_40_407 ();
 b15zdnd11an1n04x5 FILLER_40_415 ();
 b15zdnd00an1n02x5 FILLER_40_419 ();
 b15zdnd00an1n01x5 FILLER_40_421 ();
 b15zdnd11an1n08x5 FILLER_40_429 ();
 b15zdnd11an1n04x5 FILLER_40_437 ();
 b15zdnd00an1n01x5 FILLER_40_441 ();
 b15zdnd11an1n32x5 FILLER_40_457 ();
 b15zdnd00an1n01x5 FILLER_40_489 ();
 b15zdnd11an1n16x5 FILLER_40_506 ();
 b15zdnd11an1n08x5 FILLER_40_522 ();
 b15zdnd11an1n04x5 FILLER_40_530 ();
 b15zdnd00an1n01x5 FILLER_40_534 ();
 b15zdnd11an1n04x5 FILLER_40_547 ();
 b15zdnd11an1n32x5 FILLER_40_557 ();
 b15zdnd11an1n16x5 FILLER_40_589 ();
 b15zdnd11an1n08x5 FILLER_40_605 ();
 b15zdnd11an1n04x5 FILLER_40_613 ();
 b15zdnd00an1n02x5 FILLER_40_617 ();
 b15zdnd00an1n01x5 FILLER_40_619 ();
 b15zdnd11an1n08x5 FILLER_40_625 ();
 b15zdnd11an1n04x5 FILLER_40_633 ();
 b15zdnd00an1n01x5 FILLER_40_637 ();
 b15zdnd11an1n08x5 FILLER_40_651 ();
 b15zdnd11an1n04x5 FILLER_40_659 ();
 b15zdnd00an1n02x5 FILLER_40_663 ();
 b15zdnd00an1n01x5 FILLER_40_665 ();
 b15zdnd11an1n32x5 FILLER_40_680 ();
 b15zdnd11an1n04x5 FILLER_40_712 ();
 b15zdnd00an1n02x5 FILLER_40_716 ();
 b15zdnd11an1n04x5 FILLER_40_726 ();
 b15zdnd11an1n16x5 FILLER_40_737 ();
 b15zdnd00an1n01x5 FILLER_40_753 ();
 b15zdnd11an1n04x5 FILLER_40_758 ();
 b15zdnd11an1n16x5 FILLER_40_768 ();
 b15zdnd11an1n04x5 FILLER_40_784 ();
 b15zdnd00an1n02x5 FILLER_40_788 ();
 b15zdnd00an1n01x5 FILLER_40_790 ();
 b15zdnd11an1n32x5 FILLER_40_796 ();
 b15zdnd11an1n16x5 FILLER_40_828 ();
 b15zdnd11an1n32x5 FILLER_40_870 ();
 b15zdnd00an1n01x5 FILLER_40_902 ();
 b15zdnd11an1n16x5 FILLER_40_929 ();
 b15zdnd11an1n08x5 FILLER_40_945 ();
 b15zdnd11an1n08x5 FILLER_40_965 ();
 b15zdnd00an1n02x5 FILLER_40_973 ();
 b15zdnd11an1n64x5 FILLER_40_984 ();
 b15zdnd11an1n32x5 FILLER_40_1048 ();
 b15zdnd11an1n08x5 FILLER_40_1080 ();
 b15zdnd11an1n64x5 FILLER_40_1098 ();
 b15zdnd11an1n32x5 FILLER_40_1162 ();
 b15zdnd11an1n08x5 FILLER_40_1194 ();
 b15zdnd11an1n32x5 FILLER_40_1233 ();
 b15zdnd11an1n08x5 FILLER_40_1265 ();
 b15zdnd11an1n04x5 FILLER_40_1273 ();
 b15zdnd00an1n02x5 FILLER_40_1277 ();
 b15zdnd11an1n16x5 FILLER_40_1293 ();
 b15zdnd11an1n08x5 FILLER_40_1309 ();
 b15zdnd11an1n04x5 FILLER_40_1317 ();
 b15zdnd11an1n04x5 FILLER_40_1328 ();
 b15zdnd11an1n04x5 FILLER_40_1346 ();
 b15zdnd11an1n08x5 FILLER_40_1357 ();
 b15zdnd11an1n04x5 FILLER_40_1365 ();
 b15zdnd00an1n02x5 FILLER_40_1369 ();
 b15zdnd00an1n01x5 FILLER_40_1371 ();
 b15zdnd11an1n04x5 FILLER_40_1376 ();
 b15zdnd11an1n32x5 FILLER_40_1385 ();
 b15zdnd11an1n16x5 FILLER_40_1417 ();
 b15zdnd11an1n04x5 FILLER_40_1447 ();
 b15zdnd11an1n16x5 FILLER_40_1456 ();
 b15zdnd00an1n01x5 FILLER_40_1472 ();
 b15zdnd11an1n64x5 FILLER_40_1478 ();
 b15zdnd11an1n04x5 FILLER_40_1542 ();
 b15zdnd00an1n02x5 FILLER_40_1546 ();
 b15zdnd11an1n64x5 FILLER_40_1555 ();
 b15zdnd11an1n32x5 FILLER_40_1619 ();
 b15zdnd11an1n08x5 FILLER_40_1651 ();
 b15zdnd00an1n02x5 FILLER_40_1659 ();
 b15zdnd00an1n01x5 FILLER_40_1661 ();
 b15zdnd11an1n04x5 FILLER_40_1674 ();
 b15zdnd11an1n64x5 FILLER_40_1698 ();
 b15zdnd11an1n08x5 FILLER_40_1762 ();
 b15zdnd11an1n04x5 FILLER_40_1790 ();
 b15zdnd11an1n16x5 FILLER_40_1802 ();
 b15zdnd11an1n32x5 FILLER_40_1830 ();
 b15zdnd11an1n16x5 FILLER_40_1862 ();
 b15zdnd11an1n08x5 FILLER_40_1878 ();
 b15zdnd11an1n08x5 FILLER_40_1892 ();
 b15zdnd11an1n16x5 FILLER_40_1906 ();
 b15zdnd00an1n01x5 FILLER_40_1922 ();
 b15zdnd11an1n08x5 FILLER_40_1930 ();
 b15zdnd00an1n01x5 FILLER_40_1938 ();
 b15zdnd11an1n08x5 FILLER_40_1947 ();
 b15zdnd11an1n04x5 FILLER_40_1955 ();
 b15zdnd00an1n02x5 FILLER_40_1959 ();
 b15zdnd11an1n32x5 FILLER_40_1966 ();
 b15zdnd11an1n04x5 FILLER_40_1998 ();
 b15zdnd00an1n01x5 FILLER_40_2002 ();
 b15zdnd11an1n08x5 FILLER_40_2010 ();
 b15zdnd11an1n04x5 FILLER_40_2018 ();
 b15zdnd11an1n16x5 FILLER_40_2029 ();
 b15zdnd11an1n08x5 FILLER_40_2045 ();
 b15zdnd00an1n01x5 FILLER_40_2053 ();
 b15zdnd11an1n32x5 FILLER_40_2066 ();
 b15zdnd11an1n08x5 FILLER_40_2098 ();
 b15zdnd11an1n04x5 FILLER_40_2106 ();
 b15zdnd00an1n02x5 FILLER_40_2110 ();
 b15zdnd11an1n04x5 FILLER_40_2121 ();
 b15zdnd00an1n01x5 FILLER_40_2125 ();
 b15zdnd11an1n08x5 FILLER_40_2130 ();
 b15zdnd11an1n04x5 FILLER_40_2138 ();
 b15zdnd00an1n01x5 FILLER_40_2142 ();
 b15zdnd11an1n04x5 FILLER_40_2148 ();
 b15zdnd00an1n02x5 FILLER_40_2152 ();
 b15zdnd11an1n16x5 FILLER_40_2162 ();
 b15zdnd11an1n08x5 FILLER_40_2178 ();
 b15zdnd11an1n04x5 FILLER_40_2186 ();
 b15zdnd00an1n02x5 FILLER_40_2190 ();
 b15zdnd00an1n01x5 FILLER_40_2192 ();
 b15zdnd11an1n64x5 FILLER_40_2197 ();
 b15zdnd11an1n08x5 FILLER_40_2261 ();
 b15zdnd11an1n04x5 FILLER_40_2269 ();
 b15zdnd00an1n02x5 FILLER_40_2273 ();
 b15zdnd00an1n01x5 FILLER_40_2275 ();
 b15zdnd11an1n32x5 FILLER_41_0 ();
 b15zdnd11an1n16x5 FILLER_41_32 ();
 b15zdnd11an1n64x5 FILLER_41_53 ();
 b15zdnd11an1n64x5 FILLER_41_117 ();
 b15zdnd11an1n32x5 FILLER_41_181 ();
 b15zdnd11an1n16x5 FILLER_41_213 ();
 b15zdnd11an1n04x5 FILLER_41_229 ();
 b15zdnd11an1n04x5 FILLER_41_239 ();
 b15zdnd00an1n02x5 FILLER_41_243 ();
 b15zdnd11an1n64x5 FILLER_41_252 ();
 b15zdnd11an1n08x5 FILLER_41_316 ();
 b15zdnd00an1n02x5 FILLER_41_324 ();
 b15zdnd00an1n01x5 FILLER_41_326 ();
 b15zdnd11an1n04x5 FILLER_41_331 ();
 b15zdnd11an1n64x5 FILLER_41_351 ();
 b15zdnd11an1n04x5 FILLER_41_415 ();
 b15zdnd00an1n02x5 FILLER_41_419 ();
 b15zdnd11an1n16x5 FILLER_41_430 ();
 b15zdnd00an1n01x5 FILLER_41_446 ();
 b15zdnd11an1n16x5 FILLER_41_451 ();
 b15zdnd11an1n08x5 FILLER_41_467 ();
 b15zdnd00an1n02x5 FILLER_41_475 ();
 b15zdnd00an1n01x5 FILLER_41_477 ();
 b15zdnd11an1n08x5 FILLER_41_487 ();
 b15zdnd00an1n02x5 FILLER_41_495 ();
 b15zdnd00an1n01x5 FILLER_41_497 ();
 b15zdnd11an1n16x5 FILLER_41_503 ();
 b15zdnd11an1n08x5 FILLER_41_519 ();
 b15zdnd00an1n01x5 FILLER_41_527 ();
 b15zdnd11an1n04x5 FILLER_41_543 ();
 b15zdnd11an1n08x5 FILLER_41_554 ();
 b15zdnd11an1n04x5 FILLER_41_562 ();
 b15zdnd00an1n02x5 FILLER_41_566 ();
 b15zdnd11an1n32x5 FILLER_41_580 ();
 b15zdnd11an1n04x5 FILLER_41_612 ();
 b15zdnd00an1n01x5 FILLER_41_616 ();
 b15zdnd11an1n64x5 FILLER_41_630 ();
 b15zdnd11an1n04x5 FILLER_41_694 ();
 b15zdnd00an1n02x5 FILLER_41_698 ();
 b15zdnd11an1n08x5 FILLER_41_709 ();
 b15zdnd00an1n02x5 FILLER_41_717 ();
 b15zdnd00an1n01x5 FILLER_41_719 ();
 b15zdnd11an1n32x5 FILLER_41_730 ();
 b15zdnd11an1n04x5 FILLER_41_762 ();
 b15zdnd11an1n16x5 FILLER_41_775 ();
 b15zdnd11an1n08x5 FILLER_41_791 ();
 b15zdnd00an1n02x5 FILLER_41_799 ();
 b15zdnd11an1n04x5 FILLER_41_807 ();
 b15zdnd11an1n08x5 FILLER_41_827 ();
 b15zdnd11an1n04x5 FILLER_41_844 ();
 b15zdnd11an1n16x5 FILLER_41_854 ();
 b15zdnd11an1n04x5 FILLER_41_882 ();
 b15zdnd11an1n04x5 FILLER_41_896 ();
 b15zdnd11an1n64x5 FILLER_41_932 ();
 b15zdnd11an1n64x5 FILLER_41_996 ();
 b15zdnd11an1n32x5 FILLER_41_1060 ();
 b15zdnd00an1n01x5 FILLER_41_1092 ();
 b15zdnd11an1n04x5 FILLER_41_1103 ();
 b15zdnd00an1n02x5 FILLER_41_1107 ();
 b15zdnd00an1n01x5 FILLER_41_1109 ();
 b15zdnd11an1n16x5 FILLER_41_1129 ();
 b15zdnd11an1n08x5 FILLER_41_1145 ();
 b15zdnd00an1n02x5 FILLER_41_1153 ();
 b15zdnd11an1n16x5 FILLER_41_1175 ();
 b15zdnd11an1n32x5 FILLER_41_1231 ();
 b15zdnd11an1n16x5 FILLER_41_1263 ();
 b15zdnd11an1n08x5 FILLER_41_1279 ();
 b15zdnd00an1n01x5 FILLER_41_1287 ();
 b15zdnd11an1n04x5 FILLER_41_1292 ();
 b15zdnd00an1n01x5 FILLER_41_1296 ();
 b15zdnd11an1n08x5 FILLER_41_1301 ();
 b15zdnd11an1n04x5 FILLER_41_1309 ();
 b15zdnd00an1n02x5 FILLER_41_1313 ();
 b15zdnd00an1n01x5 FILLER_41_1315 ();
 b15zdnd11an1n32x5 FILLER_41_1322 ();
 b15zdnd11an1n16x5 FILLER_41_1354 ();
 b15zdnd11an1n04x5 FILLER_41_1370 ();
 b15zdnd00an1n02x5 FILLER_41_1374 ();
 b15zdnd00an1n01x5 FILLER_41_1376 ();
 b15zdnd11an1n32x5 FILLER_41_1386 ();
 b15zdnd11an1n16x5 FILLER_41_1418 ();
 b15zdnd11an1n04x5 FILLER_41_1434 ();
 b15zdnd11an1n08x5 FILLER_41_1444 ();
 b15zdnd00an1n01x5 FILLER_41_1452 ();
 b15zdnd11an1n04x5 FILLER_41_1460 ();
 b15zdnd11an1n04x5 FILLER_41_1469 ();
 b15zdnd11an1n32x5 FILLER_41_1480 ();
 b15zdnd11an1n08x5 FILLER_41_1512 ();
 b15zdnd11an1n08x5 FILLER_41_1535 ();
 b15zdnd00an1n02x5 FILLER_41_1543 ();
 b15zdnd00an1n01x5 FILLER_41_1545 ();
 b15zdnd11an1n64x5 FILLER_41_1559 ();
 b15zdnd11an1n32x5 FILLER_41_1623 ();
 b15zdnd00an1n01x5 FILLER_41_1655 ();
 b15zdnd11an1n04x5 FILLER_41_1662 ();
 b15zdnd11an1n64x5 FILLER_41_1675 ();
 b15zdnd11an1n32x5 FILLER_41_1739 ();
 b15zdnd11an1n16x5 FILLER_41_1771 ();
 b15zdnd11an1n08x5 FILLER_41_1787 ();
 b15zdnd11an1n04x5 FILLER_41_1795 ();
 b15zdnd11an1n32x5 FILLER_41_1819 ();
 b15zdnd11an1n16x5 FILLER_41_1851 ();
 b15zdnd11an1n04x5 FILLER_41_1867 ();
 b15zdnd00an1n02x5 FILLER_41_1871 ();
 b15zdnd00an1n01x5 FILLER_41_1873 ();
 b15zdnd11an1n16x5 FILLER_41_1884 ();
 b15zdnd00an1n02x5 FILLER_41_1900 ();
 b15zdnd11an1n16x5 FILLER_41_1908 ();
 b15zdnd11an1n04x5 FILLER_41_1924 ();
 b15zdnd00an1n01x5 FILLER_41_1928 ();
 b15zdnd11an1n04x5 FILLER_41_1934 ();
 b15zdnd11an1n16x5 FILLER_41_1942 ();
 b15zdnd00an1n02x5 FILLER_41_1958 ();
 b15zdnd00an1n01x5 FILLER_41_1960 ();
 b15zdnd11an1n04x5 FILLER_41_1967 ();
 b15zdnd00an1n01x5 FILLER_41_1971 ();
 b15zdnd11an1n04x5 FILLER_41_1979 ();
 b15zdnd11an1n08x5 FILLER_41_1987 ();
 b15zdnd11an1n32x5 FILLER_41_2002 ();
 b15zdnd11an1n16x5 FILLER_41_2034 ();
 b15zdnd11an1n08x5 FILLER_41_2050 ();
 b15zdnd11an1n32x5 FILLER_41_2063 ();
 b15zdnd11an1n16x5 FILLER_41_2095 ();
 b15zdnd11an1n08x5 FILLER_41_2111 ();
 b15zdnd11an1n04x5 FILLER_41_2119 ();
 b15zdnd11an1n32x5 FILLER_41_2138 ();
 b15zdnd11an1n16x5 FILLER_41_2170 ();
 b15zdnd11an1n08x5 FILLER_41_2186 ();
 b15zdnd00an1n02x5 FILLER_41_2194 ();
 b15zdnd11an1n04x5 FILLER_41_2207 ();
 b15zdnd00an1n02x5 FILLER_41_2211 ();
 b15zdnd00an1n01x5 FILLER_41_2213 ();
 b15zdnd11an1n64x5 FILLER_41_2219 ();
 b15zdnd00an1n01x5 FILLER_41_2283 ();
 b15zdnd11an1n64x5 FILLER_42_8 ();
 b15zdnd11an1n16x5 FILLER_42_72 ();
 b15zdnd11an1n08x5 FILLER_42_88 ();
 b15zdnd11an1n04x5 FILLER_42_96 ();
 b15zdnd00an1n02x5 FILLER_42_100 ();
 b15zdnd11an1n64x5 FILLER_42_123 ();
 b15zdnd11an1n64x5 FILLER_42_187 ();
 b15zdnd11an1n16x5 FILLER_42_251 ();
 b15zdnd11an1n08x5 FILLER_42_267 ();
 b15zdnd11an1n04x5 FILLER_42_275 ();
 b15zdnd00an1n02x5 FILLER_42_279 ();
 b15zdnd00an1n01x5 FILLER_42_281 ();
 b15zdnd11an1n32x5 FILLER_42_291 ();
 b15zdnd00an1n02x5 FILLER_42_323 ();
 b15zdnd00an1n01x5 FILLER_42_325 ();
 b15zdnd11an1n08x5 FILLER_42_338 ();
 b15zdnd11an1n04x5 FILLER_42_346 ();
 b15zdnd00an1n01x5 FILLER_42_350 ();
 b15zdnd11an1n64x5 FILLER_42_361 ();
 b15zdnd11an1n32x5 FILLER_42_425 ();
 b15zdnd11an1n08x5 FILLER_42_457 ();
 b15zdnd11an1n04x5 FILLER_42_465 ();
 b15zdnd00an1n02x5 FILLER_42_469 ();
 b15zdnd00an1n01x5 FILLER_42_471 ();
 b15zdnd11an1n64x5 FILLER_42_491 ();
 b15zdnd11an1n64x5 FILLER_42_555 ();
 b15zdnd11an1n16x5 FILLER_42_619 ();
 b15zdnd11an1n08x5 FILLER_42_635 ();
 b15zdnd11an1n04x5 FILLER_42_643 ();
 b15zdnd00an1n01x5 FILLER_42_647 ();
 b15zdnd11an1n04x5 FILLER_42_657 ();
 b15zdnd00an1n02x5 FILLER_42_661 ();
 b15zdnd11an1n16x5 FILLER_42_668 ();
 b15zdnd11an1n08x5 FILLER_42_684 ();
 b15zdnd11an1n04x5 FILLER_42_692 ();
 b15zdnd00an1n02x5 FILLER_42_696 ();
 b15zdnd00an1n01x5 FILLER_42_698 ();
 b15zdnd11an1n08x5 FILLER_42_706 ();
 b15zdnd11an1n04x5 FILLER_42_714 ();
 b15zdnd11an1n64x5 FILLER_42_726 ();
 b15zdnd11an1n08x5 FILLER_42_790 ();
 b15zdnd11an1n04x5 FILLER_42_798 ();
 b15zdnd00an1n01x5 FILLER_42_802 ();
 b15zdnd11an1n64x5 FILLER_42_808 ();
 b15zdnd11an1n16x5 FILLER_42_872 ();
 b15zdnd00an1n02x5 FILLER_42_888 ();
 b15zdnd11an1n16x5 FILLER_42_894 ();
 b15zdnd00an1n02x5 FILLER_42_910 ();
 b15zdnd11an1n64x5 FILLER_42_938 ();
 b15zdnd11an1n64x5 FILLER_42_1002 ();
 b15zdnd11an1n16x5 FILLER_42_1066 ();
 b15zdnd11an1n04x5 FILLER_42_1082 ();
 b15zdnd11an1n16x5 FILLER_42_1095 ();
 b15zdnd11an1n04x5 FILLER_42_1111 ();
 b15zdnd00an1n02x5 FILLER_42_1115 ();
 b15zdnd11an1n04x5 FILLER_42_1148 ();
 b15zdnd11an1n64x5 FILLER_42_1157 ();
 b15zdnd11an1n64x5 FILLER_42_1221 ();
 b15zdnd11an1n32x5 FILLER_42_1285 ();
 b15zdnd11an1n04x5 FILLER_42_1317 ();
 b15zdnd00an1n02x5 FILLER_42_1321 ();
 b15zdnd00an1n01x5 FILLER_42_1323 ();
 b15zdnd11an1n04x5 FILLER_42_1336 ();
 b15zdnd11an1n04x5 FILLER_42_1349 ();
 b15zdnd11an1n16x5 FILLER_42_1360 ();
 b15zdnd00an1n01x5 FILLER_42_1376 ();
 b15zdnd11an1n64x5 FILLER_42_1381 ();
 b15zdnd11an1n08x5 FILLER_42_1445 ();
 b15zdnd11an1n32x5 FILLER_42_1459 ();
 b15zdnd11an1n16x5 FILLER_42_1491 ();
 b15zdnd11an1n08x5 FILLER_42_1507 ();
 b15zdnd11an1n04x5 FILLER_42_1515 ();
 b15zdnd00an1n02x5 FILLER_42_1519 ();
 b15zdnd11an1n16x5 FILLER_42_1525 ();
 b15zdnd11an1n08x5 FILLER_42_1541 ();
 b15zdnd11an1n04x5 FILLER_42_1549 ();
 b15zdnd11an1n04x5 FILLER_42_1559 ();
 b15zdnd00an1n02x5 FILLER_42_1563 ();
 b15zdnd11an1n16x5 FILLER_42_1584 ();
 b15zdnd11an1n08x5 FILLER_42_1600 ();
 b15zdnd00an1n02x5 FILLER_42_1608 ();
 b15zdnd11an1n04x5 FILLER_42_1618 ();
 b15zdnd11an1n64x5 FILLER_42_1631 ();
 b15zdnd11an1n08x5 FILLER_42_1695 ();
 b15zdnd00an1n02x5 FILLER_42_1703 ();
 b15zdnd00an1n01x5 FILLER_42_1705 ();
 b15zdnd11an1n64x5 FILLER_42_1732 ();
 b15zdnd11an1n04x5 FILLER_42_1796 ();
 b15zdnd00an1n02x5 FILLER_42_1800 ();
 b15zdnd00an1n01x5 FILLER_42_1802 ();
 b15zdnd11an1n16x5 FILLER_42_1817 ();
 b15zdnd11an1n08x5 FILLER_42_1833 ();
 b15zdnd00an1n02x5 FILLER_42_1841 ();
 b15zdnd00an1n01x5 FILLER_42_1843 ();
 b15zdnd11an1n16x5 FILLER_42_1858 ();
 b15zdnd11an1n04x5 FILLER_42_1874 ();
 b15zdnd11an1n32x5 FILLER_42_1883 ();
 b15zdnd00an1n01x5 FILLER_42_1915 ();
 b15zdnd11an1n64x5 FILLER_42_1936 ();
 b15zdnd11an1n32x5 FILLER_42_2000 ();
 b15zdnd11an1n16x5 FILLER_42_2032 ();
 b15zdnd00an1n02x5 FILLER_42_2048 ();
 b15zdnd00an1n01x5 FILLER_42_2050 ();
 b15zdnd11an1n32x5 FILLER_42_2064 ();
 b15zdnd11an1n16x5 FILLER_42_2096 ();
 b15zdnd11an1n04x5 FILLER_42_2112 ();
 b15zdnd11an1n16x5 FILLER_42_2132 ();
 b15zdnd11an1n04x5 FILLER_42_2148 ();
 b15zdnd00an1n02x5 FILLER_42_2152 ();
 b15zdnd11an1n32x5 FILLER_42_2162 ();
 b15zdnd00an1n01x5 FILLER_42_2194 ();
 b15zdnd11an1n64x5 FILLER_42_2212 ();
 b15zdnd11an1n32x5 FILLER_43_0 ();
 b15zdnd11an1n16x5 FILLER_43_32 ();
 b15zdnd11an1n08x5 FILLER_43_48 ();
 b15zdnd00an1n02x5 FILLER_43_56 ();
 b15zdnd00an1n01x5 FILLER_43_58 ();
 b15zdnd11an1n16x5 FILLER_43_75 ();
 b15zdnd11an1n04x5 FILLER_43_91 ();
 b15zdnd00an1n01x5 FILLER_43_95 ();
 b15zdnd11an1n16x5 FILLER_43_108 ();
 b15zdnd11an1n08x5 FILLER_43_124 ();
 b15zdnd00an1n02x5 FILLER_43_132 ();
 b15zdnd11an1n64x5 FILLER_43_149 ();
 b15zdnd11an1n08x5 FILLER_43_213 ();
 b15zdnd11an1n04x5 FILLER_43_221 ();
 b15zdnd00an1n01x5 FILLER_43_225 ();
 b15zdnd11an1n32x5 FILLER_43_230 ();
 b15zdnd11an1n08x5 FILLER_43_262 ();
 b15zdnd11an1n04x5 FILLER_43_270 ();
 b15zdnd11an1n16x5 FILLER_43_280 ();
 b15zdnd11an1n08x5 FILLER_43_296 ();
 b15zdnd00an1n02x5 FILLER_43_304 ();
 b15zdnd00an1n01x5 FILLER_43_306 ();
 b15zdnd11an1n64x5 FILLER_43_312 ();
 b15zdnd11an1n32x5 FILLER_43_376 ();
 b15zdnd11an1n16x5 FILLER_43_408 ();
 b15zdnd11an1n08x5 FILLER_43_424 ();
 b15zdnd11an1n04x5 FILLER_43_432 ();
 b15zdnd00an1n02x5 FILLER_43_436 ();
 b15zdnd00an1n01x5 FILLER_43_438 ();
 b15zdnd11an1n32x5 FILLER_43_451 ();
 b15zdnd11an1n16x5 FILLER_43_483 ();
 b15zdnd11an1n04x5 FILLER_43_499 ();
 b15zdnd11an1n16x5 FILLER_43_507 ();
 b15zdnd11an1n08x5 FILLER_43_523 ();
 b15zdnd11an1n04x5 FILLER_43_531 ();
 b15zdnd00an1n01x5 FILLER_43_535 ();
 b15zdnd11an1n08x5 FILLER_43_544 ();
 b15zdnd11an1n04x5 FILLER_43_552 ();
 b15zdnd00an1n02x5 FILLER_43_556 ();
 b15zdnd00an1n01x5 FILLER_43_558 ();
 b15zdnd11an1n08x5 FILLER_43_563 ();
 b15zdnd11an1n16x5 FILLER_43_587 ();
 b15zdnd11an1n04x5 FILLER_43_603 ();
 b15zdnd00an1n02x5 FILLER_43_607 ();
 b15zdnd11an1n16x5 FILLER_43_623 ();
 b15zdnd11an1n04x5 FILLER_43_639 ();
 b15zdnd00an1n02x5 FILLER_43_643 ();
 b15zdnd11an1n08x5 FILLER_43_650 ();
 b15zdnd11an1n04x5 FILLER_43_658 ();
 b15zdnd00an1n02x5 FILLER_43_662 ();
 b15zdnd00an1n01x5 FILLER_43_664 ();
 b15zdnd11an1n16x5 FILLER_43_670 ();
 b15zdnd11an1n08x5 FILLER_43_686 ();
 b15zdnd11an1n04x5 FILLER_43_694 ();
 b15zdnd00an1n02x5 FILLER_43_698 ();
 b15zdnd11an1n04x5 FILLER_43_712 ();
 b15zdnd11an1n04x5 FILLER_43_736 ();
 b15zdnd00an1n02x5 FILLER_43_740 ();
 b15zdnd00an1n01x5 FILLER_43_742 ();
 b15zdnd11an1n32x5 FILLER_43_761 ();
 b15zdnd11an1n16x5 FILLER_43_793 ();
 b15zdnd11an1n08x5 FILLER_43_809 ();
 b15zdnd00an1n01x5 FILLER_43_817 ();
 b15zdnd11an1n64x5 FILLER_43_832 ();
 b15zdnd11an1n32x5 FILLER_43_896 ();
 b15zdnd11an1n16x5 FILLER_43_928 ();
 b15zdnd11an1n08x5 FILLER_43_944 ();
 b15zdnd00an1n02x5 FILLER_43_952 ();
 b15zdnd11an1n32x5 FILLER_43_963 ();
 b15zdnd11an1n16x5 FILLER_43_995 ();
 b15zdnd11an1n04x5 FILLER_43_1011 ();
 b15zdnd00an1n02x5 FILLER_43_1015 ();
 b15zdnd00an1n01x5 FILLER_43_1017 ();
 b15zdnd11an1n04x5 FILLER_43_1023 ();
 b15zdnd11an1n04x5 FILLER_43_1031 ();
 b15zdnd11an1n16x5 FILLER_43_1053 ();
 b15zdnd00an1n01x5 FILLER_43_1069 ();
 b15zdnd11an1n64x5 FILLER_43_1080 ();
 b15zdnd11an1n32x5 FILLER_43_1144 ();
 b15zdnd11an1n08x5 FILLER_43_1176 ();
 b15zdnd11an1n04x5 FILLER_43_1184 ();
 b15zdnd11an1n64x5 FILLER_43_1192 ();
 b15zdnd11an1n32x5 FILLER_43_1256 ();
 b15zdnd11an1n04x5 FILLER_43_1288 ();
 b15zdnd11an1n32x5 FILLER_43_1298 ();
 b15zdnd11an1n04x5 FILLER_43_1330 ();
 b15zdnd11an1n04x5 FILLER_43_1348 ();
 b15zdnd11an1n64x5 FILLER_43_1362 ();
 b15zdnd11an1n32x5 FILLER_43_1426 ();
 b15zdnd11an1n16x5 FILLER_43_1458 ();
 b15zdnd11an1n04x5 FILLER_43_1474 ();
 b15zdnd00an1n01x5 FILLER_43_1478 ();
 b15zdnd11an1n16x5 FILLER_43_1489 ();
 b15zdnd00an1n02x5 FILLER_43_1505 ();
 b15zdnd00an1n01x5 FILLER_43_1507 ();
 b15zdnd11an1n04x5 FILLER_43_1520 ();
 b15zdnd11an1n16x5 FILLER_43_1545 ();
 b15zdnd11an1n08x5 FILLER_43_1561 ();
 b15zdnd11an1n32x5 FILLER_43_1589 ();
 b15zdnd11an1n08x5 FILLER_43_1621 ();
 b15zdnd00an1n02x5 FILLER_43_1629 ();
 b15zdnd11an1n08x5 FILLER_43_1635 ();
 b15zdnd11an1n16x5 FILLER_43_1648 ();
 b15zdnd11an1n08x5 FILLER_43_1664 ();
 b15zdnd11an1n04x5 FILLER_43_1672 ();
 b15zdnd00an1n01x5 FILLER_43_1676 ();
 b15zdnd11an1n32x5 FILLER_43_1689 ();
 b15zdnd11an1n16x5 FILLER_43_1721 ();
 b15zdnd11an1n08x5 FILLER_43_1737 ();
 b15zdnd11an1n04x5 FILLER_43_1745 ();
 b15zdnd00an1n02x5 FILLER_43_1749 ();
 b15zdnd11an1n16x5 FILLER_43_1769 ();
 b15zdnd11an1n04x5 FILLER_43_1785 ();
 b15zdnd11an1n32x5 FILLER_43_1802 ();
 b15zdnd11an1n16x5 FILLER_43_1834 ();
 b15zdnd00an1n02x5 FILLER_43_1850 ();
 b15zdnd00an1n01x5 FILLER_43_1852 ();
 b15zdnd11an1n64x5 FILLER_43_1859 ();
 b15zdnd11an1n16x5 FILLER_43_1923 ();
 b15zdnd00an1n01x5 FILLER_43_1939 ();
 b15zdnd11an1n64x5 FILLER_43_1944 ();
 b15zdnd00an1n02x5 FILLER_43_2008 ();
 b15zdnd11an1n04x5 FILLER_43_2022 ();
 b15zdnd00an1n02x5 FILLER_43_2026 ();
 b15zdnd11an1n16x5 FILLER_43_2038 ();
 b15zdnd00an1n01x5 FILLER_43_2054 ();
 b15zdnd11an1n08x5 FILLER_43_2075 ();
 b15zdnd11an1n04x5 FILLER_43_2083 ();
 b15zdnd00an1n02x5 FILLER_43_2087 ();
 b15zdnd00an1n01x5 FILLER_43_2089 ();
 b15zdnd11an1n16x5 FILLER_43_2098 ();
 b15zdnd11an1n04x5 FILLER_43_2114 ();
 b15zdnd00an1n02x5 FILLER_43_2118 ();
 b15zdnd00an1n01x5 FILLER_43_2120 ();
 b15zdnd11an1n32x5 FILLER_43_2130 ();
 b15zdnd11an1n16x5 FILLER_43_2162 ();
 b15zdnd11an1n08x5 FILLER_43_2178 ();
 b15zdnd11an1n04x5 FILLER_43_2191 ();
 b15zdnd11an1n04x5 FILLER_43_2204 ();
 b15zdnd11an1n64x5 FILLER_43_2215 ();
 b15zdnd11an1n04x5 FILLER_43_2279 ();
 b15zdnd00an1n01x5 FILLER_43_2283 ();
 b15zdnd11an1n32x5 FILLER_44_8 ();
 b15zdnd11an1n04x5 FILLER_44_40 ();
 b15zdnd11an1n16x5 FILLER_44_52 ();
 b15zdnd11an1n08x5 FILLER_44_68 ();
 b15zdnd00an1n01x5 FILLER_44_76 ();
 b15zdnd11an1n16x5 FILLER_44_86 ();
 b15zdnd11an1n04x5 FILLER_44_102 ();
 b15zdnd00an1n02x5 FILLER_44_106 ();
 b15zdnd11an1n16x5 FILLER_44_113 ();
 b15zdnd11an1n04x5 FILLER_44_134 ();
 b15zdnd11an1n04x5 FILLER_44_159 ();
 b15zdnd11an1n04x5 FILLER_44_175 ();
 b15zdnd11an1n08x5 FILLER_44_191 ();
 b15zdnd00an1n01x5 FILLER_44_199 ();
 b15zdnd11an1n04x5 FILLER_44_212 ();
 b15zdnd11an1n04x5 FILLER_44_226 ();
 b15zdnd11an1n04x5 FILLER_44_235 ();
 b15zdnd11an1n16x5 FILLER_44_250 ();
 b15zdnd11an1n04x5 FILLER_44_266 ();
 b15zdnd00an1n02x5 FILLER_44_270 ();
 b15zdnd11an1n32x5 FILLER_44_282 ();
 b15zdnd11an1n08x5 FILLER_44_314 ();
 b15zdnd11an1n04x5 FILLER_44_322 ();
 b15zdnd00an1n02x5 FILLER_44_326 ();
 b15zdnd11an1n04x5 FILLER_44_339 ();
 b15zdnd11an1n64x5 FILLER_44_356 ();
 b15zdnd11an1n32x5 FILLER_44_420 ();
 b15zdnd11an1n16x5 FILLER_44_452 ();
 b15zdnd11an1n04x5 FILLER_44_468 ();
 b15zdnd00an1n02x5 FILLER_44_472 ();
 b15zdnd00an1n01x5 FILLER_44_474 ();
 b15zdnd11an1n32x5 FILLER_44_489 ();
 b15zdnd11an1n08x5 FILLER_44_521 ();
 b15zdnd11an1n04x5 FILLER_44_529 ();
 b15zdnd11an1n04x5 FILLER_44_539 ();
 b15zdnd00an1n02x5 FILLER_44_543 ();
 b15zdnd00an1n01x5 FILLER_44_545 ();
 b15zdnd11an1n16x5 FILLER_44_572 ();
 b15zdnd11an1n04x5 FILLER_44_588 ();
 b15zdnd00an1n02x5 FILLER_44_592 ();
 b15zdnd00an1n01x5 FILLER_44_594 ();
 b15zdnd11an1n04x5 FILLER_44_611 ();
 b15zdnd11an1n64x5 FILLER_44_625 ();
 b15zdnd11an1n08x5 FILLER_44_689 ();
 b15zdnd11an1n04x5 FILLER_44_697 ();
 b15zdnd00an1n02x5 FILLER_44_701 ();
 b15zdnd11an1n08x5 FILLER_44_707 ();
 b15zdnd00an1n02x5 FILLER_44_715 ();
 b15zdnd00an1n01x5 FILLER_44_717 ();
 b15zdnd11an1n16x5 FILLER_44_726 ();
 b15zdnd11an1n08x5 FILLER_44_742 ();
 b15zdnd00an1n02x5 FILLER_44_750 ();
 b15zdnd00an1n01x5 FILLER_44_752 ();
 b15zdnd11an1n08x5 FILLER_44_759 ();
 b15zdnd11an1n04x5 FILLER_44_775 ();
 b15zdnd11an1n16x5 FILLER_44_785 ();
 b15zdnd00an1n02x5 FILLER_44_801 ();
 b15zdnd11an1n08x5 FILLER_44_835 ();
 b15zdnd00an1n02x5 FILLER_44_843 ();
 b15zdnd00an1n01x5 FILLER_44_845 ();
 b15zdnd11an1n04x5 FILLER_44_853 ();
 b15zdnd11an1n04x5 FILLER_44_863 ();
 b15zdnd11an1n04x5 FILLER_44_872 ();
 b15zdnd00an1n02x5 FILLER_44_876 ();
 b15zdnd11an1n32x5 FILLER_44_884 ();
 b15zdnd11an1n16x5 FILLER_44_916 ();
 b15zdnd11an1n08x5 FILLER_44_932 ();
 b15zdnd00an1n02x5 FILLER_44_940 ();
 b15zdnd00an1n01x5 FILLER_44_942 ();
 b15zdnd11an1n32x5 FILLER_44_963 ();
 b15zdnd11an1n16x5 FILLER_44_995 ();
 b15zdnd11an1n08x5 FILLER_44_1011 ();
 b15zdnd00an1n02x5 FILLER_44_1019 ();
 b15zdnd00an1n01x5 FILLER_44_1021 ();
 b15zdnd11an1n04x5 FILLER_44_1034 ();
 b15zdnd00an1n01x5 FILLER_44_1038 ();
 b15zdnd11an1n04x5 FILLER_44_1047 ();
 b15zdnd00an1n02x5 FILLER_44_1051 ();
 b15zdnd11an1n64x5 FILLER_44_1075 ();
 b15zdnd11an1n16x5 FILLER_44_1139 ();
 b15zdnd11an1n08x5 FILLER_44_1155 ();
 b15zdnd11an1n32x5 FILLER_44_1183 ();
 b15zdnd00an1n02x5 FILLER_44_1215 ();
 b15zdnd00an1n01x5 FILLER_44_1217 ();
 b15zdnd11an1n64x5 FILLER_44_1230 ();
 b15zdnd11an1n04x5 FILLER_44_1294 ();
 b15zdnd00an1n02x5 FILLER_44_1298 ();
 b15zdnd11an1n32x5 FILLER_44_1306 ();
 b15zdnd11an1n16x5 FILLER_44_1338 ();
 b15zdnd11an1n16x5 FILLER_44_1363 ();
 b15zdnd00an1n01x5 FILLER_44_1379 ();
 b15zdnd11an1n08x5 FILLER_44_1393 ();
 b15zdnd00an1n02x5 FILLER_44_1401 ();
 b15zdnd00an1n01x5 FILLER_44_1403 ();
 b15zdnd11an1n08x5 FILLER_44_1414 ();
 b15zdnd11an1n04x5 FILLER_44_1422 ();
 b15zdnd00an1n02x5 FILLER_44_1426 ();
 b15zdnd11an1n64x5 FILLER_44_1437 ();
 b15zdnd11an1n64x5 FILLER_44_1501 ();
 b15zdnd11an1n04x5 FILLER_44_1565 ();
 b15zdnd00an1n02x5 FILLER_44_1569 ();
 b15zdnd00an1n01x5 FILLER_44_1571 ();
 b15zdnd11an1n16x5 FILLER_44_1598 ();
 b15zdnd00an1n02x5 FILLER_44_1614 ();
 b15zdnd11an1n16x5 FILLER_44_1621 ();
 b15zdnd11an1n32x5 FILLER_44_1650 ();
 b15zdnd00an1n01x5 FILLER_44_1682 ();
 b15zdnd11an1n32x5 FILLER_44_1692 ();
 b15zdnd11an1n16x5 FILLER_44_1724 ();
 b15zdnd11an1n04x5 FILLER_44_1740 ();
 b15zdnd00an1n02x5 FILLER_44_1744 ();
 b15zdnd00an1n01x5 FILLER_44_1746 ();
 b15zdnd11an1n04x5 FILLER_44_1751 ();
 b15zdnd00an1n02x5 FILLER_44_1755 ();
 b15zdnd11an1n32x5 FILLER_44_1778 ();
 b15zdnd11an1n16x5 FILLER_44_1810 ();
 b15zdnd11an1n08x5 FILLER_44_1826 ();
 b15zdnd11an1n04x5 FILLER_44_1834 ();
 b15zdnd00an1n01x5 FILLER_44_1838 ();
 b15zdnd11an1n04x5 FILLER_44_1857 ();
 b15zdnd11an1n32x5 FILLER_44_1868 ();
 b15zdnd00an1n02x5 FILLER_44_1900 ();
 b15zdnd11an1n16x5 FILLER_44_1914 ();
 b15zdnd11an1n08x5 FILLER_44_1930 ();
 b15zdnd00an1n02x5 FILLER_44_1938 ();
 b15zdnd11an1n64x5 FILLER_44_1945 ();
 b15zdnd11an1n16x5 FILLER_44_2009 ();
 b15zdnd00an1n02x5 FILLER_44_2025 ();
 b15zdnd00an1n01x5 FILLER_44_2027 ();
 b15zdnd11an1n16x5 FILLER_44_2034 ();
 b15zdnd11an1n08x5 FILLER_44_2050 ();
 b15zdnd11an1n32x5 FILLER_44_2082 ();
 b15zdnd11an1n08x5 FILLER_44_2114 ();
 b15zdnd11an1n04x5 FILLER_44_2122 ();
 b15zdnd00an1n02x5 FILLER_44_2126 ();
 b15zdnd00an1n02x5 FILLER_44_2152 ();
 b15zdnd11an1n08x5 FILLER_44_2162 ();
 b15zdnd11an1n04x5 FILLER_44_2170 ();
 b15zdnd00an1n02x5 FILLER_44_2174 ();
 b15zdnd00an1n01x5 FILLER_44_2176 ();
 b15zdnd11an1n64x5 FILLER_44_2187 ();
 b15zdnd11an1n16x5 FILLER_44_2251 ();
 b15zdnd11an1n08x5 FILLER_44_2267 ();
 b15zdnd00an1n01x5 FILLER_44_2275 ();
 b15zdnd11an1n32x5 FILLER_45_0 ();
 b15zdnd11an1n04x5 FILLER_45_32 ();
 b15zdnd00an1n02x5 FILLER_45_36 ();
 b15zdnd11an1n08x5 FILLER_45_52 ();
 b15zdnd11an1n04x5 FILLER_45_60 ();
 b15zdnd11an1n04x5 FILLER_45_68 ();
 b15zdnd00an1n02x5 FILLER_45_72 ();
 b15zdnd11an1n08x5 FILLER_45_88 ();
 b15zdnd11an1n32x5 FILLER_45_117 ();
 b15zdnd11an1n08x5 FILLER_45_149 ();
 b15zdnd11an1n04x5 FILLER_45_157 ();
 b15zdnd00an1n02x5 FILLER_45_161 ();
 b15zdnd00an1n01x5 FILLER_45_163 ();
 b15zdnd11an1n64x5 FILLER_45_176 ();
 b15zdnd11an1n32x5 FILLER_45_240 ();
 b15zdnd11an1n04x5 FILLER_45_272 ();
 b15zdnd11an1n64x5 FILLER_45_286 ();
 b15zdnd11an1n64x5 FILLER_45_350 ();
 b15zdnd11an1n64x5 FILLER_45_414 ();
 b15zdnd11an1n16x5 FILLER_45_478 ();
 b15zdnd11an1n08x5 FILLER_45_506 ();
 b15zdnd00an1n01x5 FILLER_45_514 ();
 b15zdnd11an1n04x5 FILLER_45_521 ();
 b15zdnd11an1n32x5 FILLER_45_537 ();
 b15zdnd11an1n32x5 FILLER_45_580 ();
 b15zdnd11an1n04x5 FILLER_45_618 ();
 b15zdnd11an1n16x5 FILLER_45_632 ();
 b15zdnd11an1n04x5 FILLER_45_648 ();
 b15zdnd00an1n01x5 FILLER_45_652 ();
 b15zdnd11an1n04x5 FILLER_45_662 ();
 b15zdnd11an1n64x5 FILLER_45_697 ();
 b15zdnd11an1n32x5 FILLER_45_761 ();
 b15zdnd11an1n16x5 FILLER_45_793 ();
 b15zdnd11an1n08x5 FILLER_45_809 ();
 b15zdnd11an1n04x5 FILLER_45_817 ();
 b15zdnd00an1n01x5 FILLER_45_821 ();
 b15zdnd11an1n16x5 FILLER_45_827 ();
 b15zdnd11an1n08x5 FILLER_45_843 ();
 b15zdnd00an1n02x5 FILLER_45_851 ();
 b15zdnd00an1n01x5 FILLER_45_853 ();
 b15zdnd11an1n16x5 FILLER_45_861 ();
 b15zdnd11an1n08x5 FILLER_45_877 ();
 b15zdnd11an1n04x5 FILLER_45_885 ();
 b15zdnd00an1n02x5 FILLER_45_889 ();
 b15zdnd00an1n01x5 FILLER_45_891 ();
 b15zdnd11an1n08x5 FILLER_45_902 ();
 b15zdnd11an1n04x5 FILLER_45_910 ();
 b15zdnd00an1n02x5 FILLER_45_914 ();
 b15zdnd00an1n01x5 FILLER_45_916 ();
 b15zdnd11an1n64x5 FILLER_45_937 ();
 b15zdnd11an1n08x5 FILLER_45_1001 ();
 b15zdnd11an1n04x5 FILLER_45_1009 ();
 b15zdnd11an1n04x5 FILLER_45_1034 ();
 b15zdnd00an1n01x5 FILLER_45_1038 ();
 b15zdnd11an1n64x5 FILLER_45_1059 ();
 b15zdnd11an1n32x5 FILLER_45_1123 ();
 b15zdnd11an1n16x5 FILLER_45_1155 ();
 b15zdnd11an1n08x5 FILLER_45_1202 ();
 b15zdnd11an1n04x5 FILLER_45_1210 ();
 b15zdnd00an1n02x5 FILLER_45_1214 ();
 b15zdnd00an1n01x5 FILLER_45_1216 ();
 b15zdnd11an1n08x5 FILLER_45_1242 ();
 b15zdnd00an1n02x5 FILLER_45_1250 ();
 b15zdnd00an1n01x5 FILLER_45_1252 ();
 b15zdnd11an1n32x5 FILLER_45_1268 ();
 b15zdnd11an1n16x5 FILLER_45_1300 ();
 b15zdnd11an1n08x5 FILLER_45_1316 ();
 b15zdnd11an1n32x5 FILLER_45_1331 ();
 b15zdnd11an1n16x5 FILLER_45_1363 ();
 b15zdnd00an1n01x5 FILLER_45_1379 ();
 b15zdnd11an1n08x5 FILLER_45_1385 ();
 b15zdnd00an1n02x5 FILLER_45_1393 ();
 b15zdnd11an1n32x5 FILLER_45_1416 ();
 b15zdnd11an1n16x5 FILLER_45_1454 ();
 b15zdnd11an1n08x5 FILLER_45_1470 ();
 b15zdnd11an1n04x5 FILLER_45_1478 ();
 b15zdnd00an1n02x5 FILLER_45_1482 ();
 b15zdnd00an1n01x5 FILLER_45_1484 ();
 b15zdnd11an1n64x5 FILLER_45_1501 ();
 b15zdnd11an1n08x5 FILLER_45_1565 ();
 b15zdnd00an1n02x5 FILLER_45_1573 ();
 b15zdnd00an1n01x5 FILLER_45_1575 ();
 b15zdnd11an1n32x5 FILLER_45_1588 ();
 b15zdnd00an1n02x5 FILLER_45_1620 ();
 b15zdnd11an1n64x5 FILLER_45_1634 ();
 b15zdnd11an1n64x5 FILLER_45_1698 ();
 b15zdnd11an1n16x5 FILLER_45_1762 ();
 b15zdnd11an1n08x5 FILLER_45_1778 ();
 b15zdnd11an1n04x5 FILLER_45_1786 ();
 b15zdnd11an1n04x5 FILLER_45_1800 ();
 b15zdnd00an1n02x5 FILLER_45_1804 ();
 b15zdnd00an1n01x5 FILLER_45_1806 ();
 b15zdnd11an1n08x5 FILLER_45_1813 ();
 b15zdnd11an1n04x5 FILLER_45_1821 ();
 b15zdnd00an1n02x5 FILLER_45_1825 ();
 b15zdnd00an1n01x5 FILLER_45_1827 ();
 b15zdnd11an1n08x5 FILLER_45_1833 ();
 b15zdnd11an1n04x5 FILLER_45_1841 ();
 b15zdnd00an1n02x5 FILLER_45_1845 ();
 b15zdnd00an1n01x5 FILLER_45_1847 ();
 b15zdnd11an1n64x5 FILLER_45_1860 ();
 b15zdnd11an1n08x5 FILLER_45_1924 ();
 b15zdnd11an1n04x5 FILLER_45_1932 ();
 b15zdnd00an1n02x5 FILLER_45_1936 ();
 b15zdnd11an1n16x5 FILLER_45_1947 ();
 b15zdnd11an1n08x5 FILLER_45_1963 ();
 b15zdnd11an1n04x5 FILLER_45_1971 ();
 b15zdnd00an1n02x5 FILLER_45_1975 ();
 b15zdnd00an1n01x5 FILLER_45_1977 ();
 b15zdnd11an1n32x5 FILLER_45_1983 ();
 b15zdnd11an1n08x5 FILLER_45_2015 ();
 b15zdnd11an1n04x5 FILLER_45_2023 ();
 b15zdnd11an1n64x5 FILLER_45_2036 ();
 b15zdnd11an1n32x5 FILLER_45_2100 ();
 b15zdnd11an1n16x5 FILLER_45_2132 ();
 b15zdnd00an1n02x5 FILLER_45_2148 ();
 b15zdnd00an1n01x5 FILLER_45_2150 ();
 b15zdnd11an1n16x5 FILLER_45_2161 ();
 b15zdnd11an1n04x5 FILLER_45_2177 ();
 b15zdnd11an1n64x5 FILLER_45_2188 ();
 b15zdnd11an1n32x5 FILLER_45_2252 ();
 b15zdnd11an1n64x5 FILLER_46_8 ();
 b15zdnd11an1n04x5 FILLER_46_72 ();
 b15zdnd00an1n02x5 FILLER_46_76 ();
 b15zdnd00an1n01x5 FILLER_46_78 ();
 b15zdnd11an1n04x5 FILLER_46_99 ();
 b15zdnd00an1n02x5 FILLER_46_103 ();
 b15zdnd00an1n01x5 FILLER_46_105 ();
 b15zdnd11an1n64x5 FILLER_46_110 ();
 b15zdnd11an1n16x5 FILLER_46_174 ();
 b15zdnd11an1n08x5 FILLER_46_190 ();
 b15zdnd11an1n32x5 FILLER_46_203 ();
 b15zdnd11an1n04x5 FILLER_46_235 ();
 b15zdnd00an1n02x5 FILLER_46_239 ();
 b15zdnd00an1n01x5 FILLER_46_241 ();
 b15zdnd11an1n08x5 FILLER_46_268 ();
 b15zdnd11an1n04x5 FILLER_46_276 ();
 b15zdnd00an1n02x5 FILLER_46_280 ();
 b15zdnd11an1n04x5 FILLER_46_287 ();
 b15zdnd00an1n02x5 FILLER_46_291 ();
 b15zdnd00an1n01x5 FILLER_46_293 ();
 b15zdnd11an1n32x5 FILLER_46_300 ();
 b15zdnd11an1n16x5 FILLER_46_332 ();
 b15zdnd11an1n08x5 FILLER_46_348 ();
 b15zdnd11an1n04x5 FILLER_46_356 ();
 b15zdnd11an1n64x5 FILLER_46_364 ();
 b15zdnd11an1n16x5 FILLER_46_428 ();
 b15zdnd11an1n08x5 FILLER_46_449 ();
 b15zdnd00an1n02x5 FILLER_46_457 ();
 b15zdnd00an1n01x5 FILLER_46_459 ();
 b15zdnd11an1n04x5 FILLER_46_479 ();
 b15zdnd11an1n04x5 FILLER_46_490 ();
 b15zdnd11an1n04x5 FILLER_46_501 ();
 b15zdnd11an1n04x5 FILLER_46_517 ();
 b15zdnd11an1n16x5 FILLER_46_542 ();
 b15zdnd11an1n04x5 FILLER_46_558 ();
 b15zdnd11an1n04x5 FILLER_46_566 ();
 b15zdnd00an1n02x5 FILLER_46_570 ();
 b15zdnd00an1n01x5 FILLER_46_572 ();
 b15zdnd11an1n08x5 FILLER_46_578 ();
 b15zdnd00an1n01x5 FILLER_46_586 ();
 b15zdnd11an1n16x5 FILLER_46_599 ();
 b15zdnd11an1n04x5 FILLER_46_615 ();
 b15zdnd00an1n02x5 FILLER_46_619 ();
 b15zdnd00an1n01x5 FILLER_46_621 ();
 b15zdnd11an1n04x5 FILLER_46_627 ();
 b15zdnd11an1n08x5 FILLER_46_636 ();
 b15zdnd11an1n04x5 FILLER_46_644 ();
 b15zdnd00an1n02x5 FILLER_46_648 ();
 b15zdnd00an1n01x5 FILLER_46_650 ();
 b15zdnd11an1n04x5 FILLER_46_665 ();
 b15zdnd11an1n16x5 FILLER_46_690 ();
 b15zdnd11an1n08x5 FILLER_46_706 ();
 b15zdnd11an1n04x5 FILLER_46_714 ();
 b15zdnd11an1n32x5 FILLER_46_726 ();
 b15zdnd11an1n08x5 FILLER_46_758 ();
 b15zdnd11an1n04x5 FILLER_46_766 ();
 b15zdnd00an1n02x5 FILLER_46_770 ();
 b15zdnd00an1n01x5 FILLER_46_772 ();
 b15zdnd11an1n32x5 FILLER_46_787 ();
 b15zdnd00an1n01x5 FILLER_46_819 ();
 b15zdnd11an1n64x5 FILLER_46_825 ();
 b15zdnd11an1n08x5 FILLER_46_889 ();
 b15zdnd00an1n01x5 FILLER_46_897 ();
 b15zdnd11an1n64x5 FILLER_46_908 ();
 b15zdnd11an1n16x5 FILLER_46_972 ();
 b15zdnd11an1n04x5 FILLER_46_988 ();
 b15zdnd00an1n02x5 FILLER_46_992 ();
 b15zdnd00an1n01x5 FILLER_46_994 ();
 b15zdnd11an1n64x5 FILLER_46_1026 ();
 b15zdnd11an1n04x5 FILLER_46_1090 ();
 b15zdnd00an1n02x5 FILLER_46_1094 ();
 b15zdnd00an1n01x5 FILLER_46_1096 ();
 b15zdnd11an1n08x5 FILLER_46_1121 ();
 b15zdnd11an1n04x5 FILLER_46_1129 ();
 b15zdnd00an1n02x5 FILLER_46_1133 ();
 b15zdnd11an1n16x5 FILLER_46_1166 ();
 b15zdnd00an1n02x5 FILLER_46_1182 ();
 b15zdnd00an1n01x5 FILLER_46_1184 ();
 b15zdnd11an1n64x5 FILLER_46_1190 ();
 b15zdnd11an1n16x5 FILLER_46_1254 ();
 b15zdnd11an1n08x5 FILLER_46_1270 ();
 b15zdnd11an1n04x5 FILLER_46_1282 ();
 b15zdnd00an1n02x5 FILLER_46_1286 ();
 b15zdnd11an1n08x5 FILLER_46_1294 ();
 b15zdnd11an1n16x5 FILLER_46_1308 ();
 b15zdnd00an1n01x5 FILLER_46_1324 ();
 b15zdnd11an1n64x5 FILLER_46_1335 ();
 b15zdnd11an1n32x5 FILLER_46_1399 ();
 b15zdnd11an1n08x5 FILLER_46_1431 ();
 b15zdnd11an1n04x5 FILLER_46_1439 ();
 b15zdnd00an1n02x5 FILLER_46_1443 ();
 b15zdnd11an1n64x5 FILLER_46_1461 ();
 b15zdnd11an1n16x5 FILLER_46_1531 ();
 b15zdnd11an1n08x5 FILLER_46_1547 ();
 b15zdnd11an1n04x5 FILLER_46_1562 ();
 b15zdnd00an1n02x5 FILLER_46_1566 ();
 b15zdnd00an1n01x5 FILLER_46_1568 ();
 b15zdnd11an1n08x5 FILLER_46_1585 ();
 b15zdnd11an1n16x5 FILLER_46_1601 ();
 b15zdnd11an1n04x5 FILLER_46_1617 ();
 b15zdnd11an1n16x5 FILLER_46_1628 ();
 b15zdnd11an1n04x5 FILLER_46_1644 ();
 b15zdnd11an1n16x5 FILLER_46_1652 ();
 b15zdnd11an1n08x5 FILLER_46_1668 ();
 b15zdnd00an1n02x5 FILLER_46_1676 ();
 b15zdnd00an1n01x5 FILLER_46_1678 ();
 b15zdnd11an1n64x5 FILLER_46_1683 ();
 b15zdnd00an1n02x5 FILLER_46_1747 ();
 b15zdnd11an1n04x5 FILLER_46_1757 ();
 b15zdnd11an1n32x5 FILLER_46_1767 ();
 b15zdnd11an1n08x5 FILLER_46_1799 ();
 b15zdnd00an1n02x5 FILLER_46_1807 ();
 b15zdnd11an1n04x5 FILLER_46_1820 ();
 b15zdnd00an1n01x5 FILLER_46_1824 ();
 b15zdnd11an1n04x5 FILLER_46_1829 ();
 b15zdnd11an1n08x5 FILLER_46_1840 ();
 b15zdnd00an1n02x5 FILLER_46_1848 ();
 b15zdnd00an1n01x5 FILLER_46_1850 ();
 b15zdnd11an1n08x5 FILLER_46_1858 ();
 b15zdnd00an1n01x5 FILLER_46_1866 ();
 b15zdnd11an1n16x5 FILLER_46_1873 ();
 b15zdnd11an1n08x5 FILLER_46_1889 ();
 b15zdnd11an1n04x5 FILLER_46_1909 ();
 b15zdnd11an1n32x5 FILLER_46_1918 ();
 b15zdnd11an1n08x5 FILLER_46_1950 ();
 b15zdnd00an1n02x5 FILLER_46_1958 ();
 b15zdnd11an1n08x5 FILLER_46_1970 ();
 b15zdnd11an1n32x5 FILLER_46_1990 ();
 b15zdnd11an1n16x5 FILLER_46_2022 ();
 b15zdnd11an1n04x5 FILLER_46_2038 ();
 b15zdnd00an1n02x5 FILLER_46_2042 ();
 b15zdnd11an1n04x5 FILLER_46_2053 ();
 b15zdnd11an1n04x5 FILLER_46_2062 ();
 b15zdnd11an1n16x5 FILLER_46_2072 ();
 b15zdnd11an1n08x5 FILLER_46_2088 ();
 b15zdnd11an1n04x5 FILLER_46_2096 ();
 b15zdnd11an1n16x5 FILLER_46_2109 ();
 b15zdnd11an1n04x5 FILLER_46_2125 ();
 b15zdnd00an1n01x5 FILLER_46_2129 ();
 b15zdnd11an1n04x5 FILLER_46_2136 ();
 b15zdnd11an1n08x5 FILLER_46_2145 ();
 b15zdnd00an1n01x5 FILLER_46_2153 ();
 b15zdnd11an1n08x5 FILLER_46_2162 ();
 b15zdnd00an1n02x5 FILLER_46_2170 ();
 b15zdnd11an1n16x5 FILLER_46_2184 ();
 b15zdnd00an1n01x5 FILLER_46_2200 ();
 b15zdnd11an1n32x5 FILLER_46_2215 ();
 b15zdnd11an1n16x5 FILLER_46_2247 ();
 b15zdnd11an1n08x5 FILLER_46_2263 ();
 b15zdnd11an1n04x5 FILLER_46_2271 ();
 b15zdnd00an1n01x5 FILLER_46_2275 ();
 b15zdnd11an1n32x5 FILLER_47_0 ();
 b15zdnd11an1n16x5 FILLER_47_42 ();
 b15zdnd11an1n04x5 FILLER_47_58 ();
 b15zdnd00an1n02x5 FILLER_47_62 ();
 b15zdnd11an1n32x5 FILLER_47_68 ();
 b15zdnd11an1n08x5 FILLER_47_100 ();
 b15zdnd11an1n04x5 FILLER_47_108 ();
 b15zdnd11an1n04x5 FILLER_47_118 ();
 b15zdnd11an1n64x5 FILLER_47_132 ();
 b15zdnd11an1n64x5 FILLER_47_196 ();
 b15zdnd11an1n32x5 FILLER_47_260 ();
 b15zdnd11an1n08x5 FILLER_47_292 ();
 b15zdnd11an1n04x5 FILLER_47_300 ();
 b15zdnd00an1n01x5 FILLER_47_304 ();
 b15zdnd11an1n04x5 FILLER_47_318 ();
 b15zdnd00an1n01x5 FILLER_47_322 ();
 b15zdnd11an1n64x5 FILLER_47_333 ();
 b15zdnd11an1n32x5 FILLER_47_397 ();
 b15zdnd11an1n08x5 FILLER_47_429 ();
 b15zdnd00an1n02x5 FILLER_47_437 ();
 b15zdnd00an1n01x5 FILLER_47_439 ();
 b15zdnd11an1n64x5 FILLER_47_444 ();
 b15zdnd11an1n64x5 FILLER_47_508 ();
 b15zdnd11an1n08x5 FILLER_47_572 ();
 b15zdnd11an1n04x5 FILLER_47_580 ();
 b15zdnd00an1n02x5 FILLER_47_584 ();
 b15zdnd11an1n64x5 FILLER_47_591 ();
 b15zdnd11an1n64x5 FILLER_47_655 ();
 b15zdnd11an1n04x5 FILLER_47_719 ();
 b15zdnd11an1n64x5 FILLER_47_732 ();
 b15zdnd11an1n04x5 FILLER_47_796 ();
 b15zdnd00an1n01x5 FILLER_47_800 ();
 b15zdnd11an1n32x5 FILLER_47_811 ();
 b15zdnd11an1n16x5 FILLER_47_843 ();
 b15zdnd00an1n02x5 FILLER_47_859 ();
 b15zdnd11an1n64x5 FILLER_47_887 ();
 b15zdnd11an1n64x5 FILLER_47_951 ();
 b15zdnd11an1n64x5 FILLER_47_1015 ();
 b15zdnd11an1n08x5 FILLER_47_1079 ();
 b15zdnd11an1n04x5 FILLER_47_1087 ();
 b15zdnd00an1n01x5 FILLER_47_1091 ();
 b15zdnd11an1n16x5 FILLER_47_1107 ();
 b15zdnd00an1n02x5 FILLER_47_1123 ();
 b15zdnd11an1n16x5 FILLER_47_1144 ();
 b15zdnd00an1n02x5 FILLER_47_1160 ();
 b15zdnd11an1n04x5 FILLER_47_1180 ();
 b15zdnd11an1n64x5 FILLER_47_1204 ();
 b15zdnd11an1n64x5 FILLER_47_1268 ();
 b15zdnd11an1n16x5 FILLER_47_1332 ();
 b15zdnd11an1n04x5 FILLER_47_1348 ();
 b15zdnd11an1n32x5 FILLER_47_1358 ();
 b15zdnd11an1n08x5 FILLER_47_1390 ();
 b15zdnd11an1n04x5 FILLER_47_1398 ();
 b15zdnd00an1n02x5 FILLER_47_1402 ();
 b15zdnd00an1n01x5 FILLER_47_1404 ();
 b15zdnd11an1n08x5 FILLER_47_1411 ();
 b15zdnd00an1n01x5 FILLER_47_1419 ();
 b15zdnd11an1n16x5 FILLER_47_1430 ();
 b15zdnd00an1n02x5 FILLER_47_1446 ();
 b15zdnd00an1n01x5 FILLER_47_1448 ();
 b15zdnd11an1n16x5 FILLER_47_1456 ();
 b15zdnd11an1n08x5 FILLER_47_1472 ();
 b15zdnd11an1n04x5 FILLER_47_1480 ();
 b15zdnd00an1n02x5 FILLER_47_1484 ();
 b15zdnd11an1n08x5 FILLER_47_1491 ();
 b15zdnd11an1n32x5 FILLER_47_1506 ();
 b15zdnd11an1n08x5 FILLER_47_1538 ();
 b15zdnd11an1n04x5 FILLER_47_1546 ();
 b15zdnd00an1n01x5 FILLER_47_1550 ();
 b15zdnd11an1n32x5 FILLER_47_1558 ();
 b15zdnd11an1n32x5 FILLER_47_1596 ();
 b15zdnd11an1n08x5 FILLER_47_1628 ();
 b15zdnd00an1n02x5 FILLER_47_1636 ();
 b15zdnd11an1n32x5 FILLER_47_1642 ();
 b15zdnd11an1n04x5 FILLER_47_1674 ();
 b15zdnd00an1n01x5 FILLER_47_1678 ();
 b15zdnd11an1n64x5 FILLER_47_1688 ();
 b15zdnd11an1n16x5 FILLER_47_1752 ();
 b15zdnd11an1n08x5 FILLER_47_1768 ();
 b15zdnd11an1n04x5 FILLER_47_1783 ();
 b15zdnd11an1n16x5 FILLER_47_1791 ();
 b15zdnd11an1n08x5 FILLER_47_1807 ();
 b15zdnd00an1n01x5 FILLER_47_1815 ();
 b15zdnd11an1n08x5 FILLER_47_1820 ();
 b15zdnd11an1n04x5 FILLER_47_1828 ();
 b15zdnd00an1n02x5 FILLER_47_1832 ();
 b15zdnd00an1n01x5 FILLER_47_1834 ();
 b15zdnd11an1n08x5 FILLER_47_1839 ();
 b15zdnd11an1n04x5 FILLER_47_1847 ();
 b15zdnd11an1n08x5 FILLER_47_1856 ();
 b15zdnd00an1n02x5 FILLER_47_1864 ();
 b15zdnd00an1n01x5 FILLER_47_1866 ();
 b15zdnd11an1n16x5 FILLER_47_1871 ();
 b15zdnd11an1n04x5 FILLER_47_1887 ();
 b15zdnd00an1n02x5 FILLER_47_1891 ();
 b15zdnd11an1n04x5 FILLER_47_1900 ();
 b15zdnd11an1n32x5 FILLER_47_1910 ();
 b15zdnd11an1n08x5 FILLER_47_1942 ();
 b15zdnd00an1n02x5 FILLER_47_1950 ();
 b15zdnd00an1n01x5 FILLER_47_1952 ();
 b15zdnd11an1n08x5 FILLER_47_1974 ();
 b15zdnd11an1n16x5 FILLER_47_1988 ();
 b15zdnd11an1n04x5 FILLER_47_2004 ();
 b15zdnd00an1n02x5 FILLER_47_2008 ();
 b15zdnd11an1n16x5 FILLER_47_2019 ();
 b15zdnd00an1n01x5 FILLER_47_2035 ();
 b15zdnd11an1n64x5 FILLER_47_2046 ();
 b15zdnd11an1n16x5 FILLER_47_2110 ();
 b15zdnd11an1n04x5 FILLER_47_2126 ();
 b15zdnd00an1n01x5 FILLER_47_2130 ();
 b15zdnd11an1n32x5 FILLER_47_2143 ();
 b15zdnd11an1n16x5 FILLER_47_2175 ();
 b15zdnd00an1n01x5 FILLER_47_2191 ();
 b15zdnd11an1n64x5 FILLER_47_2202 ();
 b15zdnd11an1n16x5 FILLER_47_2266 ();
 b15zdnd00an1n02x5 FILLER_47_2282 ();
 b15zdnd11an1n32x5 FILLER_48_8 ();
 b15zdnd11an1n04x5 FILLER_48_40 ();
 b15zdnd00an1n02x5 FILLER_48_44 ();
 b15zdnd11an1n64x5 FILLER_48_60 ();
 b15zdnd11an1n08x5 FILLER_48_124 ();
 b15zdnd11an1n04x5 FILLER_48_132 ();
 b15zdnd11an1n04x5 FILLER_48_141 ();
 b15zdnd00an1n02x5 FILLER_48_145 ();
 b15zdnd00an1n01x5 FILLER_48_147 ();
 b15zdnd11an1n08x5 FILLER_48_153 ();
 b15zdnd00an1n02x5 FILLER_48_161 ();
 b15zdnd11an1n08x5 FILLER_48_173 ();
 b15zdnd00an1n02x5 FILLER_48_181 ();
 b15zdnd11an1n08x5 FILLER_48_190 ();
 b15zdnd11an1n64x5 FILLER_48_203 ();
 b15zdnd11an1n16x5 FILLER_48_267 ();
 b15zdnd11an1n08x5 FILLER_48_283 ();
 b15zdnd11an1n08x5 FILLER_48_300 ();
 b15zdnd11an1n04x5 FILLER_48_308 ();
 b15zdnd00an1n01x5 FILLER_48_312 ();
 b15zdnd11an1n16x5 FILLER_48_329 ();
 b15zdnd11an1n04x5 FILLER_48_345 ();
 b15zdnd00an1n02x5 FILLER_48_349 ();
 b15zdnd11an1n04x5 FILLER_48_355 ();
 b15zdnd11an1n64x5 FILLER_48_371 ();
 b15zdnd11an1n16x5 FILLER_48_435 ();
 b15zdnd11an1n08x5 FILLER_48_451 ();
 b15zdnd11an1n04x5 FILLER_48_459 ();
 b15zdnd00an1n02x5 FILLER_48_463 ();
 b15zdnd11an1n64x5 FILLER_48_477 ();
 b15zdnd11an1n04x5 FILLER_48_541 ();
 b15zdnd11an1n64x5 FILLER_48_551 ();
 b15zdnd11an1n32x5 FILLER_48_615 ();
 b15zdnd11an1n08x5 FILLER_48_647 ();
 b15zdnd00an1n02x5 FILLER_48_655 ();
 b15zdnd11an1n08x5 FILLER_48_667 ();
 b15zdnd11an1n04x5 FILLER_48_675 ();
 b15zdnd00an1n02x5 FILLER_48_679 ();
 b15zdnd00an1n01x5 FILLER_48_681 ();
 b15zdnd11an1n08x5 FILLER_48_686 ();
 b15zdnd11an1n04x5 FILLER_48_694 ();
 b15zdnd11an1n08x5 FILLER_48_708 ();
 b15zdnd00an1n02x5 FILLER_48_716 ();
 b15zdnd00an1n02x5 FILLER_48_726 ();
 b15zdnd11an1n04x5 FILLER_48_738 ();
 b15zdnd11an1n16x5 FILLER_48_746 ();
 b15zdnd00an1n01x5 FILLER_48_762 ();
 b15zdnd11an1n16x5 FILLER_48_769 ();
 b15zdnd11an1n08x5 FILLER_48_806 ();
 b15zdnd11an1n04x5 FILLER_48_814 ();
 b15zdnd00an1n02x5 FILLER_48_818 ();
 b15zdnd11an1n64x5 FILLER_48_831 ();
 b15zdnd11an1n08x5 FILLER_48_895 ();
 b15zdnd00an1n01x5 FILLER_48_903 ();
 b15zdnd11an1n08x5 FILLER_48_930 ();
 b15zdnd11an1n04x5 FILLER_48_938 ();
 b15zdnd00an1n02x5 FILLER_48_942 ();
 b15zdnd00an1n01x5 FILLER_48_944 ();
 b15zdnd11an1n08x5 FILLER_48_957 ();
 b15zdnd11an1n04x5 FILLER_48_965 ();
 b15zdnd11an1n16x5 FILLER_48_973 ();
 b15zdnd11an1n04x5 FILLER_48_989 ();
 b15zdnd11an1n16x5 FILLER_48_1002 ();
 b15zdnd11an1n08x5 FILLER_48_1018 ();
 b15zdnd11an1n04x5 FILLER_48_1026 ();
 b15zdnd11an1n64x5 FILLER_48_1061 ();
 b15zdnd11an1n32x5 FILLER_48_1125 ();
 b15zdnd11an1n08x5 FILLER_48_1157 ();
 b15zdnd00an1n02x5 FILLER_48_1165 ();
 b15zdnd00an1n01x5 FILLER_48_1167 ();
 b15zdnd11an1n64x5 FILLER_48_1180 ();
 b15zdnd11an1n32x5 FILLER_48_1244 ();
 b15zdnd11an1n16x5 FILLER_48_1276 ();
 b15zdnd11an1n08x5 FILLER_48_1292 ();
 b15zdnd00an1n02x5 FILLER_48_1300 ();
 b15zdnd11an1n16x5 FILLER_48_1314 ();
 b15zdnd11an1n08x5 FILLER_48_1330 ();
 b15zdnd00an1n02x5 FILLER_48_1338 ();
 b15zdnd00an1n01x5 FILLER_48_1340 ();
 b15zdnd11an1n64x5 FILLER_48_1355 ();
 b15zdnd11an1n08x5 FILLER_48_1419 ();
 b15zdnd11an1n16x5 FILLER_48_1432 ();
 b15zdnd00an1n01x5 FILLER_48_1448 ();
 b15zdnd11an1n08x5 FILLER_48_1458 ();
 b15zdnd11an1n04x5 FILLER_48_1466 ();
 b15zdnd00an1n02x5 FILLER_48_1470 ();
 b15zdnd00an1n01x5 FILLER_48_1472 ();
 b15zdnd11an1n08x5 FILLER_48_1478 ();
 b15zdnd00an1n02x5 FILLER_48_1486 ();
 b15zdnd00an1n01x5 FILLER_48_1488 ();
 b15zdnd11an1n16x5 FILLER_48_1501 ();
 b15zdnd11an1n04x5 FILLER_48_1517 ();
 b15zdnd00an1n02x5 FILLER_48_1521 ();
 b15zdnd00an1n01x5 FILLER_48_1523 ();
 b15zdnd11an1n16x5 FILLER_48_1534 ();
 b15zdnd11an1n64x5 FILLER_48_1562 ();
 b15zdnd11an1n08x5 FILLER_48_1626 ();
 b15zdnd00an1n02x5 FILLER_48_1634 ();
 b15zdnd11an1n04x5 FILLER_48_1645 ();
 b15zdnd00an1n02x5 FILLER_48_1649 ();
 b15zdnd11an1n08x5 FILLER_48_1655 ();
 b15zdnd11an1n04x5 FILLER_48_1663 ();
 b15zdnd11an1n64x5 FILLER_48_1693 ();
 b15zdnd11an1n32x5 FILLER_48_1757 ();
 b15zdnd11an1n16x5 FILLER_48_1789 ();
 b15zdnd11an1n04x5 FILLER_48_1805 ();
 b15zdnd00an1n02x5 FILLER_48_1809 ();
 b15zdnd11an1n64x5 FILLER_48_1818 ();
 b15zdnd11an1n32x5 FILLER_48_1882 ();
 b15zdnd11an1n04x5 FILLER_48_1914 ();
 b15zdnd11an1n32x5 FILLER_48_1928 ();
 b15zdnd11an1n16x5 FILLER_48_1960 ();
 b15zdnd11an1n04x5 FILLER_48_1976 ();
 b15zdnd00an1n02x5 FILLER_48_1980 ();
 b15zdnd11an1n32x5 FILLER_48_1986 ();
 b15zdnd11an1n08x5 FILLER_48_2018 ();
 b15zdnd00an1n01x5 FILLER_48_2026 ();
 b15zdnd11an1n04x5 FILLER_48_2041 ();
 b15zdnd11an1n64x5 FILLER_48_2056 ();
 b15zdnd11an1n32x5 FILLER_48_2120 ();
 b15zdnd00an1n02x5 FILLER_48_2152 ();
 b15zdnd11an1n64x5 FILLER_48_2162 ();
 b15zdnd11an1n32x5 FILLER_48_2226 ();
 b15zdnd11an1n16x5 FILLER_48_2258 ();
 b15zdnd00an1n02x5 FILLER_48_2274 ();
 b15zdnd11an1n32x5 FILLER_49_0 ();
 b15zdnd11an1n08x5 FILLER_49_32 ();
 b15zdnd11an1n08x5 FILLER_49_50 ();
 b15zdnd11an1n04x5 FILLER_49_58 ();
 b15zdnd11an1n32x5 FILLER_49_75 ();
 b15zdnd11an1n08x5 FILLER_49_107 ();
 b15zdnd11an1n04x5 FILLER_49_115 ();
 b15zdnd11an1n32x5 FILLER_49_128 ();
 b15zdnd11an1n64x5 FILLER_49_164 ();
 b15zdnd11an1n16x5 FILLER_49_228 ();
 b15zdnd00an1n02x5 FILLER_49_244 ();
 b15zdnd00an1n01x5 FILLER_49_246 ();
 b15zdnd11an1n04x5 FILLER_49_256 ();
 b15zdnd11an1n08x5 FILLER_49_273 ();
 b15zdnd00an1n02x5 FILLER_49_281 ();
 b15zdnd11an1n16x5 FILLER_49_297 ();
 b15zdnd11an1n08x5 FILLER_49_339 ();
 b15zdnd11an1n04x5 FILLER_49_367 ();
 b15zdnd11an1n32x5 FILLER_49_392 ();
 b15zdnd11an1n08x5 FILLER_49_424 ();
 b15zdnd00an1n02x5 FILLER_49_432 ();
 b15zdnd00an1n01x5 FILLER_49_434 ();
 b15zdnd11an1n64x5 FILLER_49_451 ();
 b15zdnd11an1n64x5 FILLER_49_515 ();
 b15zdnd11an1n64x5 FILLER_49_579 ();
 b15zdnd00an1n02x5 FILLER_49_643 ();
 b15zdnd00an1n01x5 FILLER_49_645 ();
 b15zdnd11an1n04x5 FILLER_49_672 ();
 b15zdnd11an1n32x5 FILLER_49_690 ();
 b15zdnd00an1n02x5 FILLER_49_722 ();
 b15zdnd00an1n01x5 FILLER_49_724 ();
 b15zdnd11an1n04x5 FILLER_49_730 ();
 b15zdnd00an1n02x5 FILLER_49_734 ();
 b15zdnd00an1n01x5 FILLER_49_736 ();
 b15zdnd11an1n16x5 FILLER_49_741 ();
 b15zdnd00an1n01x5 FILLER_49_757 ();
 b15zdnd11an1n32x5 FILLER_49_762 ();
 b15zdnd11an1n16x5 FILLER_49_794 ();
 b15zdnd11an1n08x5 FILLER_49_810 ();
 b15zdnd00an1n02x5 FILLER_49_818 ();
 b15zdnd11an1n32x5 FILLER_49_827 ();
 b15zdnd11an1n16x5 FILLER_49_859 ();
 b15zdnd11an1n08x5 FILLER_49_875 ();
 b15zdnd00an1n02x5 FILLER_49_883 ();
 b15zdnd00an1n01x5 FILLER_49_885 ();
 b15zdnd11an1n64x5 FILLER_49_890 ();
 b15zdnd11an1n16x5 FILLER_49_954 ();
 b15zdnd11an1n08x5 FILLER_49_970 ();
 b15zdnd00an1n02x5 FILLER_49_978 ();
 b15zdnd00an1n01x5 FILLER_49_980 ();
 b15zdnd11an1n08x5 FILLER_49_1002 ();
 b15zdnd11an1n04x5 FILLER_49_1025 ();
 b15zdnd11an1n32x5 FILLER_49_1047 ();
 b15zdnd11an1n04x5 FILLER_49_1079 ();
 b15zdnd00an1n02x5 FILLER_49_1083 ();
 b15zdnd11an1n16x5 FILLER_49_1103 ();
 b15zdnd11an1n04x5 FILLER_49_1119 ();
 b15zdnd11an1n32x5 FILLER_49_1154 ();
 b15zdnd11an1n16x5 FILLER_49_1186 ();
 b15zdnd11an1n04x5 FILLER_49_1202 ();
 b15zdnd00an1n02x5 FILLER_49_1206 ();
 b15zdnd00an1n01x5 FILLER_49_1208 ();
 b15zdnd11an1n32x5 FILLER_49_1218 ();
 b15zdnd11an1n16x5 FILLER_49_1250 ();
 b15zdnd11an1n08x5 FILLER_49_1266 ();
 b15zdnd11an1n04x5 FILLER_49_1274 ();
 b15zdnd00an1n02x5 FILLER_49_1278 ();
 b15zdnd00an1n01x5 FILLER_49_1280 ();
 b15zdnd11an1n32x5 FILLER_49_1297 ();
 b15zdnd11an1n16x5 FILLER_49_1329 ();
 b15zdnd00an1n01x5 FILLER_49_1345 ();
 b15zdnd11an1n04x5 FILLER_49_1356 ();
 b15zdnd11an1n32x5 FILLER_49_1367 ();
 b15zdnd11an1n16x5 FILLER_49_1399 ();
 b15zdnd11an1n04x5 FILLER_49_1415 ();
 b15zdnd00an1n02x5 FILLER_49_1419 ();
 b15zdnd11an1n32x5 FILLER_49_1428 ();
 b15zdnd11an1n08x5 FILLER_49_1460 ();
 b15zdnd00an1n02x5 FILLER_49_1468 ();
 b15zdnd00an1n01x5 FILLER_49_1470 ();
 b15zdnd11an1n16x5 FILLER_49_1483 ();
 b15zdnd11an1n08x5 FILLER_49_1499 ();
 b15zdnd11an1n04x5 FILLER_49_1507 ();
 b15zdnd00an1n01x5 FILLER_49_1511 ();
 b15zdnd11an1n08x5 FILLER_49_1519 ();
 b15zdnd11an1n04x5 FILLER_49_1527 ();
 b15zdnd00an1n01x5 FILLER_49_1531 ();
 b15zdnd11an1n04x5 FILLER_49_1546 ();
 b15zdnd00an1n02x5 FILLER_49_1550 ();
 b15zdnd11an1n04x5 FILLER_49_1558 ();
 b15zdnd00an1n01x5 FILLER_49_1562 ();
 b15zdnd11an1n32x5 FILLER_49_1575 ();
 b15zdnd11an1n04x5 FILLER_49_1607 ();
 b15zdnd11an1n04x5 FILLER_49_1625 ();
 b15zdnd00an1n02x5 FILLER_49_1629 ();
 b15zdnd11an1n16x5 FILLER_49_1643 ();
 b15zdnd11an1n04x5 FILLER_49_1659 ();
 b15zdnd00an1n02x5 FILLER_49_1663 ();
 b15zdnd11an1n64x5 FILLER_49_1675 ();
 b15zdnd11an1n08x5 FILLER_49_1739 ();
 b15zdnd11an1n64x5 FILLER_49_1756 ();
 b15zdnd11an1n64x5 FILLER_49_1820 ();
 b15zdnd11an1n64x5 FILLER_49_1884 ();
 b15zdnd11an1n32x5 FILLER_49_1948 ();
 b15zdnd11an1n16x5 FILLER_49_1980 ();
 b15zdnd11an1n08x5 FILLER_49_1996 ();
 b15zdnd11an1n04x5 FILLER_49_2021 ();
 b15zdnd11an1n08x5 FILLER_49_2056 ();
 b15zdnd00an1n01x5 FILLER_49_2064 ();
 b15zdnd11an1n04x5 FILLER_49_2072 ();
 b15zdnd00an1n02x5 FILLER_49_2076 ();
 b15zdnd00an1n01x5 FILLER_49_2078 ();
 b15zdnd11an1n16x5 FILLER_49_2087 ();
 b15zdnd11an1n04x5 FILLER_49_2103 ();
 b15zdnd00an1n02x5 FILLER_49_2107 ();
 b15zdnd00an1n01x5 FILLER_49_2109 ();
 b15zdnd11an1n64x5 FILLER_49_2120 ();
 b15zdnd11an1n08x5 FILLER_49_2184 ();
 b15zdnd00an1n02x5 FILLER_49_2192 ();
 b15zdnd11an1n64x5 FILLER_49_2201 ();
 b15zdnd11an1n16x5 FILLER_49_2265 ();
 b15zdnd00an1n02x5 FILLER_49_2281 ();
 b15zdnd00an1n01x5 FILLER_49_2283 ();
 b15zdnd11an1n64x5 FILLER_50_8 ();
 b15zdnd11an1n04x5 FILLER_50_72 ();
 b15zdnd00an1n02x5 FILLER_50_76 ();
 b15zdnd11an1n32x5 FILLER_50_88 ();
 b15zdnd00an1n02x5 FILLER_50_120 ();
 b15zdnd00an1n01x5 FILLER_50_122 ();
 b15zdnd11an1n32x5 FILLER_50_134 ();
 b15zdnd11an1n16x5 FILLER_50_166 ();
 b15zdnd11an1n08x5 FILLER_50_182 ();
 b15zdnd11an1n04x5 FILLER_50_190 ();
 b15zdnd00an1n02x5 FILLER_50_194 ();
 b15zdnd11an1n04x5 FILLER_50_203 ();
 b15zdnd11an1n04x5 FILLER_50_223 ();
 b15zdnd11an1n16x5 FILLER_50_233 ();
 b15zdnd00an1n02x5 FILLER_50_249 ();
 b15zdnd00an1n01x5 FILLER_50_251 ();
 b15zdnd11an1n04x5 FILLER_50_258 ();
 b15zdnd11an1n64x5 FILLER_50_282 ();
 b15zdnd11an1n08x5 FILLER_50_346 ();
 b15zdnd11an1n04x5 FILLER_50_354 ();
 b15zdnd11an1n04x5 FILLER_50_362 ();
 b15zdnd11an1n32x5 FILLER_50_379 ();
 b15zdnd11an1n16x5 FILLER_50_411 ();
 b15zdnd11an1n08x5 FILLER_50_427 ();
 b15zdnd11an1n04x5 FILLER_50_435 ();
 b15zdnd00an1n02x5 FILLER_50_439 ();
 b15zdnd00an1n01x5 FILLER_50_441 ();
 b15zdnd11an1n32x5 FILLER_50_451 ();
 b15zdnd11an1n16x5 FILLER_50_483 ();
 b15zdnd11an1n08x5 FILLER_50_499 ();
 b15zdnd00an1n02x5 FILLER_50_507 ();
 b15zdnd00an1n01x5 FILLER_50_509 ();
 b15zdnd11an1n32x5 FILLER_50_522 ();
 b15zdnd11an1n16x5 FILLER_50_554 ();
 b15zdnd00an1n02x5 FILLER_50_570 ();
 b15zdnd00an1n01x5 FILLER_50_572 ();
 b15zdnd11an1n08x5 FILLER_50_584 ();
 b15zdnd00an1n01x5 FILLER_50_592 ();
 b15zdnd11an1n04x5 FILLER_50_606 ();
 b15zdnd00an1n02x5 FILLER_50_610 ();
 b15zdnd00an1n01x5 FILLER_50_612 ();
 b15zdnd11an1n08x5 FILLER_50_619 ();
 b15zdnd11an1n04x5 FILLER_50_627 ();
 b15zdnd11an1n04x5 FILLER_50_636 ();
 b15zdnd11an1n08x5 FILLER_50_651 ();
 b15zdnd00an1n02x5 FILLER_50_659 ();
 b15zdnd00an1n01x5 FILLER_50_661 ();
 b15zdnd11an1n16x5 FILLER_50_667 ();
 b15zdnd11an1n08x5 FILLER_50_683 ();
 b15zdnd11an1n04x5 FILLER_50_691 ();
 b15zdnd00an1n02x5 FILLER_50_695 ();
 b15zdnd11an1n08x5 FILLER_50_708 ();
 b15zdnd00an1n02x5 FILLER_50_716 ();
 b15zdnd11an1n32x5 FILLER_50_726 ();
 b15zdnd11an1n16x5 FILLER_50_764 ();
 b15zdnd11an1n08x5 FILLER_50_780 ();
 b15zdnd00an1n01x5 FILLER_50_788 ();
 b15zdnd11an1n16x5 FILLER_50_794 ();
 b15zdnd11an1n08x5 FILLER_50_810 ();
 b15zdnd11an1n04x5 FILLER_50_818 ();
 b15zdnd00an1n01x5 FILLER_50_822 ();
 b15zdnd11an1n08x5 FILLER_50_829 ();
 b15zdnd11an1n04x5 FILLER_50_837 ();
 b15zdnd11an1n08x5 FILLER_50_856 ();
 b15zdnd11an1n04x5 FILLER_50_864 ();
 b15zdnd00an1n02x5 FILLER_50_868 ();
 b15zdnd11an1n64x5 FILLER_50_875 ();
 b15zdnd11an1n64x5 FILLER_50_939 ();
 b15zdnd11an1n64x5 FILLER_50_1003 ();
 b15zdnd11an1n32x5 FILLER_50_1067 ();
 b15zdnd11an1n08x5 FILLER_50_1099 ();
 b15zdnd11an1n64x5 FILLER_50_1138 ();
 b15zdnd11an1n08x5 FILLER_50_1202 ();
 b15zdnd11an1n04x5 FILLER_50_1210 ();
 b15zdnd00an1n01x5 FILLER_50_1214 ();
 b15zdnd11an1n08x5 FILLER_50_1225 ();
 b15zdnd11an1n64x5 FILLER_50_1248 ();
 b15zdnd11an1n16x5 FILLER_50_1312 ();
 b15zdnd11an1n04x5 FILLER_50_1328 ();
 b15zdnd00an1n01x5 FILLER_50_1332 ();
 b15zdnd11an1n04x5 FILLER_50_1340 ();
 b15zdnd11an1n04x5 FILLER_50_1364 ();
 b15zdnd11an1n32x5 FILLER_50_1382 ();
 b15zdnd00an1n02x5 FILLER_50_1414 ();
 b15zdnd11an1n16x5 FILLER_50_1428 ();
 b15zdnd11an1n04x5 FILLER_50_1444 ();
 b15zdnd00an1n01x5 FILLER_50_1448 ();
 b15zdnd11an1n64x5 FILLER_50_1454 ();
 b15zdnd00an1n01x5 FILLER_50_1518 ();
 b15zdnd11an1n64x5 FILLER_50_1529 ();
 b15zdnd11an1n16x5 FILLER_50_1593 ();
 b15zdnd11an1n04x5 FILLER_50_1609 ();
 b15zdnd00an1n02x5 FILLER_50_1613 ();
 b15zdnd00an1n01x5 FILLER_50_1615 ();
 b15zdnd11an1n04x5 FILLER_50_1626 ();
 b15zdnd11an1n16x5 FILLER_50_1642 ();
 b15zdnd11an1n08x5 FILLER_50_1658 ();
 b15zdnd11an1n04x5 FILLER_50_1666 ();
 b15zdnd11an1n32x5 FILLER_50_1696 ();
 b15zdnd11an1n16x5 FILLER_50_1728 ();
 b15zdnd11an1n08x5 FILLER_50_1744 ();
 b15zdnd00an1n01x5 FILLER_50_1752 ();
 b15zdnd11an1n16x5 FILLER_50_1765 ();
 b15zdnd00an1n01x5 FILLER_50_1781 ();
 b15zdnd11an1n16x5 FILLER_50_1787 ();
 b15zdnd00an1n02x5 FILLER_50_1803 ();
 b15zdnd11an1n32x5 FILLER_50_1811 ();
 b15zdnd11an1n16x5 FILLER_50_1852 ();
 b15zdnd11an1n32x5 FILLER_50_1878 ();
 b15zdnd11an1n08x5 FILLER_50_1910 ();
 b15zdnd00an1n01x5 FILLER_50_1918 ();
 b15zdnd11an1n08x5 FILLER_50_1925 ();
 b15zdnd00an1n02x5 FILLER_50_1933 ();
 b15zdnd11an1n64x5 FILLER_50_1949 ();
 b15zdnd11an1n32x5 FILLER_50_2013 ();
 b15zdnd11an1n16x5 FILLER_50_2045 ();
 b15zdnd11an1n08x5 FILLER_50_2061 ();
 b15zdnd11an1n16x5 FILLER_50_2075 ();
 b15zdnd00an1n01x5 FILLER_50_2091 ();
 b15zdnd11an1n04x5 FILLER_50_2108 ();
 b15zdnd11an1n32x5 FILLER_50_2122 ();
 b15zdnd11an1n04x5 FILLER_50_2162 ();
 b15zdnd00an1n02x5 FILLER_50_2166 ();
 b15zdnd11an1n16x5 FILLER_50_2173 ();
 b15zdnd11an1n08x5 FILLER_50_2189 ();
 b15zdnd00an1n01x5 FILLER_50_2197 ();
 b15zdnd11an1n64x5 FILLER_50_2205 ();
 b15zdnd11an1n04x5 FILLER_50_2269 ();
 b15zdnd00an1n02x5 FILLER_50_2273 ();
 b15zdnd00an1n01x5 FILLER_50_2275 ();
 b15zdnd11an1n32x5 FILLER_51_0 ();
 b15zdnd11an1n08x5 FILLER_51_32 ();
 b15zdnd11an1n08x5 FILLER_51_61 ();
 b15zdnd11an1n04x5 FILLER_51_69 ();
 b15zdnd00an1n01x5 FILLER_51_73 ();
 b15zdnd11an1n04x5 FILLER_51_90 ();
 b15zdnd11an1n64x5 FILLER_51_106 ();
 b15zdnd11an1n16x5 FILLER_51_170 ();
 b15zdnd11an1n08x5 FILLER_51_186 ();
 b15zdnd11an1n04x5 FILLER_51_194 ();
 b15zdnd00an1n02x5 FILLER_51_198 ();
 b15zdnd11an1n04x5 FILLER_51_205 ();
 b15zdnd11an1n08x5 FILLER_51_214 ();
 b15zdnd11an1n04x5 FILLER_51_222 ();
 b15zdnd00an1n01x5 FILLER_51_226 ();
 b15zdnd11an1n16x5 FILLER_51_233 ();
 b15zdnd11an1n08x5 FILLER_51_249 ();
 b15zdnd00an1n02x5 FILLER_51_257 ();
 b15zdnd00an1n01x5 FILLER_51_259 ();
 b15zdnd11an1n64x5 FILLER_51_276 ();
 b15zdnd11an1n64x5 FILLER_51_340 ();
 b15zdnd11an1n64x5 FILLER_51_404 ();
 b15zdnd00an1n02x5 FILLER_51_468 ();
 b15zdnd00an1n01x5 FILLER_51_470 ();
 b15zdnd11an1n16x5 FILLER_51_490 ();
 b15zdnd00an1n02x5 FILLER_51_506 ();
 b15zdnd11an1n08x5 FILLER_51_520 ();
 b15zdnd00an1n02x5 FILLER_51_528 ();
 b15zdnd11an1n16x5 FILLER_51_535 ();
 b15zdnd11an1n04x5 FILLER_51_551 ();
 b15zdnd11an1n08x5 FILLER_51_564 ();
 b15zdnd11an1n04x5 FILLER_51_572 ();
 b15zdnd00an1n02x5 FILLER_51_576 ();
 b15zdnd11an1n04x5 FILLER_51_598 ();
 b15zdnd11an1n08x5 FILLER_51_617 ();
 b15zdnd11an1n04x5 FILLER_51_625 ();
 b15zdnd00an1n01x5 FILLER_51_629 ();
 b15zdnd11an1n16x5 FILLER_51_642 ();
 b15zdnd11an1n08x5 FILLER_51_658 ();
 b15zdnd00an1n02x5 FILLER_51_666 ();
 b15zdnd00an1n01x5 FILLER_51_668 ();
 b15zdnd11an1n64x5 FILLER_51_686 ();
 b15zdnd11an1n08x5 FILLER_51_750 ();
 b15zdnd11an1n32x5 FILLER_51_766 ();
 b15zdnd11an1n16x5 FILLER_51_798 ();
 b15zdnd11an1n04x5 FILLER_51_814 ();
 b15zdnd00an1n02x5 FILLER_51_818 ();
 b15zdnd00an1n01x5 FILLER_51_820 ();
 b15zdnd11an1n16x5 FILLER_51_825 ();
 b15zdnd11an1n08x5 FILLER_51_841 ();
 b15zdnd11an1n04x5 FILLER_51_849 ();
 b15zdnd00an1n02x5 FILLER_51_853 ();
 b15zdnd00an1n01x5 FILLER_51_855 ();
 b15zdnd11an1n04x5 FILLER_51_862 ();
 b15zdnd11an1n04x5 FILLER_51_874 ();
 b15zdnd00an1n01x5 FILLER_51_878 ();
 b15zdnd11an1n64x5 FILLER_51_899 ();
 b15zdnd11an1n32x5 FILLER_51_963 ();
 b15zdnd11an1n16x5 FILLER_51_995 ();
 b15zdnd11an1n08x5 FILLER_51_1011 ();
 b15zdnd11an1n04x5 FILLER_51_1019 ();
 b15zdnd11an1n04x5 FILLER_51_1033 ();
 b15zdnd11an1n08x5 FILLER_51_1047 ();
 b15zdnd00an1n01x5 FILLER_51_1055 ();
 b15zdnd11an1n64x5 FILLER_51_1067 ();
 b15zdnd11an1n64x5 FILLER_51_1131 ();
 b15zdnd11an1n16x5 FILLER_51_1195 ();
 b15zdnd11an1n08x5 FILLER_51_1211 ();
 b15zdnd11an1n04x5 FILLER_51_1219 ();
 b15zdnd00an1n01x5 FILLER_51_1223 ();
 b15zdnd11an1n32x5 FILLER_51_1252 ();
 b15zdnd11an1n08x5 FILLER_51_1284 ();
 b15zdnd00an1n02x5 FILLER_51_1292 ();
 b15zdnd11an1n32x5 FILLER_51_1298 ();
 b15zdnd11an1n04x5 FILLER_51_1330 ();
 b15zdnd00an1n02x5 FILLER_51_1334 ();
 b15zdnd11an1n04x5 FILLER_51_1342 ();
 b15zdnd11an1n32x5 FILLER_51_1352 ();
 b15zdnd11an1n16x5 FILLER_51_1384 ();
 b15zdnd00an1n02x5 FILLER_51_1400 ();
 b15zdnd00an1n01x5 FILLER_51_1402 ();
 b15zdnd11an1n64x5 FILLER_51_1412 ();
 b15zdnd11an1n32x5 FILLER_51_1476 ();
 b15zdnd11an1n08x5 FILLER_51_1508 ();
 b15zdnd00an1n02x5 FILLER_51_1516 ();
 b15zdnd11an1n64x5 FILLER_51_1523 ();
 b15zdnd11an1n04x5 FILLER_51_1587 ();
 b15zdnd00an1n01x5 FILLER_51_1591 ();
 b15zdnd11an1n64x5 FILLER_51_1598 ();
 b15zdnd11an1n16x5 FILLER_51_1662 ();
 b15zdnd00an1n01x5 FILLER_51_1678 ();
 b15zdnd11an1n64x5 FILLER_51_1688 ();
 b15zdnd11an1n04x5 FILLER_51_1752 ();
 b15zdnd11an1n04x5 FILLER_51_1772 ();
 b15zdnd11an1n16x5 FILLER_51_1784 ();
 b15zdnd00an1n02x5 FILLER_51_1800 ();
 b15zdnd11an1n64x5 FILLER_51_1811 ();
 b15zdnd00an1n02x5 FILLER_51_1875 ();
 b15zdnd11an1n04x5 FILLER_51_1883 ();
 b15zdnd11an1n16x5 FILLER_51_1902 ();
 b15zdnd11an1n08x5 FILLER_51_1925 ();
 b15zdnd11an1n04x5 FILLER_51_1933 ();
 b15zdnd00an1n02x5 FILLER_51_1937 ();
 b15zdnd00an1n01x5 FILLER_51_1939 ();
 b15zdnd11an1n08x5 FILLER_51_1947 ();
 b15zdnd11an1n04x5 FILLER_51_1955 ();
 b15zdnd00an1n02x5 FILLER_51_1959 ();
 b15zdnd00an1n01x5 FILLER_51_1961 ();
 b15zdnd11an1n08x5 FILLER_51_1968 ();
 b15zdnd00an1n02x5 FILLER_51_1976 ();
 b15zdnd00an1n01x5 FILLER_51_1978 ();
 b15zdnd11an1n32x5 FILLER_51_1986 ();
 b15zdnd11an1n08x5 FILLER_51_2018 ();
 b15zdnd11an1n04x5 FILLER_51_2026 ();
 b15zdnd00an1n02x5 FILLER_51_2030 ();
 b15zdnd11an1n16x5 FILLER_51_2040 ();
 b15zdnd00an1n02x5 FILLER_51_2056 ();
 b15zdnd11an1n64x5 FILLER_51_2063 ();
 b15zdnd00an1n02x5 FILLER_51_2127 ();
 b15zdnd00an1n01x5 FILLER_51_2129 ();
 b15zdnd11an1n04x5 FILLER_51_2140 ();
 b15zdnd00an1n02x5 FILLER_51_2144 ();
 b15zdnd11an1n16x5 FILLER_51_2153 ();
 b15zdnd11an1n08x5 FILLER_51_2175 ();
 b15zdnd11an1n04x5 FILLER_51_2183 ();
 b15zdnd00an1n02x5 FILLER_51_2187 ();
 b15zdnd00an1n01x5 FILLER_51_2189 ();
 b15zdnd11an1n64x5 FILLER_51_2195 ();
 b15zdnd11an1n16x5 FILLER_51_2259 ();
 b15zdnd11an1n08x5 FILLER_51_2275 ();
 b15zdnd00an1n01x5 FILLER_51_2283 ();
 b15zdnd11an1n64x5 FILLER_52_8 ();
 b15zdnd11an1n32x5 FILLER_52_72 ();
 b15zdnd11an1n08x5 FILLER_52_104 ();
 b15zdnd11an1n04x5 FILLER_52_112 ();
 b15zdnd11an1n08x5 FILLER_52_127 ();
 b15zdnd11an1n04x5 FILLER_52_135 ();
 b15zdnd00an1n01x5 FILLER_52_139 ();
 b15zdnd11an1n16x5 FILLER_52_146 ();
 b15zdnd11an1n04x5 FILLER_52_162 ();
 b15zdnd00an1n02x5 FILLER_52_166 ();
 b15zdnd00an1n01x5 FILLER_52_168 ();
 b15zdnd11an1n64x5 FILLER_52_185 ();
 b15zdnd11an1n08x5 FILLER_52_249 ();
 b15zdnd00an1n02x5 FILLER_52_257 ();
 b15zdnd11an1n16x5 FILLER_52_266 ();
 b15zdnd11an1n08x5 FILLER_52_282 ();
 b15zdnd11an1n04x5 FILLER_52_290 ();
 b15zdnd00an1n02x5 FILLER_52_294 ();
 b15zdnd11an1n16x5 FILLER_52_306 ();
 b15zdnd00an1n02x5 FILLER_52_322 ();
 b15zdnd11an1n64x5 FILLER_52_356 ();
 b15zdnd11an1n08x5 FILLER_52_420 ();
 b15zdnd00an1n01x5 FILLER_52_428 ();
 b15zdnd11an1n32x5 FILLER_52_441 ();
 b15zdnd00an1n02x5 FILLER_52_473 ();
 b15zdnd11an1n08x5 FILLER_52_490 ();
 b15zdnd00an1n02x5 FILLER_52_498 ();
 b15zdnd11an1n32x5 FILLER_52_510 ();
 b15zdnd11an1n08x5 FILLER_52_542 ();
 b15zdnd11an1n04x5 FILLER_52_550 ();
 b15zdnd00an1n02x5 FILLER_52_554 ();
 b15zdnd00an1n01x5 FILLER_52_556 ();
 b15zdnd11an1n16x5 FILLER_52_567 ();
 b15zdnd11an1n08x5 FILLER_52_583 ();
 b15zdnd11an1n04x5 FILLER_52_604 ();
 b15zdnd11an1n08x5 FILLER_52_614 ();
 b15zdnd11an1n32x5 FILLER_52_627 ();
 b15zdnd11an1n08x5 FILLER_52_659 ();
 b15zdnd11an1n16x5 FILLER_52_680 ();
 b15zdnd00an1n02x5 FILLER_52_696 ();
 b15zdnd11an1n04x5 FILLER_52_703 ();
 b15zdnd00an1n02x5 FILLER_52_707 ();
 b15zdnd00an1n02x5 FILLER_52_716 ();
 b15zdnd11an1n16x5 FILLER_52_726 ();
 b15zdnd11an1n08x5 FILLER_52_742 ();
 b15zdnd11an1n04x5 FILLER_52_750 ();
 b15zdnd00an1n01x5 FILLER_52_754 ();
 b15zdnd11an1n16x5 FILLER_52_760 ();
 b15zdnd00an1n02x5 FILLER_52_776 ();
 b15zdnd11an1n64x5 FILLER_52_790 ();
 b15zdnd11an1n04x5 FILLER_52_854 ();
 b15zdnd00an1n01x5 FILLER_52_858 ();
 b15zdnd11an1n08x5 FILLER_52_863 ();
 b15zdnd11an1n04x5 FILLER_52_871 ();
 b15zdnd11an1n04x5 FILLER_52_891 ();
 b15zdnd11an1n04x5 FILLER_52_921 ();
 b15zdnd11an1n64x5 FILLER_52_945 ();
 b15zdnd11an1n16x5 FILLER_52_1009 ();
 b15zdnd11an1n08x5 FILLER_52_1025 ();
 b15zdnd11an1n04x5 FILLER_52_1033 ();
 b15zdnd11an1n08x5 FILLER_52_1046 ();
 b15zdnd11an1n04x5 FILLER_52_1054 ();
 b15zdnd00an1n02x5 FILLER_52_1058 ();
 b15zdnd11an1n32x5 FILLER_52_1070 ();
 b15zdnd00an1n02x5 FILLER_52_1102 ();
 b15zdnd00an1n01x5 FILLER_52_1104 ();
 b15zdnd11an1n32x5 FILLER_52_1114 ();
 b15zdnd11an1n04x5 FILLER_52_1146 ();
 b15zdnd00an1n02x5 FILLER_52_1150 ();
 b15zdnd00an1n01x5 FILLER_52_1152 ();
 b15zdnd11an1n08x5 FILLER_52_1162 ();
 b15zdnd11an1n04x5 FILLER_52_1182 ();
 b15zdnd11an1n64x5 FILLER_52_1196 ();
 b15zdnd11an1n32x5 FILLER_52_1260 ();
 b15zdnd11an1n04x5 FILLER_52_1296 ();
 b15zdnd11an1n64x5 FILLER_52_1313 ();
 b15zdnd11an1n04x5 FILLER_52_1377 ();
 b15zdnd00an1n02x5 FILLER_52_1381 ();
 b15zdnd00an1n01x5 FILLER_52_1383 ();
 b15zdnd11an1n64x5 FILLER_52_1389 ();
 b15zdnd11an1n16x5 FILLER_52_1453 ();
 b15zdnd00an1n02x5 FILLER_52_1469 ();
 b15zdnd00an1n01x5 FILLER_52_1471 ();
 b15zdnd11an1n64x5 FILLER_52_1476 ();
 b15zdnd11an1n16x5 FILLER_52_1540 ();
 b15zdnd11an1n08x5 FILLER_52_1556 ();
 b15zdnd11an1n04x5 FILLER_52_1564 ();
 b15zdnd00an1n02x5 FILLER_52_1568 ();
 b15zdnd11an1n08x5 FILLER_52_1579 ();
 b15zdnd11an1n04x5 FILLER_52_1587 ();
 b15zdnd00an1n01x5 FILLER_52_1591 ();
 b15zdnd11an1n64x5 FILLER_52_1596 ();
 b15zdnd11an1n16x5 FILLER_52_1660 ();
 b15zdnd11an1n08x5 FILLER_52_1676 ();
 b15zdnd00an1n01x5 FILLER_52_1684 ();
 b15zdnd11an1n64x5 FILLER_52_1689 ();
 b15zdnd11an1n64x5 FILLER_52_1753 ();
 b15zdnd11an1n04x5 FILLER_52_1817 ();
 b15zdnd00an1n01x5 FILLER_52_1821 ();
 b15zdnd11an1n04x5 FILLER_52_1835 ();
 b15zdnd11an1n04x5 FILLER_52_1857 ();
 b15zdnd11an1n08x5 FILLER_52_1879 ();
 b15zdnd11an1n04x5 FILLER_52_1887 ();
 b15zdnd00an1n02x5 FILLER_52_1891 ();
 b15zdnd00an1n01x5 FILLER_52_1893 ();
 b15zdnd11an1n04x5 FILLER_52_1901 ();
 b15zdnd11an1n64x5 FILLER_52_1917 ();
 b15zdnd11an1n04x5 FILLER_52_1981 ();
 b15zdnd11an1n32x5 FILLER_52_1989 ();
 b15zdnd11an1n08x5 FILLER_52_2021 ();
 b15zdnd00an1n02x5 FILLER_52_2029 ();
 b15zdnd00an1n01x5 FILLER_52_2031 ();
 b15zdnd11an1n08x5 FILLER_52_2047 ();
 b15zdnd00an1n01x5 FILLER_52_2055 ();
 b15zdnd11an1n32x5 FILLER_52_2063 ();
 b15zdnd11an1n08x5 FILLER_52_2095 ();
 b15zdnd00an1n01x5 FILLER_52_2103 ();
 b15zdnd11an1n08x5 FILLER_52_2116 ();
 b15zdnd11an1n04x5 FILLER_52_2124 ();
 b15zdnd00an1n02x5 FILLER_52_2128 ();
 b15zdnd11an1n16x5 FILLER_52_2136 ();
 b15zdnd00an1n02x5 FILLER_52_2152 ();
 b15zdnd11an1n16x5 FILLER_52_2162 ();
 b15zdnd11an1n08x5 FILLER_52_2178 ();
 b15zdnd11an1n04x5 FILLER_52_2186 ();
 b15zdnd11an1n04x5 FILLER_52_2199 ();
 b15zdnd11an1n04x5 FILLER_52_2207 ();
 b15zdnd11an1n32x5 FILLER_52_2221 ();
 b15zdnd11an1n16x5 FILLER_52_2253 ();
 b15zdnd11an1n04x5 FILLER_52_2269 ();
 b15zdnd00an1n02x5 FILLER_52_2273 ();
 b15zdnd00an1n01x5 FILLER_52_2275 ();
 b15zdnd11an1n32x5 FILLER_53_0 ();
 b15zdnd11an1n16x5 FILLER_53_32 ();
 b15zdnd00an1n01x5 FILLER_53_48 ();
 b15zdnd11an1n64x5 FILLER_53_58 ();
 b15zdnd11an1n04x5 FILLER_53_122 ();
 b15zdnd11an1n08x5 FILLER_53_140 ();
 b15zdnd11an1n04x5 FILLER_53_148 ();
 b15zdnd00an1n01x5 FILLER_53_152 ();
 b15zdnd11an1n64x5 FILLER_53_165 ();
 b15zdnd11an1n32x5 FILLER_53_229 ();
 b15zdnd11an1n08x5 FILLER_53_261 ();
 b15zdnd11an1n04x5 FILLER_53_269 ();
 b15zdnd11an1n16x5 FILLER_53_277 ();
 b15zdnd11an1n08x5 FILLER_53_293 ();
 b15zdnd00an1n01x5 FILLER_53_301 ();
 b15zdnd11an1n16x5 FILLER_53_314 ();
 b15zdnd11an1n04x5 FILLER_53_330 ();
 b15zdnd00an1n02x5 FILLER_53_334 ();
 b15zdnd11an1n04x5 FILLER_53_345 ();
 b15zdnd00an1n02x5 FILLER_53_349 ();
 b15zdnd11an1n04x5 FILLER_53_355 ();
 b15zdnd11an1n64x5 FILLER_53_363 ();
 b15zdnd11an1n16x5 FILLER_53_427 ();
 b15zdnd11an1n08x5 FILLER_53_443 ();
 b15zdnd00an1n02x5 FILLER_53_451 ();
 b15zdnd11an1n16x5 FILLER_53_474 ();
 b15zdnd11an1n08x5 FILLER_53_490 ();
 b15zdnd00an1n02x5 FILLER_53_498 ();
 b15zdnd00an1n01x5 FILLER_53_500 ();
 b15zdnd11an1n64x5 FILLER_53_509 ();
 b15zdnd11an1n16x5 FILLER_53_573 ();
 b15zdnd00an1n02x5 FILLER_53_589 ();
 b15zdnd11an1n16x5 FILLER_53_599 ();
 b15zdnd11an1n04x5 FILLER_53_615 ();
 b15zdnd00an1n02x5 FILLER_53_619 ();
 b15zdnd00an1n01x5 FILLER_53_621 ();
 b15zdnd11an1n16x5 FILLER_53_631 ();
 b15zdnd11an1n08x5 FILLER_53_647 ();
 b15zdnd11an1n04x5 FILLER_53_655 ();
 b15zdnd00an1n02x5 FILLER_53_659 ();
 b15zdnd00an1n01x5 FILLER_53_661 ();
 b15zdnd11an1n16x5 FILLER_53_674 ();
 b15zdnd11an1n08x5 FILLER_53_690 ();
 b15zdnd00an1n01x5 FILLER_53_698 ();
 b15zdnd11an1n16x5 FILLER_53_712 ();
 b15zdnd11an1n04x5 FILLER_53_728 ();
 b15zdnd00an1n02x5 FILLER_53_732 ();
 b15zdnd11an1n16x5 FILLER_53_752 ();
 b15zdnd00an1n02x5 FILLER_53_768 ();
 b15zdnd00an1n01x5 FILLER_53_770 ();
 b15zdnd11an1n04x5 FILLER_53_777 ();
 b15zdnd00an1n01x5 FILLER_53_781 ();
 b15zdnd11an1n64x5 FILLER_53_797 ();
 b15zdnd11an1n64x5 FILLER_53_861 ();
 b15zdnd11an1n08x5 FILLER_53_925 ();
 b15zdnd00an1n02x5 FILLER_53_933 ();
 b15zdnd00an1n01x5 FILLER_53_935 ();
 b15zdnd11an1n08x5 FILLER_53_962 ();
 b15zdnd00an1n01x5 FILLER_53_970 ();
 b15zdnd11an1n64x5 FILLER_53_989 ();
 b15zdnd11an1n16x5 FILLER_53_1053 ();
 b15zdnd00an1n02x5 FILLER_53_1069 ();
 b15zdnd11an1n04x5 FILLER_53_1082 ();
 b15zdnd00an1n01x5 FILLER_53_1086 ();
 b15zdnd11an1n04x5 FILLER_53_1096 ();
 b15zdnd11an1n32x5 FILLER_53_1110 ();
 b15zdnd11an1n16x5 FILLER_53_1142 ();
 b15zdnd11an1n08x5 FILLER_53_1158 ();
 b15zdnd11an1n04x5 FILLER_53_1166 ();
 b15zdnd00an1n01x5 FILLER_53_1170 ();
 b15zdnd11an1n64x5 FILLER_53_1191 ();
 b15zdnd11an1n32x5 FILLER_53_1255 ();
 b15zdnd11an1n08x5 FILLER_53_1287 ();
 b15zdnd00an1n01x5 FILLER_53_1295 ();
 b15zdnd11an1n16x5 FILLER_53_1303 ();
 b15zdnd11an1n08x5 FILLER_53_1319 ();
 b15zdnd00an1n02x5 FILLER_53_1327 ();
 b15zdnd11an1n08x5 FILLER_53_1338 ();
 b15zdnd11an1n08x5 FILLER_53_1353 ();
 b15zdnd11an1n04x5 FILLER_53_1361 ();
 b15zdnd11an1n08x5 FILLER_53_1377 ();
 b15zdnd11an1n32x5 FILLER_53_1392 ();
 b15zdnd11an1n04x5 FILLER_53_1424 ();
 b15zdnd00an1n02x5 FILLER_53_1428 ();
 b15zdnd11an1n04x5 FILLER_53_1436 ();
 b15zdnd11an1n16x5 FILLER_53_1465 ();
 b15zdnd11an1n04x5 FILLER_53_1481 ();
 b15zdnd00an1n02x5 FILLER_53_1485 ();
 b15zdnd00an1n01x5 FILLER_53_1487 ();
 b15zdnd11an1n32x5 FILLER_53_1494 ();
 b15zdnd11an1n08x5 FILLER_53_1526 ();
 b15zdnd11an1n04x5 FILLER_53_1534 ();
 b15zdnd00an1n02x5 FILLER_53_1538 ();
 b15zdnd11an1n08x5 FILLER_53_1546 ();
 b15zdnd11an1n04x5 FILLER_53_1554 ();
 b15zdnd00an1n02x5 FILLER_53_1558 ();
 b15zdnd00an1n01x5 FILLER_53_1560 ();
 b15zdnd11an1n04x5 FILLER_53_1581 ();
 b15zdnd11an1n16x5 FILLER_53_1605 ();
 b15zdnd00an1n02x5 FILLER_53_1621 ();
 b15zdnd11an1n32x5 FILLER_53_1628 ();
 b15zdnd11an1n16x5 FILLER_53_1660 ();
 b15zdnd11an1n04x5 FILLER_53_1676 ();
 b15zdnd00an1n02x5 FILLER_53_1680 ();
 b15zdnd11an1n64x5 FILLER_53_1694 ();
 b15zdnd11an1n64x5 FILLER_53_1758 ();
 b15zdnd11an1n08x5 FILLER_53_1822 ();
 b15zdnd00an1n02x5 FILLER_53_1830 ();
 b15zdnd11an1n32x5 FILLER_53_1838 ();
 b15zdnd11an1n08x5 FILLER_53_1870 ();
 b15zdnd11an1n04x5 FILLER_53_1878 ();
 b15zdnd00an1n01x5 FILLER_53_1882 ();
 b15zdnd11an1n64x5 FILLER_53_1893 ();
 b15zdnd11an1n16x5 FILLER_53_1957 ();
 b15zdnd11an1n04x5 FILLER_53_1973 ();
 b15zdnd00an1n02x5 FILLER_53_1977 ();
 b15zdnd11an1n04x5 FILLER_53_1986 ();
 b15zdnd00an1n01x5 FILLER_53_1990 ();
 b15zdnd11an1n32x5 FILLER_53_2001 ();
 b15zdnd00an1n02x5 FILLER_53_2033 ();
 b15zdnd11an1n04x5 FILLER_53_2047 ();
 b15zdnd11an1n04x5 FILLER_53_2057 ();
 b15zdnd00an1n02x5 FILLER_53_2061 ();
 b15zdnd11an1n32x5 FILLER_53_2079 ();
 b15zdnd11an1n04x5 FILLER_53_2111 ();
 b15zdnd00an1n02x5 FILLER_53_2115 ();
 b15zdnd00an1n01x5 FILLER_53_2117 ();
 b15zdnd11an1n64x5 FILLER_53_2133 ();
 b15zdnd11an1n64x5 FILLER_53_2197 ();
 b15zdnd11an1n16x5 FILLER_53_2261 ();
 b15zdnd11an1n04x5 FILLER_53_2277 ();
 b15zdnd00an1n02x5 FILLER_53_2281 ();
 b15zdnd00an1n01x5 FILLER_53_2283 ();
 b15zdnd11an1n32x5 FILLER_54_8 ();
 b15zdnd11an1n16x5 FILLER_54_40 ();
 b15zdnd00an1n02x5 FILLER_54_56 ();
 b15zdnd11an1n32x5 FILLER_54_62 ();
 b15zdnd11an1n16x5 FILLER_54_94 ();
 b15zdnd11an1n04x5 FILLER_54_110 ();
 b15zdnd00an1n02x5 FILLER_54_114 ();
 b15zdnd11an1n32x5 FILLER_54_121 ();
 b15zdnd11an1n16x5 FILLER_54_153 ();
 b15zdnd11an1n08x5 FILLER_54_169 ();
 b15zdnd11an1n04x5 FILLER_54_177 ();
 b15zdnd00an1n02x5 FILLER_54_181 ();
 b15zdnd00an1n01x5 FILLER_54_183 ();
 b15zdnd11an1n04x5 FILLER_54_189 ();
 b15zdnd11an1n32x5 FILLER_54_207 ();
 b15zdnd11an1n16x5 FILLER_54_239 ();
 b15zdnd11an1n04x5 FILLER_54_255 ();
 b15zdnd11an1n32x5 FILLER_54_273 ();
 b15zdnd11an1n16x5 FILLER_54_305 ();
 b15zdnd11an1n08x5 FILLER_54_321 ();
 b15zdnd00an1n02x5 FILLER_54_329 ();
 b15zdnd00an1n01x5 FILLER_54_331 ();
 b15zdnd11an1n64x5 FILLER_54_345 ();
 b15zdnd11an1n16x5 FILLER_54_409 ();
 b15zdnd11an1n04x5 FILLER_54_425 ();
 b15zdnd00an1n02x5 FILLER_54_429 ();
 b15zdnd00an1n01x5 FILLER_54_431 ();
 b15zdnd11an1n08x5 FILLER_54_440 ();
 b15zdnd00an1n02x5 FILLER_54_448 ();
 b15zdnd11an1n64x5 FILLER_54_469 ();
 b15zdnd11an1n16x5 FILLER_54_533 ();
 b15zdnd11an1n04x5 FILLER_54_549 ();
 b15zdnd00an1n02x5 FILLER_54_553 ();
 b15zdnd00an1n01x5 FILLER_54_555 ();
 b15zdnd11an1n64x5 FILLER_54_580 ();
 b15zdnd11an1n64x5 FILLER_54_644 ();
 b15zdnd11an1n08x5 FILLER_54_708 ();
 b15zdnd00an1n02x5 FILLER_54_716 ();
 b15zdnd11an1n16x5 FILLER_54_726 ();
 b15zdnd11an1n08x5 FILLER_54_742 ();
 b15zdnd11an1n32x5 FILLER_54_766 ();
 b15zdnd11an1n04x5 FILLER_54_798 ();
 b15zdnd00an1n01x5 FILLER_54_802 ();
 b15zdnd11an1n32x5 FILLER_54_811 ();
 b15zdnd11an1n16x5 FILLER_54_843 ();
 b15zdnd11an1n04x5 FILLER_54_859 ();
 b15zdnd00an1n02x5 FILLER_54_863 ();
 b15zdnd00an1n01x5 FILLER_54_865 ();
 b15zdnd11an1n32x5 FILLER_54_872 ();
 b15zdnd11an1n08x5 FILLER_54_904 ();
 b15zdnd11an1n04x5 FILLER_54_912 ();
 b15zdnd11an1n16x5 FILLER_54_942 ();
 b15zdnd11an1n08x5 FILLER_54_958 ();
 b15zdnd00an1n02x5 FILLER_54_966 ();
 b15zdnd11an1n16x5 FILLER_54_978 ();
 b15zdnd11an1n04x5 FILLER_54_994 ();
 b15zdnd00an1n02x5 FILLER_54_998 ();
 b15zdnd11an1n04x5 FILLER_54_1026 ();
 b15zdnd11an1n64x5 FILLER_54_1045 ();
 b15zdnd11an1n32x5 FILLER_54_1109 ();
 b15zdnd11an1n08x5 FILLER_54_1141 ();
 b15zdnd11an1n04x5 FILLER_54_1149 ();
 b15zdnd11an1n16x5 FILLER_54_1171 ();
 b15zdnd11an1n04x5 FILLER_54_1187 ();
 b15zdnd00an1n01x5 FILLER_54_1191 ();
 b15zdnd11an1n04x5 FILLER_54_1217 ();
 b15zdnd11an1n64x5 FILLER_54_1246 ();
 b15zdnd11an1n08x5 FILLER_54_1310 ();
 b15zdnd11an1n04x5 FILLER_54_1318 ();
 b15zdnd00an1n02x5 FILLER_54_1322 ();
 b15zdnd11an1n08x5 FILLER_54_1339 ();
 b15zdnd00an1n02x5 FILLER_54_1347 ();
 b15zdnd11an1n08x5 FILLER_54_1356 ();
 b15zdnd11an1n04x5 FILLER_54_1364 ();
 b15zdnd00an1n02x5 FILLER_54_1368 ();
 b15zdnd11an1n32x5 FILLER_54_1401 ();
 b15zdnd11an1n04x5 FILLER_54_1441 ();
 b15zdnd11an1n08x5 FILLER_54_1449 ();
 b15zdnd00an1n02x5 FILLER_54_1457 ();
 b15zdnd11an1n04x5 FILLER_54_1471 ();
 b15zdnd11an1n04x5 FILLER_54_1481 ();
 b15zdnd00an1n01x5 FILLER_54_1485 ();
 b15zdnd11an1n64x5 FILLER_54_1499 ();
 b15zdnd11an1n08x5 FILLER_54_1563 ();
 b15zdnd00an1n02x5 FILLER_54_1571 ();
 b15zdnd11an1n08x5 FILLER_54_1584 ();
 b15zdnd11an1n08x5 FILLER_54_1598 ();
 b15zdnd00an1n01x5 FILLER_54_1606 ();
 b15zdnd11an1n08x5 FILLER_54_1612 ();
 b15zdnd00an1n02x5 FILLER_54_1620 ();
 b15zdnd11an1n08x5 FILLER_54_1634 ();
 b15zdnd11an1n04x5 FILLER_54_1642 ();
 b15zdnd00an1n02x5 FILLER_54_1646 ();
 b15zdnd00an1n01x5 FILLER_54_1648 ();
 b15zdnd11an1n16x5 FILLER_54_1656 ();
 b15zdnd11an1n04x5 FILLER_54_1672 ();
 b15zdnd00an1n01x5 FILLER_54_1676 ();
 b15zdnd11an1n64x5 FILLER_54_1683 ();
 b15zdnd11an1n16x5 FILLER_54_1747 ();
 b15zdnd11an1n04x5 FILLER_54_1763 ();
 b15zdnd00an1n02x5 FILLER_54_1767 ();
 b15zdnd11an1n64x5 FILLER_54_1777 ();
 b15zdnd11an1n64x5 FILLER_54_1841 ();
 b15zdnd11an1n64x5 FILLER_54_1905 ();
 b15zdnd11an1n64x5 FILLER_54_1969 ();
 b15zdnd11an1n16x5 FILLER_54_2033 ();
 b15zdnd00an1n02x5 FILLER_54_2049 ();
 b15zdnd11an1n32x5 FILLER_54_2055 ();
 b15zdnd11an1n08x5 FILLER_54_2087 ();
 b15zdnd11an1n04x5 FILLER_54_2095 ();
 b15zdnd00an1n02x5 FILLER_54_2099 ();
 b15zdnd11an1n16x5 FILLER_54_2106 ();
 b15zdnd11an1n08x5 FILLER_54_2122 ();
 b15zdnd00an1n02x5 FILLER_54_2152 ();
 b15zdnd11an1n64x5 FILLER_54_2162 ();
 b15zdnd11an1n32x5 FILLER_54_2226 ();
 b15zdnd11an1n16x5 FILLER_54_2258 ();
 b15zdnd00an1n02x5 FILLER_54_2274 ();
 b15zdnd11an1n32x5 FILLER_55_0 ();
 b15zdnd11an1n04x5 FILLER_55_32 ();
 b15zdnd00an1n01x5 FILLER_55_36 ();
 b15zdnd11an1n04x5 FILLER_55_46 ();
 b15zdnd11an1n32x5 FILLER_55_64 ();
 b15zdnd11an1n08x5 FILLER_55_106 ();
 b15zdnd11an1n04x5 FILLER_55_114 ();
 b15zdnd00an1n01x5 FILLER_55_118 ();
 b15zdnd11an1n04x5 FILLER_55_131 ();
 b15zdnd11an1n32x5 FILLER_55_161 ();
 b15zdnd11an1n08x5 FILLER_55_193 ();
 b15zdnd11an1n16x5 FILLER_55_207 ();
 b15zdnd11an1n04x5 FILLER_55_223 ();
 b15zdnd00an1n02x5 FILLER_55_227 ();
 b15zdnd00an1n01x5 FILLER_55_229 ();
 b15zdnd11an1n04x5 FILLER_55_234 ();
 b15zdnd11an1n08x5 FILLER_55_247 ();
 b15zdnd11an1n04x5 FILLER_55_255 ();
 b15zdnd11an1n16x5 FILLER_55_264 ();
 b15zdnd00an1n02x5 FILLER_55_280 ();
 b15zdnd00an1n01x5 FILLER_55_282 ();
 b15zdnd11an1n08x5 FILLER_55_299 ();
 b15zdnd11an1n04x5 FILLER_55_307 ();
 b15zdnd11an1n16x5 FILLER_55_319 ();
 b15zdnd11an1n04x5 FILLER_55_335 ();
 b15zdnd11an1n64x5 FILLER_55_347 ();
 b15zdnd11an1n16x5 FILLER_55_411 ();
 b15zdnd11an1n08x5 FILLER_55_427 ();
 b15zdnd11an1n04x5 FILLER_55_435 ();
 b15zdnd11an1n32x5 FILLER_55_449 ();
 b15zdnd11an1n08x5 FILLER_55_481 ();
 b15zdnd00an1n02x5 FILLER_55_489 ();
 b15zdnd11an1n64x5 FILLER_55_507 ();
 b15zdnd11an1n16x5 FILLER_55_571 ();
 b15zdnd11an1n08x5 FILLER_55_587 ();
 b15zdnd11an1n04x5 FILLER_55_595 ();
 b15zdnd00an1n02x5 FILLER_55_599 ();
 b15zdnd11an1n64x5 FILLER_55_606 ();
 b15zdnd11an1n64x5 FILLER_55_670 ();
 b15zdnd11an1n04x5 FILLER_55_734 ();
 b15zdnd00an1n02x5 FILLER_55_738 ();
 b15zdnd00an1n01x5 FILLER_55_740 ();
 b15zdnd11an1n04x5 FILLER_55_750 ();
 b15zdnd11an1n08x5 FILLER_55_758 ();
 b15zdnd11an1n04x5 FILLER_55_766 ();
 b15zdnd00an1n02x5 FILLER_55_770 ();
 b15zdnd11an1n08x5 FILLER_55_792 ();
 b15zdnd11an1n04x5 FILLER_55_800 ();
 b15zdnd00an1n01x5 FILLER_55_804 ();
 b15zdnd11an1n16x5 FILLER_55_809 ();
 b15zdnd00an1n02x5 FILLER_55_825 ();
 b15zdnd00an1n01x5 FILLER_55_827 ();
 b15zdnd11an1n08x5 FILLER_55_833 ();
 b15zdnd00an1n01x5 FILLER_55_841 ();
 b15zdnd11an1n04x5 FILLER_55_848 ();
 b15zdnd11an1n32x5 FILLER_55_857 ();
 b15zdnd11an1n04x5 FILLER_55_889 ();
 b15zdnd00an1n02x5 FILLER_55_893 ();
 b15zdnd00an1n01x5 FILLER_55_895 ();
 b15zdnd11an1n16x5 FILLER_55_919 ();
 b15zdnd11an1n08x5 FILLER_55_935 ();
 b15zdnd11an1n04x5 FILLER_55_943 ();
 b15zdnd00an1n02x5 FILLER_55_947 ();
 b15zdnd00an1n01x5 FILLER_55_949 ();
 b15zdnd11an1n64x5 FILLER_55_968 ();
 b15zdnd11an1n32x5 FILLER_55_1032 ();
 b15zdnd11an1n16x5 FILLER_55_1064 ();
 b15zdnd00an1n02x5 FILLER_55_1080 ();
 b15zdnd00an1n01x5 FILLER_55_1082 ();
 b15zdnd11an1n64x5 FILLER_55_1106 ();
 b15zdnd11an1n64x5 FILLER_55_1170 ();
 b15zdnd11an1n64x5 FILLER_55_1234 ();
 b15zdnd00an1n01x5 FILLER_55_1298 ();
 b15zdnd11an1n04x5 FILLER_55_1310 ();
 b15zdnd00an1n02x5 FILLER_55_1314 ();
 b15zdnd11an1n08x5 FILLER_55_1322 ();
 b15zdnd00an1n01x5 FILLER_55_1330 ();
 b15zdnd11an1n64x5 FILLER_55_1337 ();
 b15zdnd11an1n16x5 FILLER_55_1401 ();
 b15zdnd11an1n08x5 FILLER_55_1417 ();
 b15zdnd00an1n02x5 FILLER_55_1425 ();
 b15zdnd11an1n08x5 FILLER_55_1434 ();
 b15zdnd11an1n04x5 FILLER_55_1442 ();
 b15zdnd00an1n01x5 FILLER_55_1446 ();
 b15zdnd11an1n32x5 FILLER_55_1453 ();
 b15zdnd11an1n08x5 FILLER_55_1485 ();
 b15zdnd00an1n01x5 FILLER_55_1493 ();
 b15zdnd11an1n08x5 FILLER_55_1507 ();
 b15zdnd11an1n04x5 FILLER_55_1515 ();
 b15zdnd11an1n04x5 FILLER_55_1529 ();
 b15zdnd11an1n32x5 FILLER_55_1548 ();
 b15zdnd00an1n01x5 FILLER_55_1580 ();
 b15zdnd11an1n16x5 FILLER_55_1586 ();
 b15zdnd11an1n08x5 FILLER_55_1602 ();
 b15zdnd00an1n01x5 FILLER_55_1610 ();
 b15zdnd11an1n16x5 FILLER_55_1632 ();
 b15zdnd11an1n04x5 FILLER_55_1648 ();
 b15zdnd11an1n64x5 FILLER_55_1656 ();
 b15zdnd11an1n16x5 FILLER_55_1720 ();
 b15zdnd11an1n08x5 FILLER_55_1736 ();
 b15zdnd00an1n02x5 FILLER_55_1744 ();
 b15zdnd11an1n16x5 FILLER_55_1756 ();
 b15zdnd00an1n02x5 FILLER_55_1772 ();
 b15zdnd00an1n01x5 FILLER_55_1774 ();
 b15zdnd11an1n64x5 FILLER_55_1781 ();
 b15zdnd11an1n64x5 FILLER_55_1845 ();
 b15zdnd11an1n08x5 FILLER_55_1909 ();
 b15zdnd11an1n04x5 FILLER_55_1924 ();
 b15zdnd00an1n02x5 FILLER_55_1928 ();
 b15zdnd00an1n01x5 FILLER_55_1930 ();
 b15zdnd11an1n64x5 FILLER_55_1945 ();
 b15zdnd11an1n64x5 FILLER_55_2009 ();
 b15zdnd11an1n08x5 FILLER_55_2073 ();
 b15zdnd11an1n04x5 FILLER_55_2081 ();
 b15zdnd11an1n64x5 FILLER_55_2095 ();
 b15zdnd11an1n16x5 FILLER_55_2159 ();
 b15zdnd11an1n08x5 FILLER_55_2175 ();
 b15zdnd11an1n04x5 FILLER_55_2183 ();
 b15zdnd00an1n01x5 FILLER_55_2187 ();
 b15zdnd11an1n04x5 FILLER_55_2193 ();
 b15zdnd00an1n01x5 FILLER_55_2197 ();
 b15zdnd11an1n64x5 FILLER_55_2203 ();
 b15zdnd11an1n16x5 FILLER_55_2267 ();
 b15zdnd00an1n01x5 FILLER_55_2283 ();
 b15zdnd11an1n64x5 FILLER_56_8 ();
 b15zdnd11an1n16x5 FILLER_56_72 ();
 b15zdnd11an1n04x5 FILLER_56_88 ();
 b15zdnd00an1n01x5 FILLER_56_92 ();
 b15zdnd11an1n16x5 FILLER_56_107 ();
 b15zdnd00an1n02x5 FILLER_56_123 ();
 b15zdnd00an1n01x5 FILLER_56_125 ();
 b15zdnd11an1n04x5 FILLER_56_132 ();
 b15zdnd11an1n32x5 FILLER_56_160 ();
 b15zdnd11an1n08x5 FILLER_56_192 ();
 b15zdnd00an1n02x5 FILLER_56_200 ();
 b15zdnd00an1n01x5 FILLER_56_202 ();
 b15zdnd11an1n16x5 FILLER_56_209 ();
 b15zdnd11an1n32x5 FILLER_56_253 ();
 b15zdnd11an1n16x5 FILLER_56_285 ();
 b15zdnd11an1n04x5 FILLER_56_306 ();
 b15zdnd00an1n01x5 FILLER_56_310 ();
 b15zdnd11an1n04x5 FILLER_56_315 ();
 b15zdnd00an1n01x5 FILLER_56_319 ();
 b15zdnd11an1n04x5 FILLER_56_332 ();
 b15zdnd11an1n04x5 FILLER_56_348 ();
 b15zdnd11an1n04x5 FILLER_56_358 ();
 b15zdnd11an1n64x5 FILLER_56_366 ();
 b15zdnd11an1n32x5 FILLER_56_430 ();
 b15zdnd11an1n16x5 FILLER_56_462 ();
 b15zdnd11an1n08x5 FILLER_56_478 ();
 b15zdnd11an1n04x5 FILLER_56_486 ();
 b15zdnd00an1n02x5 FILLER_56_490 ();
 b15zdnd00an1n01x5 FILLER_56_492 ();
 b15zdnd11an1n64x5 FILLER_56_507 ();
 b15zdnd00an1n02x5 FILLER_56_571 ();
 b15zdnd11an1n08x5 FILLER_56_582 ();
 b15zdnd11an1n04x5 FILLER_56_590 ();
 b15zdnd00an1n01x5 FILLER_56_594 ();
 b15zdnd11an1n08x5 FILLER_56_608 ();
 b15zdnd11an1n04x5 FILLER_56_616 ();
 b15zdnd11an1n04x5 FILLER_56_626 ();
 b15zdnd11an1n04x5 FILLER_56_638 ();
 b15zdnd11an1n32x5 FILLER_56_651 ();
 b15zdnd11an1n08x5 FILLER_56_683 ();
 b15zdnd11an1n04x5 FILLER_56_691 ();
 b15zdnd00an1n01x5 FILLER_56_695 ();
 b15zdnd00an1n02x5 FILLER_56_716 ();
 b15zdnd11an1n16x5 FILLER_56_726 ();
 b15zdnd11an1n08x5 FILLER_56_742 ();
 b15zdnd11an1n04x5 FILLER_56_750 ();
 b15zdnd00an1n02x5 FILLER_56_754 ();
 b15zdnd00an1n01x5 FILLER_56_756 ();
 b15zdnd11an1n64x5 FILLER_56_763 ();
 b15zdnd11an1n08x5 FILLER_56_827 ();
 b15zdnd00an1n02x5 FILLER_56_835 ();
 b15zdnd00an1n01x5 FILLER_56_837 ();
 b15zdnd11an1n04x5 FILLER_56_843 ();
 b15zdnd11an1n04x5 FILLER_56_856 ();
 b15zdnd11an1n64x5 FILLER_56_866 ();
 b15zdnd11an1n16x5 FILLER_56_930 ();
 b15zdnd11an1n04x5 FILLER_56_946 ();
 b15zdnd11an1n64x5 FILLER_56_962 ();
 b15zdnd11an1n04x5 FILLER_56_1026 ();
 b15zdnd00an1n02x5 FILLER_56_1030 ();
 b15zdnd11an1n08x5 FILLER_56_1063 ();
 b15zdnd00an1n02x5 FILLER_56_1071 ();
 b15zdnd00an1n01x5 FILLER_56_1073 ();
 b15zdnd11an1n64x5 FILLER_56_1099 ();
 b15zdnd11an1n08x5 FILLER_56_1163 ();
 b15zdnd11an1n04x5 FILLER_56_1171 ();
 b15zdnd00an1n02x5 FILLER_56_1175 ();
 b15zdnd11an1n04x5 FILLER_56_1203 ();
 b15zdnd11an1n64x5 FILLER_56_1216 ();
 b15zdnd11an1n32x5 FILLER_56_1280 ();
 b15zdnd11an1n08x5 FILLER_56_1312 ();
 b15zdnd11an1n16x5 FILLER_56_1327 ();
 b15zdnd11an1n08x5 FILLER_56_1343 ();
 b15zdnd11an1n04x5 FILLER_56_1351 ();
 b15zdnd00an1n02x5 FILLER_56_1355 ();
 b15zdnd11an1n64x5 FILLER_56_1363 ();
 b15zdnd11an1n08x5 FILLER_56_1436 ();
 b15zdnd11an1n04x5 FILLER_56_1444 ();
 b15zdnd00an1n02x5 FILLER_56_1448 ();
 b15zdnd00an1n01x5 FILLER_56_1450 ();
 b15zdnd11an1n32x5 FILLER_56_1482 ();
 b15zdnd11an1n08x5 FILLER_56_1514 ();
 b15zdnd11an1n04x5 FILLER_56_1522 ();
 b15zdnd11an1n32x5 FILLER_56_1535 ();
 b15zdnd11an1n16x5 FILLER_56_1567 ();
 b15zdnd11an1n08x5 FILLER_56_1583 ();
 b15zdnd00an1n02x5 FILLER_56_1591 ();
 b15zdnd00an1n01x5 FILLER_56_1593 ();
 b15zdnd11an1n64x5 FILLER_56_1599 ();
 b15zdnd11an1n64x5 FILLER_56_1663 ();
 b15zdnd11an1n08x5 FILLER_56_1727 ();
 b15zdnd00an1n02x5 FILLER_56_1735 ();
 b15zdnd00an1n01x5 FILLER_56_1737 ();
 b15zdnd11an1n04x5 FILLER_56_1745 ();
 b15zdnd11an1n08x5 FILLER_56_1756 ();
 b15zdnd11an1n04x5 FILLER_56_1764 ();
 b15zdnd00an1n02x5 FILLER_56_1768 ();
 b15zdnd00an1n01x5 FILLER_56_1770 ();
 b15zdnd11an1n16x5 FILLER_56_1780 ();
 b15zdnd11an1n08x5 FILLER_56_1796 ();
 b15zdnd11an1n32x5 FILLER_56_1813 ();
 b15zdnd11an1n08x5 FILLER_56_1845 ();
 b15zdnd11an1n04x5 FILLER_56_1853 ();
 b15zdnd00an1n01x5 FILLER_56_1857 ();
 b15zdnd11an1n04x5 FILLER_56_1865 ();
 b15zdnd11an1n32x5 FILLER_56_1873 ();
 b15zdnd11an1n08x5 FILLER_56_1905 ();
 b15zdnd11an1n04x5 FILLER_56_1913 ();
 b15zdnd00an1n02x5 FILLER_56_1917 ();
 b15zdnd11an1n04x5 FILLER_56_1923 ();
 b15zdnd11an1n16x5 FILLER_56_1938 ();
 b15zdnd11an1n04x5 FILLER_56_1954 ();
 b15zdnd00an1n02x5 FILLER_56_1958 ();
 b15zdnd11an1n32x5 FILLER_56_1972 ();
 b15zdnd11an1n16x5 FILLER_56_2004 ();
 b15zdnd00an1n02x5 FILLER_56_2020 ();
 b15zdnd11an1n64x5 FILLER_56_2035 ();
 b15zdnd11an1n16x5 FILLER_56_2099 ();
 b15zdnd00an1n02x5 FILLER_56_2115 ();
 b15zdnd11an1n16x5 FILLER_56_2137 ();
 b15zdnd00an1n01x5 FILLER_56_2153 ();
 b15zdnd11an1n16x5 FILLER_56_2162 ();
 b15zdnd11an1n08x5 FILLER_56_2178 ();
 b15zdnd00an1n02x5 FILLER_56_2186 ();
 b15zdnd00an1n01x5 FILLER_56_2188 ();
 b15zdnd11an1n64x5 FILLER_56_2196 ();
 b15zdnd11an1n16x5 FILLER_56_2260 ();
 b15zdnd11an1n64x5 FILLER_57_0 ();
 b15zdnd11an1n08x5 FILLER_57_64 ();
 b15zdnd11an1n04x5 FILLER_57_72 ();
 b15zdnd00an1n02x5 FILLER_57_76 ();
 b15zdnd00an1n01x5 FILLER_57_78 ();
 b15zdnd11an1n64x5 FILLER_57_102 ();
 b15zdnd00an1n01x5 FILLER_57_166 ();
 b15zdnd11an1n16x5 FILLER_57_177 ();
 b15zdnd00an1n02x5 FILLER_57_193 ();
 b15zdnd11an1n16x5 FILLER_57_205 ();
 b15zdnd11an1n08x5 FILLER_57_221 ();
 b15zdnd00an1n02x5 FILLER_57_229 ();
 b15zdnd00an1n01x5 FILLER_57_231 ();
 b15zdnd11an1n64x5 FILLER_57_240 ();
 b15zdnd11an1n64x5 FILLER_57_304 ();
 b15zdnd11an1n64x5 FILLER_57_368 ();
 b15zdnd11an1n32x5 FILLER_57_432 ();
 b15zdnd00an1n02x5 FILLER_57_464 ();
 b15zdnd00an1n01x5 FILLER_57_466 ();
 b15zdnd11an1n08x5 FILLER_57_480 ();
 b15zdnd00an1n01x5 FILLER_57_488 ();
 b15zdnd11an1n04x5 FILLER_57_498 ();
 b15zdnd11an1n16x5 FILLER_57_510 ();
 b15zdnd11an1n04x5 FILLER_57_526 ();
 b15zdnd11an1n16x5 FILLER_57_546 ();
 b15zdnd11an1n04x5 FILLER_57_577 ();
 b15zdnd11an1n08x5 FILLER_57_586 ();
 b15zdnd11an1n16x5 FILLER_57_599 ();
 b15zdnd11an1n08x5 FILLER_57_615 ();
 b15zdnd11an1n04x5 FILLER_57_623 ();
 b15zdnd00an1n02x5 FILLER_57_627 ();
 b15zdnd00an1n01x5 FILLER_57_629 ();
 b15zdnd11an1n16x5 FILLER_57_638 ();
 b15zdnd11an1n08x5 FILLER_57_654 ();
 b15zdnd11an1n04x5 FILLER_57_662 ();
 b15zdnd00an1n02x5 FILLER_57_666 ();
 b15zdnd11an1n16x5 FILLER_57_674 ();
 b15zdnd11an1n64x5 FILLER_57_695 ();
 b15zdnd11an1n32x5 FILLER_57_759 ();
 b15zdnd00an1n02x5 FILLER_57_791 ();
 b15zdnd00an1n01x5 FILLER_57_793 ();
 b15zdnd11an1n32x5 FILLER_57_806 ();
 b15zdnd11an1n16x5 FILLER_57_838 ();
 b15zdnd11an1n32x5 FILLER_57_860 ();
 b15zdnd11an1n04x5 FILLER_57_892 ();
 b15zdnd11an1n32x5 FILLER_57_927 ();
 b15zdnd11an1n16x5 FILLER_57_959 ();
 b15zdnd11an1n08x5 FILLER_57_975 ();
 b15zdnd11an1n04x5 FILLER_57_983 ();
 b15zdnd00an1n02x5 FILLER_57_987 ();
 b15zdnd00an1n01x5 FILLER_57_989 ();
 b15zdnd11an1n64x5 FILLER_57_1047 ();
 b15zdnd11an1n16x5 FILLER_57_1111 ();
 b15zdnd11an1n08x5 FILLER_57_1127 ();
 b15zdnd11an1n32x5 FILLER_57_1150 ();
 b15zdnd11an1n16x5 FILLER_57_1182 ();
 b15zdnd11an1n08x5 FILLER_57_1198 ();
 b15zdnd00an1n02x5 FILLER_57_1206 ();
 b15zdnd00an1n01x5 FILLER_57_1208 ();
 b15zdnd11an1n32x5 FILLER_57_1230 ();
 b15zdnd00an1n01x5 FILLER_57_1262 ();
 b15zdnd11an1n04x5 FILLER_57_1294 ();
 b15zdnd00an1n01x5 FILLER_57_1298 ();
 b15zdnd11an1n32x5 FILLER_57_1303 ();
 b15zdnd11an1n16x5 FILLER_57_1335 ();
 b15zdnd11an1n08x5 FILLER_57_1351 ();
 b15zdnd00an1n02x5 FILLER_57_1359 ();
 b15zdnd11an1n04x5 FILLER_57_1368 ();
 b15zdnd11an1n64x5 FILLER_57_1378 ();
 b15zdnd11an1n64x5 FILLER_57_1442 ();
 b15zdnd11an1n32x5 FILLER_57_1506 ();
 b15zdnd00an1n02x5 FILLER_57_1538 ();
 b15zdnd11an1n32x5 FILLER_57_1544 ();
 b15zdnd11an1n16x5 FILLER_57_1576 ();
 b15zdnd11an1n64x5 FILLER_57_1602 ();
 b15zdnd11an1n64x5 FILLER_57_1666 ();
 b15zdnd11an1n64x5 FILLER_57_1730 ();
 b15zdnd00an1n02x5 FILLER_57_1794 ();
 b15zdnd00an1n01x5 FILLER_57_1796 ();
 b15zdnd11an1n04x5 FILLER_57_1812 ();
 b15zdnd11an1n08x5 FILLER_57_1826 ();
 b15zdnd11an1n04x5 FILLER_57_1840 ();
 b15zdnd11an1n16x5 FILLER_57_1869 ();
 b15zdnd11an1n04x5 FILLER_57_1885 ();
 b15zdnd00an1n02x5 FILLER_57_1889 ();
 b15zdnd11an1n64x5 FILLER_57_1896 ();
 b15zdnd00an1n02x5 FILLER_57_1960 ();
 b15zdnd11an1n04x5 FILLER_57_1967 ();
 b15zdnd11an1n32x5 FILLER_57_1975 ();
 b15zdnd11an1n08x5 FILLER_57_2007 ();
 b15zdnd11an1n04x5 FILLER_57_2015 ();
 b15zdnd00an1n02x5 FILLER_57_2019 ();
 b15zdnd00an1n01x5 FILLER_57_2021 ();
 b15zdnd11an1n16x5 FILLER_57_2029 ();
 b15zdnd11an1n08x5 FILLER_57_2045 ();
 b15zdnd00an1n02x5 FILLER_57_2053 ();
 b15zdnd11an1n04x5 FILLER_57_2059 ();
 b15zdnd11an1n16x5 FILLER_57_2069 ();
 b15zdnd00an1n01x5 FILLER_57_2085 ();
 b15zdnd11an1n04x5 FILLER_57_2101 ();
 b15zdnd11an1n08x5 FILLER_57_2110 ();
 b15zdnd00an1n01x5 FILLER_57_2118 ();
 b15zdnd11an1n08x5 FILLER_57_2127 ();
 b15zdnd00an1n02x5 FILLER_57_2135 ();
 b15zdnd00an1n01x5 FILLER_57_2137 ();
 b15zdnd11an1n04x5 FILLER_57_2150 ();
 b15zdnd11an1n08x5 FILLER_57_2176 ();
 b15zdnd00an1n02x5 FILLER_57_2184 ();
 b15zdnd00an1n01x5 FILLER_57_2186 ();
 b15zdnd11an1n64x5 FILLER_57_2203 ();
 b15zdnd11an1n16x5 FILLER_57_2267 ();
 b15zdnd00an1n01x5 FILLER_57_2283 ();
 b15zdnd11an1n32x5 FILLER_58_8 ();
 b15zdnd11an1n04x5 FILLER_58_40 ();
 b15zdnd00an1n01x5 FILLER_58_44 ();
 b15zdnd11an1n04x5 FILLER_58_49 ();
 b15zdnd00an1n02x5 FILLER_58_53 ();
 b15zdnd11an1n32x5 FILLER_58_65 ();
 b15zdnd11an1n16x5 FILLER_58_97 ();
 b15zdnd00an1n02x5 FILLER_58_113 ();
 b15zdnd11an1n32x5 FILLER_58_120 ();
 b15zdnd11an1n16x5 FILLER_58_152 ();
 b15zdnd00an1n01x5 FILLER_58_168 ();
 b15zdnd11an1n16x5 FILLER_58_174 ();
 b15zdnd11an1n08x5 FILLER_58_190 ();
 b15zdnd00an1n01x5 FILLER_58_198 ();
 b15zdnd11an1n16x5 FILLER_58_209 ();
 b15zdnd11an1n08x5 FILLER_58_225 ();
 b15zdnd00an1n02x5 FILLER_58_233 ();
 b15zdnd00an1n01x5 FILLER_58_235 ();
 b15zdnd11an1n64x5 FILLER_58_255 ();
 b15zdnd11an1n64x5 FILLER_58_319 ();
 b15zdnd11an1n32x5 FILLER_58_383 ();
 b15zdnd11an1n08x5 FILLER_58_415 ();
 b15zdnd11an1n08x5 FILLER_58_439 ();
 b15zdnd11an1n04x5 FILLER_58_447 ();
 b15zdnd11an1n16x5 FILLER_58_459 ();
 b15zdnd11an1n04x5 FILLER_58_475 ();
 b15zdnd00an1n01x5 FILLER_58_479 ();
 b15zdnd11an1n32x5 FILLER_58_486 ();
 b15zdnd11an1n16x5 FILLER_58_518 ();
 b15zdnd11an1n08x5 FILLER_58_534 ();
 b15zdnd00an1n01x5 FILLER_58_542 ();
 b15zdnd11an1n16x5 FILLER_58_552 ();
 b15zdnd00an1n02x5 FILLER_58_568 ();
 b15zdnd11an1n04x5 FILLER_58_586 ();
 b15zdnd11an1n64x5 FILLER_58_604 ();
 b15zdnd11an1n08x5 FILLER_58_668 ();
 b15zdnd11an1n04x5 FILLER_58_676 ();
 b15zdnd00an1n02x5 FILLER_58_680 ();
 b15zdnd11an1n04x5 FILLER_58_694 ();
 b15zdnd00an1n02x5 FILLER_58_698 ();
 b15zdnd00an1n01x5 FILLER_58_700 ();
 b15zdnd00an1n02x5 FILLER_58_715 ();
 b15zdnd00an1n01x5 FILLER_58_717 ();
 b15zdnd11an1n08x5 FILLER_58_726 ();
 b15zdnd11an1n04x5 FILLER_58_734 ();
 b15zdnd00an1n02x5 FILLER_58_738 ();
 b15zdnd11an1n64x5 FILLER_58_748 ();
 b15zdnd11an1n32x5 FILLER_58_812 ();
 b15zdnd11an1n08x5 FILLER_58_844 ();
 b15zdnd11an1n32x5 FILLER_58_858 ();
 b15zdnd11an1n08x5 FILLER_58_890 ();
 b15zdnd00an1n02x5 FILLER_58_898 ();
 b15zdnd00an1n01x5 FILLER_58_900 ();
 b15zdnd11an1n64x5 FILLER_58_905 ();
 b15zdnd11an1n04x5 FILLER_58_969 ();
 b15zdnd00an1n02x5 FILLER_58_973 ();
 b15zdnd00an1n01x5 FILLER_58_975 ();
 b15zdnd11an1n04x5 FILLER_58_980 ();
 b15zdnd11an1n04x5 FILLER_58_1006 ();
 b15zdnd11an1n64x5 FILLER_58_1036 ();
 b15zdnd00an1n02x5 FILLER_58_1100 ();
 b15zdnd00an1n01x5 FILLER_58_1102 ();
 b15zdnd11an1n04x5 FILLER_58_1134 ();
 b15zdnd11an1n16x5 FILLER_58_1157 ();
 b15zdnd11an1n08x5 FILLER_58_1173 ();
 b15zdnd11an1n04x5 FILLER_58_1199 ();
 b15zdnd11an1n64x5 FILLER_58_1213 ();
 b15zdnd11an1n16x5 FILLER_58_1277 ();
 b15zdnd00an1n01x5 FILLER_58_1293 ();
 b15zdnd11an1n32x5 FILLER_58_1305 ();
 b15zdnd11an1n08x5 FILLER_58_1337 ();
 b15zdnd11an1n04x5 FILLER_58_1345 ();
 b15zdnd11an1n04x5 FILLER_58_1354 ();
 b15zdnd11an1n04x5 FILLER_58_1363 ();
 b15zdnd00an1n02x5 FILLER_58_1367 ();
 b15zdnd11an1n16x5 FILLER_58_1382 ();
 b15zdnd11an1n04x5 FILLER_58_1398 ();
 b15zdnd00an1n02x5 FILLER_58_1402 ();
 b15zdnd11an1n32x5 FILLER_58_1410 ();
 b15zdnd11an1n16x5 FILLER_58_1442 ();
 b15zdnd11an1n08x5 FILLER_58_1458 ();
 b15zdnd11an1n04x5 FILLER_58_1466 ();
 b15zdnd00an1n01x5 FILLER_58_1470 ();
 b15zdnd11an1n08x5 FILLER_58_1477 ();
 b15zdnd11an1n64x5 FILLER_58_1495 ();
 b15zdnd11an1n16x5 FILLER_58_1559 ();
 b15zdnd00an1n01x5 FILLER_58_1575 ();
 b15zdnd11an1n04x5 FILLER_58_1590 ();
 b15zdnd11an1n32x5 FILLER_58_1599 ();
 b15zdnd11an1n04x5 FILLER_58_1631 ();
 b15zdnd00an1n02x5 FILLER_58_1635 ();
 b15zdnd11an1n16x5 FILLER_58_1650 ();
 b15zdnd11an1n08x5 FILLER_58_1666 ();
 b15zdnd00an1n01x5 FILLER_58_1674 ();
 b15zdnd11an1n16x5 FILLER_58_1682 ();
 b15zdnd11an1n04x5 FILLER_58_1698 ();
 b15zdnd00an1n02x5 FILLER_58_1702 ();
 b15zdnd11an1n64x5 FILLER_58_1722 ();
 b15zdnd11an1n04x5 FILLER_58_1786 ();
 b15zdnd00an1n02x5 FILLER_58_1790 ();
 b15zdnd00an1n01x5 FILLER_58_1792 ();
 b15zdnd11an1n04x5 FILLER_58_1799 ();
 b15zdnd11an1n04x5 FILLER_58_1829 ();
 b15zdnd11an1n08x5 FILLER_58_1839 ();
 b15zdnd11an1n04x5 FILLER_58_1847 ();
 b15zdnd00an1n02x5 FILLER_58_1851 ();
 b15zdnd00an1n01x5 FILLER_58_1853 ();
 b15zdnd11an1n32x5 FILLER_58_1861 ();
 b15zdnd00an1n01x5 FILLER_58_1893 ();
 b15zdnd11an1n16x5 FILLER_58_1899 ();
 b15zdnd11an1n08x5 FILLER_58_1915 ();
 b15zdnd11an1n04x5 FILLER_58_1923 ();
 b15zdnd00an1n02x5 FILLER_58_1927 ();
 b15zdnd00an1n01x5 FILLER_58_1929 ();
 b15zdnd11an1n32x5 FILLER_58_1936 ();
 b15zdnd11an1n16x5 FILLER_58_1973 ();
 b15zdnd00an1n01x5 FILLER_58_1989 ();
 b15zdnd11an1n04x5 FILLER_58_1996 ();
 b15zdnd11an1n32x5 FILLER_58_2012 ();
 b15zdnd00an1n01x5 FILLER_58_2044 ();
 b15zdnd11an1n04x5 FILLER_58_2050 ();
 b15zdnd00an1n02x5 FILLER_58_2054 ();
 b15zdnd00an1n01x5 FILLER_58_2056 ();
 b15zdnd11an1n16x5 FILLER_58_2063 ();
 b15zdnd11an1n04x5 FILLER_58_2079 ();
 b15zdnd00an1n02x5 FILLER_58_2083 ();
 b15zdnd11an1n08x5 FILLER_58_2095 ();
 b15zdnd00an1n01x5 FILLER_58_2103 ();
 b15zdnd11an1n16x5 FILLER_58_2110 ();
 b15zdnd11an1n08x5 FILLER_58_2126 ();
 b15zdnd00an1n01x5 FILLER_58_2134 ();
 b15zdnd11an1n04x5 FILLER_58_2148 ();
 b15zdnd00an1n02x5 FILLER_58_2152 ();
 b15zdnd11an1n64x5 FILLER_58_2162 ();
 b15zdnd11an1n32x5 FILLER_58_2226 ();
 b15zdnd11an1n16x5 FILLER_58_2258 ();
 b15zdnd00an1n02x5 FILLER_58_2274 ();
 b15zdnd11an1n16x5 FILLER_59_0 ();
 b15zdnd11an1n08x5 FILLER_59_16 ();
 b15zdnd11an1n04x5 FILLER_59_24 ();
 b15zdnd00an1n02x5 FILLER_59_28 ();
 b15zdnd11an1n04x5 FILLER_59_42 ();
 b15zdnd11an1n16x5 FILLER_59_56 ();
 b15zdnd11an1n08x5 FILLER_59_72 ();
 b15zdnd00an1n02x5 FILLER_59_80 ();
 b15zdnd11an1n16x5 FILLER_59_92 ();
 b15zdnd11an1n08x5 FILLER_59_108 ();
 b15zdnd11an1n04x5 FILLER_59_123 ();
 b15zdnd11an1n16x5 FILLER_59_132 ();
 b15zdnd11an1n08x5 FILLER_59_148 ();
 b15zdnd11an1n04x5 FILLER_59_156 ();
 b15zdnd00an1n02x5 FILLER_59_160 ();
 b15zdnd00an1n01x5 FILLER_59_162 ();
 b15zdnd11an1n04x5 FILLER_59_170 ();
 b15zdnd11an1n04x5 FILLER_59_184 ();
 b15zdnd00an1n02x5 FILLER_59_188 ();
 b15zdnd11an1n32x5 FILLER_59_204 ();
 b15zdnd11an1n08x5 FILLER_59_236 ();
 b15zdnd11an1n04x5 FILLER_59_256 ();
 b15zdnd11an1n04x5 FILLER_59_281 ();
 b15zdnd11an1n04x5 FILLER_59_294 ();
 b15zdnd11an1n32x5 FILLER_59_311 ();
 b15zdnd00an1n02x5 FILLER_59_343 ();
 b15zdnd00an1n01x5 FILLER_59_345 ();
 b15zdnd11an1n08x5 FILLER_59_356 ();
 b15zdnd11an1n64x5 FILLER_59_371 ();
 b15zdnd11an1n04x5 FILLER_59_435 ();
 b15zdnd11an1n04x5 FILLER_59_444 ();
 b15zdnd11an1n04x5 FILLER_59_455 ();
 b15zdnd00an1n02x5 FILLER_59_459 ();
 b15zdnd00an1n01x5 FILLER_59_461 ();
 b15zdnd11an1n04x5 FILLER_59_476 ();
 b15zdnd11an1n04x5 FILLER_59_486 ();
 b15zdnd11an1n32x5 FILLER_59_503 ();
 b15zdnd11an1n04x5 FILLER_59_535 ();
 b15zdnd00an1n01x5 FILLER_59_539 ();
 b15zdnd11an1n64x5 FILLER_59_547 ();
 b15zdnd11an1n16x5 FILLER_59_611 ();
 b15zdnd00an1n02x5 FILLER_59_627 ();
 b15zdnd11an1n16x5 FILLER_59_641 ();
 b15zdnd11an1n08x5 FILLER_59_657 ();
 b15zdnd11an1n04x5 FILLER_59_665 ();
 b15zdnd00an1n01x5 FILLER_59_669 ();
 b15zdnd11an1n04x5 FILLER_59_679 ();
 b15zdnd11an1n16x5 FILLER_59_694 ();
 b15zdnd11an1n04x5 FILLER_59_710 ();
 b15zdnd11an1n08x5 FILLER_59_724 ();
 b15zdnd00an1n02x5 FILLER_59_732 ();
 b15zdnd11an1n16x5 FILLER_59_741 ();
 b15zdnd11an1n04x5 FILLER_59_757 ();
 b15zdnd00an1n01x5 FILLER_59_761 ();
 b15zdnd11an1n08x5 FILLER_59_778 ();
 b15zdnd00an1n02x5 FILLER_59_786 ();
 b15zdnd11an1n64x5 FILLER_59_802 ();
 b15zdnd11an1n64x5 FILLER_59_866 ();
 b15zdnd11an1n16x5 FILLER_59_930 ();
 b15zdnd11an1n08x5 FILLER_59_946 ();
 b15zdnd11an1n04x5 FILLER_59_954 ();
 b15zdnd00an1n02x5 FILLER_59_958 ();
 b15zdnd11an1n04x5 FILLER_59_969 ();
 b15zdnd11an1n64x5 FILLER_59_978 ();
 b15zdnd11an1n64x5 FILLER_59_1042 ();
 b15zdnd11an1n64x5 FILLER_59_1106 ();
 b15zdnd11an1n64x5 FILLER_59_1170 ();
 b15zdnd11an1n64x5 FILLER_59_1234 ();
 b15zdnd11an1n64x5 FILLER_59_1298 ();
 b15zdnd11an1n32x5 FILLER_59_1362 ();
 b15zdnd11an1n04x5 FILLER_59_1394 ();
 b15zdnd00an1n02x5 FILLER_59_1398 ();
 b15zdnd11an1n16x5 FILLER_59_1406 ();
 b15zdnd11an1n08x5 FILLER_59_1422 ();
 b15zdnd11an1n04x5 FILLER_59_1430 ();
 b15zdnd11an1n32x5 FILLER_59_1450 ();
 b15zdnd00an1n02x5 FILLER_59_1482 ();
 b15zdnd00an1n01x5 FILLER_59_1484 ();
 b15zdnd11an1n08x5 FILLER_59_1492 ();
 b15zdnd00an1n02x5 FILLER_59_1500 ();
 b15zdnd00an1n01x5 FILLER_59_1502 ();
 b15zdnd11an1n08x5 FILLER_59_1507 ();
 b15zdnd11an1n04x5 FILLER_59_1515 ();
 b15zdnd11an1n32x5 FILLER_59_1531 ();
 b15zdnd00an1n02x5 FILLER_59_1563 ();
 b15zdnd11an1n64x5 FILLER_59_1580 ();
 b15zdnd11an1n04x5 FILLER_59_1644 ();
 b15zdnd00an1n02x5 FILLER_59_1648 ();
 b15zdnd11an1n08x5 FILLER_59_1670 ();
 b15zdnd11an1n04x5 FILLER_59_1683 ();
 b15zdnd11an1n64x5 FILLER_59_1691 ();
 b15zdnd11an1n16x5 FILLER_59_1755 ();
 b15zdnd00an1n02x5 FILLER_59_1771 ();
 b15zdnd11an1n32x5 FILLER_59_1779 ();
 b15zdnd11an1n16x5 FILLER_59_1811 ();
 b15zdnd11an1n08x5 FILLER_59_1827 ();
 b15zdnd00an1n01x5 FILLER_59_1835 ();
 b15zdnd11an1n04x5 FILLER_59_1847 ();
 b15zdnd11an1n08x5 FILLER_59_1861 ();
 b15zdnd11an1n04x5 FILLER_59_1869 ();
 b15zdnd00an1n02x5 FILLER_59_1873 ();
 b15zdnd11an1n08x5 FILLER_59_1881 ();
 b15zdnd11an1n04x5 FILLER_59_1889 ();
 b15zdnd00an1n01x5 FILLER_59_1893 ();
 b15zdnd11an1n16x5 FILLER_59_1901 ();
 b15zdnd11an1n08x5 FILLER_59_1917 ();
 b15zdnd00an1n02x5 FILLER_59_1925 ();
 b15zdnd00an1n01x5 FILLER_59_1927 ();
 b15zdnd11an1n32x5 FILLER_59_1935 ();
 b15zdnd11an1n32x5 FILLER_59_1978 ();
 b15zdnd11an1n08x5 FILLER_59_2010 ();
 b15zdnd11an1n04x5 FILLER_59_2018 ();
 b15zdnd00an1n02x5 FILLER_59_2022 ();
 b15zdnd11an1n08x5 FILLER_59_2029 ();
 b15zdnd00an1n02x5 FILLER_59_2037 ();
 b15zdnd00an1n01x5 FILLER_59_2039 ();
 b15zdnd11an1n04x5 FILLER_59_2052 ();
 b15zdnd11an1n64x5 FILLER_59_2068 ();
 b15zdnd11an1n64x5 FILLER_59_2132 ();
 b15zdnd11an1n64x5 FILLER_59_2196 ();
 b15zdnd11an1n16x5 FILLER_59_2260 ();
 b15zdnd11an1n08x5 FILLER_59_2276 ();
 b15zdnd11an1n32x5 FILLER_60_8 ();
 b15zdnd11an1n16x5 FILLER_60_40 ();
 b15zdnd11an1n04x5 FILLER_60_56 ();
 b15zdnd00an1n01x5 FILLER_60_60 ();
 b15zdnd11an1n08x5 FILLER_60_65 ();
 b15zdnd11an1n04x5 FILLER_60_73 ();
 b15zdnd00an1n02x5 FILLER_60_77 ();
 b15zdnd11an1n08x5 FILLER_60_89 ();
 b15zdnd11an1n04x5 FILLER_60_97 ();
 b15zdnd00an1n01x5 FILLER_60_101 ();
 b15zdnd11an1n04x5 FILLER_60_107 ();
 b15zdnd00an1n02x5 FILLER_60_111 ();
 b15zdnd11an1n08x5 FILLER_60_128 ();
 b15zdnd11an1n04x5 FILLER_60_148 ();
 b15zdnd11an1n32x5 FILLER_60_161 ();
 b15zdnd00an1n01x5 FILLER_60_193 ();
 b15zdnd11an1n16x5 FILLER_60_198 ();
 b15zdnd11an1n08x5 FILLER_60_214 ();
 b15zdnd11an1n04x5 FILLER_60_222 ();
 b15zdnd11an1n08x5 FILLER_60_233 ();
 b15zdnd11an1n04x5 FILLER_60_241 ();
 b15zdnd00an1n02x5 FILLER_60_245 ();
 b15zdnd11an1n32x5 FILLER_60_256 ();
 b15zdnd11an1n16x5 FILLER_60_288 ();
 b15zdnd11an1n04x5 FILLER_60_304 ();
 b15zdnd00an1n01x5 FILLER_60_308 ();
 b15zdnd11an1n16x5 FILLER_60_324 ();
 b15zdnd11an1n04x5 FILLER_60_344 ();
 b15zdnd11an1n08x5 FILLER_60_354 ();
 b15zdnd00an1n02x5 FILLER_60_362 ();
 b15zdnd00an1n01x5 FILLER_60_364 ();
 b15zdnd11an1n08x5 FILLER_60_372 ();
 b15zdnd11an1n04x5 FILLER_60_380 ();
 b15zdnd11an1n64x5 FILLER_60_403 ();
 b15zdnd11an1n32x5 FILLER_60_467 ();
 b15zdnd11an1n16x5 FILLER_60_499 ();
 b15zdnd11an1n08x5 FILLER_60_515 ();
 b15zdnd11an1n04x5 FILLER_60_523 ();
 b15zdnd00an1n02x5 FILLER_60_527 ();
 b15zdnd11an1n64x5 FILLER_60_550 ();
 b15zdnd11an1n32x5 FILLER_60_614 ();
 b15zdnd11an1n16x5 FILLER_60_646 ();
 b15zdnd11an1n04x5 FILLER_60_662 ();
 b15zdnd11an1n16x5 FILLER_60_671 ();
 b15zdnd11an1n08x5 FILLER_60_687 ();
 b15zdnd11an1n04x5 FILLER_60_695 ();
 b15zdnd00an1n01x5 FILLER_60_699 ();
 b15zdnd00an1n02x5 FILLER_60_716 ();
 b15zdnd11an1n08x5 FILLER_60_726 ();
 b15zdnd11an1n16x5 FILLER_60_739 ();
 b15zdnd11an1n08x5 FILLER_60_755 ();
 b15zdnd00an1n02x5 FILLER_60_763 ();
 b15zdnd00an1n01x5 FILLER_60_765 ();
 b15zdnd11an1n04x5 FILLER_60_770 ();
 b15zdnd11an1n04x5 FILLER_60_780 ();
 b15zdnd11an1n16x5 FILLER_60_790 ();
 b15zdnd11an1n04x5 FILLER_60_806 ();
 b15zdnd11an1n32x5 FILLER_60_826 ();
 b15zdnd11an1n16x5 FILLER_60_890 ();
 b15zdnd00an1n01x5 FILLER_60_906 ();
 b15zdnd11an1n04x5 FILLER_60_912 ();
 b15zdnd11an1n32x5 FILLER_60_936 ();
 b15zdnd11an1n16x5 FILLER_60_968 ();
 b15zdnd00an1n01x5 FILLER_60_984 ();
 b15zdnd11an1n64x5 FILLER_60_994 ();
 b15zdnd11an1n64x5 FILLER_60_1058 ();
 b15zdnd11an1n64x5 FILLER_60_1122 ();
 b15zdnd11an1n08x5 FILLER_60_1186 ();
 b15zdnd11an1n32x5 FILLER_60_1214 ();
 b15zdnd11an1n08x5 FILLER_60_1246 ();
 b15zdnd00an1n01x5 FILLER_60_1254 ();
 b15zdnd11an1n04x5 FILLER_60_1286 ();
 b15zdnd11an1n16x5 FILLER_60_1297 ();
 b15zdnd11an1n08x5 FILLER_60_1313 ();
 b15zdnd00an1n02x5 FILLER_60_1321 ();
 b15zdnd00an1n01x5 FILLER_60_1323 ();
 b15zdnd11an1n16x5 FILLER_60_1339 ();
 b15zdnd11an1n08x5 FILLER_60_1355 ();
 b15zdnd11an1n04x5 FILLER_60_1363 ();
 b15zdnd11an1n16x5 FILLER_60_1379 ();
 b15zdnd11an1n08x5 FILLER_60_1395 ();
 b15zdnd00an1n02x5 FILLER_60_1403 ();
 b15zdnd00an1n01x5 FILLER_60_1405 ();
 b15zdnd11an1n08x5 FILLER_60_1412 ();
 b15zdnd00an1n01x5 FILLER_60_1420 ();
 b15zdnd11an1n04x5 FILLER_60_1429 ();
 b15zdnd11an1n08x5 FILLER_60_1438 ();
 b15zdnd00an1n01x5 FILLER_60_1446 ();
 b15zdnd11an1n16x5 FILLER_60_1459 ();
 b15zdnd11an1n08x5 FILLER_60_1475 ();
 b15zdnd00an1n01x5 FILLER_60_1483 ();
 b15zdnd11an1n32x5 FILLER_60_1490 ();
 b15zdnd00an1n02x5 FILLER_60_1522 ();
 b15zdnd11an1n08x5 FILLER_60_1530 ();
 b15zdnd11an1n04x5 FILLER_60_1538 ();
 b15zdnd00an1n01x5 FILLER_60_1542 ();
 b15zdnd11an1n32x5 FILLER_60_1553 ();
 b15zdnd11an1n08x5 FILLER_60_1585 ();
 b15zdnd00an1n02x5 FILLER_60_1593 ();
 b15zdnd00an1n01x5 FILLER_60_1595 ();
 b15zdnd11an1n04x5 FILLER_60_1607 ();
 b15zdnd11an1n32x5 FILLER_60_1617 ();
 b15zdnd00an1n02x5 FILLER_60_1649 ();
 b15zdnd00an1n01x5 FILLER_60_1651 ();
 b15zdnd11an1n08x5 FILLER_60_1662 ();
 b15zdnd11an1n64x5 FILLER_60_1674 ();
 b15zdnd11an1n64x5 FILLER_60_1738 ();
 b15zdnd11an1n64x5 FILLER_60_1802 ();
 b15zdnd11an1n16x5 FILLER_60_1866 ();
 b15zdnd11an1n08x5 FILLER_60_1882 ();
 b15zdnd00an1n01x5 FILLER_60_1890 ();
 b15zdnd11an1n32x5 FILLER_60_1896 ();
 b15zdnd11an1n64x5 FILLER_60_1933 ();
 b15zdnd11an1n64x5 FILLER_60_1997 ();
 b15zdnd11an1n32x5 FILLER_60_2061 ();
 b15zdnd11an1n16x5 FILLER_60_2093 ();
 b15zdnd11an1n08x5 FILLER_60_2109 ();
 b15zdnd11an1n04x5 FILLER_60_2117 ();
 b15zdnd00an1n01x5 FILLER_60_2121 ();
 b15zdnd11an1n16x5 FILLER_60_2127 ();
 b15zdnd11an1n08x5 FILLER_60_2143 ();
 b15zdnd00an1n02x5 FILLER_60_2151 ();
 b15zdnd00an1n01x5 FILLER_60_2153 ();
 b15zdnd11an1n64x5 FILLER_60_2162 ();
 b15zdnd11an1n32x5 FILLER_60_2226 ();
 b15zdnd11an1n16x5 FILLER_60_2258 ();
 b15zdnd00an1n02x5 FILLER_60_2274 ();
 b15zdnd11an1n32x5 FILLER_61_0 ();
 b15zdnd11an1n08x5 FILLER_61_32 ();
 b15zdnd11an1n04x5 FILLER_61_40 ();
 b15zdnd00an1n02x5 FILLER_61_44 ();
 b15zdnd00an1n01x5 FILLER_61_46 ();
 b15zdnd11an1n16x5 FILLER_61_52 ();
 b15zdnd00an1n02x5 FILLER_61_68 ();
 b15zdnd00an1n01x5 FILLER_61_70 ();
 b15zdnd11an1n08x5 FILLER_61_76 ();
 b15zdnd00an1n01x5 FILLER_61_84 ();
 b15zdnd11an1n64x5 FILLER_61_90 ();
 b15zdnd11an1n16x5 FILLER_61_154 ();
 b15zdnd11an1n04x5 FILLER_61_170 ();
 b15zdnd00an1n02x5 FILLER_61_174 ();
 b15zdnd00an1n01x5 FILLER_61_176 ();
 b15zdnd11an1n16x5 FILLER_61_186 ();
 b15zdnd11an1n08x5 FILLER_61_202 ();
 b15zdnd11an1n04x5 FILLER_61_210 ();
 b15zdnd00an1n02x5 FILLER_61_214 ();
 b15zdnd11an1n64x5 FILLER_61_228 ();
 b15zdnd11an1n32x5 FILLER_61_292 ();
 b15zdnd00an1n02x5 FILLER_61_324 ();
 b15zdnd00an1n01x5 FILLER_61_326 ();
 b15zdnd11an1n64x5 FILLER_61_340 ();
 b15zdnd11an1n32x5 FILLER_61_404 ();
 b15zdnd11an1n16x5 FILLER_61_436 ();
 b15zdnd11an1n08x5 FILLER_61_452 ();
 b15zdnd00an1n02x5 FILLER_61_460 ();
 b15zdnd00an1n01x5 FILLER_61_462 ();
 b15zdnd11an1n16x5 FILLER_61_477 ();
 b15zdnd11an1n04x5 FILLER_61_493 ();
 b15zdnd11an1n04x5 FILLER_61_503 ();
 b15zdnd11an1n32x5 FILLER_61_516 ();
 b15zdnd11an1n08x5 FILLER_61_548 ();
 b15zdnd00an1n02x5 FILLER_61_556 ();
 b15zdnd00an1n01x5 FILLER_61_558 ();
 b15zdnd11an1n32x5 FILLER_61_565 ();
 b15zdnd11an1n16x5 FILLER_61_597 ();
 b15zdnd00an1n01x5 FILLER_61_613 ();
 b15zdnd11an1n32x5 FILLER_61_618 ();
 b15zdnd11an1n16x5 FILLER_61_650 ();
 b15zdnd11an1n64x5 FILLER_61_671 ();
 b15zdnd11an1n64x5 FILLER_61_735 ();
 b15zdnd11an1n04x5 FILLER_61_799 ();
 b15zdnd00an1n02x5 FILLER_61_803 ();
 b15zdnd11an1n04x5 FILLER_61_810 ();
 b15zdnd11an1n32x5 FILLER_61_819 ();
 b15zdnd11an1n04x5 FILLER_61_882 ();
 b15zdnd11an1n32x5 FILLER_61_918 ();
 b15zdnd11an1n16x5 FILLER_61_950 ();
 b15zdnd11an1n08x5 FILLER_61_966 ();
 b15zdnd11an1n04x5 FILLER_61_974 ();
 b15zdnd11an1n16x5 FILLER_61_998 ();
 b15zdnd11an1n08x5 FILLER_61_1014 ();
 b15zdnd11an1n08x5 FILLER_61_1047 ();
 b15zdnd11an1n08x5 FILLER_61_1081 ();
 b15zdnd00an1n02x5 FILLER_61_1089 ();
 b15zdnd11an1n16x5 FILLER_61_1104 ();
 b15zdnd00an1n02x5 FILLER_61_1120 ();
 b15zdnd00an1n01x5 FILLER_61_1122 ();
 b15zdnd11an1n16x5 FILLER_61_1154 ();
 b15zdnd11an1n04x5 FILLER_61_1170 ();
 b15zdnd00an1n02x5 FILLER_61_1174 ();
 b15zdnd00an1n01x5 FILLER_61_1176 ();
 b15zdnd11an1n04x5 FILLER_61_1202 ();
 b15zdnd11an1n32x5 FILLER_61_1230 ();
 b15zdnd11an1n16x5 FILLER_61_1262 ();
 b15zdnd11an1n08x5 FILLER_61_1278 ();
 b15zdnd11an1n04x5 FILLER_61_1291 ();
 b15zdnd11an1n04x5 FILLER_61_1306 ();
 b15zdnd00an1n02x5 FILLER_61_1310 ();
 b15zdnd11an1n08x5 FILLER_61_1316 ();
 b15zdnd00an1n01x5 FILLER_61_1324 ();
 b15zdnd11an1n04x5 FILLER_61_1341 ();
 b15zdnd11an1n16x5 FILLER_61_1351 ();
 b15zdnd11an1n08x5 FILLER_61_1367 ();
 b15zdnd11an1n32x5 FILLER_61_1400 ();
 b15zdnd11an1n04x5 FILLER_61_1432 ();
 b15zdnd00an1n02x5 FILLER_61_1436 ();
 b15zdnd00an1n01x5 FILLER_61_1438 ();
 b15zdnd11an1n32x5 FILLER_61_1451 ();
 b15zdnd11an1n16x5 FILLER_61_1483 ();
 b15zdnd11an1n08x5 FILLER_61_1499 ();
 b15zdnd11an1n04x5 FILLER_61_1507 ();
 b15zdnd00an1n02x5 FILLER_61_1511 ();
 b15zdnd00an1n01x5 FILLER_61_1513 ();
 b15zdnd11an1n16x5 FILLER_61_1520 ();
 b15zdnd11an1n08x5 FILLER_61_1541 ();
 b15zdnd11an1n04x5 FILLER_61_1549 ();
 b15zdnd11an1n16x5 FILLER_61_1569 ();
 b15zdnd11an1n04x5 FILLER_61_1585 ();
 b15zdnd11an1n16x5 FILLER_61_1596 ();
 b15zdnd11an1n04x5 FILLER_61_1612 ();
 b15zdnd00an1n01x5 FILLER_61_1616 ();
 b15zdnd11an1n64x5 FILLER_61_1628 ();
 b15zdnd11an1n64x5 FILLER_61_1692 ();
 b15zdnd11an1n04x5 FILLER_61_1756 ();
 b15zdnd00an1n02x5 FILLER_61_1760 ();
 b15zdnd00an1n01x5 FILLER_61_1762 ();
 b15zdnd11an1n04x5 FILLER_61_1769 ();
 b15zdnd11an1n64x5 FILLER_61_1778 ();
 b15zdnd11an1n08x5 FILLER_61_1842 ();
 b15zdnd11an1n04x5 FILLER_61_1850 ();
 b15zdnd11an1n64x5 FILLER_61_1859 ();
 b15zdnd11an1n32x5 FILLER_61_1923 ();
 b15zdnd11an1n16x5 FILLER_61_1955 ();
 b15zdnd11an1n04x5 FILLER_61_1971 ();
 b15zdnd11an1n64x5 FILLER_61_1980 ();
 b15zdnd11an1n08x5 FILLER_61_2044 ();
 b15zdnd00an1n02x5 FILLER_61_2052 ();
 b15zdnd00an1n01x5 FILLER_61_2054 ();
 b15zdnd11an1n16x5 FILLER_61_2065 ();
 b15zdnd11an1n04x5 FILLER_61_2081 ();
 b15zdnd11an1n08x5 FILLER_61_2101 ();
 b15zdnd11an1n04x5 FILLER_61_2109 ();
 b15zdnd00an1n02x5 FILLER_61_2113 ();
 b15zdnd11an1n16x5 FILLER_61_2121 ();
 b15zdnd11an1n08x5 FILLER_61_2137 ();
 b15zdnd11an1n04x5 FILLER_61_2145 ();
 b15zdnd00an1n02x5 FILLER_61_2149 ();
 b15zdnd11an1n64x5 FILLER_61_2169 ();
 b15zdnd11an1n32x5 FILLER_61_2233 ();
 b15zdnd11an1n16x5 FILLER_61_2265 ();
 b15zdnd00an1n02x5 FILLER_61_2281 ();
 b15zdnd00an1n01x5 FILLER_61_2283 ();
 b15zdnd11an1n64x5 FILLER_62_8 ();
 b15zdnd11an1n32x5 FILLER_62_72 ();
 b15zdnd11an1n04x5 FILLER_62_104 ();
 b15zdnd00an1n01x5 FILLER_62_108 ();
 b15zdnd11an1n08x5 FILLER_62_114 ();
 b15zdnd11an1n04x5 FILLER_62_122 ();
 b15zdnd00an1n02x5 FILLER_62_126 ();
 b15zdnd00an1n01x5 FILLER_62_128 ();
 b15zdnd11an1n32x5 FILLER_62_139 ();
 b15zdnd11an1n08x5 FILLER_62_171 ();
 b15zdnd00an1n01x5 FILLER_62_179 ();
 b15zdnd11an1n08x5 FILLER_62_200 ();
 b15zdnd00an1n02x5 FILLER_62_208 ();
 b15zdnd00an1n01x5 FILLER_62_210 ();
 b15zdnd11an1n04x5 FILLER_62_215 ();
 b15zdnd11an1n32x5 FILLER_62_236 ();
 b15zdnd11an1n16x5 FILLER_62_268 ();
 b15zdnd00an1n02x5 FILLER_62_284 ();
 b15zdnd00an1n01x5 FILLER_62_286 ();
 b15zdnd11an1n32x5 FILLER_62_297 ();
 b15zdnd11an1n64x5 FILLER_62_360 ();
 b15zdnd11an1n32x5 FILLER_62_424 ();
 b15zdnd00an1n01x5 FILLER_62_456 ();
 b15zdnd11an1n04x5 FILLER_62_467 ();
 b15zdnd11an1n32x5 FILLER_62_487 ();
 b15zdnd11an1n04x5 FILLER_62_519 ();
 b15zdnd00an1n02x5 FILLER_62_523 ();
 b15zdnd00an1n01x5 FILLER_62_525 ();
 b15zdnd11an1n04x5 FILLER_62_542 ();
 b15zdnd11an1n04x5 FILLER_62_557 ();
 b15zdnd11an1n16x5 FILLER_62_575 ();
 b15zdnd11an1n08x5 FILLER_62_591 ();
 b15zdnd11an1n04x5 FILLER_62_599 ();
 b15zdnd00an1n02x5 FILLER_62_603 ();
 b15zdnd00an1n01x5 FILLER_62_605 ();
 b15zdnd11an1n08x5 FILLER_62_615 ();
 b15zdnd00an1n02x5 FILLER_62_623 ();
 b15zdnd11an1n64x5 FILLER_62_632 ();
 b15zdnd11an1n16x5 FILLER_62_696 ();
 b15zdnd11an1n04x5 FILLER_62_712 ();
 b15zdnd00an1n02x5 FILLER_62_716 ();
 b15zdnd11an1n64x5 FILLER_62_726 ();
 b15zdnd11an1n08x5 FILLER_62_790 ();
 b15zdnd11an1n04x5 FILLER_62_798 ();
 b15zdnd00an1n01x5 FILLER_62_802 ();
 b15zdnd11an1n16x5 FILLER_62_815 ();
 b15zdnd11an1n04x5 FILLER_62_831 ();
 b15zdnd00an1n02x5 FILLER_62_835 ();
 b15zdnd00an1n01x5 FILLER_62_837 ();
 b15zdnd11an1n16x5 FILLER_62_864 ();
 b15zdnd11an1n08x5 FILLER_62_880 ();
 b15zdnd11an1n64x5 FILLER_62_906 ();
 b15zdnd11an1n64x5 FILLER_62_970 ();
 b15zdnd11an1n08x5 FILLER_62_1043 ();
 b15zdnd00an1n01x5 FILLER_62_1051 ();
 b15zdnd11an1n16x5 FILLER_62_1070 ();
 b15zdnd11an1n04x5 FILLER_62_1086 ();
 b15zdnd00an1n02x5 FILLER_62_1090 ();
 b15zdnd11an1n16x5 FILLER_62_1101 ();
 b15zdnd11an1n08x5 FILLER_62_1117 ();
 b15zdnd11an1n04x5 FILLER_62_1125 ();
 b15zdnd00an1n02x5 FILLER_62_1129 ();
 b15zdnd00an1n01x5 FILLER_62_1131 ();
 b15zdnd11an1n04x5 FILLER_62_1142 ();
 b15zdnd11an1n04x5 FILLER_62_1203 ();
 b15zdnd00an1n01x5 FILLER_62_1207 ();
 b15zdnd11an1n64x5 FILLER_62_1226 ();
 b15zdnd11an1n08x5 FILLER_62_1290 ();
 b15zdnd11an1n04x5 FILLER_62_1298 ();
 b15zdnd00an1n02x5 FILLER_62_1302 ();
 b15zdnd00an1n01x5 FILLER_62_1304 ();
 b15zdnd11an1n16x5 FILLER_62_1311 ();
 b15zdnd11an1n64x5 FILLER_62_1333 ();
 b15zdnd11an1n32x5 FILLER_62_1397 ();
 b15zdnd11an1n16x5 FILLER_62_1429 ();
 b15zdnd11an1n08x5 FILLER_62_1445 ();
 b15zdnd11an1n04x5 FILLER_62_1453 ();
 b15zdnd00an1n02x5 FILLER_62_1457 ();
 b15zdnd00an1n01x5 FILLER_62_1459 ();
 b15zdnd11an1n08x5 FILLER_62_1471 ();
 b15zdnd00an1n02x5 FILLER_62_1479 ();
 b15zdnd11an1n16x5 FILLER_62_1487 ();
 b15zdnd11an1n08x5 FILLER_62_1503 ();
 b15zdnd11an1n04x5 FILLER_62_1511 ();
 b15zdnd00an1n01x5 FILLER_62_1515 ();
 b15zdnd11an1n32x5 FILLER_62_1530 ();
 b15zdnd00an1n01x5 FILLER_62_1562 ();
 b15zdnd11an1n16x5 FILLER_62_1567 ();
 b15zdnd11an1n08x5 FILLER_62_1583 ();
 b15zdnd11an1n04x5 FILLER_62_1591 ();
 b15zdnd11an1n16x5 FILLER_62_1600 ();
 b15zdnd11an1n04x5 FILLER_62_1616 ();
 b15zdnd00an1n01x5 FILLER_62_1620 ();
 b15zdnd11an1n32x5 FILLER_62_1629 ();
 b15zdnd11an1n08x5 FILLER_62_1661 ();
 b15zdnd11an1n04x5 FILLER_62_1681 ();
 b15zdnd00an1n02x5 FILLER_62_1685 ();
 b15zdnd00an1n01x5 FILLER_62_1687 ();
 b15zdnd11an1n04x5 FILLER_62_1693 ();
 b15zdnd11an1n32x5 FILLER_62_1700 ();
 b15zdnd11an1n16x5 FILLER_62_1732 ();
 b15zdnd11an1n04x5 FILLER_62_1748 ();
 b15zdnd11an1n08x5 FILLER_62_1758 ();
 b15zdnd11an1n04x5 FILLER_62_1766 ();
 b15zdnd00an1n02x5 FILLER_62_1770 ();
 b15zdnd11an1n32x5 FILLER_62_1787 ();
 b15zdnd11an1n16x5 FILLER_62_1819 ();
 b15zdnd00an1n02x5 FILLER_62_1835 ();
 b15zdnd11an1n04x5 FILLER_62_1849 ();
 b15zdnd11an1n32x5 FILLER_62_1860 ();
 b15zdnd00an1n02x5 FILLER_62_1892 ();
 b15zdnd11an1n32x5 FILLER_62_1901 ();
 b15zdnd00an1n01x5 FILLER_62_1933 ();
 b15zdnd11an1n08x5 FILLER_62_1946 ();
 b15zdnd11an1n04x5 FILLER_62_1954 ();
 b15zdnd00an1n02x5 FILLER_62_1958 ();
 b15zdnd11an1n04x5 FILLER_62_1965 ();
 b15zdnd00an1n01x5 FILLER_62_1969 ();
 b15zdnd11an1n08x5 FILLER_62_1974 ();
 b15zdnd11an1n04x5 FILLER_62_1982 ();
 b15zdnd11an1n08x5 FILLER_62_1991 ();
 b15zdnd11an1n04x5 FILLER_62_1999 ();
 b15zdnd00an1n02x5 FILLER_62_2003 ();
 b15zdnd00an1n01x5 FILLER_62_2005 ();
 b15zdnd11an1n08x5 FILLER_62_2027 ();
 b15zdnd11an1n04x5 FILLER_62_2035 ();
 b15zdnd00an1n02x5 FILLER_62_2039 ();
 b15zdnd00an1n01x5 FILLER_62_2041 ();
 b15zdnd11an1n16x5 FILLER_62_2063 ();
 b15zdnd11an1n08x5 FILLER_62_2079 ();
 b15zdnd11an1n08x5 FILLER_62_2103 ();
 b15zdnd11an1n04x5 FILLER_62_2111 ();
 b15zdnd11an1n16x5 FILLER_62_2124 ();
 b15zdnd11an1n08x5 FILLER_62_2140 ();
 b15zdnd11an1n04x5 FILLER_62_2148 ();
 b15zdnd00an1n02x5 FILLER_62_2152 ();
 b15zdnd11an1n16x5 FILLER_62_2162 ();
 b15zdnd11an1n04x5 FILLER_62_2186 ();
 b15zdnd11an1n64x5 FILLER_62_2204 ();
 b15zdnd11an1n08x5 FILLER_62_2268 ();
 b15zdnd11an1n32x5 FILLER_63_0 ();
 b15zdnd11an1n16x5 FILLER_63_32 ();
 b15zdnd11an1n04x5 FILLER_63_48 ();
 b15zdnd00an1n01x5 FILLER_63_52 ();
 b15zdnd11an1n32x5 FILLER_63_68 ();
 b15zdnd11an1n16x5 FILLER_63_100 ();
 b15zdnd00an1n02x5 FILLER_63_116 ();
 b15zdnd11an1n64x5 FILLER_63_127 ();
 b15zdnd11an1n32x5 FILLER_63_191 ();
 b15zdnd11an1n16x5 FILLER_63_223 ();
 b15zdnd11an1n04x5 FILLER_63_239 ();
 b15zdnd11an1n32x5 FILLER_63_253 ();
 b15zdnd00an1n02x5 FILLER_63_285 ();
 b15zdnd11an1n04x5 FILLER_63_299 ();
 b15zdnd11an1n16x5 FILLER_63_310 ();
 b15zdnd11an1n08x5 FILLER_63_326 ();
 b15zdnd11an1n04x5 FILLER_63_334 ();
 b15zdnd00an1n02x5 FILLER_63_338 ();
 b15zdnd00an1n01x5 FILLER_63_340 ();
 b15zdnd11an1n64x5 FILLER_63_355 ();
 b15zdnd11an1n16x5 FILLER_63_419 ();
 b15zdnd11an1n04x5 FILLER_63_435 ();
 b15zdnd00an1n02x5 FILLER_63_439 ();
 b15zdnd11an1n04x5 FILLER_63_459 ();
 b15zdnd11an1n16x5 FILLER_63_470 ();
 b15zdnd00an1n02x5 FILLER_63_486 ();
 b15zdnd11an1n32x5 FILLER_63_498 ();
 b15zdnd11an1n16x5 FILLER_63_530 ();
 b15zdnd11an1n08x5 FILLER_63_546 ();
 b15zdnd11an1n04x5 FILLER_63_554 ();
 b15zdnd00an1n02x5 FILLER_63_558 ();
 b15zdnd00an1n01x5 FILLER_63_560 ();
 b15zdnd11an1n32x5 FILLER_63_565 ();
 b15zdnd11an1n16x5 FILLER_63_597 ();
 b15zdnd11an1n04x5 FILLER_63_613 ();
 b15zdnd00an1n01x5 FILLER_63_617 ();
 b15zdnd11an1n04x5 FILLER_63_624 ();
 b15zdnd11an1n08x5 FILLER_63_644 ();
 b15zdnd00an1n01x5 FILLER_63_652 ();
 b15zdnd11an1n08x5 FILLER_63_661 ();
 b15zdnd11an1n04x5 FILLER_63_669 ();
 b15zdnd00an1n01x5 FILLER_63_673 ();
 b15zdnd11an1n04x5 FILLER_63_688 ();
 b15zdnd11an1n32x5 FILLER_63_697 ();
 b15zdnd11an1n16x5 FILLER_63_729 ();
 b15zdnd11an1n04x5 FILLER_63_745 ();
 b15zdnd11an1n04x5 FILLER_63_758 ();
 b15zdnd11an1n16x5 FILLER_63_775 ();
 b15zdnd11an1n08x5 FILLER_63_791 ();
 b15zdnd11an1n04x5 FILLER_63_799 ();
 b15zdnd00an1n02x5 FILLER_63_803 ();
 b15zdnd11an1n16x5 FILLER_63_825 ();
 b15zdnd11an1n16x5 FILLER_63_851 ();
 b15zdnd11an1n04x5 FILLER_63_867 ();
 b15zdnd00an1n01x5 FILLER_63_871 ();
 b15zdnd11an1n64x5 FILLER_63_886 ();
 b15zdnd11an1n32x5 FILLER_63_950 ();
 b15zdnd11an1n04x5 FILLER_63_982 ();
 b15zdnd00an1n02x5 FILLER_63_986 ();
 b15zdnd11an1n32x5 FILLER_63_997 ();
 b15zdnd11an1n16x5 FILLER_63_1029 ();
 b15zdnd11an1n08x5 FILLER_63_1045 ();
 b15zdnd00an1n02x5 FILLER_63_1053 ();
 b15zdnd00an1n01x5 FILLER_63_1055 ();
 b15zdnd11an1n64x5 FILLER_63_1081 ();
 b15zdnd11an1n32x5 FILLER_63_1145 ();
 b15zdnd11an1n04x5 FILLER_63_1208 ();
 b15zdnd11an1n32x5 FILLER_63_1230 ();
 b15zdnd11an1n16x5 FILLER_63_1262 ();
 b15zdnd11an1n04x5 FILLER_63_1278 ();
 b15zdnd00an1n02x5 FILLER_63_1282 ();
 b15zdnd00an1n01x5 FILLER_63_1284 ();
 b15zdnd11an1n32x5 FILLER_63_1291 ();
 b15zdnd11an1n16x5 FILLER_63_1323 ();
 b15zdnd11an1n08x5 FILLER_63_1339 ();
 b15zdnd00an1n01x5 FILLER_63_1347 ();
 b15zdnd11an1n64x5 FILLER_63_1353 ();
 b15zdnd11an1n32x5 FILLER_63_1417 ();
 b15zdnd11an1n08x5 FILLER_63_1449 ();
 b15zdnd00an1n02x5 FILLER_63_1457 ();
 b15zdnd00an1n01x5 FILLER_63_1459 ();
 b15zdnd11an1n04x5 FILLER_63_1470 ();
 b15zdnd00an1n02x5 FILLER_63_1474 ();
 b15zdnd00an1n01x5 FILLER_63_1476 ();
 b15zdnd11an1n64x5 FILLER_63_1490 ();
 b15zdnd11an1n08x5 FILLER_63_1554 ();
 b15zdnd00an1n02x5 FILLER_63_1562 ();
 b15zdnd00an1n01x5 FILLER_63_1564 ();
 b15zdnd11an1n64x5 FILLER_63_1577 ();
 b15zdnd11an1n08x5 FILLER_63_1641 ();
 b15zdnd11an1n04x5 FILLER_63_1649 ();
 b15zdnd00an1n01x5 FILLER_63_1653 ();
 b15zdnd11an1n16x5 FILLER_63_1660 ();
 b15zdnd11an1n08x5 FILLER_63_1676 ();
 b15zdnd00an1n02x5 FILLER_63_1684 ();
 b15zdnd00an1n01x5 FILLER_63_1686 ();
 b15zdnd11an1n32x5 FILLER_63_1707 ();
 b15zdnd11an1n08x5 FILLER_63_1739 ();
 b15zdnd11an1n04x5 FILLER_63_1747 ();
 b15zdnd00an1n02x5 FILLER_63_1751 ();
 b15zdnd11an1n04x5 FILLER_63_1785 ();
 b15zdnd11an1n04x5 FILLER_63_1820 ();
 b15zdnd11an1n04x5 FILLER_63_1850 ();
 b15zdnd11an1n04x5 FILLER_63_1870 ();
 b15zdnd00an1n02x5 FILLER_63_1874 ();
 b15zdnd00an1n01x5 FILLER_63_1876 ();
 b15zdnd11an1n04x5 FILLER_63_1883 ();
 b15zdnd11an1n04x5 FILLER_63_1898 ();
 b15zdnd11an1n04x5 FILLER_63_1912 ();
 b15zdnd11an1n16x5 FILLER_63_1924 ();
 b15zdnd11an1n04x5 FILLER_63_1940 ();
 b15zdnd11an1n08x5 FILLER_63_1950 ();
 b15zdnd11an1n04x5 FILLER_63_1958 ();
 b15zdnd00an1n02x5 FILLER_63_1962 ();
 b15zdnd11an1n16x5 FILLER_63_1971 ();
 b15zdnd00an1n01x5 FILLER_63_1987 ();
 b15zdnd11an1n16x5 FILLER_63_1995 ();
 b15zdnd11an1n32x5 FILLER_63_2016 ();
 b15zdnd11an1n04x5 FILLER_63_2048 ();
 b15zdnd11an1n04x5 FILLER_63_2060 ();
 b15zdnd11an1n16x5 FILLER_63_2096 ();
 b15zdnd11an1n04x5 FILLER_63_2112 ();
 b15zdnd00an1n02x5 FILLER_63_2116 ();
 b15zdnd11an1n04x5 FILLER_63_2123 ();
 b15zdnd00an1n01x5 FILLER_63_2127 ();
 b15zdnd11an1n16x5 FILLER_63_2160 ();
 b15zdnd11an1n08x5 FILLER_63_2176 ();
 b15zdnd11an1n08x5 FILLER_63_2188 ();
 b15zdnd11an1n04x5 FILLER_63_2196 ();
 b15zdnd11an1n08x5 FILLER_63_2204 ();
 b15zdnd00an1n02x5 FILLER_63_2212 ();
 b15zdnd00an1n01x5 FILLER_63_2214 ();
 b15zdnd11an1n32x5 FILLER_63_2237 ();
 b15zdnd11an1n08x5 FILLER_63_2269 ();
 b15zdnd11an1n04x5 FILLER_63_2277 ();
 b15zdnd00an1n02x5 FILLER_63_2281 ();
 b15zdnd00an1n01x5 FILLER_63_2283 ();
 b15zdnd11an1n16x5 FILLER_64_8 ();
 b15zdnd11an1n04x5 FILLER_64_24 ();
 b15zdnd11an1n08x5 FILLER_64_42 ();
 b15zdnd00an1n01x5 FILLER_64_50 ();
 b15zdnd11an1n08x5 FILLER_64_59 ();
 b15zdnd11an1n04x5 FILLER_64_67 ();
 b15zdnd00an1n02x5 FILLER_64_71 ();
 b15zdnd00an1n01x5 FILLER_64_73 ();
 b15zdnd11an1n32x5 FILLER_64_81 ();
 b15zdnd11an1n16x5 FILLER_64_113 ();
 b15zdnd11an1n32x5 FILLER_64_135 ();
 b15zdnd11an1n16x5 FILLER_64_167 ();
 b15zdnd11an1n08x5 FILLER_64_183 ();
 b15zdnd11an1n64x5 FILLER_64_196 ();
 b15zdnd11an1n32x5 FILLER_64_260 ();
 b15zdnd11an1n16x5 FILLER_64_292 ();
 b15zdnd00an1n02x5 FILLER_64_308 ();
 b15zdnd11an1n04x5 FILLER_64_316 ();
 b15zdnd11an1n32x5 FILLER_64_326 ();
 b15zdnd11an1n08x5 FILLER_64_358 ();
 b15zdnd11an1n04x5 FILLER_64_381 ();
 b15zdnd11an1n64x5 FILLER_64_389 ();
 b15zdnd11an1n64x5 FILLER_64_453 ();
 b15zdnd11an1n08x5 FILLER_64_517 ();
 b15zdnd00an1n02x5 FILLER_64_525 ();
 b15zdnd00an1n01x5 FILLER_64_527 ();
 b15zdnd11an1n16x5 FILLER_64_532 ();
 b15zdnd11an1n08x5 FILLER_64_548 ();
 b15zdnd00an1n02x5 FILLER_64_556 ();
 b15zdnd11an1n16x5 FILLER_64_564 ();
 b15zdnd11an1n08x5 FILLER_64_580 ();
 b15zdnd11an1n04x5 FILLER_64_588 ();
 b15zdnd00an1n02x5 FILLER_64_592 ();
 b15zdnd00an1n01x5 FILLER_64_594 ();
 b15zdnd11an1n08x5 FILLER_64_612 ();
 b15zdnd11an1n04x5 FILLER_64_620 ();
 b15zdnd11an1n16x5 FILLER_64_636 ();
 b15zdnd00an1n02x5 FILLER_64_652 ();
 b15zdnd00an1n01x5 FILLER_64_654 ();
 b15zdnd11an1n16x5 FILLER_64_664 ();
 b15zdnd11an1n08x5 FILLER_64_680 ();
 b15zdnd11an1n04x5 FILLER_64_688 ();
 b15zdnd00an1n02x5 FILLER_64_692 ();
 b15zdnd00an1n01x5 FILLER_64_694 ();
 b15zdnd11an1n16x5 FILLER_64_701 ();
 b15zdnd00an1n01x5 FILLER_64_717 ();
 b15zdnd11an1n08x5 FILLER_64_726 ();
 b15zdnd00an1n02x5 FILLER_64_734 ();
 b15zdnd00an1n01x5 FILLER_64_736 ();
 b15zdnd11an1n32x5 FILLER_64_742 ();
 b15zdnd11an1n16x5 FILLER_64_774 ();
 b15zdnd11an1n08x5 FILLER_64_790 ();
 b15zdnd00an1n02x5 FILLER_64_798 ();
 b15zdnd00an1n01x5 FILLER_64_800 ();
 b15zdnd11an1n16x5 FILLER_64_817 ();
 b15zdnd11an1n64x5 FILLER_64_851 ();
 b15zdnd11an1n64x5 FILLER_64_915 ();
 b15zdnd11an1n08x5 FILLER_64_979 ();
 b15zdnd00an1n01x5 FILLER_64_987 ();
 b15zdnd11an1n64x5 FILLER_64_997 ();
 b15zdnd11an1n64x5 FILLER_64_1061 ();
 b15zdnd11an1n32x5 FILLER_64_1125 ();
 b15zdnd11an1n08x5 FILLER_64_1157 ();
 b15zdnd11an1n16x5 FILLER_64_1183 ();
 b15zdnd11an1n64x5 FILLER_64_1227 ();
 b15zdnd11an1n16x5 FILLER_64_1291 ();
 b15zdnd11an1n08x5 FILLER_64_1307 ();
 b15zdnd11an1n04x5 FILLER_64_1315 ();
 b15zdnd00an1n02x5 FILLER_64_1319 ();
 b15zdnd00an1n01x5 FILLER_64_1321 ();
 b15zdnd11an1n08x5 FILLER_64_1331 ();
 b15zdnd00an1n02x5 FILLER_64_1339 ();
 b15zdnd00an1n01x5 FILLER_64_1341 ();
 b15zdnd11an1n04x5 FILLER_64_1349 ();
 b15zdnd11an1n64x5 FILLER_64_1360 ();
 b15zdnd00an1n01x5 FILLER_64_1424 ();
 b15zdnd11an1n04x5 FILLER_64_1442 ();
 b15zdnd11an1n64x5 FILLER_64_1456 ();
 b15zdnd11an1n32x5 FILLER_64_1520 ();
 b15zdnd11an1n08x5 FILLER_64_1552 ();
 b15zdnd11an1n04x5 FILLER_64_1560 ();
 b15zdnd00an1n01x5 FILLER_64_1564 ();
 b15zdnd11an1n64x5 FILLER_64_1581 ();
 b15zdnd11an1n08x5 FILLER_64_1645 ();
 b15zdnd00an1n02x5 FILLER_64_1653 ();
 b15zdnd11an1n64x5 FILLER_64_1668 ();
 b15zdnd11an1n64x5 FILLER_64_1732 ();
 b15zdnd11an1n16x5 FILLER_64_1796 ();
 b15zdnd11an1n04x5 FILLER_64_1812 ();
 b15zdnd00an1n02x5 FILLER_64_1816 ();
 b15zdnd11an1n08x5 FILLER_64_1829 ();
 b15zdnd11an1n04x5 FILLER_64_1856 ();
 b15zdnd00an1n02x5 FILLER_64_1860 ();
 b15zdnd00an1n01x5 FILLER_64_1862 ();
 b15zdnd11an1n04x5 FILLER_64_1879 ();
 b15zdnd11an1n64x5 FILLER_64_1889 ();
 b15zdnd11an1n08x5 FILLER_64_1953 ();
 b15zdnd00an1n01x5 FILLER_64_1961 ();
 b15zdnd11an1n32x5 FILLER_64_1974 ();
 b15zdnd11an1n04x5 FILLER_64_2006 ();
 b15zdnd00an1n02x5 FILLER_64_2010 ();
 b15zdnd11an1n64x5 FILLER_64_2018 ();
 b15zdnd11an1n64x5 FILLER_64_2082 ();
 b15zdnd11an1n08x5 FILLER_64_2146 ();
 b15zdnd11an1n16x5 FILLER_64_2162 ();
 b15zdnd00an1n02x5 FILLER_64_2178 ();
 b15zdnd00an1n01x5 FILLER_64_2180 ();
 b15zdnd11an1n64x5 FILLER_64_2195 ();
 b15zdnd11an1n16x5 FILLER_64_2259 ();
 b15zdnd00an1n01x5 FILLER_64_2275 ();
 b15zdnd11an1n64x5 FILLER_65_0 ();
 b15zdnd11an1n04x5 FILLER_65_64 ();
 b15zdnd00an1n02x5 FILLER_65_68 ();
 b15zdnd11an1n32x5 FILLER_65_82 ();
 b15zdnd11an1n16x5 FILLER_65_114 ();
 b15zdnd11an1n04x5 FILLER_65_130 ();
 b15zdnd00an1n01x5 FILLER_65_134 ();
 b15zdnd11an1n32x5 FILLER_65_141 ();
 b15zdnd11an1n16x5 FILLER_65_173 ();
 b15zdnd00an1n02x5 FILLER_65_189 ();
 b15zdnd00an1n01x5 FILLER_65_191 ();
 b15zdnd11an1n16x5 FILLER_65_198 ();
 b15zdnd00an1n01x5 FILLER_65_214 ();
 b15zdnd11an1n64x5 FILLER_65_222 ();
 b15zdnd11an1n64x5 FILLER_65_290 ();
 b15zdnd11an1n64x5 FILLER_65_354 ();
 b15zdnd11an1n64x5 FILLER_65_418 ();
 b15zdnd11an1n04x5 FILLER_65_482 ();
 b15zdnd00an1n02x5 FILLER_65_486 ();
 b15zdnd11an1n16x5 FILLER_65_499 ();
 b15zdnd11an1n08x5 FILLER_65_515 ();
 b15zdnd00an1n02x5 FILLER_65_523 ();
 b15zdnd11an1n64x5 FILLER_65_540 ();
 b15zdnd11an1n64x5 FILLER_65_604 ();
 b15zdnd11an1n16x5 FILLER_65_668 ();
 b15zdnd11an1n04x5 FILLER_65_684 ();
 b15zdnd00an1n02x5 FILLER_65_688 ();
 b15zdnd00an1n01x5 FILLER_65_690 ();
 b15zdnd11an1n32x5 FILLER_65_698 ();
 b15zdnd11an1n08x5 FILLER_65_730 ();
 b15zdnd11an1n16x5 FILLER_65_750 ();
 b15zdnd11an1n04x5 FILLER_65_766 ();
 b15zdnd11an1n64x5 FILLER_65_791 ();
 b15zdnd00an1n02x5 FILLER_65_855 ();
 b15zdnd00an1n01x5 FILLER_65_857 ();
 b15zdnd11an1n04x5 FILLER_65_862 ();
 b15zdnd00an1n02x5 FILLER_65_866 ();
 b15zdnd00an1n01x5 FILLER_65_868 ();
 b15zdnd11an1n64x5 FILLER_65_895 ();
 b15zdnd11an1n64x5 FILLER_65_959 ();
 b15zdnd11an1n32x5 FILLER_65_1023 ();
 b15zdnd11an1n16x5 FILLER_65_1055 ();
 b15zdnd11an1n08x5 FILLER_65_1071 ();
 b15zdnd11an1n04x5 FILLER_65_1079 ();
 b15zdnd11an1n04x5 FILLER_65_1087 ();
 b15zdnd11an1n32x5 FILLER_65_1100 ();
 b15zdnd00an1n01x5 FILLER_65_1132 ();
 b15zdnd11an1n32x5 FILLER_65_1159 ();
 b15zdnd00an1n01x5 FILLER_65_1191 ();
 b15zdnd11an1n32x5 FILLER_65_1217 ();
 b15zdnd11an1n16x5 FILLER_65_1249 ();
 b15zdnd11an1n08x5 FILLER_65_1265 ();
 b15zdnd11an1n04x5 FILLER_65_1273 ();
 b15zdnd00an1n01x5 FILLER_65_1277 ();
 b15zdnd11an1n04x5 FILLER_65_1285 ();
 b15zdnd11an1n32x5 FILLER_65_1298 ();
 b15zdnd11an1n16x5 FILLER_65_1330 ();
 b15zdnd11an1n04x5 FILLER_65_1346 ();
 b15zdnd00an1n02x5 FILLER_65_1350 ();
 b15zdnd00an1n01x5 FILLER_65_1352 ();
 b15zdnd11an1n32x5 FILLER_65_1358 ();
 b15zdnd11an1n08x5 FILLER_65_1390 ();
 b15zdnd11an1n04x5 FILLER_65_1398 ();
 b15zdnd00an1n01x5 FILLER_65_1402 ();
 b15zdnd11an1n32x5 FILLER_65_1418 ();
 b15zdnd11an1n16x5 FILLER_65_1462 ();
 b15zdnd11an1n08x5 FILLER_65_1478 ();
 b15zdnd00an1n01x5 FILLER_65_1486 ();
 b15zdnd11an1n32x5 FILLER_65_1492 ();
 b15zdnd11an1n16x5 FILLER_65_1524 ();
 b15zdnd11an1n08x5 FILLER_65_1540 ();
 b15zdnd00an1n02x5 FILLER_65_1548 ();
 b15zdnd11an1n64x5 FILLER_65_1562 ();
 b15zdnd11an1n16x5 FILLER_65_1626 ();
 b15zdnd11an1n08x5 FILLER_65_1642 ();
 b15zdnd00an1n01x5 FILLER_65_1650 ();
 b15zdnd11an1n64x5 FILLER_65_1665 ();
 b15zdnd11an1n64x5 FILLER_65_1729 ();
 b15zdnd11an1n64x5 FILLER_65_1793 ();
 b15zdnd11an1n16x5 FILLER_65_1857 ();
 b15zdnd11an1n04x5 FILLER_65_1873 ();
 b15zdnd00an1n02x5 FILLER_65_1877 ();
 b15zdnd11an1n64x5 FILLER_65_1895 ();
 b15zdnd11an1n64x5 FILLER_65_1959 ();
 b15zdnd11an1n64x5 FILLER_65_2023 ();
 b15zdnd11an1n64x5 FILLER_65_2087 ();
 b15zdnd11an1n64x5 FILLER_65_2151 ();
 b15zdnd11an1n64x5 FILLER_65_2215 ();
 b15zdnd11an1n04x5 FILLER_65_2279 ();
 b15zdnd00an1n01x5 FILLER_65_2283 ();
 b15zdnd11an1n64x5 FILLER_66_8 ();
 b15zdnd11an1n32x5 FILLER_66_72 ();
 b15zdnd11an1n08x5 FILLER_66_104 ();
 b15zdnd11an1n16x5 FILLER_66_136 ();
 b15zdnd00an1n02x5 FILLER_66_152 ();
 b15zdnd00an1n01x5 FILLER_66_154 ();
 b15zdnd11an1n08x5 FILLER_66_161 ();
 b15zdnd00an1n02x5 FILLER_66_169 ();
 b15zdnd11an1n16x5 FILLER_66_176 ();
 b15zdnd11an1n08x5 FILLER_66_199 ();
 b15zdnd11an1n04x5 FILLER_66_207 ();
 b15zdnd00an1n02x5 FILLER_66_211 ();
 b15zdnd00an1n01x5 FILLER_66_213 ();
 b15zdnd11an1n08x5 FILLER_66_226 ();
 b15zdnd11an1n04x5 FILLER_66_234 ();
 b15zdnd11an1n08x5 FILLER_66_244 ();
 b15zdnd11an1n04x5 FILLER_66_252 ();
 b15zdnd00an1n02x5 FILLER_66_256 ();
 b15zdnd00an1n01x5 FILLER_66_258 ();
 b15zdnd11an1n04x5 FILLER_66_266 ();
 b15zdnd11an1n04x5 FILLER_66_286 ();
 b15zdnd00an1n02x5 FILLER_66_290 ();
 b15zdnd00an1n01x5 FILLER_66_292 ();
 b15zdnd11an1n32x5 FILLER_66_297 ();
 b15zdnd11an1n16x5 FILLER_66_329 ();
 b15zdnd11an1n08x5 FILLER_66_345 ();
 b15zdnd11an1n04x5 FILLER_66_353 ();
 b15zdnd00an1n02x5 FILLER_66_357 ();
 b15zdnd00an1n01x5 FILLER_66_359 ();
 b15zdnd11an1n04x5 FILLER_66_367 ();
 b15zdnd00an1n02x5 FILLER_66_371 ();
 b15zdnd00an1n01x5 FILLER_66_373 ();
 b15zdnd11an1n04x5 FILLER_66_380 ();
 b15zdnd11an1n64x5 FILLER_66_388 ();
 b15zdnd11an1n32x5 FILLER_66_452 ();
 b15zdnd11an1n04x5 FILLER_66_484 ();
 b15zdnd11an1n16x5 FILLER_66_506 ();
 b15zdnd11an1n04x5 FILLER_66_522 ();
 b15zdnd00an1n02x5 FILLER_66_526 ();
 b15zdnd00an1n01x5 FILLER_66_528 ();
 b15zdnd11an1n16x5 FILLER_66_536 ();
 b15zdnd11an1n08x5 FILLER_66_552 ();
 b15zdnd00an1n02x5 FILLER_66_560 ();
 b15zdnd11an1n16x5 FILLER_66_573 ();
 b15zdnd11an1n08x5 FILLER_66_589 ();
 b15zdnd11an1n16x5 FILLER_66_613 ();
 b15zdnd11an1n04x5 FILLER_66_629 ();
 b15zdnd11an1n04x5 FILLER_66_659 ();
 b15zdnd11an1n16x5 FILLER_66_667 ();
 b15zdnd11an1n04x5 FILLER_66_683 ();
 b15zdnd00an1n01x5 FILLER_66_687 ();
 b15zdnd11an1n04x5 FILLER_66_695 ();
 b15zdnd00an1n01x5 FILLER_66_699 ();
 b15zdnd00an1n02x5 FILLER_66_716 ();
 b15zdnd11an1n04x5 FILLER_66_726 ();
 b15zdnd00an1n02x5 FILLER_66_730 ();
 b15zdnd00an1n01x5 FILLER_66_732 ();
 b15zdnd11an1n16x5 FILLER_66_738 ();
 b15zdnd00an1n02x5 FILLER_66_754 ();
 b15zdnd11an1n32x5 FILLER_66_761 ();
 b15zdnd11an1n64x5 FILLER_66_811 ();
 b15zdnd11an1n32x5 FILLER_66_875 ();
 b15zdnd00an1n01x5 FILLER_66_907 ();
 b15zdnd11an1n08x5 FILLER_66_914 ();
 b15zdnd00an1n02x5 FILLER_66_922 ();
 b15zdnd11an1n16x5 FILLER_66_949 ();
 b15zdnd11an1n08x5 FILLER_66_965 ();
 b15zdnd11an1n04x5 FILLER_66_973 ();
 b15zdnd11an1n08x5 FILLER_66_997 ();
 b15zdnd11an1n04x5 FILLER_66_1005 ();
 b15zdnd00an1n02x5 FILLER_66_1009 ();
 b15zdnd00an1n01x5 FILLER_66_1011 ();
 b15zdnd11an1n32x5 FILLER_66_1038 ();
 b15zdnd11an1n16x5 FILLER_66_1070 ();
 b15zdnd11an1n08x5 FILLER_66_1086 ();
 b15zdnd00an1n01x5 FILLER_66_1094 ();
 b15zdnd11an1n32x5 FILLER_66_1105 ();
 b15zdnd11an1n04x5 FILLER_66_1137 ();
 b15zdnd00an1n02x5 FILLER_66_1141 ();
 b15zdnd11an1n64x5 FILLER_66_1153 ();
 b15zdnd11an1n16x5 FILLER_66_1217 ();
 b15zdnd00an1n01x5 FILLER_66_1233 ();
 b15zdnd11an1n16x5 FILLER_66_1260 ();
 b15zdnd11an1n08x5 FILLER_66_1276 ();
 b15zdnd11an1n04x5 FILLER_66_1284 ();
 b15zdnd11an1n32x5 FILLER_66_1294 ();
 b15zdnd11an1n16x5 FILLER_66_1326 ();
 b15zdnd11an1n08x5 FILLER_66_1342 ();
 b15zdnd00an1n02x5 FILLER_66_1350 ();
 b15zdnd00an1n01x5 FILLER_66_1352 ();
 b15zdnd11an1n16x5 FILLER_66_1357 ();
 b15zdnd11an1n08x5 FILLER_66_1373 ();
 b15zdnd00an1n02x5 FILLER_66_1381 ();
 b15zdnd11an1n04x5 FILLER_66_1400 ();
 b15zdnd11an1n32x5 FILLER_66_1411 ();
 b15zdnd00an1n02x5 FILLER_66_1443 ();
 b15zdnd00an1n01x5 FILLER_66_1445 ();
 b15zdnd11an1n32x5 FILLER_66_1455 ();
 b15zdnd11an1n04x5 FILLER_66_1487 ();
 b15zdnd11an1n32x5 FILLER_66_1500 ();
 b15zdnd11an1n16x5 FILLER_66_1532 ();
 b15zdnd11an1n16x5 FILLER_66_1555 ();
 b15zdnd11an1n08x5 FILLER_66_1571 ();
 b15zdnd11an1n04x5 FILLER_66_1579 ();
 b15zdnd00an1n01x5 FILLER_66_1583 ();
 b15zdnd11an1n08x5 FILLER_66_1588 ();
 b15zdnd00an1n02x5 FILLER_66_1596 ();
 b15zdnd11an1n04x5 FILLER_66_1604 ();
 b15zdnd11an1n04x5 FILLER_66_1615 ();
 b15zdnd11an1n04x5 FILLER_66_1625 ();
 b15zdnd00an1n01x5 FILLER_66_1629 ();
 b15zdnd11an1n08x5 FILLER_66_1635 ();
 b15zdnd11an1n04x5 FILLER_66_1643 ();
 b15zdnd00an1n02x5 FILLER_66_1647 ();
 b15zdnd00an1n01x5 FILLER_66_1649 ();
 b15zdnd11an1n64x5 FILLER_66_1658 ();
 b15zdnd11an1n64x5 FILLER_66_1722 ();
 b15zdnd11an1n64x5 FILLER_66_1786 ();
 b15zdnd11an1n64x5 FILLER_66_1850 ();
 b15zdnd11an1n64x5 FILLER_66_1914 ();
 b15zdnd11an1n64x5 FILLER_66_1978 ();
 b15zdnd11an1n64x5 FILLER_66_2042 ();
 b15zdnd11an1n32x5 FILLER_66_2106 ();
 b15zdnd11an1n16x5 FILLER_66_2138 ();
 b15zdnd11an1n64x5 FILLER_66_2162 ();
 b15zdnd11an1n32x5 FILLER_66_2226 ();
 b15zdnd11an1n16x5 FILLER_66_2258 ();
 b15zdnd00an1n02x5 FILLER_66_2274 ();
 b15zdnd11an1n32x5 FILLER_67_0 ();
 b15zdnd11an1n04x5 FILLER_67_32 ();
 b15zdnd00an1n02x5 FILLER_67_36 ();
 b15zdnd00an1n01x5 FILLER_67_38 ();
 b15zdnd11an1n04x5 FILLER_67_43 ();
 b15zdnd00an1n02x5 FILLER_67_47 ();
 b15zdnd00an1n01x5 FILLER_67_49 ();
 b15zdnd11an1n16x5 FILLER_67_66 ();
 b15zdnd11an1n08x5 FILLER_67_82 ();
 b15zdnd00an1n01x5 FILLER_67_90 ();
 b15zdnd11an1n32x5 FILLER_67_99 ();
 b15zdnd11an1n16x5 FILLER_67_131 ();
 b15zdnd11an1n08x5 FILLER_67_147 ();
 b15zdnd11an1n16x5 FILLER_67_161 ();
 b15zdnd11an1n04x5 FILLER_67_177 ();
 b15zdnd11an1n04x5 FILLER_67_213 ();
 b15zdnd11an1n08x5 FILLER_67_224 ();
 b15zdnd11an1n04x5 FILLER_67_232 ();
 b15zdnd00an1n02x5 FILLER_67_236 ();
 b15zdnd11an1n04x5 FILLER_67_247 ();
 b15zdnd11an1n04x5 FILLER_67_256 ();
 b15zdnd11an1n04x5 FILLER_67_286 ();
 b15zdnd00an1n01x5 FILLER_67_290 ();
 b15zdnd11an1n32x5 FILLER_67_300 ();
 b15zdnd11an1n16x5 FILLER_67_332 ();
 b15zdnd11an1n08x5 FILLER_67_348 ();
 b15zdnd11an1n04x5 FILLER_67_356 ();
 b15zdnd00an1n02x5 FILLER_67_360 ();
 b15zdnd00an1n01x5 FILLER_67_362 ();
 b15zdnd11an1n04x5 FILLER_67_373 ();
 b15zdnd11an1n16x5 FILLER_67_384 ();
 b15zdnd00an1n01x5 FILLER_67_400 ();
 b15zdnd11an1n04x5 FILLER_67_407 ();
 b15zdnd11an1n32x5 FILLER_67_419 ();
 b15zdnd11an1n08x5 FILLER_67_451 ();
 b15zdnd00an1n01x5 FILLER_67_459 ();
 b15zdnd11an1n32x5 FILLER_67_483 ();
 b15zdnd11an1n16x5 FILLER_67_515 ();
 b15zdnd11an1n08x5 FILLER_67_531 ();
 b15zdnd11an1n04x5 FILLER_67_539 ();
 b15zdnd00an1n01x5 FILLER_67_543 ();
 b15zdnd11an1n16x5 FILLER_67_557 ();
 b15zdnd11an1n08x5 FILLER_67_587 ();
 b15zdnd11an1n04x5 FILLER_67_595 ();
 b15zdnd00an1n01x5 FILLER_67_599 ();
 b15zdnd11an1n32x5 FILLER_67_607 ();
 b15zdnd11an1n16x5 FILLER_67_639 ();
 b15zdnd11an1n04x5 FILLER_67_655 ();
 b15zdnd00an1n02x5 FILLER_67_659 ();
 b15zdnd00an1n01x5 FILLER_67_661 ();
 b15zdnd11an1n08x5 FILLER_67_678 ();
 b15zdnd11an1n04x5 FILLER_67_686 ();
 b15zdnd00an1n01x5 FILLER_67_690 ();
 b15zdnd11an1n16x5 FILLER_67_697 ();
 b15zdnd00an1n02x5 FILLER_67_713 ();
 b15zdnd11an1n04x5 FILLER_67_720 ();
 b15zdnd00an1n01x5 FILLER_67_724 ();
 b15zdnd11an1n64x5 FILLER_67_733 ();
 b15zdnd11an1n32x5 FILLER_67_797 ();
 b15zdnd11an1n32x5 FILLER_67_834 ();
 b15zdnd11an1n04x5 FILLER_67_866 ();
 b15zdnd00an1n02x5 FILLER_67_870 ();
 b15zdnd11an1n16x5 FILLER_67_892 ();
 b15zdnd00an1n02x5 FILLER_67_908 ();
 b15zdnd11an1n64x5 FILLER_67_930 ();
 b15zdnd11an1n32x5 FILLER_67_994 ();
 b15zdnd11an1n16x5 FILLER_67_1026 ();
 b15zdnd11an1n08x5 FILLER_67_1042 ();
 b15zdnd00an1n02x5 FILLER_67_1050 ();
 b15zdnd00an1n01x5 FILLER_67_1052 ();
 b15zdnd11an1n64x5 FILLER_67_1058 ();
 b15zdnd11an1n64x5 FILLER_67_1122 ();
 b15zdnd11an1n64x5 FILLER_67_1186 ();
 b15zdnd11an1n32x5 FILLER_67_1250 ();
 b15zdnd00an1n02x5 FILLER_67_1282 ();
 b15zdnd00an1n01x5 FILLER_67_1284 ();
 b15zdnd11an1n32x5 FILLER_67_1290 ();
 b15zdnd11an1n04x5 FILLER_67_1322 ();
 b15zdnd00an1n02x5 FILLER_67_1326 ();
 b15zdnd00an1n01x5 FILLER_67_1328 ();
 b15zdnd11an1n32x5 FILLER_67_1345 ();
 b15zdnd00an1n02x5 FILLER_67_1377 ();
 b15zdnd11an1n04x5 FILLER_67_1385 ();
 b15zdnd00an1n01x5 FILLER_67_1389 ();
 b15zdnd11an1n32x5 FILLER_67_1402 ();
 b15zdnd11an1n08x5 FILLER_67_1434 ();
 b15zdnd11an1n04x5 FILLER_67_1442 ();
 b15zdnd11an1n32x5 FILLER_67_1455 ();
 b15zdnd11an1n16x5 FILLER_67_1487 ();
 b15zdnd11an1n08x5 FILLER_67_1503 ();
 b15zdnd00an1n01x5 FILLER_67_1511 ();
 b15zdnd11an1n04x5 FILLER_67_1518 ();
 b15zdnd00an1n02x5 FILLER_67_1522 ();
 b15zdnd00an1n01x5 FILLER_67_1524 ();
 b15zdnd11an1n16x5 FILLER_67_1540 ();
 b15zdnd11an1n04x5 FILLER_67_1556 ();
 b15zdnd00an1n01x5 FILLER_67_1560 ();
 b15zdnd11an1n04x5 FILLER_67_1579 ();
 b15zdnd00an1n02x5 FILLER_67_1583 ();
 b15zdnd11an1n08x5 FILLER_67_1590 ();
 b15zdnd00an1n02x5 FILLER_67_1598 ();
 b15zdnd11an1n08x5 FILLER_67_1606 ();
 b15zdnd11an1n04x5 FILLER_67_1614 ();
 b15zdnd00an1n02x5 FILLER_67_1618 ();
 b15zdnd00an1n01x5 FILLER_67_1620 ();
 b15zdnd11an1n16x5 FILLER_67_1638 ();
 b15zdnd11an1n08x5 FILLER_67_1654 ();
 b15zdnd00an1n02x5 FILLER_67_1662 ();
 b15zdnd00an1n01x5 FILLER_67_1664 ();
 b15zdnd11an1n64x5 FILLER_67_1675 ();
 b15zdnd11an1n08x5 FILLER_67_1739 ();
 b15zdnd00an1n01x5 FILLER_67_1747 ();
 b15zdnd11an1n64x5 FILLER_67_1774 ();
 b15zdnd11an1n64x5 FILLER_67_1838 ();
 b15zdnd11an1n64x5 FILLER_67_1902 ();
 b15zdnd11an1n64x5 FILLER_67_1966 ();
 b15zdnd11an1n64x5 FILLER_67_2030 ();
 b15zdnd11an1n64x5 FILLER_67_2094 ();
 b15zdnd11an1n64x5 FILLER_67_2158 ();
 b15zdnd11an1n32x5 FILLER_67_2222 ();
 b15zdnd11an1n16x5 FILLER_67_2254 ();
 b15zdnd11an1n08x5 FILLER_67_2270 ();
 b15zdnd11an1n04x5 FILLER_67_2278 ();
 b15zdnd00an1n02x5 FILLER_67_2282 ();
 b15zdnd11an1n16x5 FILLER_68_8 ();
 b15zdnd11an1n08x5 FILLER_68_24 ();
 b15zdnd11an1n04x5 FILLER_68_32 ();
 b15zdnd00an1n02x5 FILLER_68_36 ();
 b15zdnd11an1n32x5 FILLER_68_51 ();
 b15zdnd11an1n16x5 FILLER_68_83 ();
 b15zdnd11an1n08x5 FILLER_68_99 ();
 b15zdnd00an1n01x5 FILLER_68_107 ();
 b15zdnd11an1n16x5 FILLER_68_120 ();
 b15zdnd11an1n08x5 FILLER_68_136 ();
 b15zdnd00an1n01x5 FILLER_68_144 ();
 b15zdnd11an1n64x5 FILLER_68_158 ();
 b15zdnd11an1n16x5 FILLER_68_222 ();
 b15zdnd11an1n08x5 FILLER_68_238 ();
 b15zdnd11an1n04x5 FILLER_68_246 ();
 b15zdnd00an1n02x5 FILLER_68_250 ();
 b15zdnd11an1n16x5 FILLER_68_257 ();
 b15zdnd11an1n04x5 FILLER_68_273 ();
 b15zdnd00an1n01x5 FILLER_68_277 ();
 b15zdnd11an1n08x5 FILLER_68_287 ();
 b15zdnd11an1n32x5 FILLER_68_302 ();
 b15zdnd11an1n16x5 FILLER_68_334 ();
 b15zdnd11an1n08x5 FILLER_68_350 ();
 b15zdnd00an1n01x5 FILLER_68_358 ();
 b15zdnd11an1n64x5 FILLER_68_363 ();
 b15zdnd11an1n32x5 FILLER_68_427 ();
 b15zdnd11an1n04x5 FILLER_68_459 ();
 b15zdnd00an1n02x5 FILLER_68_463 ();
 b15zdnd11an1n16x5 FILLER_68_477 ();
 b15zdnd11an1n08x5 FILLER_68_493 ();
 b15zdnd11an1n08x5 FILLER_68_517 ();
 b15zdnd00an1n02x5 FILLER_68_525 ();
 b15zdnd00an1n01x5 FILLER_68_527 ();
 b15zdnd11an1n08x5 FILLER_68_544 ();
 b15zdnd00an1n02x5 FILLER_68_552 ();
 b15zdnd11an1n04x5 FILLER_68_565 ();
 b15zdnd11an1n16x5 FILLER_68_580 ();
 b15zdnd00an1n01x5 FILLER_68_596 ();
 b15zdnd11an1n04x5 FILLER_68_603 ();
 b15zdnd11an1n16x5 FILLER_68_612 ();
 b15zdnd11an1n32x5 FILLER_68_638 ();
 b15zdnd00an1n01x5 FILLER_68_670 ();
 b15zdnd11an1n16x5 FILLER_68_687 ();
 b15zdnd11an1n08x5 FILLER_68_703 ();
 b15zdnd11an1n04x5 FILLER_68_711 ();
 b15zdnd00an1n02x5 FILLER_68_715 ();
 b15zdnd00an1n01x5 FILLER_68_717 ();
 b15zdnd11an1n64x5 FILLER_68_726 ();
 b15zdnd11an1n16x5 FILLER_68_790 ();
 b15zdnd11an1n08x5 FILLER_68_806 ();
 b15zdnd11an1n04x5 FILLER_68_814 ();
 b15zdnd00an1n02x5 FILLER_68_818 ();
 b15zdnd11an1n32x5 FILLER_68_840 ();
 b15zdnd11an1n08x5 FILLER_68_877 ();
 b15zdnd11an1n04x5 FILLER_68_885 ();
 b15zdnd11an1n16x5 FILLER_68_892 ();
 b15zdnd11an1n08x5 FILLER_68_908 ();
 b15zdnd11an1n64x5 FILLER_68_921 ();
 b15zdnd11an1n32x5 FILLER_68_997 ();
 b15zdnd00an1n02x5 FILLER_68_1029 ();
 b15zdnd00an1n01x5 FILLER_68_1031 ();
 b15zdnd11an1n04x5 FILLER_68_1052 ();
 b15zdnd11an1n64x5 FILLER_68_1059 ();
 b15zdnd11an1n16x5 FILLER_68_1123 ();
 b15zdnd11an1n04x5 FILLER_68_1139 ();
 b15zdnd00an1n02x5 FILLER_68_1143 ();
 b15zdnd00an1n01x5 FILLER_68_1145 ();
 b15zdnd11an1n04x5 FILLER_68_1164 ();
 b15zdnd11an1n16x5 FILLER_68_1193 ();
 b15zdnd11an1n64x5 FILLER_68_1221 ();
 b15zdnd00an1n02x5 FILLER_68_1285 ();
 b15zdnd00an1n01x5 FILLER_68_1287 ();
 b15zdnd11an1n16x5 FILLER_68_1293 ();
 b15zdnd11an1n08x5 FILLER_68_1309 ();
 b15zdnd00an1n02x5 FILLER_68_1317 ();
 b15zdnd00an1n01x5 FILLER_68_1319 ();
 b15zdnd11an1n04x5 FILLER_68_1330 ();
 b15zdnd11an1n32x5 FILLER_68_1352 ();
 b15zdnd11an1n32x5 FILLER_68_1390 ();
 b15zdnd11an1n16x5 FILLER_68_1422 ();
 b15zdnd00an1n02x5 FILLER_68_1438 ();
 b15zdnd11an1n08x5 FILLER_68_1447 ();
 b15zdnd11an1n04x5 FILLER_68_1455 ();
 b15zdnd00an1n02x5 FILLER_68_1459 ();
 b15zdnd11an1n04x5 FILLER_68_1472 ();
 b15zdnd00an1n02x5 FILLER_68_1476 ();
 b15zdnd00an1n01x5 FILLER_68_1478 ();
 b15zdnd11an1n16x5 FILLER_68_1493 ();
 b15zdnd11an1n16x5 FILLER_68_1521 ();
 b15zdnd11an1n08x5 FILLER_68_1537 ();
 b15zdnd11an1n04x5 FILLER_68_1545 ();
 b15zdnd00an1n02x5 FILLER_68_1549 ();
 b15zdnd11an1n16x5 FILLER_68_1563 ();
 b15zdnd11an1n04x5 FILLER_68_1579 ();
 b15zdnd00an1n02x5 FILLER_68_1583 ();
 b15zdnd00an1n01x5 FILLER_68_1585 ();
 b15zdnd11an1n32x5 FILLER_68_1599 ();
 b15zdnd11an1n04x5 FILLER_68_1631 ();
 b15zdnd00an1n02x5 FILLER_68_1635 ();
 b15zdnd11an1n32x5 FILLER_68_1658 ();
 b15zdnd11an1n08x5 FILLER_68_1690 ();
 b15zdnd11an1n04x5 FILLER_68_1698 ();
 b15zdnd00an1n01x5 FILLER_68_1702 ();
 b15zdnd11an1n64x5 FILLER_68_1709 ();
 b15zdnd11an1n64x5 FILLER_68_1773 ();
 b15zdnd11an1n64x5 FILLER_68_1837 ();
 b15zdnd11an1n64x5 FILLER_68_1901 ();
 b15zdnd11an1n64x5 FILLER_68_1965 ();
 b15zdnd11an1n16x5 FILLER_68_2029 ();
 b15zdnd11an1n08x5 FILLER_68_2045 ();
 b15zdnd00an1n01x5 FILLER_68_2053 ();
 b15zdnd11an1n64x5 FILLER_68_2063 ();
 b15zdnd11an1n16x5 FILLER_68_2127 ();
 b15zdnd11an1n08x5 FILLER_68_2143 ();
 b15zdnd00an1n02x5 FILLER_68_2151 ();
 b15zdnd00an1n01x5 FILLER_68_2153 ();
 b15zdnd11an1n64x5 FILLER_68_2162 ();
 b15zdnd11an1n32x5 FILLER_68_2226 ();
 b15zdnd11an1n16x5 FILLER_68_2258 ();
 b15zdnd00an1n02x5 FILLER_68_2274 ();
 b15zdnd11an1n32x5 FILLER_69_0 ();
 b15zdnd11an1n16x5 FILLER_69_32 ();
 b15zdnd11an1n08x5 FILLER_69_48 ();
 b15zdnd00an1n01x5 FILLER_69_56 ();
 b15zdnd11an1n16x5 FILLER_69_74 ();
 b15zdnd11an1n08x5 FILLER_69_90 ();
 b15zdnd00an1n02x5 FILLER_69_98 ();
 b15zdnd00an1n01x5 FILLER_69_100 ();
 b15zdnd11an1n04x5 FILLER_69_105 ();
 b15zdnd11an1n32x5 FILLER_69_116 ();
 b15zdnd11an1n16x5 FILLER_69_148 ();
 b15zdnd00an1n01x5 FILLER_69_164 ();
 b15zdnd11an1n64x5 FILLER_69_171 ();
 b15zdnd11an1n64x5 FILLER_69_235 ();
 b15zdnd11an1n04x5 FILLER_69_299 ();
 b15zdnd00an1n02x5 FILLER_69_303 ();
 b15zdnd00an1n01x5 FILLER_69_305 ();
 b15zdnd11an1n04x5 FILLER_69_332 ();
 b15zdnd00an1n01x5 FILLER_69_336 ();
 b15zdnd11an1n64x5 FILLER_69_347 ();
 b15zdnd11an1n64x5 FILLER_69_411 ();
 b15zdnd11an1n64x5 FILLER_69_475 ();
 b15zdnd11an1n32x5 FILLER_69_539 ();
 b15zdnd11an1n16x5 FILLER_69_571 ();
 b15zdnd11an1n08x5 FILLER_69_587 ();
 b15zdnd11an1n04x5 FILLER_69_595 ();
 b15zdnd11an1n04x5 FILLER_69_611 ();
 b15zdnd00an1n02x5 FILLER_69_615 ();
 b15zdnd11an1n64x5 FILLER_69_625 ();
 b15zdnd11an1n64x5 FILLER_69_689 ();
 b15zdnd11an1n64x5 FILLER_69_753 ();
 b15zdnd00an1n02x5 FILLER_69_817 ();
 b15zdnd00an1n01x5 FILLER_69_819 ();
 b15zdnd11an1n64x5 FILLER_69_826 ();
 b15zdnd11an1n32x5 FILLER_69_890 ();
 b15zdnd00an1n02x5 FILLER_69_922 ();
 b15zdnd00an1n01x5 FILLER_69_924 ();
 b15zdnd11an1n32x5 FILLER_69_945 ();
 b15zdnd00an1n02x5 FILLER_69_977 ();
 b15zdnd11an1n08x5 FILLER_69_989 ();
 b15zdnd00an1n01x5 FILLER_69_997 ();
 b15zdnd11an1n04x5 FILLER_69_1003 ();
 b15zdnd11an1n32x5 FILLER_69_1013 ();
 b15zdnd11an1n04x5 FILLER_69_1045 ();
 b15zdnd00an1n02x5 FILLER_69_1049 ();
 b15zdnd00an1n01x5 FILLER_69_1051 ();
 b15zdnd11an1n16x5 FILLER_69_1074 ();
 b15zdnd00an1n02x5 FILLER_69_1090 ();
 b15zdnd00an1n01x5 FILLER_69_1092 ();
 b15zdnd11an1n64x5 FILLER_69_1116 ();
 b15zdnd11an1n08x5 FILLER_69_1180 ();
 b15zdnd11an1n04x5 FILLER_69_1188 ();
 b15zdnd00an1n02x5 FILLER_69_1192 ();
 b15zdnd11an1n04x5 FILLER_69_1206 ();
 b15zdnd11an1n32x5 FILLER_69_1227 ();
 b15zdnd11an1n16x5 FILLER_69_1259 ();
 b15zdnd11an1n08x5 FILLER_69_1275 ();
 b15zdnd00an1n02x5 FILLER_69_1283 ();
 b15zdnd11an1n32x5 FILLER_69_1293 ();
 b15zdnd00an1n01x5 FILLER_69_1325 ();
 b15zdnd11an1n08x5 FILLER_69_1332 ();
 b15zdnd00an1n01x5 FILLER_69_1340 ();
 b15zdnd11an1n64x5 FILLER_69_1348 ();
 b15zdnd11an1n32x5 FILLER_69_1412 ();
 b15zdnd11an1n16x5 FILLER_69_1444 ();
 b15zdnd11an1n08x5 FILLER_69_1460 ();
 b15zdnd00an1n02x5 FILLER_69_1468 ();
 b15zdnd00an1n01x5 FILLER_69_1470 ();
 b15zdnd11an1n32x5 FILLER_69_1492 ();
 b15zdnd11an1n16x5 FILLER_69_1524 ();
 b15zdnd11an1n04x5 FILLER_69_1540 ();
 b15zdnd00an1n02x5 FILLER_69_1544 ();
 b15zdnd00an1n01x5 FILLER_69_1546 ();
 b15zdnd11an1n32x5 FILLER_69_1553 ();
 b15zdnd00an1n01x5 FILLER_69_1585 ();
 b15zdnd11an1n64x5 FILLER_69_1590 ();
 b15zdnd00an1n02x5 FILLER_69_1654 ();
 b15zdnd00an1n01x5 FILLER_69_1656 ();
 b15zdnd11an1n32x5 FILLER_69_1662 ();
 b15zdnd11an1n08x5 FILLER_69_1694 ();
 b15zdnd00an1n02x5 FILLER_69_1702 ();
 b15zdnd11an1n64x5 FILLER_69_1724 ();
 b15zdnd11an1n64x5 FILLER_69_1788 ();
 b15zdnd11an1n64x5 FILLER_69_1852 ();
 b15zdnd00an1n02x5 FILLER_69_1916 ();
 b15zdnd11an1n16x5 FILLER_69_1926 ();
 b15zdnd11an1n08x5 FILLER_69_1942 ();
 b15zdnd11an1n04x5 FILLER_69_1950 ();
 b15zdnd00an1n01x5 FILLER_69_1954 ();
 b15zdnd11an1n16x5 FILLER_69_1971 ();
 b15zdnd11an1n32x5 FILLER_69_1994 ();
 b15zdnd11an1n16x5 FILLER_69_2026 ();
 b15zdnd11an1n08x5 FILLER_69_2042 ();
 b15zdnd00an1n02x5 FILLER_69_2050 ();
 b15zdnd11an1n08x5 FILLER_69_2064 ();
 b15zdnd00an1n02x5 FILLER_69_2072 ();
 b15zdnd00an1n01x5 FILLER_69_2074 ();
 b15zdnd11an1n04x5 FILLER_69_2090 ();
 b15zdnd11an1n16x5 FILLER_69_2098 ();
 b15zdnd00an1n01x5 FILLER_69_2114 ();
 b15zdnd11an1n04x5 FILLER_69_2120 ();
 b15zdnd11an1n04x5 FILLER_69_2130 ();
 b15zdnd11an1n32x5 FILLER_69_2143 ();
 b15zdnd11an1n08x5 FILLER_69_2175 ();
 b15zdnd00an1n01x5 FILLER_69_2183 ();
 b15zdnd11an1n64x5 FILLER_69_2192 ();
 b15zdnd11an1n16x5 FILLER_69_2256 ();
 b15zdnd11an1n08x5 FILLER_69_2272 ();
 b15zdnd11an1n04x5 FILLER_69_2280 ();
 b15zdnd11an1n32x5 FILLER_70_8 ();
 b15zdnd11an1n16x5 FILLER_70_40 ();
 b15zdnd11an1n04x5 FILLER_70_56 ();
 b15zdnd00an1n01x5 FILLER_70_60 ();
 b15zdnd11an1n16x5 FILLER_70_67 ();
 b15zdnd11an1n08x5 FILLER_70_83 ();
 b15zdnd11an1n04x5 FILLER_70_91 ();
 b15zdnd00an1n01x5 FILLER_70_95 ();
 b15zdnd11an1n64x5 FILLER_70_112 ();
 b15zdnd11an1n08x5 FILLER_70_176 ();
 b15zdnd11an1n04x5 FILLER_70_184 ();
 b15zdnd11an1n32x5 FILLER_70_193 ();
 b15zdnd11an1n08x5 FILLER_70_225 ();
 b15zdnd11an1n04x5 FILLER_70_233 ();
 b15zdnd00an1n02x5 FILLER_70_237 ();
 b15zdnd00an1n01x5 FILLER_70_239 ();
 b15zdnd11an1n64x5 FILLER_70_245 ();
 b15zdnd11an1n16x5 FILLER_70_309 ();
 b15zdnd11an1n08x5 FILLER_70_325 ();
 b15zdnd11an1n04x5 FILLER_70_333 ();
 b15zdnd00an1n01x5 FILLER_70_337 ();
 b15zdnd11an1n08x5 FILLER_70_356 ();
 b15zdnd11an1n04x5 FILLER_70_364 ();
 b15zdnd00an1n01x5 FILLER_70_368 ();
 b15zdnd11an1n64x5 FILLER_70_377 ();
 b15zdnd11an1n64x5 FILLER_70_441 ();
 b15zdnd11an1n64x5 FILLER_70_505 ();
 b15zdnd11an1n64x5 FILLER_70_569 ();
 b15zdnd11an1n64x5 FILLER_70_633 ();
 b15zdnd11an1n16x5 FILLER_70_697 ();
 b15zdnd11an1n04x5 FILLER_70_713 ();
 b15zdnd00an1n01x5 FILLER_70_717 ();
 b15zdnd11an1n64x5 FILLER_70_726 ();
 b15zdnd11an1n64x5 FILLER_70_790 ();
 b15zdnd11an1n64x5 FILLER_70_854 ();
 b15zdnd11an1n32x5 FILLER_70_918 ();
 b15zdnd11an1n08x5 FILLER_70_950 ();
 b15zdnd11an1n04x5 FILLER_70_958 ();
 b15zdnd00an1n02x5 FILLER_70_962 ();
 b15zdnd00an1n01x5 FILLER_70_964 ();
 b15zdnd11an1n04x5 FILLER_70_976 ();
 b15zdnd00an1n02x5 FILLER_70_980 ();
 b15zdnd11an1n64x5 FILLER_70_1002 ();
 b15zdnd11an1n32x5 FILLER_70_1066 ();
 b15zdnd11an1n08x5 FILLER_70_1098 ();
 b15zdnd11an1n04x5 FILLER_70_1106 ();
 b15zdnd00an1n02x5 FILLER_70_1110 ();
 b15zdnd11an1n16x5 FILLER_70_1116 ();
 b15zdnd00an1n01x5 FILLER_70_1132 ();
 b15zdnd11an1n04x5 FILLER_70_1142 ();
 b15zdnd11an1n16x5 FILLER_70_1172 ();
 b15zdnd11an1n08x5 FILLER_70_1188 ();
 b15zdnd00an1n02x5 FILLER_70_1196 ();
 b15zdnd11an1n64x5 FILLER_70_1208 ();
 b15zdnd11an1n32x5 FILLER_70_1272 ();
 b15zdnd11an1n04x5 FILLER_70_1304 ();
 b15zdnd00an1n02x5 FILLER_70_1308 ();
 b15zdnd00an1n01x5 FILLER_70_1310 ();
 b15zdnd11an1n32x5 FILLER_70_1327 ();
 b15zdnd00an1n02x5 FILLER_70_1359 ();
 b15zdnd00an1n01x5 FILLER_70_1361 ();
 b15zdnd11an1n04x5 FILLER_70_1370 ();
 b15zdnd11an1n08x5 FILLER_70_1381 ();
 b15zdnd00an1n02x5 FILLER_70_1389 ();
 b15zdnd00an1n01x5 FILLER_70_1391 ();
 b15zdnd11an1n64x5 FILLER_70_1396 ();
 b15zdnd11an1n16x5 FILLER_70_1472 ();
 b15zdnd11an1n04x5 FILLER_70_1488 ();
 b15zdnd00an1n02x5 FILLER_70_1492 ();
 b15zdnd00an1n01x5 FILLER_70_1494 ();
 b15zdnd11an1n16x5 FILLER_70_1505 ();
 b15zdnd11an1n08x5 FILLER_70_1521 ();
 b15zdnd00an1n02x5 FILLER_70_1529 ();
 b15zdnd11an1n64x5 FILLER_70_1541 ();
 b15zdnd11an1n32x5 FILLER_70_1605 ();
 b15zdnd11an1n04x5 FILLER_70_1637 ();
 b15zdnd00an1n02x5 FILLER_70_1641 ();
 b15zdnd11an1n32x5 FILLER_70_1653 ();
 b15zdnd11an1n08x5 FILLER_70_1685 ();
 b15zdnd00an1n02x5 FILLER_70_1693 ();
 b15zdnd11an1n08x5 FILLER_70_1699 ();
 b15zdnd11an1n04x5 FILLER_70_1707 ();
 b15zdnd00an1n01x5 FILLER_70_1711 ();
 b15zdnd11an1n32x5 FILLER_70_1717 ();
 b15zdnd11an1n16x5 FILLER_70_1749 ();
 b15zdnd11an1n04x5 FILLER_70_1765 ();
 b15zdnd11an1n16x5 FILLER_70_1792 ();
 b15zdnd11an1n16x5 FILLER_70_1834 ();
 b15zdnd11an1n04x5 FILLER_70_1850 ();
 b15zdnd11an1n16x5 FILLER_70_1860 ();
 b15zdnd11an1n08x5 FILLER_70_1876 ();
 b15zdnd11an1n04x5 FILLER_70_1884 ();
 b15zdnd00an1n02x5 FILLER_70_1888 ();
 b15zdnd00an1n01x5 FILLER_70_1890 ();
 b15zdnd11an1n04x5 FILLER_70_1899 ();
 b15zdnd11an1n08x5 FILLER_70_1915 ();
 b15zdnd00an1n01x5 FILLER_70_1923 ();
 b15zdnd11an1n08x5 FILLER_70_1934 ();
 b15zdnd11an1n04x5 FILLER_70_1942 ();
 b15zdnd00an1n02x5 FILLER_70_1946 ();
 b15zdnd00an1n01x5 FILLER_70_1948 ();
 b15zdnd11an1n04x5 FILLER_70_1965 ();
 b15zdnd11an1n08x5 FILLER_70_1990 ();
 b15zdnd11an1n04x5 FILLER_70_1998 ();
 b15zdnd00an1n02x5 FILLER_70_2002 ();
 b15zdnd11an1n04x5 FILLER_70_2011 ();
 b15zdnd11an1n04x5 FILLER_70_2022 ();
 b15zdnd00an1n02x5 FILLER_70_2026 ();
 b15zdnd00an1n01x5 FILLER_70_2028 ();
 b15zdnd11an1n08x5 FILLER_70_2044 ();
 b15zdnd00an1n01x5 FILLER_70_2052 ();
 b15zdnd11an1n16x5 FILLER_70_2057 ();
 b15zdnd11an1n04x5 FILLER_70_2073 ();
 b15zdnd00an1n01x5 FILLER_70_2077 ();
 b15zdnd11an1n04x5 FILLER_70_2091 ();
 b15zdnd11an1n08x5 FILLER_70_2101 ();
 b15zdnd00an1n02x5 FILLER_70_2109 ();
 b15zdnd11an1n04x5 FILLER_70_2124 ();
 b15zdnd11an1n04x5 FILLER_70_2133 ();
 b15zdnd00an1n01x5 FILLER_70_2137 ();
 b15zdnd11an1n08x5 FILLER_70_2146 ();
 b15zdnd11an1n08x5 FILLER_70_2162 ();
 b15zdnd11an1n04x5 FILLER_70_2170 ();
 b15zdnd00an1n02x5 FILLER_70_2174 ();
 b15zdnd11an1n04x5 FILLER_70_2180 ();
 b15zdnd11an1n64x5 FILLER_70_2195 ();
 b15zdnd11an1n16x5 FILLER_70_2259 ();
 b15zdnd00an1n01x5 FILLER_70_2275 ();
 b15zdnd11an1n64x5 FILLER_71_0 ();
 b15zdnd11an1n16x5 FILLER_71_64 ();
 b15zdnd11an1n04x5 FILLER_71_80 ();
 b15zdnd00an1n02x5 FILLER_71_84 ();
 b15zdnd11an1n16x5 FILLER_71_97 ();
 b15zdnd11an1n08x5 FILLER_71_113 ();
 b15zdnd00an1n02x5 FILLER_71_121 ();
 b15zdnd00an1n01x5 FILLER_71_123 ();
 b15zdnd11an1n04x5 FILLER_71_130 ();
 b15zdnd11an1n32x5 FILLER_71_139 ();
 b15zdnd11an1n08x5 FILLER_71_171 ();
 b15zdnd11an1n04x5 FILLER_71_179 ();
 b15zdnd00an1n02x5 FILLER_71_183 ();
 b15zdnd00an1n01x5 FILLER_71_185 ();
 b15zdnd11an1n08x5 FILLER_71_190 ();
 b15zdnd11an1n04x5 FILLER_71_198 ();
 b15zdnd00an1n02x5 FILLER_71_202 ();
 b15zdnd00an1n01x5 FILLER_71_204 ();
 b15zdnd11an1n08x5 FILLER_71_217 ();
 b15zdnd00an1n02x5 FILLER_71_225 ();
 b15zdnd11an1n04x5 FILLER_71_239 ();
 b15zdnd11an1n08x5 FILLER_71_248 ();
 b15zdnd00an1n01x5 FILLER_71_256 ();
 b15zdnd11an1n04x5 FILLER_71_273 ();
 b15zdnd11an1n04x5 FILLER_71_283 ();
 b15zdnd11an1n32x5 FILLER_71_293 ();
 b15zdnd11an1n16x5 FILLER_71_325 ();
 b15zdnd11an1n08x5 FILLER_71_341 ();
 b15zdnd00an1n02x5 FILLER_71_349 ();
 b15zdnd00an1n01x5 FILLER_71_351 ();
 b15zdnd11an1n16x5 FILLER_71_361 ();
 b15zdnd11an1n08x5 FILLER_71_377 ();
 b15zdnd00an1n01x5 FILLER_71_385 ();
 b15zdnd11an1n04x5 FILLER_71_399 ();
 b15zdnd11an1n64x5 FILLER_71_408 ();
 b15zdnd11an1n64x5 FILLER_71_472 ();
 b15zdnd11an1n64x5 FILLER_71_536 ();
 b15zdnd11an1n64x5 FILLER_71_600 ();
 b15zdnd11an1n64x5 FILLER_71_664 ();
 b15zdnd11an1n32x5 FILLER_71_728 ();
 b15zdnd11an1n16x5 FILLER_71_760 ();
 b15zdnd00an1n01x5 FILLER_71_776 ();
 b15zdnd11an1n32x5 FILLER_71_797 ();
 b15zdnd11an1n08x5 FILLER_71_829 ();
 b15zdnd00an1n02x5 FILLER_71_837 ();
 b15zdnd00an1n01x5 FILLER_71_839 ();
 b15zdnd11an1n32x5 FILLER_71_852 ();
 b15zdnd11an1n04x5 FILLER_71_884 ();
 b15zdnd00an1n01x5 FILLER_71_888 ();
 b15zdnd11an1n16x5 FILLER_71_897 ();
 b15zdnd11an1n04x5 FILLER_71_913 ();
 b15zdnd11an1n64x5 FILLER_71_929 ();
 b15zdnd11an1n64x5 FILLER_71_993 ();
 b15zdnd11an1n32x5 FILLER_71_1057 ();
 b15zdnd11an1n16x5 FILLER_71_1089 ();
 b15zdnd11an1n08x5 FILLER_71_1105 ();
 b15zdnd11an1n04x5 FILLER_71_1113 ();
 b15zdnd11an1n64x5 FILLER_71_1127 ();
 b15zdnd11an1n64x5 FILLER_71_1191 ();
 b15zdnd11an1n32x5 FILLER_71_1255 ();
 b15zdnd11an1n16x5 FILLER_71_1287 ();
 b15zdnd11an1n64x5 FILLER_71_1319 ();
 b15zdnd00an1n01x5 FILLER_71_1383 ();
 b15zdnd11an1n04x5 FILLER_71_1389 ();
 b15zdnd11an1n08x5 FILLER_71_1407 ();
 b15zdnd00an1n01x5 FILLER_71_1415 ();
 b15zdnd11an1n04x5 FILLER_71_1431 ();
 b15zdnd11an1n08x5 FILLER_71_1447 ();
 b15zdnd11an1n08x5 FILLER_71_1470 ();
 b15zdnd00an1n02x5 FILLER_71_1478 ();
 b15zdnd11an1n16x5 FILLER_71_1488 ();
 b15zdnd11an1n08x5 FILLER_71_1504 ();
 b15zdnd11an1n64x5 FILLER_71_1520 ();
 b15zdnd11an1n32x5 FILLER_71_1584 ();
 b15zdnd11an1n04x5 FILLER_71_1616 ();
 b15zdnd00an1n02x5 FILLER_71_1620 ();
 b15zdnd00an1n01x5 FILLER_71_1622 ();
 b15zdnd11an1n16x5 FILLER_71_1628 ();
 b15zdnd11an1n04x5 FILLER_71_1644 ();
 b15zdnd11an1n64x5 FILLER_71_1653 ();
 b15zdnd11an1n32x5 FILLER_71_1717 ();
 b15zdnd11an1n08x5 FILLER_71_1749 ();
 b15zdnd11an1n04x5 FILLER_71_1757 ();
 b15zdnd00an1n02x5 FILLER_71_1761 ();
 b15zdnd11an1n08x5 FILLER_71_1781 ();
 b15zdnd00an1n02x5 FILLER_71_1789 ();
 b15zdnd00an1n01x5 FILLER_71_1791 ();
 b15zdnd11an1n08x5 FILLER_71_1804 ();
 b15zdnd00an1n02x5 FILLER_71_1812 ();
 b15zdnd11an1n16x5 FILLER_71_1845 ();
 b15zdnd11an1n08x5 FILLER_71_1861 ();
 b15zdnd11an1n08x5 FILLER_71_1885 ();
 b15zdnd00an1n02x5 FILLER_71_1893 ();
 b15zdnd00an1n01x5 FILLER_71_1895 ();
 b15zdnd11an1n32x5 FILLER_71_1903 ();
 b15zdnd11an1n16x5 FILLER_71_1935 ();
 b15zdnd11an1n04x5 FILLER_71_1951 ();
 b15zdnd11an1n16x5 FILLER_71_1960 ();
 b15zdnd11an1n04x5 FILLER_71_1976 ();
 b15zdnd11an1n16x5 FILLER_71_1985 ();
 b15zdnd11an1n08x5 FILLER_71_2001 ();
 b15zdnd11an1n32x5 FILLER_71_2014 ();
 b15zdnd11an1n16x5 FILLER_71_2046 ();
 b15zdnd11an1n08x5 FILLER_71_2062 ();
 b15zdnd11an1n04x5 FILLER_71_2070 ();
 b15zdnd00an1n02x5 FILLER_71_2074 ();
 b15zdnd11an1n32x5 FILLER_71_2083 ();
 b15zdnd11an1n08x5 FILLER_71_2115 ();
 b15zdnd11an1n08x5 FILLER_71_2129 ();
 b15zdnd00an1n02x5 FILLER_71_2137 ();
 b15zdnd00an1n01x5 FILLER_71_2139 ();
 b15zdnd11an1n16x5 FILLER_71_2146 ();
 b15zdnd11an1n08x5 FILLER_71_2162 ();
 b15zdnd11an1n04x5 FILLER_71_2170 ();
 b15zdnd00an1n02x5 FILLER_71_2174 ();
 b15zdnd00an1n01x5 FILLER_71_2176 ();
 b15zdnd11an1n04x5 FILLER_71_2183 ();
 b15zdnd00an1n01x5 FILLER_71_2187 ();
 b15zdnd11an1n04x5 FILLER_71_2193 ();
 b15zdnd11an1n64x5 FILLER_71_2215 ();
 b15zdnd11an1n04x5 FILLER_71_2279 ();
 b15zdnd00an1n01x5 FILLER_71_2283 ();
 b15zdnd11an1n32x5 FILLER_72_8 ();
 b15zdnd11an1n08x5 FILLER_72_40 ();
 b15zdnd11an1n04x5 FILLER_72_48 ();
 b15zdnd00an1n01x5 FILLER_72_52 ();
 b15zdnd11an1n32x5 FILLER_72_67 ();
 b15zdnd11an1n16x5 FILLER_72_99 ();
 b15zdnd11an1n08x5 FILLER_72_115 ();
 b15zdnd11an1n04x5 FILLER_72_123 ();
 b15zdnd00an1n02x5 FILLER_72_127 ();
 b15zdnd00an1n01x5 FILLER_72_129 ();
 b15zdnd11an1n32x5 FILLER_72_137 ();
 b15zdnd00an1n02x5 FILLER_72_169 ();
 b15zdnd00an1n01x5 FILLER_72_171 ();
 b15zdnd11an1n04x5 FILLER_72_180 ();
 b15zdnd11an1n04x5 FILLER_72_198 ();
 b15zdnd00an1n01x5 FILLER_72_202 ();
 b15zdnd11an1n16x5 FILLER_72_231 ();
 b15zdnd11an1n08x5 FILLER_72_247 ();
 b15zdnd11an1n04x5 FILLER_72_255 ();
 b15zdnd00an1n02x5 FILLER_72_259 ();
 b15zdnd11an1n16x5 FILLER_72_268 ();
 b15zdnd11an1n08x5 FILLER_72_284 ();
 b15zdnd00an1n01x5 FILLER_72_292 ();
 b15zdnd11an1n16x5 FILLER_72_301 ();
 b15zdnd11an1n04x5 FILLER_72_317 ();
 b15zdnd00an1n01x5 FILLER_72_321 ();
 b15zdnd11an1n04x5 FILLER_72_331 ();
 b15zdnd11an1n08x5 FILLER_72_339 ();
 b15zdnd11an1n04x5 FILLER_72_354 ();
 b15zdnd11an1n16x5 FILLER_72_384 ();
 b15zdnd00an1n01x5 FILLER_72_400 ();
 b15zdnd11an1n04x5 FILLER_72_407 ();
 b15zdnd11an1n64x5 FILLER_72_418 ();
 b15zdnd11an1n64x5 FILLER_72_482 ();
 b15zdnd11an1n64x5 FILLER_72_546 ();
 b15zdnd11an1n64x5 FILLER_72_610 ();
 b15zdnd11an1n32x5 FILLER_72_674 ();
 b15zdnd11an1n08x5 FILLER_72_706 ();
 b15zdnd11an1n04x5 FILLER_72_714 ();
 b15zdnd11an1n32x5 FILLER_72_726 ();
 b15zdnd11an1n16x5 FILLER_72_758 ();
 b15zdnd00an1n01x5 FILLER_72_774 ();
 b15zdnd11an1n64x5 FILLER_72_801 ();
 b15zdnd11an1n16x5 FILLER_72_865 ();
 b15zdnd11an1n04x5 FILLER_72_881 ();
 b15zdnd00an1n01x5 FILLER_72_885 ();
 b15zdnd11an1n08x5 FILLER_72_890 ();
 b15zdnd00an1n02x5 FILLER_72_898 ();
 b15zdnd00an1n01x5 FILLER_72_900 ();
 b15zdnd11an1n64x5 FILLER_72_926 ();
 b15zdnd11an1n64x5 FILLER_72_990 ();
 b15zdnd11an1n16x5 FILLER_72_1054 ();
 b15zdnd11an1n08x5 FILLER_72_1070 ();
 b15zdnd11an1n32x5 FILLER_72_1082 ();
 b15zdnd11an1n16x5 FILLER_72_1114 ();
 b15zdnd11an1n08x5 FILLER_72_1130 ();
 b15zdnd11an1n04x5 FILLER_72_1138 ();
 b15zdnd11an1n64x5 FILLER_72_1168 ();
 b15zdnd11an1n16x5 FILLER_72_1232 ();
 b15zdnd11an1n08x5 FILLER_72_1248 ();
 b15zdnd11an1n04x5 FILLER_72_1256 ();
 b15zdnd00an1n01x5 FILLER_72_1260 ();
 b15zdnd11an1n04x5 FILLER_72_1292 ();
 b15zdnd11an1n04x5 FILLER_72_1328 ();
 b15zdnd11an1n08x5 FILLER_72_1340 ();
 b15zdnd11an1n04x5 FILLER_72_1348 ();
 b15zdnd00an1n01x5 FILLER_72_1352 ();
 b15zdnd11an1n32x5 FILLER_72_1367 ();
 b15zdnd11an1n04x5 FILLER_72_1399 ();
 b15zdnd00an1n02x5 FILLER_72_1403 ();
 b15zdnd00an1n01x5 FILLER_72_1405 ();
 b15zdnd11an1n04x5 FILLER_72_1418 ();
 b15zdnd11an1n16x5 FILLER_72_1427 ();
 b15zdnd11an1n08x5 FILLER_72_1443 ();
 b15zdnd11an1n04x5 FILLER_72_1451 ();
 b15zdnd00an1n02x5 FILLER_72_1455 ();
 b15zdnd11an1n16x5 FILLER_72_1464 ();
 b15zdnd00an1n01x5 FILLER_72_1480 ();
 b15zdnd11an1n16x5 FILLER_72_1488 ();
 b15zdnd11an1n04x5 FILLER_72_1504 ();
 b15zdnd00an1n01x5 FILLER_72_1508 ();
 b15zdnd11an1n32x5 FILLER_72_1522 ();
 b15zdnd11an1n08x5 FILLER_72_1554 ();
 b15zdnd00an1n01x5 FILLER_72_1562 ();
 b15zdnd11an1n04x5 FILLER_72_1572 ();
 b15zdnd11an1n08x5 FILLER_72_1593 ();
 b15zdnd11an1n04x5 FILLER_72_1601 ();
 b15zdnd00an1n02x5 FILLER_72_1605 ();
 b15zdnd00an1n01x5 FILLER_72_1607 ();
 b15zdnd11an1n08x5 FILLER_72_1614 ();
 b15zdnd00an1n01x5 FILLER_72_1622 ();
 b15zdnd11an1n04x5 FILLER_72_1635 ();
 b15zdnd11an1n64x5 FILLER_72_1660 ();
 b15zdnd11an1n64x5 FILLER_72_1724 ();
 b15zdnd11an1n08x5 FILLER_72_1788 ();
 b15zdnd00an1n02x5 FILLER_72_1796 ();
 b15zdnd11an1n04x5 FILLER_72_1816 ();
 b15zdnd00an1n01x5 FILLER_72_1820 ();
 b15zdnd11an1n08x5 FILLER_72_1839 ();
 b15zdnd11an1n16x5 FILLER_72_1859 ();
 b15zdnd11an1n04x5 FILLER_72_1875 ();
 b15zdnd00an1n02x5 FILLER_72_1879 ();
 b15zdnd00an1n01x5 FILLER_72_1881 ();
 b15zdnd11an1n64x5 FILLER_72_1900 ();
 b15zdnd11an1n32x5 FILLER_72_1964 ();
 b15zdnd11an1n08x5 FILLER_72_1996 ();
 b15zdnd11an1n32x5 FILLER_72_2015 ();
 b15zdnd11an1n08x5 FILLER_72_2047 ();
 b15zdnd11an1n04x5 FILLER_72_2055 ();
 b15zdnd00an1n01x5 FILLER_72_2059 ();
 b15zdnd11an1n64x5 FILLER_72_2064 ();
 b15zdnd11an1n16x5 FILLER_72_2128 ();
 b15zdnd11an1n08x5 FILLER_72_2144 ();
 b15zdnd00an1n02x5 FILLER_72_2152 ();
 b15zdnd11an1n64x5 FILLER_72_2162 ();
 b15zdnd11an1n32x5 FILLER_72_2226 ();
 b15zdnd11an1n16x5 FILLER_72_2258 ();
 b15zdnd00an1n02x5 FILLER_72_2274 ();
 b15zdnd11an1n32x5 FILLER_73_0 ();
 b15zdnd11an1n04x5 FILLER_73_32 ();
 b15zdnd11an1n04x5 FILLER_73_42 ();
 b15zdnd11an1n08x5 FILLER_73_60 ();
 b15zdnd00an1n02x5 FILLER_73_68 ();
 b15zdnd00an1n01x5 FILLER_73_70 ();
 b15zdnd11an1n08x5 FILLER_73_89 ();
 b15zdnd11an1n16x5 FILLER_73_108 ();
 b15zdnd11an1n08x5 FILLER_73_124 ();
 b15zdnd00an1n01x5 FILLER_73_132 ();
 b15zdnd11an1n16x5 FILLER_73_138 ();
 b15zdnd11an1n08x5 FILLER_73_154 ();
 b15zdnd11an1n04x5 FILLER_73_162 ();
 b15zdnd00an1n02x5 FILLER_73_166 ();
 b15zdnd00an1n01x5 FILLER_73_168 ();
 b15zdnd11an1n32x5 FILLER_73_175 ();
 b15zdnd11an1n04x5 FILLER_73_207 ();
 b15zdnd00an1n02x5 FILLER_73_211 ();
 b15zdnd00an1n01x5 FILLER_73_213 ();
 b15zdnd11an1n16x5 FILLER_73_222 ();
 b15zdnd11an1n08x5 FILLER_73_238 ();
 b15zdnd00an1n02x5 FILLER_73_246 ();
 b15zdnd00an1n01x5 FILLER_73_248 ();
 b15zdnd11an1n04x5 FILLER_73_263 ();
 b15zdnd11an1n32x5 FILLER_73_273 ();
 b15zdnd11an1n16x5 FILLER_73_305 ();
 b15zdnd11an1n08x5 FILLER_73_321 ();
 b15zdnd00an1n02x5 FILLER_73_329 ();
 b15zdnd00an1n01x5 FILLER_73_331 ();
 b15zdnd11an1n32x5 FILLER_73_339 ();
 b15zdnd11an1n08x5 FILLER_73_371 ();
 b15zdnd11an1n04x5 FILLER_73_379 ();
 b15zdnd00an1n02x5 FILLER_73_383 ();
 b15zdnd11an1n08x5 FILLER_73_394 ();
 b15zdnd00an1n01x5 FILLER_73_402 ();
 b15zdnd11an1n64x5 FILLER_73_409 ();
 b15zdnd11an1n08x5 FILLER_73_473 ();
 b15zdnd11an1n04x5 FILLER_73_481 ();
 b15zdnd00an1n01x5 FILLER_73_485 ();
 b15zdnd11an1n04x5 FILLER_73_504 ();
 b15zdnd11an1n64x5 FILLER_73_524 ();
 b15zdnd11an1n64x5 FILLER_73_588 ();
 b15zdnd11an1n32x5 FILLER_73_652 ();
 b15zdnd11an1n16x5 FILLER_73_684 ();
 b15zdnd11an1n08x5 FILLER_73_700 ();
 b15zdnd11an1n04x5 FILLER_73_708 ();
 b15zdnd11an1n04x5 FILLER_73_717 ();
 b15zdnd11an1n08x5 FILLER_73_729 ();
 b15zdnd11an1n04x5 FILLER_73_737 ();
 b15zdnd00an1n02x5 FILLER_73_741 ();
 b15zdnd11an1n64x5 FILLER_73_748 ();
 b15zdnd11an1n32x5 FILLER_73_812 ();
 b15zdnd11an1n16x5 FILLER_73_844 ();
 b15zdnd11an1n04x5 FILLER_73_860 ();
 b15zdnd00an1n02x5 FILLER_73_864 ();
 b15zdnd11an1n04x5 FILLER_73_877 ();
 b15zdnd00an1n02x5 FILLER_73_881 ();
 b15zdnd00an1n01x5 FILLER_73_883 ();
 b15zdnd11an1n04x5 FILLER_73_889 ();
 b15zdnd11an1n64x5 FILLER_73_913 ();
 b15zdnd11an1n64x5 FILLER_73_977 ();
 b15zdnd11an1n04x5 FILLER_73_1041 ();
 b15zdnd00an1n02x5 FILLER_73_1045 ();
 b15zdnd11an1n04x5 FILLER_73_1067 ();
 b15zdnd11an1n16x5 FILLER_73_1076 ();
 b15zdnd00an1n02x5 FILLER_73_1092 ();
 b15zdnd11an1n04x5 FILLER_73_1098 ();
 b15zdnd11an1n04x5 FILLER_73_1133 ();
 b15zdnd11an1n32x5 FILLER_73_1149 ();
 b15zdnd11an1n08x5 FILLER_73_1181 ();
 b15zdnd11an1n64x5 FILLER_73_1208 ();
 b15zdnd11an1n16x5 FILLER_73_1272 ();
 b15zdnd11an1n08x5 FILLER_73_1288 ();
 b15zdnd11an1n04x5 FILLER_73_1296 ();
 b15zdnd00an1n02x5 FILLER_73_1300 ();
 b15zdnd11an1n08x5 FILLER_73_1318 ();
 b15zdnd11an1n04x5 FILLER_73_1326 ();
 b15zdnd00an1n01x5 FILLER_73_1330 ();
 b15zdnd11an1n04x5 FILLER_73_1337 ();
 b15zdnd11an1n64x5 FILLER_73_1353 ();
 b15zdnd00an1n02x5 FILLER_73_1417 ();
 b15zdnd00an1n01x5 FILLER_73_1419 ();
 b15zdnd11an1n16x5 FILLER_73_1432 ();
 b15zdnd11an1n08x5 FILLER_73_1448 ();
 b15zdnd11an1n32x5 FILLER_73_1476 ();
 b15zdnd11an1n04x5 FILLER_73_1508 ();
 b15zdnd11an1n32x5 FILLER_73_1516 ();
 b15zdnd00an1n01x5 FILLER_73_1548 ();
 b15zdnd11an1n04x5 FILLER_73_1554 ();
 b15zdnd11an1n04x5 FILLER_73_1576 ();
 b15zdnd00an1n02x5 FILLER_73_1580 ();
 b15zdnd00an1n01x5 FILLER_73_1582 ();
 b15zdnd11an1n16x5 FILLER_73_1599 ();
 b15zdnd11an1n08x5 FILLER_73_1615 ();
 b15zdnd11an1n16x5 FILLER_73_1630 ();
 b15zdnd00an1n02x5 FILLER_73_1646 ();
 b15zdnd00an1n01x5 FILLER_73_1648 ();
 b15zdnd11an1n16x5 FILLER_73_1669 ();
 b15zdnd11an1n08x5 FILLER_73_1685 ();
 b15zdnd00an1n02x5 FILLER_73_1693 ();
 b15zdnd11an1n04x5 FILLER_73_1700 ();
 b15zdnd00an1n02x5 FILLER_73_1704 ();
 b15zdnd11an1n32x5 FILLER_73_1710 ();
 b15zdnd00an1n02x5 FILLER_73_1742 ();
 b15zdnd00an1n01x5 FILLER_73_1744 ();
 b15zdnd11an1n04x5 FILLER_73_1765 ();
 b15zdnd11an1n04x5 FILLER_73_1792 ();
 b15zdnd00an1n01x5 FILLER_73_1796 ();
 b15zdnd11an1n64x5 FILLER_73_1803 ();
 b15zdnd11an1n16x5 FILLER_73_1867 ();
 b15zdnd11an1n08x5 FILLER_73_1883 ();
 b15zdnd11an1n04x5 FILLER_73_1895 ();
 b15zdnd00an1n02x5 FILLER_73_1899 ();
 b15zdnd11an1n08x5 FILLER_73_1906 ();
 b15zdnd11an1n04x5 FILLER_73_1914 ();
 b15zdnd00an1n01x5 FILLER_73_1918 ();
 b15zdnd11an1n04x5 FILLER_73_1929 ();
 b15zdnd11an1n04x5 FILLER_73_1937 ();
 b15zdnd00an1n01x5 FILLER_73_1941 ();
 b15zdnd11an1n16x5 FILLER_73_1952 ();
 b15zdnd11an1n08x5 FILLER_73_1968 ();
 b15zdnd11an1n04x5 FILLER_73_1976 ();
 b15zdnd00an1n02x5 FILLER_73_1980 ();
 b15zdnd00an1n01x5 FILLER_73_1982 ();
 b15zdnd11an1n16x5 FILLER_73_1991 ();
 b15zdnd11an1n04x5 FILLER_73_2007 ();
 b15zdnd00an1n01x5 FILLER_73_2011 ();
 b15zdnd11an1n04x5 FILLER_73_2017 ();
 b15zdnd11an1n08x5 FILLER_73_2034 ();
 b15zdnd11an1n04x5 FILLER_73_2042 ();
 b15zdnd00an1n02x5 FILLER_73_2046 ();
 b15zdnd00an1n01x5 FILLER_73_2048 ();
 b15zdnd11an1n04x5 FILLER_73_2058 ();
 b15zdnd11an1n04x5 FILLER_73_2066 ();
 b15zdnd11an1n16x5 FILLER_73_2082 ();
 b15zdnd00an1n01x5 FILLER_73_2098 ();
 b15zdnd11an1n64x5 FILLER_73_2107 ();
 b15zdnd11an1n16x5 FILLER_73_2187 ();
 b15zdnd00an1n02x5 FILLER_73_2203 ();
 b15zdnd11an1n64x5 FILLER_73_2209 ();
 b15zdnd11an1n08x5 FILLER_73_2273 ();
 b15zdnd00an1n02x5 FILLER_73_2281 ();
 b15zdnd00an1n01x5 FILLER_73_2283 ();
 b15zdnd11an1n32x5 FILLER_74_8 ();
 b15zdnd11an1n04x5 FILLER_74_40 ();
 b15zdnd11an1n16x5 FILLER_74_49 ();
 b15zdnd11an1n04x5 FILLER_74_65 ();
 b15zdnd11an1n16x5 FILLER_74_78 ();
 b15zdnd00an1n01x5 FILLER_74_94 ();
 b15zdnd11an1n64x5 FILLER_74_106 ();
 b15zdnd00an1n01x5 FILLER_74_170 ();
 b15zdnd11an1n64x5 FILLER_74_176 ();
 b15zdnd11an1n32x5 FILLER_74_240 ();
 b15zdnd11an1n16x5 FILLER_74_272 ();
 b15zdnd11an1n08x5 FILLER_74_288 ();
 b15zdnd11an1n04x5 FILLER_74_296 ();
 b15zdnd11an1n32x5 FILLER_74_310 ();
 b15zdnd00an1n01x5 FILLER_74_342 ();
 b15zdnd11an1n16x5 FILLER_74_355 ();
 b15zdnd11an1n08x5 FILLER_74_371 ();
 b15zdnd11an1n04x5 FILLER_74_379 ();
 b15zdnd00an1n02x5 FILLER_74_383 ();
 b15zdnd11an1n64x5 FILLER_74_400 ();
 b15zdnd11an1n08x5 FILLER_74_464 ();
 b15zdnd11an1n08x5 FILLER_74_503 ();
 b15zdnd11an1n04x5 FILLER_74_511 ();
 b15zdnd00an1n02x5 FILLER_74_515 ();
 b15zdnd11an1n04x5 FILLER_74_524 ();
 b15zdnd11an1n04x5 FILLER_74_540 ();
 b15zdnd11an1n16x5 FILLER_74_556 ();
 b15zdnd00an1n02x5 FILLER_74_572 ();
 b15zdnd11an1n16x5 FILLER_74_584 ();
 b15zdnd11an1n08x5 FILLER_74_600 ();
 b15zdnd00an1n01x5 FILLER_74_608 ();
 b15zdnd11an1n04x5 FILLER_74_619 ();
 b15zdnd11an1n08x5 FILLER_74_628 ();
 b15zdnd00an1n01x5 FILLER_74_636 ();
 b15zdnd11an1n04x5 FILLER_74_644 ();
 b15zdnd11an1n04x5 FILLER_74_670 ();
 b15zdnd11an1n16x5 FILLER_74_682 ();
 b15zdnd00an1n01x5 FILLER_74_698 ();
 b15zdnd11an1n04x5 FILLER_74_704 ();
 b15zdnd00an1n02x5 FILLER_74_715 ();
 b15zdnd00an1n01x5 FILLER_74_717 ();
 b15zdnd11an1n04x5 FILLER_74_726 ();
 b15zdnd00an1n02x5 FILLER_74_730 ();
 b15zdnd11an1n04x5 FILLER_74_739 ();
 b15zdnd00an1n02x5 FILLER_74_743 ();
 b15zdnd00an1n01x5 FILLER_74_745 ();
 b15zdnd11an1n08x5 FILLER_74_756 ();
 b15zdnd11an1n04x5 FILLER_74_764 ();
 b15zdnd00an1n02x5 FILLER_74_768 ();
 b15zdnd11an1n04x5 FILLER_74_791 ();
 b15zdnd11an1n04x5 FILLER_74_807 ();
 b15zdnd11an1n32x5 FILLER_74_830 ();
 b15zdnd11an1n04x5 FILLER_74_862 ();
 b15zdnd00an1n02x5 FILLER_74_866 ();
 b15zdnd00an1n01x5 FILLER_74_868 ();
 b15zdnd11an1n08x5 FILLER_74_884 ();
 b15zdnd11an1n04x5 FILLER_74_892 ();
 b15zdnd00an1n02x5 FILLER_74_896 ();
 b15zdnd00an1n01x5 FILLER_74_898 ();
 b15zdnd11an1n64x5 FILLER_74_902 ();
 b15zdnd00an1n01x5 FILLER_74_966 ();
 b15zdnd11an1n04x5 FILLER_74_987 ();
 b15zdnd11an1n64x5 FILLER_74_1022 ();
 b15zdnd11an1n64x5 FILLER_74_1086 ();
 b15zdnd11an1n32x5 FILLER_74_1150 ();
 b15zdnd11an1n16x5 FILLER_74_1182 ();
 b15zdnd11an1n04x5 FILLER_74_1198 ();
 b15zdnd00an1n02x5 FILLER_74_1202 ();
 b15zdnd00an1n01x5 FILLER_74_1204 ();
 b15zdnd11an1n64x5 FILLER_74_1209 ();
 b15zdnd11an1n64x5 FILLER_74_1273 ();
 b15zdnd11an1n04x5 FILLER_74_1342 ();
 b15zdnd11an1n64x5 FILLER_74_1354 ();
 b15zdnd11an1n32x5 FILLER_74_1418 ();
 b15zdnd11an1n16x5 FILLER_74_1450 ();
 b15zdnd11an1n08x5 FILLER_74_1466 ();
 b15zdnd11an1n04x5 FILLER_74_1474 ();
 b15zdnd00an1n02x5 FILLER_74_1478 ();
 b15zdnd00an1n01x5 FILLER_74_1480 ();
 b15zdnd11an1n32x5 FILLER_74_1487 ();
 b15zdnd11an1n16x5 FILLER_74_1519 ();
 b15zdnd11an1n08x5 FILLER_74_1535 ();
 b15zdnd11an1n04x5 FILLER_74_1543 ();
 b15zdnd00an1n02x5 FILLER_74_1547 ();
 b15zdnd11an1n04x5 FILLER_74_1561 ();
 b15zdnd11an1n16x5 FILLER_74_1585 ();
 b15zdnd11an1n08x5 FILLER_74_1601 ();
 b15zdnd00an1n02x5 FILLER_74_1609 ();
 b15zdnd11an1n32x5 FILLER_74_1631 ();
 b15zdnd11an1n16x5 FILLER_74_1663 ();
 b15zdnd11an1n08x5 FILLER_74_1679 ();
 b15zdnd11an1n04x5 FILLER_74_1687 ();
 b15zdnd00an1n01x5 FILLER_74_1691 ();
 b15zdnd11an1n64x5 FILLER_74_1712 ();
 b15zdnd11an1n16x5 FILLER_74_1776 ();
 b15zdnd11an1n04x5 FILLER_74_1792 ();
 b15zdnd00an1n02x5 FILLER_74_1796 ();
 b15zdnd11an1n64x5 FILLER_74_1803 ();
 b15zdnd11an1n16x5 FILLER_74_1867 ();
 b15zdnd11an1n08x5 FILLER_74_1883 ();
 b15zdnd00an1n02x5 FILLER_74_1891 ();
 b15zdnd00an1n01x5 FILLER_74_1893 ();
 b15zdnd11an1n08x5 FILLER_74_1904 ();
 b15zdnd11an1n04x5 FILLER_74_1912 ();
 b15zdnd00an1n02x5 FILLER_74_1916 ();
 b15zdnd11an1n16x5 FILLER_74_1923 ();
 b15zdnd00an1n02x5 FILLER_74_1939 ();
 b15zdnd11an1n64x5 FILLER_74_1955 ();
 b15zdnd11an1n32x5 FILLER_74_2019 ();
 b15zdnd11an1n16x5 FILLER_74_2051 ();
 b15zdnd11an1n64x5 FILLER_74_2073 ();
 b15zdnd11an1n16x5 FILLER_74_2137 ();
 b15zdnd00an1n01x5 FILLER_74_2153 ();
 b15zdnd11an1n08x5 FILLER_74_2162 ();
 b15zdnd11an1n04x5 FILLER_74_2170 ();
 b15zdnd00an1n02x5 FILLER_74_2174 ();
 b15zdnd11an1n08x5 FILLER_74_2191 ();
 b15zdnd11an1n04x5 FILLER_74_2199 ();
 b15zdnd00an1n02x5 FILLER_74_2203 ();
 b15zdnd00an1n01x5 FILLER_74_2205 ();
 b15zdnd11an1n32x5 FILLER_74_2220 ();
 b15zdnd11an1n16x5 FILLER_74_2252 ();
 b15zdnd11an1n08x5 FILLER_74_2268 ();
 b15zdnd11an1n64x5 FILLER_75_0 ();
 b15zdnd11an1n16x5 FILLER_75_64 ();
 b15zdnd11an1n08x5 FILLER_75_80 ();
 b15zdnd11an1n04x5 FILLER_75_88 ();
 b15zdnd00an1n01x5 FILLER_75_92 ();
 b15zdnd11an1n32x5 FILLER_75_102 ();
 b15zdnd11an1n04x5 FILLER_75_134 ();
 b15zdnd00an1n02x5 FILLER_75_138 ();
 b15zdnd11an1n16x5 FILLER_75_146 ();
 b15zdnd11an1n04x5 FILLER_75_162 ();
 b15zdnd00an1n02x5 FILLER_75_166 ();
 b15zdnd00an1n01x5 FILLER_75_168 ();
 b15zdnd11an1n08x5 FILLER_75_176 ();
 b15zdnd11an1n64x5 FILLER_75_190 ();
 b15zdnd11an1n08x5 FILLER_75_254 ();
 b15zdnd00an1n02x5 FILLER_75_262 ();
 b15zdnd00an1n01x5 FILLER_75_264 ();
 b15zdnd11an1n64x5 FILLER_75_273 ();
 b15zdnd11an1n64x5 FILLER_75_337 ();
 b15zdnd11an1n32x5 FILLER_75_401 ();
 b15zdnd00an1n02x5 FILLER_75_433 ();
 b15zdnd11an1n64x5 FILLER_75_449 ();
 b15zdnd11an1n16x5 FILLER_75_513 ();
 b15zdnd11an1n04x5 FILLER_75_529 ();
 b15zdnd00an1n02x5 FILLER_75_533 ();
 b15zdnd11an1n32x5 FILLER_75_550 ();
 b15zdnd11an1n08x5 FILLER_75_582 ();
 b15zdnd00an1n02x5 FILLER_75_590 ();
 b15zdnd00an1n01x5 FILLER_75_592 ();
 b15zdnd11an1n04x5 FILLER_75_611 ();
 b15zdnd11an1n04x5 FILLER_75_629 ();
 b15zdnd11an1n16x5 FILLER_75_643 ();
 b15zdnd11an1n32x5 FILLER_75_663 ();
 b15zdnd00an1n01x5 FILLER_75_695 ();
 b15zdnd11an1n08x5 FILLER_75_704 ();
 b15zdnd00an1n02x5 FILLER_75_712 ();
 b15zdnd00an1n01x5 FILLER_75_714 ();
 b15zdnd11an1n32x5 FILLER_75_720 ();
 b15zdnd11an1n16x5 FILLER_75_752 ();
 b15zdnd11an1n32x5 FILLER_75_774 ();
 b15zdnd11an1n04x5 FILLER_75_806 ();
 b15zdnd00an1n01x5 FILLER_75_810 ();
 b15zdnd11an1n16x5 FILLER_75_817 ();
 b15zdnd11an1n08x5 FILLER_75_833 ();
 b15zdnd11an1n04x5 FILLER_75_841 ();
 b15zdnd11an1n32x5 FILLER_75_858 ();
 b15zdnd11an1n08x5 FILLER_75_890 ();
 b15zdnd11an1n04x5 FILLER_75_898 ();
 b15zdnd00an1n02x5 FILLER_75_902 ();
 b15zdnd11an1n64x5 FILLER_75_927 ();
 b15zdnd11an1n64x5 FILLER_75_991 ();
 b15zdnd11an1n04x5 FILLER_75_1055 ();
 b15zdnd00an1n01x5 FILLER_75_1059 ();
 b15zdnd11an1n04x5 FILLER_75_1070 ();
 b15zdnd11an1n04x5 FILLER_75_1083 ();
 b15zdnd11an1n64x5 FILLER_75_1092 ();
 b15zdnd11an1n08x5 FILLER_75_1156 ();
 b15zdnd00an1n02x5 FILLER_75_1164 ();
 b15zdnd00an1n01x5 FILLER_75_1166 ();
 b15zdnd11an1n08x5 FILLER_75_1175 ();
 b15zdnd11an1n04x5 FILLER_75_1183 ();
 b15zdnd00an1n02x5 FILLER_75_1187 ();
 b15zdnd00an1n01x5 FILLER_75_1189 ();
 b15zdnd11an1n64x5 FILLER_75_1195 ();
 b15zdnd11an1n08x5 FILLER_75_1259 ();
 b15zdnd00an1n01x5 FILLER_75_1267 ();
 b15zdnd11an1n32x5 FILLER_75_1294 ();
 b15zdnd11an1n16x5 FILLER_75_1326 ();
 b15zdnd00an1n02x5 FILLER_75_1342 ();
 b15zdnd00an1n01x5 FILLER_75_1344 ();
 b15zdnd11an1n32x5 FILLER_75_1359 ();
 b15zdnd00an1n02x5 FILLER_75_1391 ();
 b15zdnd11an1n64x5 FILLER_75_1410 ();
 b15zdnd11an1n64x5 FILLER_75_1474 ();
 b15zdnd11an1n08x5 FILLER_75_1553 ();
 b15zdnd11an1n04x5 FILLER_75_1561 ();
 b15zdnd00an1n02x5 FILLER_75_1565 ();
 b15zdnd11an1n16x5 FILLER_75_1576 ();
 b15zdnd00an1n01x5 FILLER_75_1592 ();
 b15zdnd11an1n32x5 FILLER_75_1613 ();
 b15zdnd11an1n16x5 FILLER_75_1645 ();
 b15zdnd11an1n08x5 FILLER_75_1661 ();
 b15zdnd00an1n01x5 FILLER_75_1669 ();
 b15zdnd11an1n32x5 FILLER_75_1688 ();
 b15zdnd11an1n16x5 FILLER_75_1720 ();
 b15zdnd11an1n04x5 FILLER_75_1736 ();
 b15zdnd00an1n02x5 FILLER_75_1740 ();
 b15zdnd11an1n04x5 FILLER_75_1756 ();
 b15zdnd11an1n32x5 FILLER_75_1791 ();
 b15zdnd11an1n16x5 FILLER_75_1823 ();
 b15zdnd11an1n04x5 FILLER_75_1859 ();
 b15zdnd11an1n64x5 FILLER_75_1868 ();
 b15zdnd11an1n32x5 FILLER_75_1932 ();
 b15zdnd11an1n16x5 FILLER_75_1964 ();
 b15zdnd00an1n01x5 FILLER_75_1980 ();
 b15zdnd11an1n64x5 FILLER_75_1989 ();
 b15zdnd11an1n16x5 FILLER_75_2053 ();
 b15zdnd11an1n32x5 FILLER_75_2074 ();
 b15zdnd11an1n04x5 FILLER_75_2106 ();
 b15zdnd00an1n02x5 FILLER_75_2110 ();
 b15zdnd00an1n01x5 FILLER_75_2112 ();
 b15zdnd11an1n16x5 FILLER_75_2123 ();
 b15zdnd00an1n02x5 FILLER_75_2139 ();
 b15zdnd00an1n01x5 FILLER_75_2141 ();
 b15zdnd11an1n16x5 FILLER_75_2148 ();
 b15zdnd11an1n04x5 FILLER_75_2164 ();
 b15zdnd00an1n01x5 FILLER_75_2168 ();
 b15zdnd11an1n64x5 FILLER_75_2187 ();
 b15zdnd11an1n32x5 FILLER_75_2251 ();
 b15zdnd00an1n01x5 FILLER_75_2283 ();
 b15zdnd11an1n32x5 FILLER_76_8 ();
 b15zdnd00an1n01x5 FILLER_76_40 ();
 b15zdnd11an1n08x5 FILLER_76_58 ();
 b15zdnd11an1n04x5 FILLER_76_66 ();
 b15zdnd00an1n01x5 FILLER_76_70 ();
 b15zdnd11an1n32x5 FILLER_76_77 ();
 b15zdnd11an1n16x5 FILLER_76_109 ();
 b15zdnd00an1n01x5 FILLER_76_125 ();
 b15zdnd11an1n04x5 FILLER_76_138 ();
 b15zdnd11an1n32x5 FILLER_76_154 ();
 b15zdnd00an1n02x5 FILLER_76_186 ();
 b15zdnd11an1n32x5 FILLER_76_194 ();
 b15zdnd11an1n04x5 FILLER_76_226 ();
 b15zdnd00an1n01x5 FILLER_76_230 ();
 b15zdnd11an1n04x5 FILLER_76_235 ();
 b15zdnd00an1n01x5 FILLER_76_239 ();
 b15zdnd11an1n16x5 FILLER_76_245 ();
 b15zdnd11an1n08x5 FILLER_76_261 ();
 b15zdnd00an1n02x5 FILLER_76_269 ();
 b15zdnd00an1n01x5 FILLER_76_271 ();
 b15zdnd11an1n04x5 FILLER_76_284 ();
 b15zdnd11an1n16x5 FILLER_76_309 ();
 b15zdnd11an1n04x5 FILLER_76_325 ();
 b15zdnd00an1n02x5 FILLER_76_329 ();
 b15zdnd00an1n01x5 FILLER_76_331 ();
 b15zdnd11an1n32x5 FILLER_76_338 ();
 b15zdnd11an1n08x5 FILLER_76_370 ();
 b15zdnd00an1n01x5 FILLER_76_378 ();
 b15zdnd11an1n64x5 FILLER_76_385 ();
 b15zdnd11an1n64x5 FILLER_76_449 ();
 b15zdnd11an1n16x5 FILLER_76_513 ();
 b15zdnd11an1n08x5 FILLER_76_529 ();
 b15zdnd00an1n01x5 FILLER_76_537 ();
 b15zdnd11an1n08x5 FILLER_76_550 ();
 b15zdnd11an1n04x5 FILLER_76_558 ();
 b15zdnd00an1n02x5 FILLER_76_562 ();
 b15zdnd11an1n08x5 FILLER_76_570 ();
 b15zdnd11an1n04x5 FILLER_76_578 ();
 b15zdnd00an1n02x5 FILLER_76_582 ();
 b15zdnd11an1n04x5 FILLER_76_597 ();
 b15zdnd11an1n64x5 FILLER_76_606 ();
 b15zdnd11an1n32x5 FILLER_76_670 ();
 b15zdnd11an1n16x5 FILLER_76_702 ();
 b15zdnd11an1n32x5 FILLER_76_726 ();
 b15zdnd11an1n04x5 FILLER_76_758 ();
 b15zdnd11an1n64x5 FILLER_76_766 ();
 b15zdnd11an1n64x5 FILLER_76_830 ();
 b15zdnd11an1n64x5 FILLER_76_894 ();
 b15zdnd11an1n32x5 FILLER_76_958 ();
 b15zdnd11an1n16x5 FILLER_76_990 ();
 b15zdnd11an1n08x5 FILLER_76_1006 ();
 b15zdnd00an1n02x5 FILLER_76_1014 ();
 b15zdnd00an1n01x5 FILLER_76_1016 ();
 b15zdnd11an1n64x5 FILLER_76_1021 ();
 b15zdnd11an1n64x5 FILLER_76_1085 ();
 b15zdnd11an1n04x5 FILLER_76_1149 ();
 b15zdnd00an1n02x5 FILLER_76_1153 ();
 b15zdnd00an1n01x5 FILLER_76_1155 ();
 b15zdnd11an1n16x5 FILLER_76_1160 ();
 b15zdnd11an1n08x5 FILLER_76_1176 ();
 b15zdnd11an1n64x5 FILLER_76_1215 ();
 b15zdnd11an1n16x5 FILLER_76_1279 ();
 b15zdnd11an1n04x5 FILLER_76_1295 ();
 b15zdnd11an1n04x5 FILLER_76_1322 ();
 b15zdnd00an1n02x5 FILLER_76_1326 ();
 b15zdnd11an1n32x5 FILLER_76_1340 ();
 b15zdnd11an1n08x5 FILLER_76_1372 ();
 b15zdnd11an1n04x5 FILLER_76_1380 ();
 b15zdnd00an1n02x5 FILLER_76_1384 ();
 b15zdnd11an1n32x5 FILLER_76_1416 ();
 b15zdnd00an1n02x5 FILLER_76_1448 ();
 b15zdnd11an1n64x5 FILLER_76_1454 ();
 b15zdnd11an1n08x5 FILLER_76_1544 ();
 b15zdnd00an1n02x5 FILLER_76_1552 ();
 b15zdnd11an1n08x5 FILLER_76_1567 ();
 b15zdnd11an1n32x5 FILLER_76_1601 ();
 b15zdnd11an1n08x5 FILLER_76_1633 ();
 b15zdnd11an1n04x5 FILLER_76_1641 ();
 b15zdnd00an1n02x5 FILLER_76_1645 ();
 b15zdnd11an1n04x5 FILLER_76_1663 ();
 b15zdnd11an1n64x5 FILLER_76_1687 ();
 b15zdnd11an1n04x5 FILLER_76_1751 ();
 b15zdnd00an1n02x5 FILLER_76_1755 ();
 b15zdnd11an1n16x5 FILLER_76_1788 ();
 b15zdnd11an1n04x5 FILLER_76_1804 ();
 b15zdnd00an1n01x5 FILLER_76_1808 ();
 b15zdnd11an1n32x5 FILLER_76_1813 ();
 b15zdnd11an1n08x5 FILLER_76_1845 ();
 b15zdnd00an1n02x5 FILLER_76_1853 ();
 b15zdnd00an1n01x5 FILLER_76_1855 ();
 b15zdnd11an1n16x5 FILLER_76_1868 ();
 b15zdnd00an1n02x5 FILLER_76_1884 ();
 b15zdnd11an1n32x5 FILLER_76_1893 ();
 b15zdnd11an1n16x5 FILLER_76_1925 ();
 b15zdnd11an1n04x5 FILLER_76_1941 ();
 b15zdnd00an1n02x5 FILLER_76_1945 ();
 b15zdnd11an1n16x5 FILLER_76_1953 ();
 b15zdnd11an1n08x5 FILLER_76_1969 ();
 b15zdnd00an1n02x5 FILLER_76_1977 ();
 b15zdnd11an1n64x5 FILLER_76_1983 ();
 b15zdnd11an1n64x5 FILLER_76_2047 ();
 b15zdnd11an1n08x5 FILLER_76_2111 ();
 b15zdnd11an1n04x5 FILLER_76_2119 ();
 b15zdnd00an1n01x5 FILLER_76_2123 ();
 b15zdnd11an1n08x5 FILLER_76_2129 ();
 b15zdnd00an1n01x5 FILLER_76_2137 ();
 b15zdnd00an1n02x5 FILLER_76_2152 ();
 b15zdnd11an1n32x5 FILLER_76_2162 ();
 b15zdnd11an1n08x5 FILLER_76_2194 ();
 b15zdnd11an1n04x5 FILLER_76_2202 ();
 b15zdnd00an1n01x5 FILLER_76_2206 ();
 b15zdnd11an1n04x5 FILLER_76_2211 ();
 b15zdnd11an1n32x5 FILLER_76_2235 ();
 b15zdnd11an1n08x5 FILLER_76_2267 ();
 b15zdnd00an1n01x5 FILLER_76_2275 ();
 b15zdnd11an1n32x5 FILLER_77_0 ();
 b15zdnd11an1n04x5 FILLER_77_32 ();
 b15zdnd00an1n02x5 FILLER_77_36 ();
 b15zdnd11an1n08x5 FILLER_77_48 ();
 b15zdnd00an1n02x5 FILLER_77_56 ();
 b15zdnd00an1n01x5 FILLER_77_58 ();
 b15zdnd11an1n16x5 FILLER_77_63 ();
 b15zdnd11an1n08x5 FILLER_77_79 ();
 b15zdnd00an1n02x5 FILLER_77_87 ();
 b15zdnd11an1n16x5 FILLER_77_96 ();
 b15zdnd11an1n08x5 FILLER_77_112 ();
 b15zdnd11an1n64x5 FILLER_77_132 ();
 b15zdnd11an1n08x5 FILLER_77_196 ();
 b15zdnd00an1n02x5 FILLER_77_204 ();
 b15zdnd00an1n01x5 FILLER_77_206 ();
 b15zdnd11an1n04x5 FILLER_77_218 ();
 b15zdnd00an1n02x5 FILLER_77_222 ();
 b15zdnd11an1n04x5 FILLER_77_231 ();
 b15zdnd11an1n04x5 FILLER_77_242 ();
 b15zdnd11an1n08x5 FILLER_77_258 ();
 b15zdnd00an1n02x5 FILLER_77_266 ();
 b15zdnd11an1n64x5 FILLER_77_272 ();
 b15zdnd00an1n02x5 FILLER_77_336 ();
 b15zdnd00an1n01x5 FILLER_77_338 ();
 b15zdnd11an1n04x5 FILLER_77_359 ();
 b15zdnd11an1n04x5 FILLER_77_372 ();
 b15zdnd11an1n32x5 FILLER_77_380 ();
 b15zdnd11an1n16x5 FILLER_77_412 ();
 b15zdnd11an1n08x5 FILLER_77_428 ();
 b15zdnd11an1n04x5 FILLER_77_436 ();
 b15zdnd00an1n02x5 FILLER_77_440 ();
 b15zdnd00an1n01x5 FILLER_77_442 ();
 b15zdnd11an1n16x5 FILLER_77_475 ();
 b15zdnd00an1n01x5 FILLER_77_491 ();
 b15zdnd11an1n04x5 FILLER_77_508 ();
 b15zdnd00an1n02x5 FILLER_77_512 ();
 b15zdnd00an1n01x5 FILLER_77_514 ();
 b15zdnd11an1n04x5 FILLER_77_547 ();
 b15zdnd00an1n02x5 FILLER_77_551 ();
 b15zdnd11an1n04x5 FILLER_77_561 ();
 b15zdnd11an1n16x5 FILLER_77_596 ();
 b15zdnd11an1n04x5 FILLER_77_612 ();
 b15zdnd00an1n01x5 FILLER_77_616 ();
 b15zdnd11an1n16x5 FILLER_77_638 ();
 b15zdnd00an1n02x5 FILLER_77_654 ();
 b15zdnd11an1n32x5 FILLER_77_666 ();
 b15zdnd11an1n04x5 FILLER_77_698 ();
 b15zdnd00an1n02x5 FILLER_77_702 ();
 b15zdnd00an1n01x5 FILLER_77_704 ();
 b15zdnd11an1n64x5 FILLER_77_711 ();
 b15zdnd11an1n32x5 FILLER_77_775 ();
 b15zdnd11an1n08x5 FILLER_77_807 ();
 b15zdnd11an1n04x5 FILLER_77_815 ();
 b15zdnd00an1n01x5 FILLER_77_819 ();
 b15zdnd11an1n32x5 FILLER_77_828 ();
 b15zdnd11an1n16x5 FILLER_77_860 ();
 b15zdnd11an1n08x5 FILLER_77_876 ();
 b15zdnd11an1n04x5 FILLER_77_884 ();
 b15zdnd00an1n02x5 FILLER_77_888 ();
 b15zdnd11an1n16x5 FILLER_77_904 ();
 b15zdnd11an1n04x5 FILLER_77_920 ();
 b15zdnd11an1n04x5 FILLER_77_935 ();
 b15zdnd00an1n02x5 FILLER_77_939 ();
 b15zdnd11an1n16x5 FILLER_77_950 ();
 b15zdnd11an1n08x5 FILLER_77_966 ();
 b15zdnd00an1n01x5 FILLER_77_974 ();
 b15zdnd11an1n08x5 FILLER_77_1000 ();
 b15zdnd11an1n04x5 FILLER_77_1008 ();
 b15zdnd00an1n01x5 FILLER_77_1012 ();
 b15zdnd11an1n32x5 FILLER_77_1033 ();
 b15zdnd11an1n16x5 FILLER_77_1065 ();
 b15zdnd00an1n02x5 FILLER_77_1081 ();
 b15zdnd00an1n01x5 FILLER_77_1083 ();
 b15zdnd11an1n64x5 FILLER_77_1104 ();
 b15zdnd11an1n32x5 FILLER_77_1168 ();
 b15zdnd11an1n16x5 FILLER_77_1200 ();
 b15zdnd11an1n08x5 FILLER_77_1216 ();
 b15zdnd00an1n02x5 FILLER_77_1224 ();
 b15zdnd11an1n04x5 FILLER_77_1257 ();
 b15zdnd11an1n16x5 FILLER_77_1265 ();
 b15zdnd11an1n08x5 FILLER_77_1281 ();
 b15zdnd00an1n02x5 FILLER_77_1289 ();
 b15zdnd11an1n04x5 FILLER_77_1322 ();
 b15zdnd11an1n16x5 FILLER_77_1342 ();
 b15zdnd00an1n01x5 FILLER_77_1358 ();
 b15zdnd11an1n16x5 FILLER_77_1365 ();
 b15zdnd00an1n02x5 FILLER_77_1381 ();
 b15zdnd11an1n16x5 FILLER_77_1392 ();
 b15zdnd11an1n04x5 FILLER_77_1408 ();
 b15zdnd11an1n08x5 FILLER_77_1427 ();
 b15zdnd00an1n02x5 FILLER_77_1435 ();
 b15zdnd11an1n08x5 FILLER_77_1452 ();
 b15zdnd00an1n02x5 FILLER_77_1460 ();
 b15zdnd11an1n08x5 FILLER_77_1468 ();
 b15zdnd00an1n02x5 FILLER_77_1476 ();
 b15zdnd11an1n04x5 FILLER_77_1484 ();
 b15zdnd11an1n16x5 FILLER_77_1499 ();
 b15zdnd11an1n08x5 FILLER_77_1520 ();
 b15zdnd00an1n02x5 FILLER_77_1528 ();
 b15zdnd11an1n04x5 FILLER_77_1540 ();
 b15zdnd11an1n16x5 FILLER_77_1550 ();
 b15zdnd11an1n08x5 FILLER_77_1566 ();
 b15zdnd00an1n01x5 FILLER_77_1574 ();
 b15zdnd11an1n08x5 FILLER_77_1586 ();
 b15zdnd11an1n04x5 FILLER_77_1594 ();
 b15zdnd00an1n01x5 FILLER_77_1598 ();
 b15zdnd11an1n04x5 FILLER_77_1604 ();
 b15zdnd11an1n04x5 FILLER_77_1614 ();
 b15zdnd11an1n08x5 FILLER_77_1623 ();
 b15zdnd00an1n02x5 FILLER_77_1631 ();
 b15zdnd11an1n08x5 FILLER_77_1646 ();
 b15zdnd11an1n04x5 FILLER_77_1654 ();
 b15zdnd00an1n01x5 FILLER_77_1658 ();
 b15zdnd11an1n04x5 FILLER_77_1677 ();
 b15zdnd11an1n64x5 FILLER_77_1701 ();
 b15zdnd11an1n08x5 FILLER_77_1765 ();
 b15zdnd11an1n04x5 FILLER_77_1773 ();
 b15zdnd00an1n01x5 FILLER_77_1777 ();
 b15zdnd11an1n16x5 FILLER_77_1787 ();
 b15zdnd11an1n04x5 FILLER_77_1803 ();
 b15zdnd00an1n02x5 FILLER_77_1807 ();
 b15zdnd11an1n32x5 FILLER_77_1814 ();
 b15zdnd11an1n08x5 FILLER_77_1846 ();
 b15zdnd00an1n02x5 FILLER_77_1854 ();
 b15zdnd11an1n16x5 FILLER_77_1868 ();
 b15zdnd11an1n04x5 FILLER_77_1884 ();
 b15zdnd11an1n32x5 FILLER_77_1894 ();
 b15zdnd11an1n16x5 FILLER_77_1926 ();
 b15zdnd11an1n08x5 FILLER_77_1942 ();
 b15zdnd11an1n04x5 FILLER_77_1950 ();
 b15zdnd00an1n02x5 FILLER_77_1954 ();
 b15zdnd11an1n04x5 FILLER_77_1974 ();
 b15zdnd11an1n16x5 FILLER_77_1984 ();
 b15zdnd11an1n08x5 FILLER_77_2000 ();
 b15zdnd00an1n01x5 FILLER_77_2008 ();
 b15zdnd11an1n04x5 FILLER_77_2022 ();
 b15zdnd11an1n08x5 FILLER_77_2033 ();
 b15zdnd11an1n04x5 FILLER_77_2041 ();
 b15zdnd00an1n02x5 FILLER_77_2045 ();
 b15zdnd11an1n16x5 FILLER_77_2051 ();
 b15zdnd11an1n08x5 FILLER_77_2067 ();
 b15zdnd00an1n02x5 FILLER_77_2075 ();
 b15zdnd00an1n01x5 FILLER_77_2077 ();
 b15zdnd11an1n04x5 FILLER_77_2087 ();
 b15zdnd11an1n16x5 FILLER_77_2099 ();
 b15zdnd11an1n08x5 FILLER_77_2133 ();
 b15zdnd00an1n01x5 FILLER_77_2141 ();
 b15zdnd11an1n08x5 FILLER_77_2147 ();
 b15zdnd11an1n04x5 FILLER_77_2155 ();
 b15zdnd11an1n04x5 FILLER_77_2165 ();
 b15zdnd11an1n64x5 FILLER_77_2189 ();
 b15zdnd11an1n16x5 FILLER_77_2253 ();
 b15zdnd11an1n08x5 FILLER_77_2269 ();
 b15zdnd11an1n04x5 FILLER_77_2277 ();
 b15zdnd00an1n02x5 FILLER_77_2281 ();
 b15zdnd00an1n01x5 FILLER_77_2283 ();
 b15zdnd11an1n32x5 FILLER_78_8 ();
 b15zdnd00an1n02x5 FILLER_78_40 ();
 b15zdnd11an1n04x5 FILLER_78_59 ();
 b15zdnd11an1n08x5 FILLER_78_81 ();
 b15zdnd00an1n02x5 FILLER_78_89 ();
 b15zdnd00an1n01x5 FILLER_78_91 ();
 b15zdnd11an1n04x5 FILLER_78_118 ();
 b15zdnd11an1n64x5 FILLER_78_129 ();
 b15zdnd11an1n64x5 FILLER_78_193 ();
 b15zdnd00an1n02x5 FILLER_78_257 ();
 b15zdnd00an1n01x5 FILLER_78_259 ();
 b15zdnd11an1n16x5 FILLER_78_266 ();
 b15zdnd00an1n02x5 FILLER_78_282 ();
 b15zdnd11an1n04x5 FILLER_78_289 ();
 b15zdnd11an1n16x5 FILLER_78_308 ();
 b15zdnd11an1n08x5 FILLER_78_324 ();
 b15zdnd00an1n01x5 FILLER_78_332 ();
 b15zdnd11an1n32x5 FILLER_78_341 ();
 b15zdnd00an1n01x5 FILLER_78_373 ();
 b15zdnd11an1n32x5 FILLER_78_379 ();
 b15zdnd11an1n16x5 FILLER_78_411 ();
 b15zdnd11an1n04x5 FILLER_78_427 ();
 b15zdnd00an1n01x5 FILLER_78_431 ();
 b15zdnd11an1n04x5 FILLER_78_448 ();
 b15zdnd11an1n16x5 FILLER_78_478 ();
 b15zdnd11an1n08x5 FILLER_78_494 ();
 b15zdnd00an1n01x5 FILLER_78_502 ();
 b15zdnd11an1n16x5 FILLER_78_535 ();
 b15zdnd00an1n01x5 FILLER_78_551 ();
 b15zdnd11an1n04x5 FILLER_78_560 ();
 b15zdnd00an1n02x5 FILLER_78_564 ();
 b15zdnd00an1n01x5 FILLER_78_566 ();
 b15zdnd11an1n64x5 FILLER_78_583 ();
 b15zdnd11an1n64x5 FILLER_78_647 ();
 b15zdnd11an1n04x5 FILLER_78_711 ();
 b15zdnd00an1n02x5 FILLER_78_715 ();
 b15zdnd00an1n01x5 FILLER_78_717 ();
 b15zdnd11an1n16x5 FILLER_78_726 ();
 b15zdnd00an1n02x5 FILLER_78_742 ();
 b15zdnd00an1n01x5 FILLER_78_744 ();
 b15zdnd11an1n04x5 FILLER_78_761 ();
 b15zdnd11an1n32x5 FILLER_78_774 ();
 b15zdnd11an1n08x5 FILLER_78_806 ();
 b15zdnd11an1n04x5 FILLER_78_814 ();
 b15zdnd00an1n02x5 FILLER_78_818 ();
 b15zdnd00an1n01x5 FILLER_78_820 ();
 b15zdnd11an1n16x5 FILLER_78_825 ();
 b15zdnd11an1n08x5 FILLER_78_841 ();
 b15zdnd11an1n04x5 FILLER_78_849 ();
 b15zdnd00an1n01x5 FILLER_78_853 ();
 b15zdnd11an1n32x5 FILLER_78_860 ();
 b15zdnd00an1n02x5 FILLER_78_892 ();
 b15zdnd00an1n01x5 FILLER_78_894 ();
 b15zdnd11an1n32x5 FILLER_78_909 ();
 b15zdnd00an1n02x5 FILLER_78_941 ();
 b15zdnd00an1n01x5 FILLER_78_943 ();
 b15zdnd11an1n08x5 FILLER_78_964 ();
 b15zdnd11an1n04x5 FILLER_78_972 ();
 b15zdnd00an1n01x5 FILLER_78_976 ();
 b15zdnd11an1n04x5 FILLER_78_1008 ();
 b15zdnd00an1n02x5 FILLER_78_1012 ();
 b15zdnd11an1n08x5 FILLER_78_1019 ();
 b15zdnd00an1n01x5 FILLER_78_1027 ();
 b15zdnd11an1n64x5 FILLER_78_1032 ();
 b15zdnd11an1n32x5 FILLER_78_1096 ();
 b15zdnd11an1n16x5 FILLER_78_1128 ();
 b15zdnd11an1n16x5 FILLER_78_1149 ();
 b15zdnd11an1n08x5 FILLER_78_1165 ();
 b15zdnd00an1n02x5 FILLER_78_1173 ();
 b15zdnd11an1n32x5 FILLER_78_1195 ();
 b15zdnd11an1n16x5 FILLER_78_1227 ();
 b15zdnd11an1n08x5 FILLER_78_1243 ();
 b15zdnd11an1n04x5 FILLER_78_1251 ();
 b15zdnd00an1n02x5 FILLER_78_1255 ();
 b15zdnd11an1n64x5 FILLER_78_1262 ();
 b15zdnd11an1n04x5 FILLER_78_1326 ();
 b15zdnd00an1n02x5 FILLER_78_1330 ();
 b15zdnd00an1n01x5 FILLER_78_1332 ();
 b15zdnd11an1n32x5 FILLER_78_1344 ();
 b15zdnd11an1n08x5 FILLER_78_1376 ();
 b15zdnd11an1n04x5 FILLER_78_1390 ();
 b15zdnd00an1n02x5 FILLER_78_1394 ();
 b15zdnd00an1n01x5 FILLER_78_1396 ();
 b15zdnd11an1n04x5 FILLER_78_1407 ();
 b15zdnd11an1n08x5 FILLER_78_1426 ();
 b15zdnd00an1n01x5 FILLER_78_1434 ();
 b15zdnd11an1n08x5 FILLER_78_1448 ();
 b15zdnd11an1n04x5 FILLER_78_1456 ();
 b15zdnd00an1n01x5 FILLER_78_1460 ();
 b15zdnd11an1n08x5 FILLER_78_1467 ();
 b15zdnd11an1n04x5 FILLER_78_1489 ();
 b15zdnd11an1n04x5 FILLER_78_1499 ();
 b15zdnd00an1n01x5 FILLER_78_1503 ();
 b15zdnd11an1n08x5 FILLER_78_1509 ();
 b15zdnd11an1n64x5 FILLER_78_1525 ();
 b15zdnd11an1n64x5 FILLER_78_1589 ();
 b15zdnd11an1n64x5 FILLER_78_1653 ();
 b15zdnd11an1n64x5 FILLER_78_1717 ();
 b15zdnd11an1n16x5 FILLER_78_1781 ();
 b15zdnd11an1n08x5 FILLER_78_1797 ();
 b15zdnd00an1n02x5 FILLER_78_1805 ();
 b15zdnd00an1n01x5 FILLER_78_1807 ();
 b15zdnd11an1n32x5 FILLER_78_1821 ();
 b15zdnd11an1n16x5 FILLER_78_1853 ();
 b15zdnd11an1n04x5 FILLER_78_1869 ();
 b15zdnd00an1n02x5 FILLER_78_1873 ();
 b15zdnd11an1n04x5 FILLER_78_1880 ();
 b15zdnd00an1n01x5 FILLER_78_1884 ();
 b15zdnd11an1n08x5 FILLER_78_1900 ();
 b15zdnd11an1n04x5 FILLER_78_1908 ();
 b15zdnd00an1n01x5 FILLER_78_1912 ();
 b15zdnd11an1n32x5 FILLER_78_1919 ();
 b15zdnd11an1n16x5 FILLER_78_1951 ();
 b15zdnd11an1n08x5 FILLER_78_1967 ();
 b15zdnd11an1n04x5 FILLER_78_1975 ();
 b15zdnd00an1n02x5 FILLER_78_1979 ();
 b15zdnd11an1n16x5 FILLER_78_1993 ();
 b15zdnd11an1n08x5 FILLER_78_2009 ();
 b15zdnd00an1n02x5 FILLER_78_2017 ();
 b15zdnd11an1n32x5 FILLER_78_2023 ();
 b15zdnd11an1n16x5 FILLER_78_2055 ();
 b15zdnd00an1n01x5 FILLER_78_2071 ();
 b15zdnd11an1n04x5 FILLER_78_2088 ();
 b15zdnd11an1n32x5 FILLER_78_2099 ();
 b15zdnd11an1n16x5 FILLER_78_2131 ();
 b15zdnd11an1n04x5 FILLER_78_2147 ();
 b15zdnd00an1n02x5 FILLER_78_2151 ();
 b15zdnd00an1n01x5 FILLER_78_2153 ();
 b15zdnd11an1n64x5 FILLER_78_2162 ();
 b15zdnd11an1n32x5 FILLER_78_2226 ();
 b15zdnd11an1n16x5 FILLER_78_2258 ();
 b15zdnd00an1n02x5 FILLER_78_2274 ();
 b15zdnd11an1n64x5 FILLER_79_0 ();
 b15zdnd11an1n08x5 FILLER_79_64 ();
 b15zdnd11an1n04x5 FILLER_79_84 ();
 b15zdnd11an1n16x5 FILLER_79_97 ();
 b15zdnd11an1n08x5 FILLER_79_113 ();
 b15zdnd11an1n16x5 FILLER_79_128 ();
 b15zdnd11an1n08x5 FILLER_79_144 ();
 b15zdnd00an1n02x5 FILLER_79_152 ();
 b15zdnd11an1n08x5 FILLER_79_160 ();
 b15zdnd11an1n16x5 FILLER_79_175 ();
 b15zdnd11an1n08x5 FILLER_79_191 ();
 b15zdnd00an1n01x5 FILLER_79_199 ();
 b15zdnd11an1n32x5 FILLER_79_212 ();
 b15zdnd11an1n08x5 FILLER_79_244 ();
 b15zdnd11an1n04x5 FILLER_79_252 ();
 b15zdnd00an1n02x5 FILLER_79_256 ();
 b15zdnd11an1n64x5 FILLER_79_264 ();
 b15zdnd11an1n16x5 FILLER_79_328 ();
 b15zdnd11an1n08x5 FILLER_79_344 ();
 b15zdnd11an1n04x5 FILLER_79_352 ();
 b15zdnd00an1n01x5 FILLER_79_356 ();
 b15zdnd11an1n16x5 FILLER_79_364 ();
 b15zdnd11an1n08x5 FILLER_79_380 ();
 b15zdnd11an1n32x5 FILLER_79_397 ();
 b15zdnd11an1n04x5 FILLER_79_429 ();
 b15zdnd11an1n04x5 FILLER_79_454 ();
 b15zdnd11an1n32x5 FILLER_79_474 ();
 b15zdnd11an1n04x5 FILLER_79_506 ();
 b15zdnd11an1n32x5 FILLER_79_526 ();
 b15zdnd11an1n08x5 FILLER_79_558 ();
 b15zdnd11an1n64x5 FILLER_79_577 ();
 b15zdnd11an1n08x5 FILLER_79_641 ();
 b15zdnd11an1n04x5 FILLER_79_649 ();
 b15zdnd00an1n02x5 FILLER_79_653 ();
 b15zdnd00an1n01x5 FILLER_79_655 ();
 b15zdnd11an1n32x5 FILLER_79_661 ();
 b15zdnd11an1n04x5 FILLER_79_705 ();
 b15zdnd00an1n01x5 FILLER_79_709 ();
 b15zdnd11an1n16x5 FILLER_79_715 ();
 b15zdnd11an1n32x5 FILLER_79_738 ();
 b15zdnd11an1n04x5 FILLER_79_770 ();
 b15zdnd11an1n08x5 FILLER_79_780 ();
 b15zdnd11an1n16x5 FILLER_79_794 ();
 b15zdnd00an1n02x5 FILLER_79_810 ();
 b15zdnd00an1n01x5 FILLER_79_812 ();
 b15zdnd11an1n04x5 FILLER_79_826 ();
 b15zdnd11an1n32x5 FILLER_79_843 ();
 b15zdnd00an1n01x5 FILLER_79_875 ();
 b15zdnd11an1n04x5 FILLER_79_907 ();
 b15zdnd11an1n16x5 FILLER_79_936 ();
 b15zdnd11an1n08x5 FILLER_79_952 ();
 b15zdnd00an1n02x5 FILLER_79_960 ();
 b15zdnd00an1n01x5 FILLER_79_962 ();
 b15zdnd11an1n64x5 FILLER_79_983 ();
 b15zdnd11an1n08x5 FILLER_79_1047 ();
 b15zdnd11an1n04x5 FILLER_79_1055 ();
 b15zdnd11an1n16x5 FILLER_79_1070 ();
 b15zdnd11an1n08x5 FILLER_79_1086 ();
 b15zdnd11an1n04x5 FILLER_79_1094 ();
 b15zdnd00an1n02x5 FILLER_79_1098 ();
 b15zdnd11an1n08x5 FILLER_79_1104 ();
 b15zdnd11an1n04x5 FILLER_79_1112 ();
 b15zdnd11an1n04x5 FILLER_79_1136 ();
 b15zdnd11an1n64x5 FILLER_79_1160 ();
 b15zdnd00an1n01x5 FILLER_79_1224 ();
 b15zdnd11an1n04x5 FILLER_79_1251 ();
 b15zdnd11an1n64x5 FILLER_79_1275 ();
 b15zdnd00an1n02x5 FILLER_79_1339 ();
 b15zdnd11an1n04x5 FILLER_79_1346 ();
 b15zdnd11an1n64x5 FILLER_79_1359 ();
 b15zdnd11an1n04x5 FILLER_79_1432 ();
 b15zdnd11an1n64x5 FILLER_79_1445 ();
 b15zdnd11an1n64x5 FILLER_79_1509 ();
 b15zdnd11an1n64x5 FILLER_79_1573 ();
 b15zdnd11an1n04x5 FILLER_79_1637 ();
 b15zdnd00an1n02x5 FILLER_79_1641 ();
 b15zdnd00an1n01x5 FILLER_79_1643 ();
 b15zdnd11an1n32x5 FILLER_79_1660 ();
 b15zdnd11an1n16x5 FILLER_79_1692 ();
 b15zdnd11an1n04x5 FILLER_79_1708 ();
 b15zdnd00an1n02x5 FILLER_79_1712 ();
 b15zdnd11an1n32x5 FILLER_79_1726 ();
 b15zdnd11an1n16x5 FILLER_79_1758 ();
 b15zdnd00an1n02x5 FILLER_79_1774 ();
 b15zdnd00an1n01x5 FILLER_79_1776 ();
 b15zdnd11an1n32x5 FILLER_79_1782 ();
 b15zdnd11an1n16x5 FILLER_79_1814 ();
 b15zdnd11an1n08x5 FILLER_79_1830 ();
 b15zdnd11an1n04x5 FILLER_79_1838 ();
 b15zdnd00an1n02x5 FILLER_79_1842 ();
 b15zdnd00an1n01x5 FILLER_79_1844 ();
 b15zdnd11an1n08x5 FILLER_79_1858 ();
 b15zdnd00an1n02x5 FILLER_79_1866 ();
 b15zdnd11an1n16x5 FILLER_79_1880 ();
 b15zdnd11an1n04x5 FILLER_79_1896 ();
 b15zdnd11an1n08x5 FILLER_79_1905 ();
 b15zdnd11an1n32x5 FILLER_79_1925 ();
 b15zdnd11an1n08x5 FILLER_79_1957 ();
 b15zdnd11an1n04x5 FILLER_79_1974 ();
 b15zdnd11an1n32x5 FILLER_79_1983 ();
 b15zdnd11an1n08x5 FILLER_79_2015 ();
 b15zdnd00an1n01x5 FILLER_79_2023 ();
 b15zdnd11an1n04x5 FILLER_79_2029 ();
 b15zdnd00an1n01x5 FILLER_79_2033 ();
 b15zdnd11an1n04x5 FILLER_79_2044 ();
 b15zdnd11an1n08x5 FILLER_79_2067 ();
 b15zdnd11an1n32x5 FILLER_79_2084 ();
 b15zdnd11an1n04x5 FILLER_79_2116 ();
 b15zdnd00an1n01x5 FILLER_79_2120 ();
 b15zdnd11an1n64x5 FILLER_79_2142 ();
 b15zdnd00an1n01x5 FILLER_79_2206 ();
 b15zdnd11an1n32x5 FILLER_79_2223 ();
 b15zdnd11an1n16x5 FILLER_79_2255 ();
 b15zdnd11an1n08x5 FILLER_79_2271 ();
 b15zdnd11an1n04x5 FILLER_79_2279 ();
 b15zdnd00an1n01x5 FILLER_79_2283 ();
 b15zdnd11an1n32x5 FILLER_80_8 ();
 b15zdnd11an1n04x5 FILLER_80_40 ();
 b15zdnd00an1n02x5 FILLER_80_44 ();
 b15zdnd00an1n01x5 FILLER_80_46 ();
 b15zdnd11an1n64x5 FILLER_80_67 ();
 b15zdnd11an1n16x5 FILLER_80_131 ();
 b15zdnd11an1n08x5 FILLER_80_147 ();
 b15zdnd11an1n04x5 FILLER_80_163 ();
 b15zdnd00an1n02x5 FILLER_80_167 ();
 b15zdnd11an1n64x5 FILLER_80_177 ();
 b15zdnd11an1n32x5 FILLER_80_241 ();
 b15zdnd11an1n16x5 FILLER_80_273 ();
 b15zdnd11an1n04x5 FILLER_80_289 ();
 b15zdnd11an1n04x5 FILLER_80_305 ();
 b15zdnd11an1n32x5 FILLER_80_320 ();
 b15zdnd00an1n02x5 FILLER_80_352 ();
 b15zdnd11an1n64x5 FILLER_80_360 ();
 b15zdnd11an1n64x5 FILLER_80_424 ();
 b15zdnd11an1n04x5 FILLER_80_488 ();
 b15zdnd00an1n02x5 FILLER_80_492 ();
 b15zdnd11an1n04x5 FILLER_80_510 ();
 b15zdnd11an1n32x5 FILLER_80_546 ();
 b15zdnd11an1n16x5 FILLER_80_578 ();
 b15zdnd00an1n01x5 FILLER_80_594 ();
 b15zdnd11an1n32x5 FILLER_80_600 ();
 b15zdnd11an1n16x5 FILLER_80_632 ();
 b15zdnd11an1n08x5 FILLER_80_648 ();
 b15zdnd11an1n04x5 FILLER_80_656 ();
 b15zdnd00an1n02x5 FILLER_80_660 ();
 b15zdnd11an1n04x5 FILLER_80_672 ();
 b15zdnd11an1n16x5 FILLER_80_680 ();
 b15zdnd00an1n01x5 FILLER_80_696 ();
 b15zdnd11an1n04x5 FILLER_80_701 ();
 b15zdnd00an1n02x5 FILLER_80_705 ();
 b15zdnd00an1n02x5 FILLER_80_716 ();
 b15zdnd11an1n32x5 FILLER_80_726 ();
 b15zdnd11an1n08x5 FILLER_80_758 ();
 b15zdnd11an1n04x5 FILLER_80_766 ();
 b15zdnd11an1n04x5 FILLER_80_774 ();
 b15zdnd11an1n16x5 FILLER_80_794 ();
 b15zdnd11an1n08x5 FILLER_80_810 ();
 b15zdnd00an1n01x5 FILLER_80_818 ();
 b15zdnd11an1n16x5 FILLER_80_825 ();
 b15zdnd11an1n08x5 FILLER_80_841 ();
 b15zdnd00an1n02x5 FILLER_80_849 ();
 b15zdnd11an1n16x5 FILLER_80_855 ();
 b15zdnd11an1n08x5 FILLER_80_871 ();
 b15zdnd11an1n04x5 FILLER_80_879 ();
 b15zdnd00an1n02x5 FILLER_80_883 ();
 b15zdnd11an1n64x5 FILLER_80_911 ();
 b15zdnd11an1n64x5 FILLER_80_975 ();
 b15zdnd11an1n64x5 FILLER_80_1039 ();
 b15zdnd11an1n64x5 FILLER_80_1103 ();
 b15zdnd11an1n08x5 FILLER_80_1167 ();
 b15zdnd00an1n02x5 FILLER_80_1175 ();
 b15zdnd11an1n64x5 FILLER_80_1197 ();
 b15zdnd11an1n32x5 FILLER_80_1261 ();
 b15zdnd11an1n04x5 FILLER_80_1293 ();
 b15zdnd00an1n02x5 FILLER_80_1297 ();
 b15zdnd11an1n04x5 FILLER_80_1331 ();
 b15zdnd11an1n32x5 FILLER_80_1345 ();
 b15zdnd11an1n08x5 FILLER_80_1377 ();
 b15zdnd11an1n04x5 FILLER_80_1385 ();
 b15zdnd00an1n01x5 FILLER_80_1389 ();
 b15zdnd11an1n64x5 FILLER_80_1397 ();
 b15zdnd11an1n64x5 FILLER_80_1461 ();
 b15zdnd11an1n04x5 FILLER_80_1525 ();
 b15zdnd00an1n01x5 FILLER_80_1529 ();
 b15zdnd11an1n04x5 FILLER_80_1535 ();
 b15zdnd11an1n04x5 FILLER_80_1552 ();
 b15zdnd11an1n04x5 FILLER_80_1562 ();
 b15zdnd11an1n32x5 FILLER_80_1587 ();
 b15zdnd11an1n08x5 FILLER_80_1619 ();
 b15zdnd11an1n04x5 FILLER_80_1627 ();
 b15zdnd11an1n32x5 FILLER_80_1643 ();
 b15zdnd11an1n08x5 FILLER_80_1675 ();
 b15zdnd11an1n08x5 FILLER_80_1703 ();
 b15zdnd00an1n02x5 FILLER_80_1711 ();
 b15zdnd00an1n01x5 FILLER_80_1713 ();
 b15zdnd11an1n32x5 FILLER_80_1723 ();
 b15zdnd00an1n02x5 FILLER_80_1755 ();
 b15zdnd11an1n32x5 FILLER_80_1773 ();
 b15zdnd11an1n04x5 FILLER_80_1828 ();
 b15zdnd11an1n16x5 FILLER_80_1845 ();
 b15zdnd11an1n08x5 FILLER_80_1861 ();
 b15zdnd00an1n01x5 FILLER_80_1869 ();
 b15zdnd11an1n16x5 FILLER_80_1878 ();
 b15zdnd11an1n08x5 FILLER_80_1894 ();
 b15zdnd11an1n04x5 FILLER_80_1902 ();
 b15zdnd00an1n01x5 FILLER_80_1906 ();
 b15zdnd11an1n04x5 FILLER_80_1916 ();
 b15zdnd11an1n64x5 FILLER_80_1928 ();
 b15zdnd11an1n64x5 FILLER_80_1992 ();
 b15zdnd11an1n64x5 FILLER_80_2056 ();
 b15zdnd11an1n08x5 FILLER_80_2120 ();
 b15zdnd11an1n04x5 FILLER_80_2128 ();
 b15zdnd00an1n01x5 FILLER_80_2132 ();
 b15zdnd11an1n16x5 FILLER_80_2137 ();
 b15zdnd00an1n01x5 FILLER_80_2153 ();
 b15zdnd11an1n08x5 FILLER_80_2162 ();
 b15zdnd11an1n04x5 FILLER_80_2170 ();
 b15zdnd00an1n02x5 FILLER_80_2174 ();
 b15zdnd11an1n64x5 FILLER_80_2182 ();
 b15zdnd11an1n16x5 FILLER_80_2246 ();
 b15zdnd11an1n08x5 FILLER_80_2262 ();
 b15zdnd11an1n04x5 FILLER_80_2270 ();
 b15zdnd00an1n02x5 FILLER_80_2274 ();
 b15zdnd11an1n64x5 FILLER_81_0 ();
 b15zdnd11an1n16x5 FILLER_81_64 ();
 b15zdnd11an1n08x5 FILLER_81_80 ();
 b15zdnd11an1n04x5 FILLER_81_88 ();
 b15zdnd00an1n01x5 FILLER_81_92 ();
 b15zdnd11an1n08x5 FILLER_81_111 ();
 b15zdnd11an1n04x5 FILLER_81_119 ();
 b15zdnd11an1n16x5 FILLER_81_129 ();
 b15zdnd11an1n08x5 FILLER_81_145 ();
 b15zdnd11an1n04x5 FILLER_81_153 ();
 b15zdnd00an1n01x5 FILLER_81_157 ();
 b15zdnd11an1n08x5 FILLER_81_163 ();
 b15zdnd00an1n01x5 FILLER_81_171 ();
 b15zdnd11an1n16x5 FILLER_81_192 ();
 b15zdnd11an1n04x5 FILLER_81_208 ();
 b15zdnd00an1n02x5 FILLER_81_212 ();
 b15zdnd00an1n01x5 FILLER_81_214 ();
 b15zdnd11an1n32x5 FILLER_81_220 ();
 b15zdnd11an1n04x5 FILLER_81_252 ();
 b15zdnd00an1n02x5 FILLER_81_256 ();
 b15zdnd11an1n32x5 FILLER_81_263 ();
 b15zdnd00an1n01x5 FILLER_81_295 ();
 b15zdnd11an1n64x5 FILLER_81_303 ();
 b15zdnd11an1n64x5 FILLER_81_367 ();
 b15zdnd11an1n08x5 FILLER_81_431 ();
 b15zdnd11an1n04x5 FILLER_81_439 ();
 b15zdnd00an1n02x5 FILLER_81_443 ();
 b15zdnd11an1n64x5 FILLER_81_461 ();
 b15zdnd11an1n64x5 FILLER_81_525 ();
 b15zdnd11an1n08x5 FILLER_81_589 ();
 b15zdnd00an1n02x5 FILLER_81_597 ();
 b15zdnd00an1n01x5 FILLER_81_599 ();
 b15zdnd11an1n04x5 FILLER_81_623 ();
 b15zdnd11an1n08x5 FILLER_81_632 ();
 b15zdnd00an1n01x5 FILLER_81_640 ();
 b15zdnd11an1n08x5 FILLER_81_647 ();
 b15zdnd11an1n04x5 FILLER_81_655 ();
 b15zdnd11an1n64x5 FILLER_81_669 ();
 b15zdnd11an1n08x5 FILLER_81_742 ();
 b15zdnd11an1n04x5 FILLER_81_750 ();
 b15zdnd00an1n02x5 FILLER_81_754 ();
 b15zdnd00an1n01x5 FILLER_81_756 ();
 b15zdnd11an1n32x5 FILLER_81_762 ();
 b15zdnd11an1n16x5 FILLER_81_794 ();
 b15zdnd11an1n08x5 FILLER_81_810 ();
 b15zdnd00an1n01x5 FILLER_81_818 ();
 b15zdnd11an1n32x5 FILLER_81_826 ();
 b15zdnd11an1n16x5 FILLER_81_858 ();
 b15zdnd11an1n08x5 FILLER_81_874 ();
 b15zdnd11an1n04x5 FILLER_81_882 ();
 b15zdnd00an1n02x5 FILLER_81_886 ();
 b15zdnd11an1n64x5 FILLER_81_919 ();
 b15zdnd11an1n64x5 FILLER_81_983 ();
 b15zdnd11an1n08x5 FILLER_81_1047 ();
 b15zdnd11an1n04x5 FILLER_81_1055 ();
 b15zdnd00an1n02x5 FILLER_81_1059 ();
 b15zdnd11an1n64x5 FILLER_81_1081 ();
 b15zdnd11an1n32x5 FILLER_81_1145 ();
 b15zdnd11an1n16x5 FILLER_81_1177 ();
 b15zdnd11an1n08x5 FILLER_81_1193 ();
 b15zdnd11an1n64x5 FILLER_81_1207 ();
 b15zdnd11an1n16x5 FILLER_81_1271 ();
 b15zdnd11an1n64x5 FILLER_81_1296 ();
 b15zdnd11an1n08x5 FILLER_81_1360 ();
 b15zdnd00an1n02x5 FILLER_81_1368 ();
 b15zdnd11an1n64x5 FILLER_81_1386 ();
 b15zdnd11an1n64x5 FILLER_81_1450 ();
 b15zdnd11an1n32x5 FILLER_81_1514 ();
 b15zdnd11an1n16x5 FILLER_81_1546 ();
 b15zdnd11an1n04x5 FILLER_81_1562 ();
 b15zdnd11an1n04x5 FILLER_81_1570 ();
 b15zdnd11an1n04x5 FILLER_81_1586 ();
 b15zdnd11an1n08x5 FILLER_81_1596 ();
 b15zdnd00an1n01x5 FILLER_81_1604 ();
 b15zdnd11an1n04x5 FILLER_81_1617 ();
 b15zdnd11an1n04x5 FILLER_81_1647 ();
 b15zdnd11an1n04x5 FILLER_81_1657 ();
 b15zdnd11an1n64x5 FILLER_81_1666 ();
 b15zdnd11an1n16x5 FILLER_81_1730 ();
 b15zdnd11an1n08x5 FILLER_81_1746 ();
 b15zdnd00an1n02x5 FILLER_81_1754 ();
 b15zdnd11an1n08x5 FILLER_81_1760 ();
 b15zdnd00an1n02x5 FILLER_81_1768 ();
 b15zdnd11an1n32x5 FILLER_81_1777 ();
 b15zdnd00an1n01x5 FILLER_81_1809 ();
 b15zdnd11an1n64x5 FILLER_81_1841 ();
 b15zdnd11an1n16x5 FILLER_81_1905 ();
 b15zdnd11an1n04x5 FILLER_81_1921 ();
 b15zdnd11an1n32x5 FILLER_81_1937 ();
 b15zdnd11an1n08x5 FILLER_81_1969 ();
 b15zdnd11an1n04x5 FILLER_81_1977 ();
 b15zdnd11an1n16x5 FILLER_81_1986 ();
 b15zdnd11an1n08x5 FILLER_81_2002 ();
 b15zdnd11an1n04x5 FILLER_81_2010 ();
 b15zdnd00an1n02x5 FILLER_81_2014 ();
 b15zdnd11an1n04x5 FILLER_81_2022 ();
 b15zdnd11an1n32x5 FILLER_81_2030 ();
 b15zdnd11an1n16x5 FILLER_81_2062 ();
 b15zdnd00an1n02x5 FILLER_81_2078 ();
 b15zdnd11an1n64x5 FILLER_81_2087 ();
 b15zdnd00an1n02x5 FILLER_81_2151 ();
 b15zdnd11an1n16x5 FILLER_81_2157 ();
 b15zdnd11an1n04x5 FILLER_81_2173 ();
 b15zdnd00an1n02x5 FILLER_81_2177 ();
 b15zdnd00an1n01x5 FILLER_81_2179 ();
 b15zdnd11an1n64x5 FILLER_81_2190 ();
 b15zdnd11an1n16x5 FILLER_81_2254 ();
 b15zdnd11an1n08x5 FILLER_81_2270 ();
 b15zdnd11an1n04x5 FILLER_81_2278 ();
 b15zdnd00an1n02x5 FILLER_81_2282 ();
 b15zdnd11an1n16x5 FILLER_82_8 ();
 b15zdnd11an1n08x5 FILLER_82_24 ();
 b15zdnd11an1n04x5 FILLER_82_32 ();
 b15zdnd00an1n02x5 FILLER_82_36 ();
 b15zdnd00an1n01x5 FILLER_82_38 ();
 b15zdnd11an1n08x5 FILLER_82_55 ();
 b15zdnd11an1n04x5 FILLER_82_63 ();
 b15zdnd00an1n02x5 FILLER_82_67 ();
 b15zdnd00an1n01x5 FILLER_82_69 ();
 b15zdnd11an1n04x5 FILLER_82_77 ();
 b15zdnd00an1n02x5 FILLER_82_81 ();
 b15zdnd00an1n01x5 FILLER_82_83 ();
 b15zdnd11an1n08x5 FILLER_82_89 ();
 b15zdnd11an1n04x5 FILLER_82_97 ();
 b15zdnd00an1n02x5 FILLER_82_101 ();
 b15zdnd11an1n64x5 FILLER_82_110 ();
 b15zdnd11an1n32x5 FILLER_82_174 ();
 b15zdnd11an1n04x5 FILLER_82_206 ();
 b15zdnd00an1n01x5 FILLER_82_210 ();
 b15zdnd11an1n16x5 FILLER_82_221 ();
 b15zdnd11an1n08x5 FILLER_82_237 ();
 b15zdnd00an1n02x5 FILLER_82_245 ();
 b15zdnd11an1n32x5 FILLER_82_254 ();
 b15zdnd11an1n08x5 FILLER_82_286 ();
 b15zdnd11an1n04x5 FILLER_82_294 ();
 b15zdnd00an1n02x5 FILLER_82_298 ();
 b15zdnd11an1n32x5 FILLER_82_310 ();
 b15zdnd11an1n16x5 FILLER_82_342 ();
 b15zdnd11an1n04x5 FILLER_82_365 ();
 b15zdnd11an1n04x5 FILLER_82_377 ();
 b15zdnd00an1n02x5 FILLER_82_381 ();
 b15zdnd11an1n64x5 FILLER_82_409 ();
 b15zdnd11an1n08x5 FILLER_82_473 ();
 b15zdnd11an1n04x5 FILLER_82_501 ();
 b15zdnd11an1n32x5 FILLER_82_536 ();
 b15zdnd00an1n01x5 FILLER_82_568 ();
 b15zdnd11an1n32x5 FILLER_82_574 ();
 b15zdnd11an1n08x5 FILLER_82_606 ();
 b15zdnd11an1n04x5 FILLER_82_614 ();
 b15zdnd00an1n01x5 FILLER_82_618 ();
 b15zdnd11an1n04x5 FILLER_82_632 ();
 b15zdnd11an1n16x5 FILLER_82_646 ();
 b15zdnd11an1n04x5 FILLER_82_662 ();
 b15zdnd11an1n04x5 FILLER_82_671 ();
 b15zdnd00an1n02x5 FILLER_82_675 ();
 b15zdnd11an1n16x5 FILLER_82_687 ();
 b15zdnd11an1n08x5 FILLER_82_703 ();
 b15zdnd11an1n04x5 FILLER_82_711 ();
 b15zdnd00an1n02x5 FILLER_82_715 ();
 b15zdnd00an1n01x5 FILLER_82_717 ();
 b15zdnd11an1n16x5 FILLER_82_726 ();
 b15zdnd11an1n08x5 FILLER_82_742 ();
 b15zdnd11an1n04x5 FILLER_82_750 ();
 b15zdnd00an1n02x5 FILLER_82_754 ();
 b15zdnd00an1n01x5 FILLER_82_756 ();
 b15zdnd11an1n16x5 FILLER_82_762 ();
 b15zdnd11an1n08x5 FILLER_82_778 ();
 b15zdnd11an1n04x5 FILLER_82_786 ();
 b15zdnd00an1n02x5 FILLER_82_790 ();
 b15zdnd00an1n01x5 FILLER_82_792 ();
 b15zdnd11an1n64x5 FILLER_82_797 ();
 b15zdnd11an1n64x5 FILLER_82_861 ();
 b15zdnd11an1n16x5 FILLER_82_925 ();
 b15zdnd11an1n08x5 FILLER_82_941 ();
 b15zdnd11an1n04x5 FILLER_82_949 ();
 b15zdnd00an1n02x5 FILLER_82_953 ();
 b15zdnd00an1n01x5 FILLER_82_955 ();
 b15zdnd11an1n04x5 FILLER_82_976 ();
 b15zdnd11an1n32x5 FILLER_82_989 ();
 b15zdnd11an1n04x5 FILLER_82_1021 ();
 b15zdnd00an1n01x5 FILLER_82_1025 ();
 b15zdnd11an1n32x5 FILLER_82_1030 ();
 b15zdnd11an1n04x5 FILLER_82_1062 ();
 b15zdnd11an1n08x5 FILLER_82_1084 ();
 b15zdnd11an1n04x5 FILLER_82_1092 ();
 b15zdnd00an1n01x5 FILLER_82_1096 ();
 b15zdnd11an1n32x5 FILLER_82_1102 ();
 b15zdnd00an1n02x5 FILLER_82_1134 ();
 b15zdnd11an1n32x5 FILLER_82_1161 ();
 b15zdnd11an1n64x5 FILLER_82_1213 ();
 b15zdnd11an1n04x5 FILLER_82_1277 ();
 b15zdnd00an1n02x5 FILLER_82_1281 ();
 b15zdnd00an1n01x5 FILLER_82_1283 ();
 b15zdnd11an1n04x5 FILLER_82_1298 ();
 b15zdnd11an1n04x5 FILLER_82_1320 ();
 b15zdnd00an1n02x5 FILLER_82_1324 ();
 b15zdnd00an1n01x5 FILLER_82_1326 ();
 b15zdnd11an1n16x5 FILLER_82_1345 ();
 b15zdnd00an1n01x5 FILLER_82_1361 ();
 b15zdnd11an1n08x5 FILLER_82_1368 ();
 b15zdnd11an1n04x5 FILLER_82_1376 ();
 b15zdnd00an1n02x5 FILLER_82_1380 ();
 b15zdnd11an1n04x5 FILLER_82_1403 ();
 b15zdnd00an1n02x5 FILLER_82_1407 ();
 b15zdnd11an1n32x5 FILLER_82_1418 ();
 b15zdnd11an1n08x5 FILLER_82_1450 ();
 b15zdnd11an1n04x5 FILLER_82_1458 ();
 b15zdnd11an1n04x5 FILLER_82_1467 ();
 b15zdnd00an1n01x5 FILLER_82_1471 ();
 b15zdnd11an1n08x5 FILLER_82_1478 ();
 b15zdnd11an1n04x5 FILLER_82_1486 ();
 b15zdnd00an1n02x5 FILLER_82_1490 ();
 b15zdnd00an1n01x5 FILLER_82_1492 ();
 b15zdnd11an1n64x5 FILLER_82_1507 ();
 b15zdnd11an1n16x5 FILLER_82_1571 ();
 b15zdnd11an1n08x5 FILLER_82_1587 ();
 b15zdnd11an1n04x5 FILLER_82_1595 ();
 b15zdnd11an1n32x5 FILLER_82_1625 ();
 b15zdnd11an1n08x5 FILLER_82_1657 ();
 b15zdnd00an1n01x5 FILLER_82_1665 ();
 b15zdnd11an1n64x5 FILLER_82_1692 ();
 b15zdnd11an1n32x5 FILLER_82_1756 ();
 b15zdnd11an1n08x5 FILLER_82_1788 ();
 b15zdnd11an1n04x5 FILLER_82_1796 ();
 b15zdnd00an1n02x5 FILLER_82_1800 ();
 b15zdnd11an1n64x5 FILLER_82_1809 ();
 b15zdnd11an1n32x5 FILLER_82_1873 ();
 b15zdnd11an1n16x5 FILLER_82_1905 ();
 b15zdnd11an1n08x5 FILLER_82_1921 ();
 b15zdnd11an1n16x5 FILLER_82_1946 ();
 b15zdnd11an1n08x5 FILLER_82_1962 ();
 b15zdnd00an1n01x5 FILLER_82_1970 ();
 b15zdnd11an1n16x5 FILLER_82_1985 ();
 b15zdnd11an1n08x5 FILLER_82_2001 ();
 b15zdnd11an1n04x5 FILLER_82_2009 ();
 b15zdnd11an1n32x5 FILLER_82_2022 ();
 b15zdnd00an1n01x5 FILLER_82_2054 ();
 b15zdnd11an1n64x5 FILLER_82_2061 ();
 b15zdnd11an1n08x5 FILLER_82_2131 ();
 b15zdnd11an1n04x5 FILLER_82_2139 ();
 b15zdnd00an1n01x5 FILLER_82_2143 ();
 b15zdnd00an1n02x5 FILLER_82_2152 ();
 b15zdnd11an1n16x5 FILLER_82_2162 ();
 b15zdnd11an1n04x5 FILLER_82_2192 ();
 b15zdnd11an1n64x5 FILLER_82_2206 ();
 b15zdnd11an1n04x5 FILLER_82_2270 ();
 b15zdnd00an1n02x5 FILLER_82_2274 ();
 b15zdnd11an1n64x5 FILLER_83_0 ();
 b15zdnd11an1n16x5 FILLER_83_64 ();
 b15zdnd11an1n04x5 FILLER_83_80 ();
 b15zdnd00an1n02x5 FILLER_83_84 ();
 b15zdnd00an1n01x5 FILLER_83_86 ();
 b15zdnd11an1n16x5 FILLER_83_108 ();
 b15zdnd11an1n64x5 FILLER_83_138 ();
 b15zdnd11an1n64x5 FILLER_83_202 ();
 b15zdnd11an1n08x5 FILLER_83_266 ();
 b15zdnd11an1n04x5 FILLER_83_274 ();
 b15zdnd00an1n02x5 FILLER_83_278 ();
 b15zdnd00an1n01x5 FILLER_83_280 ();
 b15zdnd11an1n32x5 FILLER_83_286 ();
 b15zdnd11an1n08x5 FILLER_83_318 ();
 b15zdnd11an1n04x5 FILLER_83_326 ();
 b15zdnd11an1n04x5 FILLER_83_356 ();
 b15zdnd11an1n32x5 FILLER_83_380 ();
 b15zdnd11an1n16x5 FILLER_83_412 ();
 b15zdnd11an1n04x5 FILLER_83_438 ();
 b15zdnd11an1n32x5 FILLER_83_458 ();
 b15zdnd11an1n08x5 FILLER_83_490 ();
 b15zdnd11an1n04x5 FILLER_83_498 ();
 b15zdnd00an1n01x5 FILLER_83_502 ();
 b15zdnd11an1n32x5 FILLER_83_512 ();
 b15zdnd11an1n16x5 FILLER_83_544 ();
 b15zdnd11an1n04x5 FILLER_83_560 ();
 b15zdnd00an1n02x5 FILLER_83_564 ();
 b15zdnd11an1n16x5 FILLER_83_576 ();
 b15zdnd00an1n02x5 FILLER_83_592 ();
 b15zdnd11an1n16x5 FILLER_83_610 ();
 b15zdnd11an1n08x5 FILLER_83_626 ();
 b15zdnd00an1n01x5 FILLER_83_634 ();
 b15zdnd11an1n32x5 FILLER_83_650 ();
 b15zdnd00an1n02x5 FILLER_83_682 ();
 b15zdnd11an1n04x5 FILLER_83_709 ();
 b15zdnd11an1n16x5 FILLER_83_723 ();
 b15zdnd11an1n08x5 FILLER_83_739 ();
 b15zdnd00an1n01x5 FILLER_83_747 ();
 b15zdnd11an1n32x5 FILLER_83_758 ();
 b15zdnd00an1n02x5 FILLER_83_790 ();
 b15zdnd11an1n16x5 FILLER_83_799 ();
 b15zdnd11an1n08x5 FILLER_83_815 ();
 b15zdnd11an1n04x5 FILLER_83_823 ();
 b15zdnd00an1n01x5 FILLER_83_827 ();
 b15zdnd11an1n08x5 FILLER_83_833 ();
 b15zdnd11an1n04x5 FILLER_83_841 ();
 b15zdnd00an1n02x5 FILLER_83_845 ();
 b15zdnd11an1n08x5 FILLER_83_852 ();
 b15zdnd00an1n02x5 FILLER_83_860 ();
 b15zdnd11an1n16x5 FILLER_83_876 ();
 b15zdnd11an1n08x5 FILLER_83_892 ();
 b15zdnd11an1n04x5 FILLER_83_900 ();
 b15zdnd11an1n64x5 FILLER_83_922 ();
 b15zdnd11an1n32x5 FILLER_83_986 ();
 b15zdnd00an1n02x5 FILLER_83_1018 ();
 b15zdnd11an1n64x5 FILLER_83_1025 ();
 b15zdnd11an1n16x5 FILLER_83_1089 ();
 b15zdnd11an1n08x5 FILLER_83_1105 ();
 b15zdnd11an1n04x5 FILLER_83_1113 ();
 b15zdnd00an1n02x5 FILLER_83_1117 ();
 b15zdnd11an1n32x5 FILLER_83_1150 ();
 b15zdnd11an1n04x5 FILLER_83_1182 ();
 b15zdnd11an1n08x5 FILLER_83_1190 ();
 b15zdnd11an1n04x5 FILLER_83_1198 ();
 b15zdnd11an1n64x5 FILLER_83_1207 ();
 b15zdnd11an1n16x5 FILLER_83_1271 ();
 b15zdnd00an1n02x5 FILLER_83_1287 ();
 b15zdnd11an1n32x5 FILLER_83_1309 ();
 b15zdnd11an1n08x5 FILLER_83_1341 ();
 b15zdnd00an1n01x5 FILLER_83_1349 ();
 b15zdnd11an1n08x5 FILLER_83_1360 ();
 b15zdnd11an1n04x5 FILLER_83_1368 ();
 b15zdnd00an1n02x5 FILLER_83_1372 ();
 b15zdnd11an1n16x5 FILLER_83_1384 ();
 b15zdnd11an1n08x5 FILLER_83_1400 ();
 b15zdnd00an1n01x5 FILLER_83_1408 ();
 b15zdnd11an1n04x5 FILLER_83_1413 ();
 b15zdnd11an1n16x5 FILLER_83_1429 ();
 b15zdnd00an1n01x5 FILLER_83_1445 ();
 b15zdnd11an1n32x5 FILLER_83_1453 ();
 b15zdnd11an1n08x5 FILLER_83_1485 ();
 b15zdnd00an1n01x5 FILLER_83_1493 ();
 b15zdnd11an1n04x5 FILLER_83_1506 ();
 b15zdnd11an1n64x5 FILLER_83_1522 ();
 b15zdnd11an1n16x5 FILLER_83_1586 ();
 b15zdnd11an1n08x5 FILLER_83_1602 ();
 b15zdnd11an1n04x5 FILLER_83_1610 ();
 b15zdnd11an1n04x5 FILLER_83_1623 ();
 b15zdnd11an1n04x5 FILLER_83_1642 ();
 b15zdnd11an1n04x5 FILLER_83_1661 ();
 b15zdnd00an1n01x5 FILLER_83_1665 ();
 b15zdnd11an1n64x5 FILLER_83_1682 ();
 b15zdnd11an1n64x5 FILLER_83_1746 ();
 b15zdnd11an1n16x5 FILLER_83_1810 ();
 b15zdnd00an1n02x5 FILLER_83_1826 ();
 b15zdnd00an1n01x5 FILLER_83_1828 ();
 b15zdnd11an1n04x5 FILLER_83_1839 ();
 b15zdnd00an1n02x5 FILLER_83_1843 ();
 b15zdnd11an1n32x5 FILLER_83_1853 ();
 b15zdnd11an1n04x5 FILLER_83_1885 ();
 b15zdnd00an1n02x5 FILLER_83_1889 ();
 b15zdnd11an1n04x5 FILLER_83_1901 ();
 b15zdnd11an1n64x5 FILLER_83_1921 ();
 b15zdnd11an1n32x5 FILLER_83_1985 ();
 b15zdnd11an1n16x5 FILLER_83_2017 ();
 b15zdnd11an1n08x5 FILLER_83_2033 ();
 b15zdnd11an1n04x5 FILLER_83_2041 ();
 b15zdnd00an1n02x5 FILLER_83_2045 ();
 b15zdnd00an1n01x5 FILLER_83_2047 ();
 b15zdnd11an1n32x5 FILLER_83_2054 ();
 b15zdnd11an1n08x5 FILLER_83_2086 ();
 b15zdnd11an1n04x5 FILLER_83_2094 ();
 b15zdnd11an1n04x5 FILLER_83_2103 ();
 b15zdnd11an1n16x5 FILLER_83_2112 ();
 b15zdnd00an1n02x5 FILLER_83_2128 ();
 b15zdnd11an1n16x5 FILLER_83_2135 ();
 b15zdnd11an1n04x5 FILLER_83_2151 ();
 b15zdnd11an1n16x5 FILLER_83_2163 ();
 b15zdnd00an1n02x5 FILLER_83_2179 ();
 b15zdnd11an1n04x5 FILLER_83_2195 ();
 b15zdnd11an1n32x5 FILLER_83_2223 ();
 b15zdnd11an1n16x5 FILLER_83_2255 ();
 b15zdnd11an1n08x5 FILLER_83_2271 ();
 b15zdnd11an1n04x5 FILLER_83_2279 ();
 b15zdnd00an1n01x5 FILLER_83_2283 ();
 b15zdnd11an1n64x5 FILLER_84_8 ();
 b15zdnd11an1n04x5 FILLER_84_72 ();
 b15zdnd00an1n02x5 FILLER_84_76 ();
 b15zdnd11an1n32x5 FILLER_84_88 ();
 b15zdnd11an1n64x5 FILLER_84_130 ();
 b15zdnd11an1n16x5 FILLER_84_194 ();
 b15zdnd11an1n04x5 FILLER_84_210 ();
 b15zdnd11an1n04x5 FILLER_84_220 ();
 b15zdnd11an1n16x5 FILLER_84_230 ();
 b15zdnd00an1n02x5 FILLER_84_246 ();
 b15zdnd00an1n01x5 FILLER_84_248 ();
 b15zdnd11an1n16x5 FILLER_84_261 ();
 b15zdnd11an1n04x5 FILLER_84_277 ();
 b15zdnd00an1n02x5 FILLER_84_281 ();
 b15zdnd11an1n04x5 FILLER_84_297 ();
 b15zdnd11an1n08x5 FILLER_84_307 ();
 b15zdnd11an1n04x5 FILLER_84_315 ();
 b15zdnd11an1n04x5 FILLER_84_329 ();
 b15zdnd11an1n04x5 FILLER_84_354 ();
 b15zdnd00an1n02x5 FILLER_84_358 ();
 b15zdnd11an1n32x5 FILLER_84_378 ();
 b15zdnd11an1n16x5 FILLER_84_410 ();
 b15zdnd11an1n08x5 FILLER_84_426 ();
 b15zdnd11an1n04x5 FILLER_84_434 ();
 b15zdnd00an1n01x5 FILLER_84_438 ();
 b15zdnd11an1n16x5 FILLER_84_452 ();
 b15zdnd11an1n08x5 FILLER_84_468 ();
 b15zdnd11an1n04x5 FILLER_84_476 ();
 b15zdnd11an1n04x5 FILLER_84_488 ();
 b15zdnd11an1n16x5 FILLER_84_508 ();
 b15zdnd11an1n08x5 FILLER_84_524 ();
 b15zdnd11an1n04x5 FILLER_84_532 ();
 b15zdnd00an1n02x5 FILLER_84_536 ();
 b15zdnd11an1n04x5 FILLER_84_544 ();
 b15zdnd00an1n01x5 FILLER_84_548 ();
 b15zdnd11an1n64x5 FILLER_84_555 ();
 b15zdnd11an1n64x5 FILLER_84_619 ();
 b15zdnd11an1n08x5 FILLER_84_683 ();
 b15zdnd00an1n02x5 FILLER_84_691 ();
 b15zdnd11an1n16x5 FILLER_84_700 ();
 b15zdnd00an1n02x5 FILLER_84_716 ();
 b15zdnd11an1n16x5 FILLER_84_726 ();
 b15zdnd00an1n01x5 FILLER_84_742 ();
 b15zdnd11an1n04x5 FILLER_84_750 ();
 b15zdnd00an1n02x5 FILLER_84_754 ();
 b15zdnd11an1n08x5 FILLER_84_768 ();
 b15zdnd11an1n04x5 FILLER_84_792 ();
 b15zdnd11an1n16x5 FILLER_84_803 ();
 b15zdnd00an1n01x5 FILLER_84_819 ();
 b15zdnd11an1n04x5 FILLER_84_841 ();
 b15zdnd00an1n01x5 FILLER_84_845 ();
 b15zdnd11an1n04x5 FILLER_84_852 ();
 b15zdnd11an1n16x5 FILLER_84_871 ();
 b15zdnd11an1n08x5 FILLER_84_887 ();
 b15zdnd00an1n02x5 FILLER_84_895 ();
 b15zdnd11an1n32x5 FILLER_84_910 ();
 b15zdnd11an1n08x5 FILLER_84_942 ();
 b15zdnd11an1n04x5 FILLER_84_950 ();
 b15zdnd00an1n02x5 FILLER_84_954 ();
 b15zdnd11an1n04x5 FILLER_84_976 ();
 b15zdnd11an1n16x5 FILLER_84_992 ();
 b15zdnd11an1n04x5 FILLER_84_1008 ();
 b15zdnd00an1n02x5 FILLER_84_1012 ();
 b15zdnd11an1n32x5 FILLER_84_1034 ();
 b15zdnd11an1n16x5 FILLER_84_1066 ();
 b15zdnd11an1n08x5 FILLER_84_1082 ();
 b15zdnd11an1n04x5 FILLER_84_1090 ();
 b15zdnd00an1n02x5 FILLER_84_1094 ();
 b15zdnd11an1n32x5 FILLER_84_1116 ();
 b15zdnd11an1n16x5 FILLER_84_1148 ();
 b15zdnd11an1n08x5 FILLER_84_1164 ();
 b15zdnd00an1n02x5 FILLER_84_1172 ();
 b15zdnd11an1n32x5 FILLER_84_1200 ();
 b15zdnd11an1n08x5 FILLER_84_1232 ();
 b15zdnd00an1n01x5 FILLER_84_1240 ();
 b15zdnd11an1n08x5 FILLER_84_1245 ();
 b15zdnd11an1n16x5 FILLER_84_1279 ();
 b15zdnd00an1n01x5 FILLER_84_1295 ();
 b15zdnd11an1n04x5 FILLER_84_1327 ();
 b15zdnd11an1n64x5 FILLER_84_1363 ();
 b15zdnd11an1n16x5 FILLER_84_1427 ();
 b15zdnd11an1n08x5 FILLER_84_1443 ();
 b15zdnd00an1n01x5 FILLER_84_1451 ();
 b15zdnd11an1n08x5 FILLER_84_1464 ();
 b15zdnd00an1n02x5 FILLER_84_1472 ();
 b15zdnd11an1n04x5 FILLER_84_1479 ();
 b15zdnd11an1n16x5 FILLER_84_1509 ();
 b15zdnd11an1n08x5 FILLER_84_1525 ();
 b15zdnd00an1n01x5 FILLER_84_1533 ();
 b15zdnd11an1n32x5 FILLER_84_1548 ();
 b15zdnd11an1n08x5 FILLER_84_1580 ();
 b15zdnd11an1n04x5 FILLER_84_1588 ();
 b15zdnd00an1n02x5 FILLER_84_1592 ();
 b15zdnd00an1n01x5 FILLER_84_1594 ();
 b15zdnd11an1n08x5 FILLER_84_1618 ();
 b15zdnd11an1n16x5 FILLER_84_1635 ();
 b15zdnd11an1n64x5 FILLER_84_1657 ();
 b15zdnd11an1n16x5 FILLER_84_1721 ();
 b15zdnd11an1n08x5 FILLER_84_1737 ();
 b15zdnd11an1n04x5 FILLER_84_1745 ();
 b15zdnd11an1n04x5 FILLER_84_1758 ();
 b15zdnd11an1n08x5 FILLER_84_1771 ();
 b15zdnd00an1n02x5 FILLER_84_1779 ();
 b15zdnd00an1n01x5 FILLER_84_1781 ();
 b15zdnd11an1n08x5 FILLER_84_1787 ();
 b15zdnd11an1n04x5 FILLER_84_1795 ();
 b15zdnd00an1n02x5 FILLER_84_1799 ();
 b15zdnd11an1n16x5 FILLER_84_1807 ();
 b15zdnd11an1n08x5 FILLER_84_1823 ();
 b15zdnd11an1n04x5 FILLER_84_1831 ();
 b15zdnd00an1n02x5 FILLER_84_1835 ();
 b15zdnd11an1n16x5 FILLER_84_1853 ();
 b15zdnd11an1n04x5 FILLER_84_1884 ();
 b15zdnd11an1n08x5 FILLER_84_1897 ();
 b15zdnd11an1n04x5 FILLER_84_1910 ();
 b15zdnd11an1n08x5 FILLER_84_1919 ();
 b15zdnd00an1n02x5 FILLER_84_1927 ();
 b15zdnd11an1n04x5 FILLER_84_1939 ();
 b15zdnd11an1n32x5 FILLER_84_1948 ();
 b15zdnd11an1n04x5 FILLER_84_1980 ();
 b15zdnd11an1n16x5 FILLER_84_1994 ();
 b15zdnd11an1n08x5 FILLER_84_2010 ();
 b15zdnd11an1n04x5 FILLER_84_2030 ();
 b15zdnd11an1n16x5 FILLER_84_2048 ();
 b15zdnd11an1n16x5 FILLER_84_2071 ();
 b15zdnd11an1n08x5 FILLER_84_2087 ();
 b15zdnd00an1n02x5 FILLER_84_2095 ();
 b15zdnd00an1n01x5 FILLER_84_2097 ();
 b15zdnd11an1n16x5 FILLER_84_2105 ();
 b15zdnd11an1n04x5 FILLER_84_2121 ();
 b15zdnd00an1n01x5 FILLER_84_2125 ();
 b15zdnd11an1n04x5 FILLER_84_2133 ();
 b15zdnd11an1n04x5 FILLER_84_2150 ();
 b15zdnd11an1n32x5 FILLER_84_2162 ();
 b15zdnd11an1n16x5 FILLER_84_2194 ();
 b15zdnd11an1n32x5 FILLER_84_2214 ();
 b15zdnd11an1n16x5 FILLER_84_2246 ();
 b15zdnd11an1n08x5 FILLER_84_2262 ();
 b15zdnd11an1n04x5 FILLER_84_2270 ();
 b15zdnd00an1n02x5 FILLER_84_2274 ();
 b15zdnd11an1n32x5 FILLER_85_0 ();
 b15zdnd11an1n16x5 FILLER_85_32 ();
 b15zdnd11an1n08x5 FILLER_85_48 ();
 b15zdnd00an1n02x5 FILLER_85_56 ();
 b15zdnd00an1n01x5 FILLER_85_58 ();
 b15zdnd11an1n04x5 FILLER_85_79 ();
 b15zdnd11an1n08x5 FILLER_85_109 ();
 b15zdnd11an1n04x5 FILLER_85_117 ();
 b15zdnd00an1n01x5 FILLER_85_121 ();
 b15zdnd11an1n16x5 FILLER_85_129 ();
 b15zdnd11an1n08x5 FILLER_85_145 ();
 b15zdnd00an1n02x5 FILLER_85_153 ();
 b15zdnd11an1n32x5 FILLER_85_164 ();
 b15zdnd00an1n01x5 FILLER_85_196 ();
 b15zdnd11an1n04x5 FILLER_85_204 ();
 b15zdnd00an1n02x5 FILLER_85_208 ();
 b15zdnd00an1n01x5 FILLER_85_210 ();
 b15zdnd11an1n32x5 FILLER_85_217 ();
 b15zdnd11an1n08x5 FILLER_85_249 ();
 b15zdnd11an1n04x5 FILLER_85_257 ();
 b15zdnd00an1n02x5 FILLER_85_261 ();
 b15zdnd00an1n01x5 FILLER_85_263 ();
 b15zdnd11an1n08x5 FILLER_85_290 ();
 b15zdnd00an1n02x5 FILLER_85_298 ();
 b15zdnd11an1n08x5 FILLER_85_320 ();
 b15zdnd11an1n04x5 FILLER_85_328 ();
 b15zdnd00an1n02x5 FILLER_85_332 ();
 b15zdnd00an1n01x5 FILLER_85_334 ();
 b15zdnd11an1n08x5 FILLER_85_361 ();
 b15zdnd11an1n04x5 FILLER_85_369 ();
 b15zdnd00an1n02x5 FILLER_85_373 ();
 b15zdnd00an1n01x5 FILLER_85_375 ();
 b15zdnd11an1n32x5 FILLER_85_402 ();
 b15zdnd11an1n16x5 FILLER_85_434 ();
 b15zdnd11an1n08x5 FILLER_85_450 ();
 b15zdnd11an1n04x5 FILLER_85_458 ();
 b15zdnd00an1n01x5 FILLER_85_462 ();
 b15zdnd11an1n16x5 FILLER_85_495 ();
 b15zdnd11an1n08x5 FILLER_85_511 ();
 b15zdnd00an1n02x5 FILLER_85_519 ();
 b15zdnd11an1n08x5 FILLER_85_527 ();
 b15zdnd00an1n02x5 FILLER_85_535 ();
 b15zdnd11an1n08x5 FILLER_85_544 ();
 b15zdnd00an1n02x5 FILLER_85_552 ();
 b15zdnd11an1n64x5 FILLER_85_561 ();
 b15zdnd11an1n08x5 FILLER_85_625 ();
 b15zdnd11an1n04x5 FILLER_85_633 ();
 b15zdnd11an1n64x5 FILLER_85_649 ();
 b15zdnd11an1n32x5 FILLER_85_713 ();
 b15zdnd11an1n16x5 FILLER_85_745 ();
 b15zdnd11an1n08x5 FILLER_85_761 ();
 b15zdnd11an1n16x5 FILLER_85_781 ();
 b15zdnd11an1n08x5 FILLER_85_797 ();
 b15zdnd11an1n04x5 FILLER_85_805 ();
 b15zdnd00an1n01x5 FILLER_85_809 ();
 b15zdnd11an1n08x5 FILLER_85_826 ();
 b15zdnd11an1n04x5 FILLER_85_834 ();
 b15zdnd00an1n01x5 FILLER_85_838 ();
 b15zdnd11an1n16x5 FILLER_85_844 ();
 b15zdnd00an1n02x5 FILLER_85_860 ();
 b15zdnd11an1n16x5 FILLER_85_868 ();
 b15zdnd00an1n02x5 FILLER_85_884 ();
 b15zdnd11an1n04x5 FILLER_85_917 ();
 b15zdnd11an1n08x5 FILLER_85_941 ();
 b15zdnd00an1n02x5 FILLER_85_949 ();
 b15zdnd11an1n08x5 FILLER_85_957 ();
 b15zdnd11an1n04x5 FILLER_85_965 ();
 b15zdnd00an1n01x5 FILLER_85_969 ();
 b15zdnd11an1n04x5 FILLER_85_975 ();
 b15zdnd00an1n02x5 FILLER_85_979 ();
 b15zdnd11an1n16x5 FILLER_85_1007 ();
 b15zdnd11an1n04x5 FILLER_85_1023 ();
 b15zdnd00an1n02x5 FILLER_85_1027 ();
 b15zdnd11an1n16x5 FILLER_85_1032 ();
 b15zdnd11an1n08x5 FILLER_85_1048 ();
 b15zdnd11an1n04x5 FILLER_85_1056 ();
 b15zdnd00an1n01x5 FILLER_85_1060 ();
 b15zdnd11an1n64x5 FILLER_85_1076 ();
 b15zdnd11an1n64x5 FILLER_85_1140 ();
 b15zdnd11an1n64x5 FILLER_85_1204 ();
 b15zdnd11an1n64x5 FILLER_85_1268 ();
 b15zdnd11an1n64x5 FILLER_85_1332 ();
 b15zdnd11an1n16x5 FILLER_85_1396 ();
 b15zdnd11an1n16x5 FILLER_85_1425 ();
 b15zdnd11an1n04x5 FILLER_85_1441 ();
 b15zdnd00an1n02x5 FILLER_85_1445 ();
 b15zdnd11an1n04x5 FILLER_85_1457 ();
 b15zdnd11an1n04x5 FILLER_85_1468 ();
 b15zdnd00an1n02x5 FILLER_85_1472 ();
 b15zdnd00an1n01x5 FILLER_85_1474 ();
 b15zdnd11an1n08x5 FILLER_85_1490 ();
 b15zdnd11an1n04x5 FILLER_85_1498 ();
 b15zdnd00an1n02x5 FILLER_85_1502 ();
 b15zdnd00an1n01x5 FILLER_85_1504 ();
 b15zdnd11an1n16x5 FILLER_85_1512 ();
 b15zdnd11an1n04x5 FILLER_85_1528 ();
 b15zdnd11an1n16x5 FILLER_85_1544 ();
 b15zdnd00an1n02x5 FILLER_85_1560 ();
 b15zdnd00an1n01x5 FILLER_85_1562 ();
 b15zdnd11an1n64x5 FILLER_85_1587 ();
 b15zdnd11an1n64x5 FILLER_85_1651 ();
 b15zdnd11an1n32x5 FILLER_85_1715 ();
 b15zdnd00an1n01x5 FILLER_85_1747 ();
 b15zdnd11an1n04x5 FILLER_85_1755 ();
 b15zdnd11an1n32x5 FILLER_85_1764 ();
 b15zdnd11an1n08x5 FILLER_85_1796 ();
 b15zdnd11an1n04x5 FILLER_85_1804 ();
 b15zdnd11an1n08x5 FILLER_85_1814 ();
 b15zdnd11an1n04x5 FILLER_85_1822 ();
 b15zdnd00an1n01x5 FILLER_85_1826 ();
 b15zdnd11an1n16x5 FILLER_85_1831 ();
 b15zdnd00an1n01x5 FILLER_85_1847 ();
 b15zdnd11an1n32x5 FILLER_85_1854 ();
 b15zdnd11an1n16x5 FILLER_85_1886 ();
 b15zdnd11an1n08x5 FILLER_85_1902 ();
 b15zdnd00an1n01x5 FILLER_85_1910 ();
 b15zdnd11an1n08x5 FILLER_85_1921 ();
 b15zdnd00an1n01x5 FILLER_85_1929 ();
 b15zdnd11an1n16x5 FILLER_85_1940 ();
 b15zdnd11an1n08x5 FILLER_85_1956 ();
 b15zdnd00an1n02x5 FILLER_85_1964 ();
 b15zdnd00an1n01x5 FILLER_85_1966 ();
 b15zdnd11an1n08x5 FILLER_85_1976 ();
 b15zdnd00an1n01x5 FILLER_85_1984 ();
 b15zdnd11an1n32x5 FILLER_85_1991 ();
 b15zdnd11an1n08x5 FILLER_85_2023 ();
 b15zdnd11an1n04x5 FILLER_85_2031 ();
 b15zdnd11an1n64x5 FILLER_85_2051 ();
 b15zdnd11an1n32x5 FILLER_85_2115 ();
 b15zdnd11an1n08x5 FILLER_85_2147 ();
 b15zdnd00an1n01x5 FILLER_85_2155 ();
 b15zdnd11an1n04x5 FILLER_85_2167 ();
 b15zdnd11an1n08x5 FILLER_85_2184 ();
 b15zdnd00an1n02x5 FILLER_85_2192 ();
 b15zdnd00an1n01x5 FILLER_85_2194 ();
 b15zdnd11an1n64x5 FILLER_85_2216 ();
 b15zdnd11an1n04x5 FILLER_85_2280 ();
 b15zdnd11an1n32x5 FILLER_86_8 ();
 b15zdnd11an1n04x5 FILLER_86_40 ();
 b15zdnd11an1n16x5 FILLER_86_52 ();
 b15zdnd00an1n02x5 FILLER_86_68 ();
 b15zdnd00an1n01x5 FILLER_86_70 ();
 b15zdnd11an1n08x5 FILLER_86_89 ();
 b15zdnd11an1n04x5 FILLER_86_97 ();
 b15zdnd00an1n02x5 FILLER_86_101 ();
 b15zdnd11an1n04x5 FILLER_86_108 ();
 b15zdnd11an1n08x5 FILLER_86_118 ();
 b15zdnd00an1n02x5 FILLER_86_126 ();
 b15zdnd11an1n16x5 FILLER_86_132 ();
 b15zdnd11an1n08x5 FILLER_86_148 ();
 b15zdnd00an1n01x5 FILLER_86_156 ();
 b15zdnd11an1n04x5 FILLER_86_171 ();
 b15zdnd00an1n02x5 FILLER_86_175 ();
 b15zdnd11an1n64x5 FILLER_86_186 ();
 b15zdnd11an1n08x5 FILLER_86_250 ();
 b15zdnd11an1n04x5 FILLER_86_282 ();
 b15zdnd11an1n04x5 FILLER_86_312 ();
 b15zdnd11an1n04x5 FILLER_86_329 ();
 b15zdnd11an1n04x5 FILLER_86_338 ();
 b15zdnd11an1n08x5 FILLER_86_347 ();
 b15zdnd00an1n02x5 FILLER_86_355 ();
 b15zdnd11an1n04x5 FILLER_86_377 ();
 b15zdnd11an1n64x5 FILLER_86_394 ();
 b15zdnd11an1n64x5 FILLER_86_458 ();
 b15zdnd00an1n02x5 FILLER_86_522 ();
 b15zdnd11an1n16x5 FILLER_86_528 ();
 b15zdnd11an1n08x5 FILLER_86_544 ();
 b15zdnd11an1n04x5 FILLER_86_552 ();
 b15zdnd00an1n02x5 FILLER_86_556 ();
 b15zdnd00an1n01x5 FILLER_86_558 ();
 b15zdnd11an1n08x5 FILLER_86_580 ();
 b15zdnd11an1n04x5 FILLER_86_588 ();
 b15zdnd00an1n01x5 FILLER_86_592 ();
 b15zdnd11an1n32x5 FILLER_86_598 ();
 b15zdnd11an1n04x5 FILLER_86_630 ();
 b15zdnd00an1n02x5 FILLER_86_634 ();
 b15zdnd00an1n01x5 FILLER_86_636 ();
 b15zdnd11an1n16x5 FILLER_86_642 ();
 b15zdnd00an1n02x5 FILLER_86_658 ();
 b15zdnd11an1n16x5 FILLER_86_678 ();
 b15zdnd11an1n16x5 FILLER_86_699 ();
 b15zdnd00an1n02x5 FILLER_86_715 ();
 b15zdnd00an1n01x5 FILLER_86_717 ();
 b15zdnd11an1n64x5 FILLER_86_726 ();
 b15zdnd11an1n32x5 FILLER_86_790 ();
 b15zdnd11an1n08x5 FILLER_86_822 ();
 b15zdnd11an1n04x5 FILLER_86_830 ();
 b15zdnd11an1n16x5 FILLER_86_846 ();
 b15zdnd00an1n02x5 FILLER_86_862 ();
 b15zdnd11an1n16x5 FILLER_86_869 ();
 b15zdnd11an1n08x5 FILLER_86_885 ();
 b15zdnd11an1n04x5 FILLER_86_893 ();
 b15zdnd11an1n64x5 FILLER_86_902 ();
 b15zdnd11an1n64x5 FILLER_86_966 ();
 b15zdnd11an1n32x5 FILLER_86_1030 ();
 b15zdnd11an1n16x5 FILLER_86_1062 ();
 b15zdnd11an1n04x5 FILLER_86_1078 ();
 b15zdnd11an1n64x5 FILLER_86_1100 ();
 b15zdnd11an1n08x5 FILLER_86_1164 ();
 b15zdnd00an1n02x5 FILLER_86_1172 ();
 b15zdnd00an1n01x5 FILLER_86_1174 ();
 b15zdnd11an1n16x5 FILLER_86_1179 ();
 b15zdnd11an1n04x5 FILLER_86_1195 ();
 b15zdnd00an1n02x5 FILLER_86_1199 ();
 b15zdnd11an1n04x5 FILLER_86_1232 ();
 b15zdnd11an1n16x5 FILLER_86_1241 ();
 b15zdnd00an1n02x5 FILLER_86_1257 ();
 b15zdnd00an1n01x5 FILLER_86_1259 ();
 b15zdnd11an1n32x5 FILLER_86_1278 ();
 b15zdnd11an1n08x5 FILLER_86_1310 ();
 b15zdnd00an1n02x5 FILLER_86_1318 ();
 b15zdnd00an1n01x5 FILLER_86_1320 ();
 b15zdnd11an1n04x5 FILLER_86_1353 ();
 b15zdnd11an1n04x5 FILLER_86_1371 ();
 b15zdnd11an1n08x5 FILLER_86_1391 ();
 b15zdnd00an1n02x5 FILLER_86_1399 ();
 b15zdnd00an1n01x5 FILLER_86_1401 ();
 b15zdnd11an1n08x5 FILLER_86_1408 ();
 b15zdnd00an1n01x5 FILLER_86_1416 ();
 b15zdnd11an1n32x5 FILLER_86_1421 ();
 b15zdnd11an1n16x5 FILLER_86_1453 ();
 b15zdnd11an1n08x5 FILLER_86_1469 ();
 b15zdnd11an1n04x5 FILLER_86_1477 ();
 b15zdnd11an1n32x5 FILLER_86_1488 ();
 b15zdnd11an1n08x5 FILLER_86_1520 ();
 b15zdnd00an1n01x5 FILLER_86_1528 ();
 b15zdnd11an1n04x5 FILLER_86_1533 ();
 b15zdnd11an1n04x5 FILLER_86_1543 ();
 b15zdnd11an1n16x5 FILLER_86_1559 ();
 b15zdnd11an1n08x5 FILLER_86_1575 ();
 b15zdnd11an1n04x5 FILLER_86_1583 ();
 b15zdnd00an1n02x5 FILLER_86_1587 ();
 b15zdnd00an1n01x5 FILLER_86_1589 ();
 b15zdnd11an1n04x5 FILLER_86_1616 ();
 b15zdnd11an1n04x5 FILLER_86_1626 ();
 b15zdnd11an1n64x5 FILLER_86_1656 ();
 b15zdnd11an1n32x5 FILLER_86_1720 ();
 b15zdnd11an1n04x5 FILLER_86_1752 ();
 b15zdnd00an1n02x5 FILLER_86_1756 ();
 b15zdnd11an1n64x5 FILLER_86_1765 ();
 b15zdnd11an1n16x5 FILLER_86_1829 ();
 b15zdnd11an1n08x5 FILLER_86_1845 ();
 b15zdnd11an1n04x5 FILLER_86_1853 ();
 b15zdnd00an1n02x5 FILLER_86_1857 ();
 b15zdnd00an1n01x5 FILLER_86_1859 ();
 b15zdnd11an1n04x5 FILLER_86_1866 ();
 b15zdnd11an1n04x5 FILLER_86_1876 ();
 b15zdnd11an1n04x5 FILLER_86_1896 ();
 b15zdnd11an1n16x5 FILLER_86_1910 ();
 b15zdnd11an1n08x5 FILLER_86_1926 ();
 b15zdnd11an1n04x5 FILLER_86_1934 ();
 b15zdnd00an1n01x5 FILLER_86_1938 ();
 b15zdnd11an1n08x5 FILLER_86_1949 ();
 b15zdnd11an1n04x5 FILLER_86_1961 ();
 b15zdnd11an1n16x5 FILLER_86_1985 ();
 b15zdnd11an1n08x5 FILLER_86_2001 ();
 b15zdnd11an1n16x5 FILLER_86_2014 ();
 b15zdnd11an1n08x5 FILLER_86_2030 ();
 b15zdnd11an1n08x5 FILLER_86_2051 ();
 b15zdnd11an1n04x5 FILLER_86_2059 ();
 b15zdnd00an1n02x5 FILLER_86_2063 ();
 b15zdnd11an1n32x5 FILLER_86_2071 ();
 b15zdnd00an1n02x5 FILLER_86_2103 ();
 b15zdnd11an1n32x5 FILLER_86_2119 ();
 b15zdnd00an1n02x5 FILLER_86_2151 ();
 b15zdnd00an1n01x5 FILLER_86_2153 ();
 b15zdnd11an1n08x5 FILLER_86_2162 ();
 b15zdnd00an1n02x5 FILLER_86_2170 ();
 b15zdnd00an1n01x5 FILLER_86_2172 ();
 b15zdnd11an1n16x5 FILLER_86_2181 ();
 b15zdnd11an1n08x5 FILLER_86_2197 ();
 b15zdnd00an1n01x5 FILLER_86_2205 ();
 b15zdnd11an1n32x5 FILLER_86_2218 ();
 b15zdnd11an1n16x5 FILLER_86_2250 ();
 b15zdnd11an1n08x5 FILLER_86_2266 ();
 b15zdnd00an1n02x5 FILLER_86_2274 ();
 b15zdnd11an1n32x5 FILLER_87_0 ();
 b15zdnd11an1n08x5 FILLER_87_32 ();
 b15zdnd00an1n01x5 FILLER_87_40 ();
 b15zdnd11an1n04x5 FILLER_87_50 ();
 b15zdnd00an1n01x5 FILLER_87_54 ();
 b15zdnd11an1n64x5 FILLER_87_65 ();
 b15zdnd11an1n04x5 FILLER_87_142 ();
 b15zdnd00an1n02x5 FILLER_87_146 ();
 b15zdnd00an1n01x5 FILLER_87_148 ();
 b15zdnd11an1n04x5 FILLER_87_159 ();
 b15zdnd00an1n01x5 FILLER_87_163 ();
 b15zdnd11an1n16x5 FILLER_87_176 ();
 b15zdnd00an1n01x5 FILLER_87_192 ();
 b15zdnd11an1n32x5 FILLER_87_203 ();
 b15zdnd11an1n08x5 FILLER_87_235 ();
 b15zdnd00an1n02x5 FILLER_87_243 ();
 b15zdnd11an1n64x5 FILLER_87_252 ();
 b15zdnd11an1n16x5 FILLER_87_316 ();
 b15zdnd11an1n08x5 FILLER_87_332 ();
 b15zdnd11an1n04x5 FILLER_87_347 ();
 b15zdnd11an1n64x5 FILLER_87_361 ();
 b15zdnd11an1n08x5 FILLER_87_425 ();
 b15zdnd11an1n04x5 FILLER_87_433 ();
 b15zdnd11an1n32x5 FILLER_87_446 ();
 b15zdnd11an1n08x5 FILLER_87_478 ();
 b15zdnd11an1n04x5 FILLER_87_486 ();
 b15zdnd11an1n04x5 FILLER_87_497 ();
 b15zdnd11an1n32x5 FILLER_87_506 ();
 b15zdnd11an1n08x5 FILLER_87_538 ();
 b15zdnd11an1n04x5 FILLER_87_546 ();
 b15zdnd11an1n08x5 FILLER_87_564 ();
 b15zdnd11an1n04x5 FILLER_87_572 ();
 b15zdnd00an1n02x5 FILLER_87_576 ();
 b15zdnd11an1n04x5 FILLER_87_584 ();
 b15zdnd00an1n01x5 FILLER_87_588 ();
 b15zdnd11an1n04x5 FILLER_87_596 ();
 b15zdnd00an1n02x5 FILLER_87_600 ();
 b15zdnd11an1n08x5 FILLER_87_608 ();
 b15zdnd11an1n04x5 FILLER_87_616 ();
 b15zdnd00an1n02x5 FILLER_87_620 ();
 b15zdnd00an1n01x5 FILLER_87_622 ();
 b15zdnd11an1n08x5 FILLER_87_634 ();
 b15zdnd00an1n02x5 FILLER_87_642 ();
 b15zdnd11an1n32x5 FILLER_87_659 ();
 b15zdnd00an1n01x5 FILLER_87_691 ();
 b15zdnd11an1n04x5 FILLER_87_705 ();
 b15zdnd00an1n02x5 FILLER_87_709 ();
 b15zdnd00an1n01x5 FILLER_87_711 ();
 b15zdnd11an1n04x5 FILLER_87_724 ();
 b15zdnd00an1n01x5 FILLER_87_728 ();
 b15zdnd11an1n04x5 FILLER_87_753 ();
 b15zdnd00an1n02x5 FILLER_87_757 ();
 b15zdnd00an1n01x5 FILLER_87_759 ();
 b15zdnd11an1n64x5 FILLER_87_767 ();
 b15zdnd11an1n32x5 FILLER_87_831 ();
 b15zdnd11an1n08x5 FILLER_87_863 ();
 b15zdnd11an1n04x5 FILLER_87_871 ();
 b15zdnd00an1n02x5 FILLER_87_875 ();
 b15zdnd11an1n08x5 FILLER_87_884 ();
 b15zdnd00an1n02x5 FILLER_87_892 ();
 b15zdnd11an1n64x5 FILLER_87_911 ();
 b15zdnd11an1n64x5 FILLER_87_975 ();
 b15zdnd11an1n32x5 FILLER_87_1039 ();
 b15zdnd11an1n08x5 FILLER_87_1071 ();
 b15zdnd11an1n04x5 FILLER_87_1079 ();
 b15zdnd00an1n02x5 FILLER_87_1083 ();
 b15zdnd00an1n01x5 FILLER_87_1085 ();
 b15zdnd11an1n64x5 FILLER_87_1090 ();
 b15zdnd11an1n16x5 FILLER_87_1154 ();
 b15zdnd11an1n04x5 FILLER_87_1170 ();
 b15zdnd00an1n01x5 FILLER_87_1174 ();
 b15zdnd11an1n32x5 FILLER_87_1200 ();
 b15zdnd11an1n04x5 FILLER_87_1232 ();
 b15zdnd00an1n01x5 FILLER_87_1236 ();
 b15zdnd11an1n16x5 FILLER_87_1255 ();
 b15zdnd11an1n08x5 FILLER_87_1271 ();
 b15zdnd00an1n02x5 FILLER_87_1279 ();
 b15zdnd00an1n01x5 FILLER_87_1281 ();
 b15zdnd11an1n04x5 FILLER_87_1292 ();
 b15zdnd11an1n64x5 FILLER_87_1307 ();
 b15zdnd11an1n08x5 FILLER_87_1371 ();
 b15zdnd11an1n04x5 FILLER_87_1379 ();
 b15zdnd00an1n02x5 FILLER_87_1383 ();
 b15zdnd00an1n01x5 FILLER_87_1385 ();
 b15zdnd11an1n32x5 FILLER_87_1393 ();
 b15zdnd11an1n16x5 FILLER_87_1425 ();
 b15zdnd00an1n02x5 FILLER_87_1441 ();
 b15zdnd00an1n01x5 FILLER_87_1443 ();
 b15zdnd11an1n16x5 FILLER_87_1453 ();
 b15zdnd11an1n04x5 FILLER_87_1469 ();
 b15zdnd00an1n02x5 FILLER_87_1473 ();
 b15zdnd11an1n64x5 FILLER_87_1486 ();
 b15zdnd11an1n16x5 FILLER_87_1550 ();
 b15zdnd11an1n08x5 FILLER_87_1566 ();
 b15zdnd11an1n04x5 FILLER_87_1574 ();
 b15zdnd11an1n16x5 FILLER_87_1591 ();
 b15zdnd11an1n08x5 FILLER_87_1607 ();
 b15zdnd00an1n02x5 FILLER_87_1615 ();
 b15zdnd00an1n01x5 FILLER_87_1617 ();
 b15zdnd11an1n32x5 FILLER_87_1629 ();
 b15zdnd11an1n08x5 FILLER_87_1661 ();
 b15zdnd11an1n04x5 FILLER_87_1669 ();
 b15zdnd11an1n32x5 FILLER_87_1677 ();
 b15zdnd11an1n16x5 FILLER_87_1709 ();
 b15zdnd11an1n32x5 FILLER_87_1756 ();
 b15zdnd11an1n08x5 FILLER_87_1788 ();
 b15zdnd11an1n64x5 FILLER_87_1803 ();
 b15zdnd11an1n64x5 FILLER_87_1867 ();
 b15zdnd11an1n64x5 FILLER_87_1931 ();
 b15zdnd11an1n08x5 FILLER_87_1995 ();
 b15zdnd11an1n04x5 FILLER_87_2003 ();
 b15zdnd11an1n04x5 FILLER_87_2016 ();
 b15zdnd00an1n01x5 FILLER_87_2020 ();
 b15zdnd11an1n32x5 FILLER_87_2037 ();
 b15zdnd00an1n02x5 FILLER_87_2069 ();
 b15zdnd00an1n01x5 FILLER_87_2071 ();
 b15zdnd11an1n16x5 FILLER_87_2081 ();
 b15zdnd11an1n08x5 FILLER_87_2097 ();
 b15zdnd00an1n02x5 FILLER_87_2105 ();
 b15zdnd00an1n01x5 FILLER_87_2107 ();
 b15zdnd11an1n32x5 FILLER_87_2118 ();
 b15zdnd11an1n16x5 FILLER_87_2150 ();
 b15zdnd11an1n08x5 FILLER_87_2166 ();
 b15zdnd11an1n64x5 FILLER_87_2179 ();
 b15zdnd11an1n32x5 FILLER_87_2243 ();
 b15zdnd11an1n08x5 FILLER_87_2275 ();
 b15zdnd00an1n01x5 FILLER_87_2283 ();
 b15zdnd11an1n64x5 FILLER_88_8 ();
 b15zdnd11an1n16x5 FILLER_88_72 ();
 b15zdnd11an1n04x5 FILLER_88_94 ();
 b15zdnd00an1n02x5 FILLER_88_98 ();
 b15zdnd00an1n01x5 FILLER_88_100 ();
 b15zdnd11an1n64x5 FILLER_88_127 ();
 b15zdnd11an1n32x5 FILLER_88_195 ();
 b15zdnd11an1n16x5 FILLER_88_227 ();
 b15zdnd11an1n04x5 FILLER_88_243 ();
 b15zdnd00an1n02x5 FILLER_88_247 ();
 b15zdnd11an1n16x5 FILLER_88_253 ();
 b15zdnd11an1n08x5 FILLER_88_269 ();
 b15zdnd00an1n02x5 FILLER_88_277 ();
 b15zdnd00an1n01x5 FILLER_88_279 ();
 b15zdnd11an1n64x5 FILLER_88_291 ();
 b15zdnd11an1n08x5 FILLER_88_355 ();
 b15zdnd11an1n04x5 FILLER_88_363 ();
 b15zdnd11an1n32x5 FILLER_88_379 ();
 b15zdnd11an1n16x5 FILLER_88_411 ();
 b15zdnd11an1n04x5 FILLER_88_427 ();
 b15zdnd00an1n02x5 FILLER_88_431 ();
 b15zdnd00an1n01x5 FILLER_88_433 ();
 b15zdnd11an1n04x5 FILLER_88_442 ();
 b15zdnd11an1n08x5 FILLER_88_467 ();
 b15zdnd11an1n04x5 FILLER_88_475 ();
 b15zdnd00an1n01x5 FILLER_88_479 ();
 b15zdnd11an1n04x5 FILLER_88_485 ();
 b15zdnd00an1n02x5 FILLER_88_489 ();
 b15zdnd11an1n32x5 FILLER_88_503 ();
 b15zdnd11an1n04x5 FILLER_88_535 ();
 b15zdnd00an1n02x5 FILLER_88_539 ();
 b15zdnd11an1n04x5 FILLER_88_548 ();
 b15zdnd00an1n02x5 FILLER_88_552 ();
 b15zdnd11an1n64x5 FILLER_88_562 ();
 b15zdnd11an1n16x5 FILLER_88_626 ();
 b15zdnd00an1n02x5 FILLER_88_642 ();
 b15zdnd00an1n01x5 FILLER_88_644 ();
 b15zdnd11an1n08x5 FILLER_88_655 ();
 b15zdnd00an1n02x5 FILLER_88_663 ();
 b15zdnd11an1n04x5 FILLER_88_673 ();
 b15zdnd11an1n04x5 FILLER_88_689 ();
 b15zdnd11an1n16x5 FILLER_88_698 ();
 b15zdnd11an1n04x5 FILLER_88_714 ();
 b15zdnd11an1n04x5 FILLER_88_726 ();
 b15zdnd00an1n01x5 FILLER_88_730 ();
 b15zdnd11an1n04x5 FILLER_88_751 ();
 b15zdnd11an1n32x5 FILLER_88_767 ();
 b15zdnd11an1n08x5 FILLER_88_799 ();
 b15zdnd11an1n04x5 FILLER_88_807 ();
 b15zdnd11an1n64x5 FILLER_88_816 ();
 b15zdnd11an1n32x5 FILLER_88_880 ();
 b15zdnd11an1n08x5 FILLER_88_912 ();
 b15zdnd11an1n04x5 FILLER_88_920 ();
 b15zdnd11an1n16x5 FILLER_88_955 ();
 b15zdnd11an1n64x5 FILLER_88_975 ();
 b15zdnd11an1n16x5 FILLER_88_1039 ();
 b15zdnd11an1n04x5 FILLER_88_1055 ();
 b15zdnd00an1n02x5 FILLER_88_1059 ();
 b15zdnd11an1n32x5 FILLER_88_1092 ();
 b15zdnd11an1n16x5 FILLER_88_1124 ();
 b15zdnd11an1n08x5 FILLER_88_1140 ();
 b15zdnd11an1n16x5 FILLER_88_1168 ();
 b15zdnd11an1n08x5 FILLER_88_1184 ();
 b15zdnd11an1n04x5 FILLER_88_1192 ();
 b15zdnd00an1n01x5 FILLER_88_1196 ();
 b15zdnd11an1n64x5 FILLER_88_1201 ();
 b15zdnd11an1n32x5 FILLER_88_1265 ();
 b15zdnd00an1n02x5 FILLER_88_1297 ();
 b15zdnd00an1n01x5 FILLER_88_1299 ();
 b15zdnd11an1n16x5 FILLER_88_1320 ();
 b15zdnd11an1n08x5 FILLER_88_1336 ();
 b15zdnd00an1n02x5 FILLER_88_1344 ();
 b15zdnd11an1n08x5 FILLER_88_1372 ();
 b15zdnd11an1n04x5 FILLER_88_1380 ();
 b15zdnd11an1n08x5 FILLER_88_1391 ();
 b15zdnd11an1n04x5 FILLER_88_1399 ();
 b15zdnd00an1n02x5 FILLER_88_1403 ();
 b15zdnd11an1n32x5 FILLER_88_1417 ();
 b15zdnd00an1n02x5 FILLER_88_1449 ();
 b15zdnd00an1n01x5 FILLER_88_1451 ();
 b15zdnd11an1n16x5 FILLER_88_1461 ();
 b15zdnd00an1n02x5 FILLER_88_1477 ();
 b15zdnd00an1n01x5 FILLER_88_1479 ();
 b15zdnd11an1n08x5 FILLER_88_1485 ();
 b15zdnd00an1n02x5 FILLER_88_1493 ();
 b15zdnd11an1n04x5 FILLER_88_1500 ();
 b15zdnd00an1n02x5 FILLER_88_1504 ();
 b15zdnd00an1n01x5 FILLER_88_1506 ();
 b15zdnd11an1n16x5 FILLER_88_1519 ();
 b15zdnd11an1n08x5 FILLER_88_1535 ();
 b15zdnd00an1n01x5 FILLER_88_1543 ();
 b15zdnd11an1n64x5 FILLER_88_1557 ();
 b15zdnd11an1n64x5 FILLER_88_1621 ();
 b15zdnd00an1n01x5 FILLER_88_1685 ();
 b15zdnd11an1n64x5 FILLER_88_1691 ();
 b15zdnd11an1n16x5 FILLER_88_1755 ();
 b15zdnd11an1n08x5 FILLER_88_1771 ();
 b15zdnd00an1n01x5 FILLER_88_1779 ();
 b15zdnd11an1n04x5 FILLER_88_1785 ();
 b15zdnd00an1n02x5 FILLER_88_1789 ();
 b15zdnd11an1n08x5 FILLER_88_1797 ();
 b15zdnd00an1n02x5 FILLER_88_1805 ();
 b15zdnd11an1n04x5 FILLER_88_1831 ();
 b15zdnd11an1n64x5 FILLER_88_1848 ();
 b15zdnd11an1n64x5 FILLER_88_1912 ();
 b15zdnd11an1n08x5 FILLER_88_1976 ();
 b15zdnd00an1n02x5 FILLER_88_1984 ();
 b15zdnd11an1n32x5 FILLER_88_2006 ();
 b15zdnd11an1n16x5 FILLER_88_2038 ();
 b15zdnd11an1n08x5 FILLER_88_2054 ();
 b15zdnd11an1n04x5 FILLER_88_2062 ();
 b15zdnd00an1n02x5 FILLER_88_2066 ();
 b15zdnd00an1n01x5 FILLER_88_2068 ();
 b15zdnd11an1n32x5 FILLER_88_2074 ();
 b15zdnd00an1n02x5 FILLER_88_2106 ();
 b15zdnd11an1n32x5 FILLER_88_2115 ();
 b15zdnd11an1n04x5 FILLER_88_2147 ();
 b15zdnd00an1n02x5 FILLER_88_2151 ();
 b15zdnd00an1n01x5 FILLER_88_2153 ();
 b15zdnd11an1n08x5 FILLER_88_2162 ();
 b15zdnd00an1n02x5 FILLER_88_2170 ();
 b15zdnd00an1n01x5 FILLER_88_2172 ();
 b15zdnd11an1n64x5 FILLER_88_2177 ();
 b15zdnd11an1n32x5 FILLER_88_2241 ();
 b15zdnd00an1n02x5 FILLER_88_2273 ();
 b15zdnd00an1n01x5 FILLER_88_2275 ();
 b15zdnd11an1n32x5 FILLER_89_0 ();
 b15zdnd11an1n16x5 FILLER_89_32 ();
 b15zdnd11an1n08x5 FILLER_89_48 ();
 b15zdnd00an1n02x5 FILLER_89_56 ();
 b15zdnd00an1n01x5 FILLER_89_58 ();
 b15zdnd11an1n64x5 FILLER_89_67 ();
 b15zdnd11an1n64x5 FILLER_89_131 ();
 b15zdnd11an1n04x5 FILLER_89_195 ();
 b15zdnd11an1n04x5 FILLER_89_214 ();
 b15zdnd11an1n04x5 FILLER_89_222 ();
 b15zdnd00an1n02x5 FILLER_89_226 ();
 b15zdnd11an1n08x5 FILLER_89_233 ();
 b15zdnd11an1n04x5 FILLER_89_241 ();
 b15zdnd11an1n08x5 FILLER_89_259 ();
 b15zdnd00an1n01x5 FILLER_89_267 ();
 b15zdnd11an1n64x5 FILLER_89_276 ();
 b15zdnd11an1n16x5 FILLER_89_340 ();
 b15zdnd11an1n04x5 FILLER_89_356 ();
 b15zdnd00an1n01x5 FILLER_89_360 ();
 b15zdnd11an1n64x5 FILLER_89_377 ();
 b15zdnd11an1n16x5 FILLER_89_441 ();
 b15zdnd11an1n04x5 FILLER_89_457 ();
 b15zdnd00an1n02x5 FILLER_89_461 ();
 b15zdnd00an1n01x5 FILLER_89_463 ();
 b15zdnd11an1n32x5 FILLER_89_469 ();
 b15zdnd11an1n04x5 FILLER_89_501 ();
 b15zdnd00an1n02x5 FILLER_89_505 ();
 b15zdnd00an1n01x5 FILLER_89_507 ();
 b15zdnd11an1n04x5 FILLER_89_528 ();
 b15zdnd00an1n02x5 FILLER_89_532 ();
 b15zdnd00an1n01x5 FILLER_89_534 ();
 b15zdnd11an1n08x5 FILLER_89_543 ();
 b15zdnd00an1n01x5 FILLER_89_551 ();
 b15zdnd11an1n64x5 FILLER_89_556 ();
 b15zdnd11an1n04x5 FILLER_89_620 ();
 b15zdnd11an1n16x5 FILLER_89_630 ();
 b15zdnd00an1n02x5 FILLER_89_646 ();
 b15zdnd11an1n04x5 FILLER_89_663 ();
 b15zdnd11an1n64x5 FILLER_89_677 ();
 b15zdnd11an1n32x5 FILLER_89_741 ();
 b15zdnd11an1n04x5 FILLER_89_773 ();
 b15zdnd00an1n01x5 FILLER_89_777 ();
 b15zdnd11an1n04x5 FILLER_89_783 ();
 b15zdnd11an1n08x5 FILLER_89_797 ();
 b15zdnd00an1n01x5 FILLER_89_805 ();
 b15zdnd11an1n04x5 FILLER_89_812 ();
 b15zdnd11an1n16x5 FILLER_89_821 ();
 b15zdnd11an1n04x5 FILLER_89_837 ();
 b15zdnd11an1n64x5 FILLER_89_847 ();
 b15zdnd11an1n64x5 FILLER_89_911 ();
 b15zdnd11an1n32x5 FILLER_89_975 ();
 b15zdnd11an1n04x5 FILLER_89_1027 ();
 b15zdnd11an1n04x5 FILLER_89_1036 ();
 b15zdnd11an1n64x5 FILLER_89_1049 ();
 b15zdnd11an1n64x5 FILLER_89_1113 ();
 b15zdnd11an1n64x5 FILLER_89_1177 ();
 b15zdnd11an1n64x5 FILLER_89_1241 ();
 b15zdnd11an1n64x5 FILLER_89_1305 ();
 b15zdnd11an1n08x5 FILLER_89_1369 ();
 b15zdnd11an1n04x5 FILLER_89_1377 ();
 b15zdnd00an1n01x5 FILLER_89_1381 ();
 b15zdnd11an1n08x5 FILLER_89_1388 ();
 b15zdnd00an1n02x5 FILLER_89_1396 ();
 b15zdnd00an1n01x5 FILLER_89_1398 ();
 b15zdnd11an1n64x5 FILLER_89_1406 ();
 b15zdnd11an1n16x5 FILLER_89_1470 ();
 b15zdnd11an1n08x5 FILLER_89_1486 ();
 b15zdnd11an1n64x5 FILLER_89_1500 ();
 b15zdnd11an1n16x5 FILLER_89_1564 ();
 b15zdnd11an1n08x5 FILLER_89_1580 ();
 b15zdnd11an1n04x5 FILLER_89_1588 ();
 b15zdnd00an1n02x5 FILLER_89_1592 ();
 b15zdnd11an1n04x5 FILLER_89_1620 ();
 b15zdnd11an1n08x5 FILLER_89_1632 ();
 b15zdnd11an1n04x5 FILLER_89_1640 ();
 b15zdnd11an1n04x5 FILLER_89_1650 ();
 b15zdnd00an1n01x5 FILLER_89_1654 ();
 b15zdnd11an1n16x5 FILLER_89_1660 ();
 b15zdnd11an1n08x5 FILLER_89_1676 ();
 b15zdnd00an1n01x5 FILLER_89_1684 ();
 b15zdnd11an1n32x5 FILLER_89_1705 ();
 b15zdnd11an1n16x5 FILLER_89_1737 ();
 b15zdnd00an1n02x5 FILLER_89_1753 ();
 b15zdnd00an1n01x5 FILLER_89_1755 ();
 b15zdnd11an1n32x5 FILLER_89_1772 ();
 b15zdnd11an1n16x5 FILLER_89_1804 ();
 b15zdnd11an1n08x5 FILLER_89_1820 ();
 b15zdnd11an1n04x5 FILLER_89_1828 ();
 b15zdnd00an1n01x5 FILLER_89_1832 ();
 b15zdnd11an1n08x5 FILLER_89_1840 ();
 b15zdnd11an1n04x5 FILLER_89_1848 ();
 b15zdnd00an1n01x5 FILLER_89_1852 ();
 b15zdnd11an1n08x5 FILLER_89_1863 ();
 b15zdnd11an1n04x5 FILLER_89_1871 ();
 b15zdnd11an1n04x5 FILLER_89_1884 ();
 b15zdnd11an1n08x5 FILLER_89_1900 ();
 b15zdnd00an1n02x5 FILLER_89_1908 ();
 b15zdnd11an1n16x5 FILLER_89_1922 ();
 b15zdnd11an1n16x5 FILLER_89_1950 ();
 b15zdnd11an1n04x5 FILLER_89_1966 ();
 b15zdnd00an1n02x5 FILLER_89_1970 ();
 b15zdnd11an1n64x5 FILLER_89_1979 ();
 b15zdnd11an1n16x5 FILLER_89_2043 ();
 b15zdnd11an1n08x5 FILLER_89_2059 ();
 b15zdnd11an1n04x5 FILLER_89_2067 ();
 b15zdnd00an1n01x5 FILLER_89_2071 ();
 b15zdnd11an1n16x5 FILLER_89_2088 ();
 b15zdnd11an1n08x5 FILLER_89_2104 ();
 b15zdnd11an1n32x5 FILLER_89_2117 ();
 b15zdnd11an1n08x5 FILLER_89_2149 ();
 b15zdnd11an1n04x5 FILLER_89_2157 ();
 b15zdnd00an1n01x5 FILLER_89_2161 ();
 b15zdnd11an1n04x5 FILLER_89_2183 ();
 b15zdnd11an1n04x5 FILLER_89_2197 ();
 b15zdnd11an1n64x5 FILLER_89_2217 ();
 b15zdnd00an1n02x5 FILLER_89_2281 ();
 b15zdnd00an1n01x5 FILLER_89_2283 ();
 b15zdnd11an1n16x5 FILLER_90_8 ();
 b15zdnd11an1n08x5 FILLER_90_24 ();
 b15zdnd00an1n02x5 FILLER_90_32 ();
 b15zdnd00an1n01x5 FILLER_90_34 ();
 b15zdnd11an1n08x5 FILLER_90_53 ();
 b15zdnd00an1n02x5 FILLER_90_61 ();
 b15zdnd11an1n16x5 FILLER_90_78 ();
 b15zdnd11an1n08x5 FILLER_90_94 ();
 b15zdnd00an1n02x5 FILLER_90_102 ();
 b15zdnd00an1n01x5 FILLER_90_104 ();
 b15zdnd11an1n32x5 FILLER_90_112 ();
 b15zdnd11an1n04x5 FILLER_90_144 ();
 b15zdnd00an1n02x5 FILLER_90_148 ();
 b15zdnd11an1n16x5 FILLER_90_156 ();
 b15zdnd11an1n08x5 FILLER_90_172 ();
 b15zdnd11an1n04x5 FILLER_90_180 ();
 b15zdnd00an1n01x5 FILLER_90_184 ();
 b15zdnd11an1n32x5 FILLER_90_195 ();
 b15zdnd11an1n16x5 FILLER_90_227 ();
 b15zdnd00an1n02x5 FILLER_90_243 ();
 b15zdnd11an1n04x5 FILLER_90_251 ();
 b15zdnd00an1n02x5 FILLER_90_255 ();
 b15zdnd11an1n16x5 FILLER_90_261 ();
 b15zdnd00an1n01x5 FILLER_90_277 ();
 b15zdnd11an1n04x5 FILLER_90_285 ();
 b15zdnd11an1n32x5 FILLER_90_315 ();
 b15zdnd11an1n08x5 FILLER_90_347 ();
 b15zdnd11an1n04x5 FILLER_90_355 ();
 b15zdnd00an1n02x5 FILLER_90_359 ();
 b15zdnd11an1n32x5 FILLER_90_371 ();
 b15zdnd11an1n16x5 FILLER_90_403 ();
 b15zdnd11an1n08x5 FILLER_90_419 ();
 b15zdnd11an1n04x5 FILLER_90_427 ();
 b15zdnd11an1n32x5 FILLER_90_447 ();
 b15zdnd11an1n16x5 FILLER_90_479 ();
 b15zdnd00an1n01x5 FILLER_90_495 ();
 b15zdnd11an1n04x5 FILLER_90_509 ();
 b15zdnd11an1n64x5 FILLER_90_518 ();
 b15zdnd11an1n64x5 FILLER_90_582 ();
 b15zdnd11an1n32x5 FILLER_90_646 ();
 b15zdnd11an1n16x5 FILLER_90_678 ();
 b15zdnd11an1n04x5 FILLER_90_694 ();
 b15zdnd00an1n02x5 FILLER_90_698 ();
 b15zdnd00an1n02x5 FILLER_90_716 ();
 b15zdnd11an1n32x5 FILLER_90_726 ();
 b15zdnd11an1n08x5 FILLER_90_758 ();
 b15zdnd00an1n02x5 FILLER_90_766 ();
 b15zdnd11an1n08x5 FILLER_90_772 ();
 b15zdnd00an1n02x5 FILLER_90_780 ();
 b15zdnd11an1n08x5 FILLER_90_794 ();
 b15zdnd11an1n04x5 FILLER_90_802 ();
 b15zdnd00an1n01x5 FILLER_90_806 ();
 b15zdnd11an1n04x5 FILLER_90_820 ();
 b15zdnd11an1n04x5 FILLER_90_844 ();
 b15zdnd00an1n02x5 FILLER_90_848 ();
 b15zdnd11an1n16x5 FILLER_90_863 ();
 b15zdnd11an1n04x5 FILLER_90_879 ();
 b15zdnd11an1n08x5 FILLER_90_887 ();
 b15zdnd00an1n02x5 FILLER_90_895 ();
 b15zdnd11an1n32x5 FILLER_90_923 ();
 b15zdnd11an1n04x5 FILLER_90_955 ();
 b15zdnd00an1n01x5 FILLER_90_959 ();
 b15zdnd11an1n64x5 FILLER_90_965 ();
 b15zdnd11an1n32x5 FILLER_90_1029 ();
 b15zdnd11an1n16x5 FILLER_90_1061 ();
 b15zdnd11an1n08x5 FILLER_90_1077 ();
 b15zdnd11an1n08x5 FILLER_90_1105 ();
 b15zdnd11an1n04x5 FILLER_90_1113 ();
 b15zdnd00an1n02x5 FILLER_90_1117 ();
 b15zdnd11an1n64x5 FILLER_90_1134 ();
 b15zdnd11an1n64x5 FILLER_90_1198 ();
 b15zdnd11an1n04x5 FILLER_90_1262 ();
 b15zdnd11an1n64x5 FILLER_90_1272 ();
 b15zdnd11an1n64x5 FILLER_90_1336 ();
 b15zdnd11an1n64x5 FILLER_90_1400 ();
 b15zdnd11an1n32x5 FILLER_90_1464 ();
 b15zdnd11an1n16x5 FILLER_90_1496 ();
 b15zdnd11an1n04x5 FILLER_90_1512 ();
 b15zdnd11an1n08x5 FILLER_90_1548 ();
 b15zdnd11an1n04x5 FILLER_90_1556 ();
 b15zdnd00an1n02x5 FILLER_90_1560 ();
 b15zdnd11an1n04x5 FILLER_90_1588 ();
 b15zdnd11an1n16x5 FILLER_90_1596 ();
 b15zdnd11an1n04x5 FILLER_90_1612 ();
 b15zdnd00an1n01x5 FILLER_90_1616 ();
 b15zdnd11an1n04x5 FILLER_90_1643 ();
 b15zdnd11an1n16x5 FILLER_90_1667 ();
 b15zdnd11an1n08x5 FILLER_90_1683 ();
 b15zdnd11an1n04x5 FILLER_90_1691 ();
 b15zdnd00an1n01x5 FILLER_90_1695 ();
 b15zdnd11an1n64x5 FILLER_90_1699 ();
 b15zdnd11an1n32x5 FILLER_90_1763 ();
 b15zdnd11an1n04x5 FILLER_90_1795 ();
 b15zdnd11an1n64x5 FILLER_90_1809 ();
 b15zdnd11an1n16x5 FILLER_90_1873 ();
 b15zdnd11an1n08x5 FILLER_90_1889 ();
 b15zdnd00an1n01x5 FILLER_90_1897 ();
 b15zdnd11an1n04x5 FILLER_90_1904 ();
 b15zdnd11an1n32x5 FILLER_90_1929 ();
 b15zdnd11an1n08x5 FILLER_90_1961 ();
 b15zdnd11an1n04x5 FILLER_90_1969 ();
 b15zdnd11an1n16x5 FILLER_90_1977 ();
 b15zdnd00an1n02x5 FILLER_90_1993 ();
 b15zdnd00an1n01x5 FILLER_90_1995 ();
 b15zdnd11an1n16x5 FILLER_90_2001 ();
 b15zdnd11an1n08x5 FILLER_90_2017 ();
 b15zdnd11an1n04x5 FILLER_90_2025 ();
 b15zdnd00an1n02x5 FILLER_90_2029 ();
 b15zdnd11an1n32x5 FILLER_90_2036 ();
 b15zdnd00an1n02x5 FILLER_90_2068 ();
 b15zdnd11an1n32x5 FILLER_90_2074 ();
 b15zdnd11an1n08x5 FILLER_90_2106 ();
 b15zdnd00an1n01x5 FILLER_90_2114 ();
 b15zdnd11an1n04x5 FILLER_90_2125 ();
 b15zdnd11an1n08x5 FILLER_90_2144 ();
 b15zdnd00an1n02x5 FILLER_90_2152 ();
 b15zdnd11an1n08x5 FILLER_90_2162 ();
 b15zdnd00an1n02x5 FILLER_90_2170 ();
 b15zdnd11an1n04x5 FILLER_90_2186 ();
 b15zdnd00an1n02x5 FILLER_90_2190 ();
 b15zdnd00an1n01x5 FILLER_90_2192 ();
 b15zdnd11an1n64x5 FILLER_90_2198 ();
 b15zdnd11an1n08x5 FILLER_90_2262 ();
 b15zdnd11an1n04x5 FILLER_90_2270 ();
 b15zdnd00an1n02x5 FILLER_90_2274 ();
 b15zdnd11an1n32x5 FILLER_91_0 ();
 b15zdnd11an1n16x5 FILLER_91_32 ();
 b15zdnd00an1n02x5 FILLER_91_48 ();
 b15zdnd00an1n01x5 FILLER_91_50 ();
 b15zdnd11an1n04x5 FILLER_91_60 ();
 b15zdnd00an1n02x5 FILLER_91_64 ();
 b15zdnd00an1n01x5 FILLER_91_66 ();
 b15zdnd11an1n16x5 FILLER_91_74 ();
 b15zdnd11an1n08x5 FILLER_91_90 ();
 b15zdnd11an1n04x5 FILLER_91_98 ();
 b15zdnd00an1n02x5 FILLER_91_102 ();
 b15zdnd11an1n08x5 FILLER_91_112 ();
 b15zdnd11an1n04x5 FILLER_91_120 ();
 b15zdnd00an1n02x5 FILLER_91_124 ();
 b15zdnd00an1n01x5 FILLER_91_126 ();
 b15zdnd11an1n08x5 FILLER_91_134 ();
 b15zdnd00an1n02x5 FILLER_91_142 ();
 b15zdnd00an1n01x5 FILLER_91_144 ();
 b15zdnd11an1n16x5 FILLER_91_155 ();
 b15zdnd11an1n08x5 FILLER_91_171 ();
 b15zdnd00an1n02x5 FILLER_91_179 ();
 b15zdnd00an1n01x5 FILLER_91_181 ();
 b15zdnd11an1n64x5 FILLER_91_194 ();
 b15zdnd11an1n08x5 FILLER_91_258 ();
 b15zdnd00an1n01x5 FILLER_91_266 ();
 b15zdnd11an1n04x5 FILLER_91_281 ();
 b15zdnd00an1n01x5 FILLER_91_285 ();
 b15zdnd11an1n08x5 FILLER_91_292 ();
 b15zdnd11an1n04x5 FILLER_91_300 ();
 b15zdnd00an1n02x5 FILLER_91_304 ();
 b15zdnd11an1n04x5 FILLER_91_313 ();
 b15zdnd11an1n32x5 FILLER_91_326 ();
 b15zdnd11an1n04x5 FILLER_91_358 ();
 b15zdnd00an1n02x5 FILLER_91_362 ();
 b15zdnd00an1n01x5 FILLER_91_364 ();
 b15zdnd11an1n64x5 FILLER_91_391 ();
 b15zdnd11an1n08x5 FILLER_91_455 ();
 b15zdnd11an1n04x5 FILLER_91_463 ();
 b15zdnd11an1n16x5 FILLER_91_472 ();
 b15zdnd11an1n08x5 FILLER_91_488 ();
 b15zdnd11an1n04x5 FILLER_91_496 ();
 b15zdnd00an1n02x5 FILLER_91_500 ();
 b15zdnd11an1n64x5 FILLER_91_511 ();
 b15zdnd11an1n64x5 FILLER_91_575 ();
 b15zdnd11an1n32x5 FILLER_91_639 ();
 b15zdnd11an1n08x5 FILLER_91_671 ();
 b15zdnd11an1n64x5 FILLER_91_693 ();
 b15zdnd11an1n04x5 FILLER_91_757 ();
 b15zdnd11an1n64x5 FILLER_91_765 ();
 b15zdnd11an1n08x5 FILLER_91_829 ();
 b15zdnd11an1n04x5 FILLER_91_837 ();
 b15zdnd00an1n02x5 FILLER_91_841 ();
 b15zdnd11an1n08x5 FILLER_91_851 ();
 b15zdnd00an1n02x5 FILLER_91_859 ();
 b15zdnd00an1n01x5 FILLER_91_861 ();
 b15zdnd11an1n16x5 FILLER_91_871 ();
 b15zdnd11an1n04x5 FILLER_91_887 ();
 b15zdnd00an1n02x5 FILLER_91_891 ();
 b15zdnd11an1n32x5 FILLER_91_919 ();
 b15zdnd00an1n02x5 FILLER_91_951 ();
 b15zdnd11an1n32x5 FILLER_91_973 ();
 b15zdnd11an1n08x5 FILLER_91_1005 ();
 b15zdnd11an1n04x5 FILLER_91_1013 ();
 b15zdnd00an1n02x5 FILLER_91_1017 ();
 b15zdnd00an1n01x5 FILLER_91_1019 ();
 b15zdnd11an1n32x5 FILLER_91_1040 ();
 b15zdnd11an1n08x5 FILLER_91_1072 ();
 b15zdnd11an1n04x5 FILLER_91_1080 ();
 b15zdnd11an1n32x5 FILLER_91_1089 ();
 b15zdnd11an1n16x5 FILLER_91_1121 ();
 b15zdnd11an1n08x5 FILLER_91_1137 ();
 b15zdnd11an1n04x5 FILLER_91_1145 ();
 b15zdnd00an1n01x5 FILLER_91_1149 ();
 b15zdnd11an1n04x5 FILLER_91_1170 ();
 b15zdnd11an1n08x5 FILLER_91_1179 ();
 b15zdnd11an1n04x5 FILLER_91_1187 ();
 b15zdnd11an1n32x5 FILLER_91_1196 ();
 b15zdnd00an1n01x5 FILLER_91_1228 ();
 b15zdnd11an1n16x5 FILLER_91_1249 ();
 b15zdnd11an1n64x5 FILLER_91_1285 ();
 b15zdnd11an1n64x5 FILLER_91_1349 ();
 b15zdnd11an1n64x5 FILLER_91_1413 ();
 b15zdnd11an1n64x5 FILLER_91_1477 ();
 b15zdnd11an1n64x5 FILLER_91_1541 ();
 b15zdnd11an1n64x5 FILLER_91_1605 ();
 b15zdnd11an1n64x5 FILLER_91_1669 ();
 b15zdnd11an1n08x5 FILLER_91_1733 ();
 b15zdnd11an1n04x5 FILLER_91_1741 ();
 b15zdnd00an1n02x5 FILLER_91_1745 ();
 b15zdnd00an1n01x5 FILLER_91_1747 ();
 b15zdnd11an1n04x5 FILLER_91_1756 ();
 b15zdnd11an1n64x5 FILLER_91_1773 ();
 b15zdnd11an1n04x5 FILLER_91_1837 ();
 b15zdnd00an1n01x5 FILLER_91_1841 ();
 b15zdnd11an1n04x5 FILLER_91_1853 ();
 b15zdnd00an1n01x5 FILLER_91_1857 ();
 b15zdnd11an1n16x5 FILLER_91_1867 ();
 b15zdnd11an1n08x5 FILLER_91_1883 ();
 b15zdnd11an1n04x5 FILLER_91_1891 ();
 b15zdnd11an1n64x5 FILLER_91_1901 ();
 b15zdnd11an1n08x5 FILLER_91_1965 ();
 b15zdnd00an1n01x5 FILLER_91_1973 ();
 b15zdnd11an1n16x5 FILLER_91_1995 ();
 b15zdnd00an1n02x5 FILLER_91_2011 ();
 b15zdnd11an1n08x5 FILLER_91_2022 ();
 b15zdnd00an1n01x5 FILLER_91_2030 ();
 b15zdnd11an1n16x5 FILLER_91_2042 ();
 b15zdnd11an1n08x5 FILLER_91_2058 ();
 b15zdnd00an1n02x5 FILLER_91_2066 ();
 b15zdnd00an1n01x5 FILLER_91_2068 ();
 b15zdnd11an1n32x5 FILLER_91_2073 ();
 b15zdnd11an1n04x5 FILLER_91_2105 ();
 b15zdnd00an1n02x5 FILLER_91_2109 ();
 b15zdnd11an1n64x5 FILLER_91_2115 ();
 b15zdnd11an1n64x5 FILLER_91_2179 ();
 b15zdnd11an1n32x5 FILLER_91_2243 ();
 b15zdnd11an1n08x5 FILLER_91_2275 ();
 b15zdnd00an1n01x5 FILLER_91_2283 ();
 b15zdnd11an1n32x5 FILLER_92_8 ();
 b15zdnd11an1n04x5 FILLER_92_40 ();
 b15zdnd11an1n08x5 FILLER_92_50 ();
 b15zdnd11an1n04x5 FILLER_92_58 ();
 b15zdnd11an1n04x5 FILLER_92_71 ();
 b15zdnd00an1n02x5 FILLER_92_75 ();
 b15zdnd11an1n16x5 FILLER_92_83 ();
 b15zdnd00an1n02x5 FILLER_92_99 ();
 b15zdnd11an1n08x5 FILLER_92_106 ();
 b15zdnd11an1n04x5 FILLER_92_120 ();
 b15zdnd00an1n02x5 FILLER_92_124 ();
 b15zdnd00an1n01x5 FILLER_92_126 ();
 b15zdnd11an1n04x5 FILLER_92_133 ();
 b15zdnd11an1n04x5 FILLER_92_142 ();
 b15zdnd11an1n32x5 FILLER_92_152 ();
 b15zdnd11an1n32x5 FILLER_92_188 ();
 b15zdnd11an1n16x5 FILLER_92_220 ();
 b15zdnd00an1n02x5 FILLER_92_236 ();
 b15zdnd11an1n64x5 FILLER_92_256 ();
 b15zdnd11an1n04x5 FILLER_92_320 ();
 b15zdnd11an1n08x5 FILLER_92_350 ();
 b15zdnd11an1n04x5 FILLER_92_358 ();
 b15zdnd11an1n32x5 FILLER_92_378 ();
 b15zdnd11an1n16x5 FILLER_92_410 ();
 b15zdnd00an1n02x5 FILLER_92_426 ();
 b15zdnd11an1n16x5 FILLER_92_432 ();
 b15zdnd11an1n08x5 FILLER_92_448 ();
 b15zdnd11an1n04x5 FILLER_92_456 ();
 b15zdnd00an1n01x5 FILLER_92_460 ();
 b15zdnd11an1n04x5 FILLER_92_471 ();
 b15zdnd11an1n32x5 FILLER_92_481 ();
 b15zdnd11an1n16x5 FILLER_92_513 ();
 b15zdnd00an1n01x5 FILLER_92_529 ();
 b15zdnd11an1n04x5 FILLER_92_537 ();
 b15zdnd11an1n16x5 FILLER_92_553 ();
 b15zdnd00an1n02x5 FILLER_92_569 ();
 b15zdnd11an1n32x5 FILLER_92_576 ();
 b15zdnd00an1n02x5 FILLER_92_608 ();
 b15zdnd11an1n04x5 FILLER_92_616 ();
 b15zdnd11an1n64x5 FILLER_92_626 ();
 b15zdnd11an1n16x5 FILLER_92_690 ();
 b15zdnd11an1n08x5 FILLER_92_706 ();
 b15zdnd11an1n04x5 FILLER_92_714 ();
 b15zdnd11an1n08x5 FILLER_92_726 ();
 b15zdnd11an1n04x5 FILLER_92_734 ();
 b15zdnd00an1n02x5 FILLER_92_738 ();
 b15zdnd00an1n01x5 FILLER_92_740 ();
 b15zdnd11an1n16x5 FILLER_92_746 ();
 b15zdnd11an1n32x5 FILLER_92_769 ();
 b15zdnd11an1n16x5 FILLER_92_801 ();
 b15zdnd11an1n04x5 FILLER_92_817 ();
 b15zdnd11an1n32x5 FILLER_92_833 ();
 b15zdnd11an1n16x5 FILLER_92_865 ();
 b15zdnd11an1n08x5 FILLER_92_881 ();
 b15zdnd11an1n04x5 FILLER_92_901 ();
 b15zdnd11an1n32x5 FILLER_92_912 ();
 b15zdnd11an1n16x5 FILLER_92_944 ();
 b15zdnd11an1n04x5 FILLER_92_960 ();
 b15zdnd00an1n01x5 FILLER_92_964 ();
 b15zdnd11an1n64x5 FILLER_92_968 ();
 b15zdnd00an1n01x5 FILLER_92_1032 ();
 b15zdnd11an1n64x5 FILLER_92_1037 ();
 b15zdnd11an1n64x5 FILLER_92_1101 ();
 b15zdnd11an1n04x5 FILLER_92_1165 ();
 b15zdnd00an1n02x5 FILLER_92_1169 ();
 b15zdnd11an1n16x5 FILLER_92_1176 ();
 b15zdnd11an1n32x5 FILLER_92_1212 ();
 b15zdnd11an1n16x5 FILLER_92_1244 ();
 b15zdnd11an1n08x5 FILLER_92_1260 ();
 b15zdnd11an1n04x5 FILLER_92_1268 ();
 b15zdnd00an1n02x5 FILLER_92_1272 ();
 b15zdnd11an1n64x5 FILLER_92_1279 ();
 b15zdnd11an1n64x5 FILLER_92_1343 ();
 b15zdnd11an1n64x5 FILLER_92_1407 ();
 b15zdnd11an1n64x5 FILLER_92_1471 ();
 b15zdnd11an1n32x5 FILLER_92_1535 ();
 b15zdnd11an1n16x5 FILLER_92_1567 ();
 b15zdnd11an1n08x5 FILLER_92_1583 ();
 b15zdnd00an1n01x5 FILLER_92_1591 ();
 b15zdnd11an1n04x5 FILLER_92_1597 ();
 b15zdnd11an1n64x5 FILLER_92_1610 ();
 b15zdnd11an1n32x5 FILLER_92_1700 ();
 b15zdnd11an1n08x5 FILLER_92_1732 ();
 b15zdnd11an1n04x5 FILLER_92_1740 ();
 b15zdnd00an1n02x5 FILLER_92_1744 ();
 b15zdnd11an1n04x5 FILLER_92_1751 ();
 b15zdnd00an1n01x5 FILLER_92_1755 ();
 b15zdnd11an1n04x5 FILLER_92_1761 ();
 b15zdnd00an1n02x5 FILLER_92_1765 ();
 b15zdnd11an1n16x5 FILLER_92_1772 ();
 b15zdnd11an1n08x5 FILLER_92_1788 ();
 b15zdnd11an1n32x5 FILLER_92_1803 ();
 b15zdnd11an1n16x5 FILLER_92_1835 ();
 b15zdnd00an1n02x5 FILLER_92_1851 ();
 b15zdnd00an1n01x5 FILLER_92_1853 ();
 b15zdnd11an1n16x5 FILLER_92_1859 ();
 b15zdnd11an1n08x5 FILLER_92_1875 ();
 b15zdnd11an1n04x5 FILLER_92_1883 ();
 b15zdnd00an1n02x5 FILLER_92_1887 ();
 b15zdnd00an1n01x5 FILLER_92_1889 ();
 b15zdnd11an1n32x5 FILLER_92_1897 ();
 b15zdnd11an1n08x5 FILLER_92_1929 ();
 b15zdnd00an1n01x5 FILLER_92_1937 ();
 b15zdnd11an1n64x5 FILLER_92_1944 ();
 b15zdnd11an1n16x5 FILLER_92_2008 ();
 b15zdnd00an1n02x5 FILLER_92_2024 ();
 b15zdnd00an1n01x5 FILLER_92_2026 ();
 b15zdnd11an1n32x5 FILLER_92_2031 ();
 b15zdnd11an1n16x5 FILLER_92_2063 ();
 b15zdnd11an1n04x5 FILLER_92_2079 ();
 b15zdnd11an1n08x5 FILLER_92_2088 ();
 b15zdnd00an1n02x5 FILLER_92_2096 ();
 b15zdnd11an1n04x5 FILLER_92_2103 ();
 b15zdnd00an1n01x5 FILLER_92_2107 ();
 b15zdnd11an1n32x5 FILLER_92_2112 ();
 b15zdnd11an1n08x5 FILLER_92_2144 ();
 b15zdnd00an1n02x5 FILLER_92_2152 ();
 b15zdnd11an1n16x5 FILLER_92_2162 ();
 b15zdnd11an1n04x5 FILLER_92_2178 ();
 b15zdnd00an1n02x5 FILLER_92_2182 ();
 b15zdnd00an1n01x5 FILLER_92_2184 ();
 b15zdnd11an1n04x5 FILLER_92_2206 ();
 b15zdnd11an1n32x5 FILLER_92_2229 ();
 b15zdnd11an1n08x5 FILLER_92_2261 ();
 b15zdnd11an1n04x5 FILLER_92_2269 ();
 b15zdnd00an1n02x5 FILLER_92_2273 ();
 b15zdnd00an1n01x5 FILLER_92_2275 ();
 b15zdnd11an1n32x5 FILLER_93_0 ();
 b15zdnd11an1n08x5 FILLER_93_32 ();
 b15zdnd00an1n02x5 FILLER_93_40 ();
 b15zdnd11an1n64x5 FILLER_93_54 ();
 b15zdnd11an1n64x5 FILLER_93_118 ();
 b15zdnd11an1n64x5 FILLER_93_182 ();
 b15zdnd11an1n32x5 FILLER_93_246 ();
 b15zdnd00an1n02x5 FILLER_93_278 ();
 b15zdnd11an1n16x5 FILLER_93_284 ();
 b15zdnd11an1n08x5 FILLER_93_300 ();
 b15zdnd11an1n08x5 FILLER_93_324 ();
 b15zdnd11an1n04x5 FILLER_93_332 ();
 b15zdnd00an1n02x5 FILLER_93_336 ();
 b15zdnd11an1n04x5 FILLER_93_358 ();
 b15zdnd11an1n32x5 FILLER_93_369 ();
 b15zdnd11an1n16x5 FILLER_93_401 ();
 b15zdnd11an1n08x5 FILLER_93_417 ();
 b15zdnd11an1n04x5 FILLER_93_425 ();
 b15zdnd00an1n02x5 FILLER_93_429 ();
 b15zdnd11an1n64x5 FILLER_93_446 ();
 b15zdnd11an1n16x5 FILLER_93_510 ();
 b15zdnd11an1n04x5 FILLER_93_526 ();
 b15zdnd11an1n16x5 FILLER_93_536 ();
 b15zdnd11an1n04x5 FILLER_93_552 ();
 b15zdnd00an1n02x5 FILLER_93_556 ();
 b15zdnd11an1n08x5 FILLER_93_565 ();
 b15zdnd00an1n02x5 FILLER_93_573 ();
 b15zdnd11an1n04x5 FILLER_93_580 ();
 b15zdnd11an1n04x5 FILLER_93_597 ();
 b15zdnd11an1n04x5 FILLER_93_610 ();
 b15zdnd11an1n16x5 FILLER_93_625 ();
 b15zdnd11an1n08x5 FILLER_93_641 ();
 b15zdnd00an1n02x5 FILLER_93_649 ();
 b15zdnd00an1n01x5 FILLER_93_651 ();
 b15zdnd11an1n16x5 FILLER_93_657 ();
 b15zdnd11an1n04x5 FILLER_93_673 ();
 b15zdnd00an1n01x5 FILLER_93_677 ();
 b15zdnd11an1n08x5 FILLER_93_683 ();
 b15zdnd00an1n02x5 FILLER_93_691 ();
 b15zdnd00an1n01x5 FILLER_93_693 ();
 b15zdnd11an1n04x5 FILLER_93_704 ();
 b15zdnd11an1n04x5 FILLER_93_716 ();
 b15zdnd11an1n04x5 FILLER_93_727 ();
 b15zdnd00an1n02x5 FILLER_93_731 ();
 b15zdnd00an1n01x5 FILLER_93_733 ();
 b15zdnd11an1n64x5 FILLER_93_744 ();
 b15zdnd11an1n08x5 FILLER_93_808 ();
 b15zdnd11an1n04x5 FILLER_93_816 ();
 b15zdnd00an1n01x5 FILLER_93_820 ();
 b15zdnd11an1n64x5 FILLER_93_827 ();
 b15zdnd11an1n04x5 FILLER_93_891 ();
 b15zdnd00an1n02x5 FILLER_93_895 ();
 b15zdnd00an1n01x5 FILLER_93_897 ();
 b15zdnd11an1n64x5 FILLER_93_908 ();
 b15zdnd11an1n64x5 FILLER_93_972 ();
 b15zdnd11an1n04x5 FILLER_93_1036 ();
 b15zdnd00an1n02x5 FILLER_93_1040 ();
 b15zdnd11an1n16x5 FILLER_93_1046 ();
 b15zdnd11an1n04x5 FILLER_93_1062 ();
 b15zdnd00an1n02x5 FILLER_93_1066 ();
 b15zdnd00an1n01x5 FILLER_93_1068 ();
 b15zdnd11an1n32x5 FILLER_93_1100 ();
 b15zdnd11an1n08x5 FILLER_93_1132 ();
 b15zdnd11an1n04x5 FILLER_93_1140 ();
 b15zdnd00an1n02x5 FILLER_93_1144 ();
 b15zdnd00an1n01x5 FILLER_93_1146 ();
 b15zdnd11an1n64x5 FILLER_93_1151 ();
 b15zdnd11an1n16x5 FILLER_93_1215 ();
 b15zdnd11an1n64x5 FILLER_93_1262 ();
 b15zdnd11an1n04x5 FILLER_93_1326 ();
 b15zdnd00an1n01x5 FILLER_93_1330 ();
 b15zdnd11an1n64x5 FILLER_93_1336 ();
 b15zdnd11an1n32x5 FILLER_93_1400 ();
 b15zdnd11an1n08x5 FILLER_93_1432 ();
 b15zdnd00an1n02x5 FILLER_93_1440 ();
 b15zdnd11an1n64x5 FILLER_93_1447 ();
 b15zdnd11an1n64x5 FILLER_93_1511 ();
 b15zdnd11an1n16x5 FILLER_93_1575 ();
 b15zdnd11an1n08x5 FILLER_93_1591 ();
 b15zdnd00an1n02x5 FILLER_93_1599 ();
 b15zdnd00an1n01x5 FILLER_93_1601 ();
 b15zdnd11an1n64x5 FILLER_93_1622 ();
 b15zdnd11an1n64x5 FILLER_93_1686 ();
 b15zdnd11an1n64x5 FILLER_93_1750 ();
 b15zdnd11an1n16x5 FILLER_93_1814 ();
 b15zdnd11an1n04x5 FILLER_93_1830 ();
 b15zdnd00an1n02x5 FILLER_93_1834 ();
 b15zdnd11an1n16x5 FILLER_93_1841 ();
 b15zdnd11an1n04x5 FILLER_93_1857 ();
 b15zdnd00an1n01x5 FILLER_93_1861 ();
 b15zdnd11an1n16x5 FILLER_93_1868 ();
 b15zdnd11an1n04x5 FILLER_93_1884 ();
 b15zdnd11an1n08x5 FILLER_93_1903 ();
 b15zdnd00an1n02x5 FILLER_93_1911 ();
 b15zdnd11an1n04x5 FILLER_93_1934 ();
 b15zdnd00an1n01x5 FILLER_93_1938 ();
 b15zdnd11an1n64x5 FILLER_93_1952 ();
 b15zdnd11an1n08x5 FILLER_93_2016 ();
 b15zdnd00an1n01x5 FILLER_93_2024 ();
 b15zdnd11an1n32x5 FILLER_93_2035 ();
 b15zdnd11an1n08x5 FILLER_93_2067 ();
 b15zdnd11an1n04x5 FILLER_93_2075 ();
 b15zdnd11an1n04x5 FILLER_93_2085 ();
 b15zdnd11an1n04x5 FILLER_93_2099 ();
 b15zdnd11an1n16x5 FILLER_93_2121 ();
 b15zdnd11an1n08x5 FILLER_93_2137 ();
 b15zdnd11an1n04x5 FILLER_93_2145 ();
 b15zdnd00an1n02x5 FILLER_93_2149 ();
 b15zdnd00an1n01x5 FILLER_93_2151 ();
 b15zdnd11an1n04x5 FILLER_93_2164 ();
 b15zdnd00an1n02x5 FILLER_93_2168 ();
 b15zdnd00an1n01x5 FILLER_93_2170 ();
 b15zdnd11an1n04x5 FILLER_93_2178 ();
 b15zdnd00an1n02x5 FILLER_93_2182 ();
 b15zdnd11an1n08x5 FILLER_93_2194 ();
 b15zdnd00an1n02x5 FILLER_93_2202 ();
 b15zdnd00an1n01x5 FILLER_93_2204 ();
 b15zdnd11an1n64x5 FILLER_93_2214 ();
 b15zdnd11an1n04x5 FILLER_93_2278 ();
 b15zdnd00an1n02x5 FILLER_93_2282 ();
 b15zdnd11an1n64x5 FILLER_94_8 ();
 b15zdnd11an1n64x5 FILLER_94_72 ();
 b15zdnd11an1n08x5 FILLER_94_136 ();
 b15zdnd11an1n04x5 FILLER_94_144 ();
 b15zdnd00an1n01x5 FILLER_94_148 ();
 b15zdnd11an1n04x5 FILLER_94_155 ();
 b15zdnd11an1n32x5 FILLER_94_165 ();
 b15zdnd11an1n16x5 FILLER_94_197 ();
 b15zdnd11an1n04x5 FILLER_94_213 ();
 b15zdnd11an1n04x5 FILLER_94_221 ();
 b15zdnd00an1n02x5 FILLER_94_225 ();
 b15zdnd00an1n01x5 FILLER_94_227 ();
 b15zdnd11an1n08x5 FILLER_94_238 ();
 b15zdnd00an1n01x5 FILLER_94_246 ();
 b15zdnd11an1n16x5 FILLER_94_257 ();
 b15zdnd11an1n08x5 FILLER_94_273 ();
 b15zdnd00an1n02x5 FILLER_94_281 ();
 b15zdnd11an1n04x5 FILLER_94_292 ();
 b15zdnd11an1n08x5 FILLER_94_321 ();
 b15zdnd11an1n04x5 FILLER_94_329 ();
 b15zdnd00an1n02x5 FILLER_94_333 ();
 b15zdnd00an1n01x5 FILLER_94_335 ();
 b15zdnd11an1n04x5 FILLER_94_350 ();
 b15zdnd00an1n01x5 FILLER_94_354 ();
 b15zdnd11an1n08x5 FILLER_94_359 ();
 b15zdnd11an1n32x5 FILLER_94_381 ();
 b15zdnd11an1n16x5 FILLER_94_413 ();
 b15zdnd11an1n04x5 FILLER_94_429 ();
 b15zdnd00an1n01x5 FILLER_94_433 ();
 b15zdnd11an1n04x5 FILLER_94_447 ();
 b15zdnd11an1n08x5 FILLER_94_467 ();
 b15zdnd00an1n02x5 FILLER_94_475 ();
 b15zdnd11an1n08x5 FILLER_94_491 ();
 b15zdnd00an1n02x5 FILLER_94_499 ();
 b15zdnd11an1n32x5 FILLER_94_527 ();
 b15zdnd11an1n08x5 FILLER_94_559 ();
 b15zdnd11an1n04x5 FILLER_94_567 ();
 b15zdnd11an1n32x5 FILLER_94_579 ();
 b15zdnd00an1n01x5 FILLER_94_611 ();
 b15zdnd11an1n16x5 FILLER_94_616 ();
 b15zdnd11an1n08x5 FILLER_94_632 ();
 b15zdnd11an1n04x5 FILLER_94_640 ();
 b15zdnd00an1n02x5 FILLER_94_644 ();
 b15zdnd00an1n01x5 FILLER_94_646 ();
 b15zdnd11an1n16x5 FILLER_94_659 ();
 b15zdnd00an1n02x5 FILLER_94_675 ();
 b15zdnd11an1n16x5 FILLER_94_690 ();
 b15zdnd11an1n08x5 FILLER_94_706 ();
 b15zdnd11an1n04x5 FILLER_94_714 ();
 b15zdnd11an1n16x5 FILLER_94_726 ();
 b15zdnd11an1n04x5 FILLER_94_742 ();
 b15zdnd00an1n02x5 FILLER_94_746 ();
 b15zdnd00an1n01x5 FILLER_94_748 ();
 b15zdnd11an1n32x5 FILLER_94_761 ();
 b15zdnd00an1n02x5 FILLER_94_793 ();
 b15zdnd00an1n01x5 FILLER_94_795 ();
 b15zdnd11an1n64x5 FILLER_94_803 ();
 b15zdnd11an1n04x5 FILLER_94_867 ();
 b15zdnd00an1n01x5 FILLER_94_871 ();
 b15zdnd11an1n08x5 FILLER_94_885 ();
 b15zdnd00an1n02x5 FILLER_94_893 ();
 b15zdnd00an1n01x5 FILLER_94_895 ();
 b15zdnd11an1n64x5 FILLER_94_909 ();
 b15zdnd11an1n64x5 FILLER_94_973 ();
 b15zdnd11an1n16x5 FILLER_94_1037 ();
 b15zdnd00an1n01x5 FILLER_94_1053 ();
 b15zdnd11an1n64x5 FILLER_94_1065 ();
 b15zdnd11an1n64x5 FILLER_94_1129 ();
 b15zdnd11an1n08x5 FILLER_94_1193 ();
 b15zdnd00an1n02x5 FILLER_94_1201 ();
 b15zdnd00an1n01x5 FILLER_94_1203 ();
 b15zdnd11an1n64x5 FILLER_94_1222 ();
 b15zdnd11an1n32x5 FILLER_94_1286 ();
 b15zdnd11an1n04x5 FILLER_94_1318 ();
 b15zdnd00an1n02x5 FILLER_94_1322 ();
 b15zdnd11an1n04x5 FILLER_94_1329 ();
 b15zdnd11an1n04x5 FILLER_94_1338 ();
 b15zdnd00an1n01x5 FILLER_94_1342 ();
 b15zdnd11an1n16x5 FILLER_94_1351 ();
 b15zdnd11an1n32x5 FILLER_94_1371 ();
 b15zdnd11an1n16x5 FILLER_94_1403 ();
 b15zdnd11an1n08x5 FILLER_94_1419 ();
 b15zdnd00an1n02x5 FILLER_94_1427 ();
 b15zdnd00an1n01x5 FILLER_94_1429 ();
 b15zdnd11an1n04x5 FILLER_94_1436 ();
 b15zdnd11an1n16x5 FILLER_94_1445 ();
 b15zdnd00an1n02x5 FILLER_94_1461 ();
 b15zdnd00an1n01x5 FILLER_94_1463 ();
 b15zdnd11an1n04x5 FILLER_94_1496 ();
 b15zdnd00an1n02x5 FILLER_94_1500 ();
 b15zdnd11an1n16x5 FILLER_94_1510 ();
 b15zdnd11an1n08x5 FILLER_94_1526 ();
 b15zdnd11an1n16x5 FILLER_94_1539 ();
 b15zdnd11an1n04x5 FILLER_94_1555 ();
 b15zdnd00an1n02x5 FILLER_94_1559 ();
 b15zdnd11an1n32x5 FILLER_94_1587 ();
 b15zdnd00an1n02x5 FILLER_94_1619 ();
 b15zdnd00an1n01x5 FILLER_94_1621 ();
 b15zdnd11an1n04x5 FILLER_94_1648 ();
 b15zdnd11an1n04x5 FILLER_94_1672 ();
 b15zdnd00an1n01x5 FILLER_94_1676 ();
 b15zdnd11an1n64x5 FILLER_94_1703 ();
 b15zdnd11an1n04x5 FILLER_94_1767 ();
 b15zdnd00an1n01x5 FILLER_94_1771 ();
 b15zdnd11an1n04x5 FILLER_94_1779 ();
 b15zdnd00an1n01x5 FILLER_94_1783 ();
 b15zdnd11an1n04x5 FILLER_94_1806 ();
 b15zdnd11an1n04x5 FILLER_94_1820 ();
 b15zdnd00an1n02x5 FILLER_94_1824 ();
 b15zdnd11an1n16x5 FILLER_94_1830 ();
 b15zdnd11an1n08x5 FILLER_94_1846 ();
 b15zdnd00an1n01x5 FILLER_94_1854 ();
 b15zdnd11an1n04x5 FILLER_94_1865 ();
 b15zdnd00an1n02x5 FILLER_94_1869 ();
 b15zdnd11an1n04x5 FILLER_94_1887 ();
 b15zdnd11an1n64x5 FILLER_94_1897 ();
 b15zdnd11an1n16x5 FILLER_94_1961 ();
 b15zdnd11an1n64x5 FILLER_94_1983 ();
 b15zdnd11an1n32x5 FILLER_94_2047 ();
 b15zdnd11an1n64x5 FILLER_94_2085 ();
 b15zdnd11an1n04x5 FILLER_94_2149 ();
 b15zdnd00an1n01x5 FILLER_94_2153 ();
 b15zdnd11an1n32x5 FILLER_94_2162 ();
 b15zdnd11an1n08x5 FILLER_94_2194 ();
 b15zdnd11an1n04x5 FILLER_94_2202 ();
 b15zdnd00an1n02x5 FILLER_94_2206 ();
 b15zdnd11an1n64x5 FILLER_94_2212 ();
 b15zdnd11an1n64x5 FILLER_95_0 ();
 b15zdnd11an1n08x5 FILLER_95_64 ();
 b15zdnd11an1n04x5 FILLER_95_72 ();
 b15zdnd00an1n02x5 FILLER_95_76 ();
 b15zdnd11an1n04x5 FILLER_95_99 ();
 b15zdnd11an1n08x5 FILLER_95_111 ();
 b15zdnd11an1n04x5 FILLER_95_119 ();
 b15zdnd11an1n16x5 FILLER_95_128 ();
 b15zdnd00an1n02x5 FILLER_95_144 ();
 b15zdnd00an1n01x5 FILLER_95_146 ();
 b15zdnd11an1n16x5 FILLER_95_152 ();
 b15zdnd11an1n08x5 FILLER_95_168 ();
 b15zdnd11an1n04x5 FILLER_95_176 ();
 b15zdnd00an1n02x5 FILLER_95_180 ();
 b15zdnd00an1n01x5 FILLER_95_182 ();
 b15zdnd11an1n16x5 FILLER_95_189 ();
 b15zdnd11an1n08x5 FILLER_95_205 ();
 b15zdnd11an1n04x5 FILLER_95_213 ();
 b15zdnd00an1n02x5 FILLER_95_217 ();
 b15zdnd11an1n08x5 FILLER_95_235 ();
 b15zdnd00an1n02x5 FILLER_95_243 ();
 b15zdnd11an1n64x5 FILLER_95_260 ();
 b15zdnd11an1n04x5 FILLER_95_324 ();
 b15zdnd00an1n02x5 FILLER_95_328 ();
 b15zdnd00an1n01x5 FILLER_95_330 ();
 b15zdnd11an1n16x5 FILLER_95_357 ();
 b15zdnd11an1n04x5 FILLER_95_373 ();
 b15zdnd00an1n02x5 FILLER_95_377 ();
 b15zdnd00an1n01x5 FILLER_95_379 ();
 b15zdnd11an1n64x5 FILLER_95_389 ();
 b15zdnd11an1n32x5 FILLER_95_459 ();
 b15zdnd11an1n16x5 FILLER_95_491 ();
 b15zdnd11an1n04x5 FILLER_95_507 ();
 b15zdnd00an1n02x5 FILLER_95_511 ();
 b15zdnd11an1n04x5 FILLER_95_533 ();
 b15zdnd11an1n64x5 FILLER_95_542 ();
 b15zdnd11an1n08x5 FILLER_95_606 ();
 b15zdnd11an1n08x5 FILLER_95_627 ();
 b15zdnd11an1n04x5 FILLER_95_635 ();
 b15zdnd00an1n02x5 FILLER_95_639 ();
 b15zdnd00an1n01x5 FILLER_95_641 ();
 b15zdnd11an1n64x5 FILLER_95_646 ();
 b15zdnd11an1n16x5 FILLER_95_710 ();
 b15zdnd11an1n32x5 FILLER_95_746 ();
 b15zdnd11an1n04x5 FILLER_95_778 ();
 b15zdnd00an1n01x5 FILLER_95_782 ();
 b15zdnd11an1n64x5 FILLER_95_798 ();
 b15zdnd11an1n16x5 FILLER_95_862 ();
 b15zdnd00an1n02x5 FILLER_95_878 ();
 b15zdnd11an1n64x5 FILLER_95_896 ();
 b15zdnd11an1n64x5 FILLER_95_960 ();
 b15zdnd11an1n32x5 FILLER_95_1024 ();
 b15zdnd11an1n16x5 FILLER_95_1076 ();
 b15zdnd11an1n08x5 FILLER_95_1092 ();
 b15zdnd11an1n04x5 FILLER_95_1120 ();
 b15zdnd11an1n32x5 FILLER_95_1129 ();
 b15zdnd11an1n16x5 FILLER_95_1161 ();
 b15zdnd11an1n04x5 FILLER_95_1177 ();
 b15zdnd00an1n02x5 FILLER_95_1181 ();
 b15zdnd11an1n64x5 FILLER_95_1214 ();
 b15zdnd11an1n32x5 FILLER_95_1278 ();
 b15zdnd11an1n16x5 FILLER_95_1310 ();
 b15zdnd11an1n04x5 FILLER_95_1326 ();
 b15zdnd00an1n02x5 FILLER_95_1330 ();
 b15zdnd11an1n04x5 FILLER_95_1338 ();
 b15zdnd00an1n02x5 FILLER_95_1342 ();
 b15zdnd00an1n01x5 FILLER_95_1344 ();
 b15zdnd11an1n08x5 FILLER_95_1349 ();
 b15zdnd11an1n04x5 FILLER_95_1357 ();
 b15zdnd00an1n01x5 FILLER_95_1361 ();
 b15zdnd11an1n32x5 FILLER_95_1375 ();
 b15zdnd11an1n16x5 FILLER_95_1407 ();
 b15zdnd11an1n04x5 FILLER_95_1423 ();
 b15zdnd00an1n02x5 FILLER_95_1427 ();
 b15zdnd00an1n01x5 FILLER_95_1429 ();
 b15zdnd11an1n16x5 FILLER_95_1444 ();
 b15zdnd11an1n04x5 FILLER_95_1460 ();
 b15zdnd11an1n16x5 FILLER_95_1469 ();
 b15zdnd11an1n08x5 FILLER_95_1485 ();
 b15zdnd00an1n02x5 FILLER_95_1493 ();
 b15zdnd00an1n01x5 FILLER_95_1495 ();
 b15zdnd11an1n04x5 FILLER_95_1527 ();
 b15zdnd00an1n02x5 FILLER_95_1531 ();
 b15zdnd11an1n32x5 FILLER_95_1545 ();
 b15zdnd11an1n16x5 FILLER_95_1577 ();
 b15zdnd11an1n08x5 FILLER_95_1593 ();
 b15zdnd11an1n04x5 FILLER_95_1601 ();
 b15zdnd11an1n16x5 FILLER_95_1630 ();
 b15zdnd11an1n04x5 FILLER_95_1646 ();
 b15zdnd11an1n16x5 FILLER_95_1659 ();
 b15zdnd11an1n08x5 FILLER_95_1675 ();
 b15zdnd11an1n04x5 FILLER_95_1683 ();
 b15zdnd00an1n02x5 FILLER_95_1687 ();
 b15zdnd00an1n01x5 FILLER_95_1689 ();
 b15zdnd11an1n32x5 FILLER_95_1701 ();
 b15zdnd11an1n04x5 FILLER_95_1733 ();
 b15zdnd00an1n01x5 FILLER_95_1737 ();
 b15zdnd11an1n16x5 FILLER_95_1750 ();
 b15zdnd11an1n08x5 FILLER_95_1766 ();
 b15zdnd00an1n02x5 FILLER_95_1774 ();
 b15zdnd00an1n01x5 FILLER_95_1776 ();
 b15zdnd11an1n08x5 FILLER_95_1781 ();
 b15zdnd11an1n04x5 FILLER_95_1789 ();
 b15zdnd00an1n02x5 FILLER_95_1793 ();
 b15zdnd11an1n64x5 FILLER_95_1801 ();
 b15zdnd00an1n02x5 FILLER_95_1865 ();
 b15zdnd00an1n01x5 FILLER_95_1867 ();
 b15zdnd11an1n16x5 FILLER_95_1872 ();
 b15zdnd11an1n08x5 FILLER_95_1888 ();
 b15zdnd11an1n04x5 FILLER_95_1896 ();
 b15zdnd11an1n16x5 FILLER_95_1905 ();
 b15zdnd11an1n04x5 FILLER_95_1921 ();
 b15zdnd11an1n32x5 FILLER_95_1933 ();
 b15zdnd00an1n02x5 FILLER_95_1965 ();
 b15zdnd00an1n01x5 FILLER_95_1967 ();
 b15zdnd11an1n04x5 FILLER_95_1973 ();
 b15zdnd11an1n32x5 FILLER_95_1986 ();
 b15zdnd11an1n08x5 FILLER_95_2018 ();
 b15zdnd00an1n02x5 FILLER_95_2026 ();
 b15zdnd11an1n32x5 FILLER_95_2032 ();
 b15zdnd11an1n08x5 FILLER_95_2064 ();
 b15zdnd11an1n04x5 FILLER_95_2072 ();
 b15zdnd00an1n01x5 FILLER_95_2076 ();
 b15zdnd11an1n16x5 FILLER_95_2083 ();
 b15zdnd00an1n02x5 FILLER_95_2099 ();
 b15zdnd11an1n16x5 FILLER_95_2107 ();
 b15zdnd00an1n02x5 FILLER_95_2123 ();
 b15zdnd11an1n04x5 FILLER_95_2130 ();
 b15zdnd11an1n64x5 FILLER_95_2142 ();
 b15zdnd11an1n64x5 FILLER_95_2206 ();
 b15zdnd11an1n08x5 FILLER_95_2270 ();
 b15zdnd00an1n02x5 FILLER_95_2282 ();
 b15zdnd11an1n64x5 FILLER_96_8 ();
 b15zdnd11an1n32x5 FILLER_96_72 ();
 b15zdnd11an1n04x5 FILLER_96_104 ();
 b15zdnd00an1n02x5 FILLER_96_108 ();
 b15zdnd11an1n04x5 FILLER_96_116 ();
 b15zdnd11an1n16x5 FILLER_96_136 ();
 b15zdnd11an1n08x5 FILLER_96_152 ();
 b15zdnd00an1n02x5 FILLER_96_160 ();
 b15zdnd00an1n01x5 FILLER_96_162 ();
 b15zdnd11an1n32x5 FILLER_96_175 ();
 b15zdnd11an1n08x5 FILLER_96_211 ();
 b15zdnd11an1n16x5 FILLER_96_228 ();
 b15zdnd11an1n08x5 FILLER_96_244 ();
 b15zdnd11an1n04x5 FILLER_96_252 ();
 b15zdnd00an1n01x5 FILLER_96_256 ();
 b15zdnd11an1n04x5 FILLER_96_261 ();
 b15zdnd00an1n02x5 FILLER_96_265 ();
 b15zdnd00an1n01x5 FILLER_96_267 ();
 b15zdnd11an1n16x5 FILLER_96_282 ();
 b15zdnd11an1n16x5 FILLER_96_314 ();
 b15zdnd11an1n04x5 FILLER_96_335 ();
 b15zdnd00an1n02x5 FILLER_96_339 ();
 b15zdnd00an1n01x5 FILLER_96_341 ();
 b15zdnd11an1n64x5 FILLER_96_352 ();
 b15zdnd11an1n64x5 FILLER_96_416 ();
 b15zdnd11an1n32x5 FILLER_96_480 ();
 b15zdnd11an1n16x5 FILLER_96_512 ();
 b15zdnd00an1n02x5 FILLER_96_528 ();
 b15zdnd00an1n01x5 FILLER_96_530 ();
 b15zdnd11an1n04x5 FILLER_96_543 ();
 b15zdnd00an1n02x5 FILLER_96_547 ();
 b15zdnd00an1n01x5 FILLER_96_549 ();
 b15zdnd11an1n64x5 FILLER_96_554 ();
 b15zdnd11an1n16x5 FILLER_96_618 ();
 b15zdnd11an1n04x5 FILLER_96_634 ();
 b15zdnd00an1n02x5 FILLER_96_638 ();
 b15zdnd11an1n04x5 FILLER_96_649 ();
 b15zdnd11an1n32x5 FILLER_96_662 ();
 b15zdnd11an1n16x5 FILLER_96_694 ();
 b15zdnd11an1n08x5 FILLER_96_710 ();
 b15zdnd11an1n32x5 FILLER_96_726 ();
 b15zdnd11an1n08x5 FILLER_96_758 ();
 b15zdnd00an1n02x5 FILLER_96_766 ();
 b15zdnd00an1n01x5 FILLER_96_768 ();
 b15zdnd11an1n04x5 FILLER_96_781 ();
 b15zdnd11an1n64x5 FILLER_96_798 ();
 b15zdnd00an1n01x5 FILLER_96_862 ();
 b15zdnd11an1n16x5 FILLER_96_875 ();
 b15zdnd11an1n04x5 FILLER_96_891 ();
 b15zdnd00an1n02x5 FILLER_96_895 ();
 b15zdnd11an1n04x5 FILLER_96_902 ();
 b15zdnd11an1n08x5 FILLER_96_912 ();
 b15zdnd11an1n04x5 FILLER_96_920 ();
 b15zdnd00an1n01x5 FILLER_96_924 ();
 b15zdnd11an1n32x5 FILLER_96_930 ();
 b15zdnd11an1n08x5 FILLER_96_962 ();
 b15zdnd00an1n01x5 FILLER_96_970 ();
 b15zdnd11an1n32x5 FILLER_96_975 ();
 b15zdnd11an1n08x5 FILLER_96_1007 ();
 b15zdnd00an1n02x5 FILLER_96_1015 ();
 b15zdnd11an1n04x5 FILLER_96_1037 ();
 b15zdnd11an1n32x5 FILLER_96_1046 ();
 b15zdnd11an1n16x5 FILLER_96_1078 ();
 b15zdnd00an1n02x5 FILLER_96_1094 ();
 b15zdnd00an1n01x5 FILLER_96_1096 ();
 b15zdnd11an1n16x5 FILLER_96_1128 ();
 b15zdnd00an1n01x5 FILLER_96_1144 ();
 b15zdnd11an1n64x5 FILLER_96_1176 ();
 b15zdnd11an1n32x5 FILLER_96_1240 ();
 b15zdnd11an1n32x5 FILLER_96_1278 ();
 b15zdnd11an1n08x5 FILLER_96_1310 ();
 b15zdnd00an1n02x5 FILLER_96_1318 ();
 b15zdnd11an1n16x5 FILLER_96_1326 ();
 b15zdnd11an1n08x5 FILLER_96_1342 ();
 b15zdnd11an1n04x5 FILLER_96_1350 ();
 b15zdnd11an1n04x5 FILLER_96_1361 ();
 b15zdnd11an1n32x5 FILLER_96_1374 ();
 b15zdnd00an1n02x5 FILLER_96_1406 ();
 b15zdnd00an1n01x5 FILLER_96_1408 ();
 b15zdnd11an1n04x5 FILLER_96_1416 ();
 b15zdnd11an1n08x5 FILLER_96_1426 ();
 b15zdnd11an1n16x5 FILLER_96_1444 ();
 b15zdnd11an1n04x5 FILLER_96_1460 ();
 b15zdnd00an1n02x5 FILLER_96_1464 ();
 b15zdnd11an1n08x5 FILLER_96_1473 ();
 b15zdnd11an1n04x5 FILLER_96_1481 ();
 b15zdnd00an1n02x5 FILLER_96_1485 ();
 b15zdnd00an1n01x5 FILLER_96_1487 ();
 b15zdnd11an1n64x5 FILLER_96_1493 ();
 b15zdnd11an1n64x5 FILLER_96_1557 ();
 b15zdnd11an1n64x5 FILLER_96_1621 ();
 b15zdnd11an1n64x5 FILLER_96_1685 ();
 b15zdnd11an1n64x5 FILLER_96_1749 ();
 b15zdnd00an1n02x5 FILLER_96_1813 ();
 b15zdnd00an1n01x5 FILLER_96_1815 ();
 b15zdnd11an1n32x5 FILLER_96_1830 ();
 b15zdnd11an1n08x5 FILLER_96_1862 ();
 b15zdnd11an1n04x5 FILLER_96_1870 ();
 b15zdnd11an1n16x5 FILLER_96_1883 ();
 b15zdnd00an1n02x5 FILLER_96_1899 ();
 b15zdnd00an1n01x5 FILLER_96_1901 ();
 b15zdnd11an1n64x5 FILLER_96_1912 ();
 b15zdnd11an1n16x5 FILLER_96_1976 ();
 b15zdnd11an1n08x5 FILLER_96_1992 ();
 b15zdnd00an1n02x5 FILLER_96_2000 ();
 b15zdnd11an1n04x5 FILLER_96_2012 ();
 b15zdnd11an1n16x5 FILLER_96_2023 ();
 b15zdnd11an1n08x5 FILLER_96_2039 ();
 b15zdnd11an1n16x5 FILLER_96_2053 ();
 b15zdnd11an1n08x5 FILLER_96_2069 ();
 b15zdnd11an1n04x5 FILLER_96_2077 ();
 b15zdnd00an1n02x5 FILLER_96_2081 ();
 b15zdnd00an1n01x5 FILLER_96_2083 ();
 b15zdnd11an1n08x5 FILLER_96_2100 ();
 b15zdnd00an1n02x5 FILLER_96_2108 ();
 b15zdnd11an1n32x5 FILLER_96_2116 ();
 b15zdnd11an1n04x5 FILLER_96_2148 ();
 b15zdnd00an1n02x5 FILLER_96_2152 ();
 b15zdnd11an1n64x5 FILLER_96_2162 ();
 b15zdnd11an1n16x5 FILLER_96_2226 ();
 b15zdnd11an1n08x5 FILLER_96_2242 ();
 b15zdnd11an1n04x5 FILLER_96_2250 ();
 b15zdnd00an1n02x5 FILLER_96_2274 ();
 b15zdnd11an1n32x5 FILLER_97_0 ();
 b15zdnd11an1n16x5 FILLER_97_32 ();
 b15zdnd11an1n04x5 FILLER_97_48 ();
 b15zdnd11an1n32x5 FILLER_97_68 ();
 b15zdnd00an1n02x5 FILLER_97_100 ();
 b15zdnd11an1n04x5 FILLER_97_110 ();
 b15zdnd11an1n64x5 FILLER_97_126 ();
 b15zdnd11an1n32x5 FILLER_97_190 ();
 b15zdnd11an1n16x5 FILLER_97_222 ();
 b15zdnd11an1n08x5 FILLER_97_238 ();
 b15zdnd11an1n04x5 FILLER_97_260 ();
 b15zdnd00an1n02x5 FILLER_97_264 ();
 b15zdnd00an1n01x5 FILLER_97_266 ();
 b15zdnd11an1n32x5 FILLER_97_287 ();
 b15zdnd11an1n08x5 FILLER_97_319 ();
 b15zdnd00an1n02x5 FILLER_97_327 ();
 b15zdnd11an1n04x5 FILLER_97_338 ();
 b15zdnd11an1n04x5 FILLER_97_350 ();
 b15zdnd00an1n01x5 FILLER_97_354 ();
 b15zdnd11an1n32x5 FILLER_97_373 ();
 b15zdnd11an1n16x5 FILLER_97_405 ();
 b15zdnd11an1n04x5 FILLER_97_421 ();
 b15zdnd00an1n02x5 FILLER_97_425 ();
 b15zdnd00an1n01x5 FILLER_97_427 ();
 b15zdnd11an1n64x5 FILLER_97_440 ();
 b15zdnd11an1n08x5 FILLER_97_504 ();
 b15zdnd11an1n08x5 FILLER_97_521 ();
 b15zdnd00an1n02x5 FILLER_97_529 ();
 b15zdnd11an1n64x5 FILLER_97_536 ();
 b15zdnd11an1n64x5 FILLER_97_612 ();
 b15zdnd11an1n08x5 FILLER_97_676 ();
 b15zdnd11an1n04x5 FILLER_97_684 ();
 b15zdnd00an1n01x5 FILLER_97_688 ();
 b15zdnd11an1n04x5 FILLER_97_701 ();
 b15zdnd11an1n64x5 FILLER_97_709 ();
 b15zdnd11an1n08x5 FILLER_97_773 ();
 b15zdnd00an1n02x5 FILLER_97_781 ();
 b15zdnd11an1n16x5 FILLER_97_792 ();
 b15zdnd00an1n02x5 FILLER_97_808 ();
 b15zdnd11an1n08x5 FILLER_97_831 ();
 b15zdnd00an1n01x5 FILLER_97_839 ();
 b15zdnd11an1n16x5 FILLER_97_846 ();
 b15zdnd11an1n04x5 FILLER_97_862 ();
 b15zdnd00an1n01x5 FILLER_97_866 ();
 b15zdnd11an1n04x5 FILLER_97_871 ();
 b15zdnd00an1n02x5 FILLER_97_875 ();
 b15zdnd11an1n32x5 FILLER_97_884 ();
 b15zdnd11an1n32x5 FILLER_97_926 ();
 b15zdnd11an1n08x5 FILLER_97_958 ();
 b15zdnd11an1n04x5 FILLER_97_966 ();
 b15zdnd00an1n01x5 FILLER_97_970 ();
 b15zdnd11an1n16x5 FILLER_97_991 ();
 b15zdnd00an1n02x5 FILLER_97_1007 ();
 b15zdnd00an1n01x5 FILLER_97_1009 ();
 b15zdnd11an1n08x5 FILLER_97_1027 ();
 b15zdnd11an1n32x5 FILLER_97_1038 ();
 b15zdnd11an1n16x5 FILLER_97_1070 ();
 b15zdnd11an1n08x5 FILLER_97_1086 ();
 b15zdnd11an1n04x5 FILLER_97_1094 ();
 b15zdnd00an1n02x5 FILLER_97_1098 ();
 b15zdnd00an1n01x5 FILLER_97_1100 ();
 b15zdnd11an1n04x5 FILLER_97_1132 ();
 b15zdnd11an1n64x5 FILLER_97_1147 ();
 b15zdnd11an1n08x5 FILLER_97_1211 ();
 b15zdnd11an1n08x5 FILLER_97_1237 ();
 b15zdnd00an1n02x5 FILLER_97_1245 ();
 b15zdnd11an1n16x5 FILLER_97_1256 ();
 b15zdnd00an1n01x5 FILLER_97_1272 ();
 b15zdnd11an1n16x5 FILLER_97_1281 ();
 b15zdnd11an1n08x5 FILLER_97_1297 ();
 b15zdnd11an1n04x5 FILLER_97_1305 ();
 b15zdnd00an1n01x5 FILLER_97_1309 ();
 b15zdnd11an1n64x5 FILLER_97_1315 ();
 b15zdnd11an1n16x5 FILLER_97_1379 ();
 b15zdnd11an1n08x5 FILLER_97_1395 ();
 b15zdnd11an1n04x5 FILLER_97_1403 ();
 b15zdnd11an1n04x5 FILLER_97_1414 ();
 b15zdnd11an1n16x5 FILLER_97_1423 ();
 b15zdnd00an1n02x5 FILLER_97_1439 ();
 b15zdnd11an1n16x5 FILLER_97_1445 ();
 b15zdnd11an1n08x5 FILLER_97_1461 ();
 b15zdnd11an1n16x5 FILLER_97_1476 ();
 b15zdnd11an1n04x5 FILLER_97_1492 ();
 b15zdnd11an1n04x5 FILLER_97_1505 ();
 b15zdnd00an1n02x5 FILLER_97_1509 ();
 b15zdnd00an1n01x5 FILLER_97_1511 ();
 b15zdnd11an1n16x5 FILLER_97_1516 ();
 b15zdnd11an1n32x5 FILLER_97_1542 ();
 b15zdnd00an1n02x5 FILLER_97_1574 ();
 b15zdnd11an1n16x5 FILLER_97_1590 ();
 b15zdnd11an1n04x5 FILLER_97_1606 ();
 b15zdnd00an1n01x5 FILLER_97_1610 ();
 b15zdnd11an1n32x5 FILLER_97_1627 ();
 b15zdnd11an1n16x5 FILLER_97_1659 ();
 b15zdnd00an1n02x5 FILLER_97_1675 ();
 b15zdnd00an1n01x5 FILLER_97_1677 ();
 b15zdnd11an1n32x5 FILLER_97_1698 ();
 b15zdnd11an1n08x5 FILLER_97_1730 ();
 b15zdnd11an1n04x5 FILLER_97_1738 ();
 b15zdnd00an1n01x5 FILLER_97_1742 ();
 b15zdnd11an1n64x5 FILLER_97_1775 ();
 b15zdnd11an1n32x5 FILLER_97_1839 ();
 b15zdnd11an1n16x5 FILLER_97_1871 ();
 b15zdnd11an1n08x5 FILLER_97_1887 ();
 b15zdnd00an1n01x5 FILLER_97_1895 ();
 b15zdnd11an1n04x5 FILLER_97_1906 ();
 b15zdnd00an1n01x5 FILLER_97_1910 ();
 b15zdnd11an1n04x5 FILLER_97_1915 ();
 b15zdnd00an1n02x5 FILLER_97_1919 ();
 b15zdnd11an1n64x5 FILLER_97_1926 ();
 b15zdnd11an1n04x5 FILLER_97_1990 ();
 b15zdnd00an1n02x5 FILLER_97_1994 ();
 b15zdnd00an1n01x5 FILLER_97_1996 ();
 b15zdnd11an1n32x5 FILLER_97_2011 ();
 b15zdnd00an1n01x5 FILLER_97_2043 ();
 b15zdnd11an1n04x5 FILLER_97_2049 ();
 b15zdnd11an1n32x5 FILLER_97_2057 ();
 b15zdnd11an1n08x5 FILLER_97_2089 ();
 b15zdnd00an1n02x5 FILLER_97_2097 ();
 b15zdnd11an1n16x5 FILLER_97_2130 ();
 b15zdnd11an1n04x5 FILLER_97_2146 ();
 b15zdnd11an1n04x5 FILLER_97_2155 ();
 b15zdnd11an1n04x5 FILLER_97_2169 ();
 b15zdnd00an1n02x5 FILLER_97_2173 ();
 b15zdnd11an1n64x5 FILLER_97_2185 ();
 b15zdnd11an1n32x5 FILLER_97_2249 ();
 b15zdnd00an1n02x5 FILLER_97_2281 ();
 b15zdnd00an1n01x5 FILLER_97_2283 ();
 b15zdnd11an1n64x5 FILLER_98_8 ();
 b15zdnd11an1n16x5 FILLER_98_72 ();
 b15zdnd11an1n08x5 FILLER_98_88 ();
 b15zdnd00an1n02x5 FILLER_98_96 ();
 b15zdnd11an1n32x5 FILLER_98_107 ();
 b15zdnd11an1n08x5 FILLER_98_139 ();
 b15zdnd00an1n02x5 FILLER_98_147 ();
 b15zdnd00an1n01x5 FILLER_98_149 ();
 b15zdnd11an1n32x5 FILLER_98_157 ();
 b15zdnd00an1n02x5 FILLER_98_189 ();
 b15zdnd00an1n01x5 FILLER_98_191 ();
 b15zdnd11an1n16x5 FILLER_98_197 ();
 b15zdnd11an1n08x5 FILLER_98_213 ();
 b15zdnd11an1n04x5 FILLER_98_221 ();
 b15zdnd00an1n02x5 FILLER_98_225 ();
 b15zdnd00an1n01x5 FILLER_98_227 ();
 b15zdnd11an1n04x5 FILLER_98_240 ();
 b15zdnd11an1n08x5 FILLER_98_250 ();
 b15zdnd11an1n04x5 FILLER_98_258 ();
 b15zdnd11an1n32x5 FILLER_98_269 ();
 b15zdnd11an1n04x5 FILLER_98_301 ();
 b15zdnd00an1n02x5 FILLER_98_305 ();
 b15zdnd00an1n01x5 FILLER_98_307 ();
 b15zdnd11an1n04x5 FILLER_98_326 ();
 b15zdnd11an1n64x5 FILLER_98_346 ();
 b15zdnd11an1n16x5 FILLER_98_410 ();
 b15zdnd11an1n08x5 FILLER_98_426 ();
 b15zdnd00an1n02x5 FILLER_98_434 ();
 b15zdnd11an1n32x5 FILLER_98_440 ();
 b15zdnd11an1n04x5 FILLER_98_472 ();
 b15zdnd00an1n02x5 FILLER_98_476 ();
 b15zdnd11an1n08x5 FILLER_98_482 ();
 b15zdnd00an1n01x5 FILLER_98_490 ();
 b15zdnd11an1n08x5 FILLER_98_498 ();
 b15zdnd11an1n04x5 FILLER_98_506 ();
 b15zdnd00an1n01x5 FILLER_98_510 ();
 b15zdnd11an1n04x5 FILLER_98_523 ();
 b15zdnd11an1n16x5 FILLER_98_534 ();
 b15zdnd11an1n04x5 FILLER_98_550 ();
 b15zdnd00an1n02x5 FILLER_98_554 ();
 b15zdnd11an1n32x5 FILLER_98_566 ();
 b15zdnd11an1n08x5 FILLER_98_598 ();
 b15zdnd00an1n01x5 FILLER_98_606 ();
 b15zdnd11an1n32x5 FILLER_98_619 ();
 b15zdnd00an1n02x5 FILLER_98_651 ();
 b15zdnd00an1n01x5 FILLER_98_653 ();
 b15zdnd11an1n08x5 FILLER_98_660 ();
 b15zdnd11an1n04x5 FILLER_98_680 ();
 b15zdnd11an1n08x5 FILLER_98_710 ();
 b15zdnd00an1n02x5 FILLER_98_726 ();
 b15zdnd11an1n04x5 FILLER_98_740 ();
 b15zdnd11an1n32x5 FILLER_98_754 ();
 b15zdnd00an1n02x5 FILLER_98_786 ();
 b15zdnd00an1n01x5 FILLER_98_788 ();
 b15zdnd11an1n32x5 FILLER_98_793 ();
 b15zdnd11an1n08x5 FILLER_98_825 ();
 b15zdnd00an1n01x5 FILLER_98_833 ();
 b15zdnd11an1n32x5 FILLER_98_843 ();
 b15zdnd11an1n16x5 FILLER_98_875 ();
 b15zdnd11an1n08x5 FILLER_98_891 ();
 b15zdnd11an1n04x5 FILLER_98_899 ();
 b15zdnd00an1n01x5 FILLER_98_903 ();
 b15zdnd11an1n16x5 FILLER_98_925 ();
 b15zdnd00an1n01x5 FILLER_98_941 ();
 b15zdnd11an1n16x5 FILLER_98_954 ();
 b15zdnd11an1n08x5 FILLER_98_975 ();
 b15zdnd11an1n04x5 FILLER_98_983 ();
 b15zdnd00an1n01x5 FILLER_98_987 ();
 b15zdnd11an1n64x5 FILLER_98_991 ();
 b15zdnd00an1n01x5 FILLER_98_1055 ();
 b15zdnd11an1n32x5 FILLER_98_1081 ();
 b15zdnd11an1n16x5 FILLER_98_1113 ();
 b15zdnd11an1n08x5 FILLER_98_1129 ();
 b15zdnd00an1n02x5 FILLER_98_1137 ();
 b15zdnd11an1n32x5 FILLER_98_1159 ();
 b15zdnd11an1n04x5 FILLER_98_1191 ();
 b15zdnd00an1n02x5 FILLER_98_1195 ();
 b15zdnd11an1n04x5 FILLER_98_1220 ();
 b15zdnd00an1n02x5 FILLER_98_1224 ();
 b15zdnd00an1n01x5 FILLER_98_1226 ();
 b15zdnd11an1n04x5 FILLER_98_1245 ();
 b15zdnd11an1n16x5 FILLER_98_1253 ();
 b15zdnd00an1n02x5 FILLER_98_1269 ();
 b15zdnd00an1n01x5 FILLER_98_1271 ();
 b15zdnd11an1n32x5 FILLER_98_1282 ();
 b15zdnd11an1n08x5 FILLER_98_1314 ();
 b15zdnd11an1n04x5 FILLER_98_1322 ();
 b15zdnd00an1n02x5 FILLER_98_1326 ();
 b15zdnd11an1n64x5 FILLER_98_1360 ();
 b15zdnd11an1n08x5 FILLER_98_1424 ();
 b15zdnd00an1n02x5 FILLER_98_1432 ();
 b15zdnd00an1n01x5 FILLER_98_1434 ();
 b15zdnd11an1n64x5 FILLER_98_1445 ();
 b15zdnd11an1n08x5 FILLER_98_1509 ();
 b15zdnd11an1n04x5 FILLER_98_1517 ();
 b15zdnd00an1n01x5 FILLER_98_1521 ();
 b15zdnd11an1n32x5 FILLER_98_1532 ();
 b15zdnd11an1n08x5 FILLER_98_1564 ();
 b15zdnd11an1n08x5 FILLER_98_1596 ();
 b15zdnd11an1n64x5 FILLER_98_1618 ();
 b15zdnd11an1n32x5 FILLER_98_1682 ();
 b15zdnd11an1n16x5 FILLER_98_1714 ();
 b15zdnd00an1n02x5 FILLER_98_1730 ();
 b15zdnd11an1n64x5 FILLER_98_1752 ();
 b15zdnd11an1n16x5 FILLER_98_1816 ();
 b15zdnd11an1n04x5 FILLER_98_1832 ();
 b15zdnd11an1n32x5 FILLER_98_1843 ();
 b15zdnd11an1n16x5 FILLER_98_1875 ();
 b15zdnd11an1n04x5 FILLER_98_1891 ();
 b15zdnd00an1n02x5 FILLER_98_1895 ();
 b15zdnd11an1n04x5 FILLER_98_1909 ();
 b15zdnd00an1n01x5 FILLER_98_1913 ();
 b15zdnd11an1n04x5 FILLER_98_1942 ();
 b15zdnd11an1n32x5 FILLER_98_1953 ();
 b15zdnd11an1n08x5 FILLER_98_1985 ();
 b15zdnd11an1n04x5 FILLER_98_1993 ();
 b15zdnd11an1n08x5 FILLER_98_2004 ();
 b15zdnd11an1n04x5 FILLER_98_2012 ();
 b15zdnd00an1n01x5 FILLER_98_2016 ();
 b15zdnd11an1n32x5 FILLER_98_2023 ();
 b15zdnd11an1n08x5 FILLER_98_2055 ();
 b15zdnd11an1n04x5 FILLER_98_2063 ();
 b15zdnd00an1n02x5 FILLER_98_2067 ();
 b15zdnd00an1n01x5 FILLER_98_2069 ();
 b15zdnd11an1n64x5 FILLER_98_2082 ();
 b15zdnd11an1n08x5 FILLER_98_2146 ();
 b15zdnd11an1n32x5 FILLER_98_2162 ();
 b15zdnd11an1n08x5 FILLER_98_2194 ();
 b15zdnd11an1n04x5 FILLER_98_2202 ();
 b15zdnd00an1n01x5 FILLER_98_2206 ();
 b15zdnd11an1n08x5 FILLER_98_2213 ();
 b15zdnd11an1n32x5 FILLER_98_2233 ();
 b15zdnd11an1n08x5 FILLER_98_2265 ();
 b15zdnd00an1n02x5 FILLER_98_2273 ();
 b15zdnd00an1n01x5 FILLER_98_2275 ();
 b15zdnd11an1n64x5 FILLER_99_0 ();
 b15zdnd11an1n64x5 FILLER_99_64 ();
 b15zdnd11an1n04x5 FILLER_99_128 ();
 b15zdnd11an1n16x5 FILLER_99_145 ();
 b15zdnd11an1n08x5 FILLER_99_161 ();
 b15zdnd00an1n01x5 FILLER_99_169 ();
 b15zdnd11an1n04x5 FILLER_99_185 ();
 b15zdnd11an1n64x5 FILLER_99_201 ();
 b15zdnd11an1n64x5 FILLER_99_265 ();
 b15zdnd11an1n64x5 FILLER_99_329 ();
 b15zdnd11an1n32x5 FILLER_99_393 ();
 b15zdnd11an1n16x5 FILLER_99_425 ();
 b15zdnd11an1n04x5 FILLER_99_441 ();
 b15zdnd00an1n02x5 FILLER_99_445 ();
 b15zdnd00an1n01x5 FILLER_99_447 ();
 b15zdnd11an1n16x5 FILLER_99_456 ();
 b15zdnd11an1n04x5 FILLER_99_472 ();
 b15zdnd11an1n08x5 FILLER_99_482 ();
 b15zdnd11an1n04x5 FILLER_99_490 ();
 b15zdnd00an1n01x5 FILLER_99_494 ();
 b15zdnd11an1n04x5 FILLER_99_499 ();
 b15zdnd11an1n08x5 FILLER_99_509 ();
 b15zdnd11an1n04x5 FILLER_99_517 ();
 b15zdnd00an1n02x5 FILLER_99_521 ();
 b15zdnd00an1n01x5 FILLER_99_523 ();
 b15zdnd11an1n16x5 FILLER_99_529 ();
 b15zdnd11an1n08x5 FILLER_99_545 ();
 b15zdnd11an1n04x5 FILLER_99_553 ();
 b15zdnd00an1n02x5 FILLER_99_557 ();
 b15zdnd00an1n01x5 FILLER_99_559 ();
 b15zdnd11an1n32x5 FILLER_99_568 ();
 b15zdnd11an1n04x5 FILLER_99_600 ();
 b15zdnd11an1n32x5 FILLER_99_617 ();
 b15zdnd11an1n16x5 FILLER_99_649 ();
 b15zdnd00an1n02x5 FILLER_99_665 ();
 b15zdnd00an1n01x5 FILLER_99_667 ();
 b15zdnd11an1n04x5 FILLER_99_694 ();
 b15zdnd11an1n04x5 FILLER_99_708 ();
 b15zdnd00an1n02x5 FILLER_99_712 ();
 b15zdnd11an1n08x5 FILLER_99_719 ();
 b15zdnd00an1n01x5 FILLER_99_727 ();
 b15zdnd11an1n32x5 FILLER_99_744 ();
 b15zdnd11an1n08x5 FILLER_99_776 ();
 b15zdnd11an1n04x5 FILLER_99_784 ();
 b15zdnd11an1n16x5 FILLER_99_802 ();
 b15zdnd00an1n02x5 FILLER_99_818 ();
 b15zdnd11an1n16x5 FILLER_99_825 ();
 b15zdnd11an1n08x5 FILLER_99_841 ();
 b15zdnd11an1n04x5 FILLER_99_849 ();
 b15zdnd00an1n02x5 FILLER_99_853 ();
 b15zdnd11an1n04x5 FILLER_99_871 ();
 b15zdnd11an1n16x5 FILLER_99_885 ();
 b15zdnd11an1n08x5 FILLER_99_901 ();
 b15zdnd00an1n02x5 FILLER_99_909 ();
 b15zdnd11an1n64x5 FILLER_99_918 ();
 b15zdnd11an1n64x5 FILLER_99_982 ();
 b15zdnd11an1n16x5 FILLER_99_1046 ();
 b15zdnd11an1n08x5 FILLER_99_1062 ();
 b15zdnd11an1n04x5 FILLER_99_1070 ();
 b15zdnd00an1n02x5 FILLER_99_1074 ();
 b15zdnd11an1n64x5 FILLER_99_1101 ();
 b15zdnd11an1n32x5 FILLER_99_1165 ();
 b15zdnd11an1n08x5 FILLER_99_1197 ();
 b15zdnd00an1n02x5 FILLER_99_1205 ();
 b15zdnd11an1n04x5 FILLER_99_1224 ();
 b15zdnd11an1n32x5 FILLER_99_1244 ();
 b15zdnd11an1n08x5 FILLER_99_1276 ();
 b15zdnd11an1n04x5 FILLER_99_1284 ();
 b15zdnd00an1n02x5 FILLER_99_1288 ();
 b15zdnd11an1n32x5 FILLER_99_1295 ();
 b15zdnd11an1n16x5 FILLER_99_1327 ();
 b15zdnd11an1n04x5 FILLER_99_1343 ();
 b15zdnd00an1n01x5 FILLER_99_1347 ();
 b15zdnd11an1n16x5 FILLER_99_1354 ();
 b15zdnd11an1n64x5 FILLER_99_1375 ();
 b15zdnd11an1n16x5 FILLER_99_1439 ();
 b15zdnd00an1n01x5 FILLER_99_1455 ();
 b15zdnd11an1n32x5 FILLER_99_1471 ();
 b15zdnd00an1n02x5 FILLER_99_1503 ();
 b15zdnd00an1n01x5 FILLER_99_1505 ();
 b15zdnd11an1n32x5 FILLER_99_1523 ();
 b15zdnd11an1n16x5 FILLER_99_1555 ();
 b15zdnd00an1n01x5 FILLER_99_1571 ();
 b15zdnd11an1n04x5 FILLER_99_1591 ();
 b15zdnd11an1n08x5 FILLER_99_1603 ();
 b15zdnd00an1n02x5 FILLER_99_1611 ();
 b15zdnd00an1n01x5 FILLER_99_1613 ();
 b15zdnd11an1n64x5 FILLER_99_1624 ();
 b15zdnd11an1n64x5 FILLER_99_1688 ();
 b15zdnd11an1n08x5 FILLER_99_1752 ();
 b15zdnd11an1n04x5 FILLER_99_1760 ();
 b15zdnd00an1n02x5 FILLER_99_1764 ();
 b15zdnd11an1n16x5 FILLER_99_1773 ();
 b15zdnd11an1n08x5 FILLER_99_1789 ();
 b15zdnd00an1n01x5 FILLER_99_1797 ();
 b15zdnd11an1n04x5 FILLER_99_1803 ();
 b15zdnd00an1n01x5 FILLER_99_1807 ();
 b15zdnd11an1n16x5 FILLER_99_1816 ();
 b15zdnd11an1n04x5 FILLER_99_1832 ();
 b15zdnd00an1n02x5 FILLER_99_1836 ();
 b15zdnd11an1n64x5 FILLER_99_1849 ();
 b15zdnd11an1n16x5 FILLER_99_1913 ();
 b15zdnd11an1n08x5 FILLER_99_1929 ();
 b15zdnd11an1n04x5 FILLER_99_1937 ();
 b15zdnd00an1n02x5 FILLER_99_1941 ();
 b15zdnd00an1n01x5 FILLER_99_1943 ();
 b15zdnd11an1n08x5 FILLER_99_1962 ();
 b15zdnd00an1n02x5 FILLER_99_1970 ();
 b15zdnd00an1n01x5 FILLER_99_1972 ();
 b15zdnd11an1n64x5 FILLER_99_1989 ();
 b15zdnd11an1n64x5 FILLER_99_2053 ();
 b15zdnd11an1n04x5 FILLER_99_2117 ();
 b15zdnd00an1n01x5 FILLER_99_2121 ();
 b15zdnd11an1n16x5 FILLER_99_2136 ();
 b15zdnd11an1n08x5 FILLER_99_2152 ();
 b15zdnd00an1n01x5 FILLER_99_2160 ();
 b15zdnd11an1n08x5 FILLER_99_2165 ();
 b15zdnd11an1n04x5 FILLER_99_2173 ();
 b15zdnd11an1n08x5 FILLER_99_2193 ();
 b15zdnd11an1n04x5 FILLER_99_2201 ();
 b15zdnd00an1n01x5 FILLER_99_2205 ();
 b15zdnd11an1n64x5 FILLER_99_2220 ();
 b15zdnd11an1n64x5 FILLER_100_8 ();
 b15zdnd11an1n32x5 FILLER_100_72 ();
 b15zdnd11an1n08x5 FILLER_100_104 ();
 b15zdnd11an1n08x5 FILLER_100_119 ();
 b15zdnd11an1n04x5 FILLER_100_127 ();
 b15zdnd00an1n01x5 FILLER_100_131 ();
 b15zdnd11an1n32x5 FILLER_100_140 ();
 b15zdnd11an1n16x5 FILLER_100_172 ();
 b15zdnd11an1n04x5 FILLER_100_188 ();
 b15zdnd00an1n02x5 FILLER_100_192 ();
 b15zdnd11an1n64x5 FILLER_100_202 ();
 b15zdnd11an1n64x5 FILLER_100_266 ();
 b15zdnd00an1n01x5 FILLER_100_330 ();
 b15zdnd11an1n64x5 FILLER_100_351 ();
 b15zdnd11an1n64x5 FILLER_100_415 ();
 b15zdnd00an1n02x5 FILLER_100_479 ();
 b15zdnd11an1n08x5 FILLER_100_487 ();
 b15zdnd11an1n04x5 FILLER_100_495 ();
 b15zdnd00an1n02x5 FILLER_100_499 ();
 b15zdnd11an1n16x5 FILLER_100_506 ();
 b15zdnd11an1n08x5 FILLER_100_522 ();
 b15zdnd11an1n04x5 FILLER_100_530 ();
 b15zdnd00an1n01x5 FILLER_100_534 ();
 b15zdnd11an1n64x5 FILLER_100_545 ();
 b15zdnd00an1n02x5 FILLER_100_609 ();
 b15zdnd11an1n04x5 FILLER_100_617 ();
 b15zdnd11an1n04x5 FILLER_100_625 ();
 b15zdnd11an1n08x5 FILLER_100_636 ();
 b15zdnd11an1n04x5 FILLER_100_644 ();
 b15zdnd00an1n02x5 FILLER_100_648 ();
 b15zdnd11an1n04x5 FILLER_100_662 ();
 b15zdnd11an1n08x5 FILLER_100_690 ();
 b15zdnd11an1n04x5 FILLER_100_698 ();
 b15zdnd00an1n02x5 FILLER_100_702 ();
 b15zdnd00an1n02x5 FILLER_100_716 ();
 b15zdnd00an1n02x5 FILLER_100_726 ();
 b15zdnd00an1n01x5 FILLER_100_728 ();
 b15zdnd11an1n08x5 FILLER_100_739 ();
 b15zdnd11an1n16x5 FILLER_100_754 ();
 b15zdnd11an1n08x5 FILLER_100_770 ();
 b15zdnd00an1n01x5 FILLER_100_778 ();
 b15zdnd11an1n32x5 FILLER_100_783 ();
 b15zdnd11an1n64x5 FILLER_100_827 ();
 b15zdnd11an1n64x5 FILLER_100_891 ();
 b15zdnd11an1n32x5 FILLER_100_955 ();
 b15zdnd11an1n16x5 FILLER_100_987 ();
 b15zdnd11an1n04x5 FILLER_100_1024 ();
 b15zdnd11an1n04x5 FILLER_100_1032 ();
 b15zdnd11an1n32x5 FILLER_100_1041 ();
 b15zdnd00an1n02x5 FILLER_100_1073 ();
 b15zdnd11an1n32x5 FILLER_100_1095 ();
 b15zdnd11an1n08x5 FILLER_100_1127 ();
 b15zdnd00an1n02x5 FILLER_100_1135 ();
 b15zdnd11an1n32x5 FILLER_100_1168 ();
 b15zdnd11an1n16x5 FILLER_100_1200 ();
 b15zdnd11an1n04x5 FILLER_100_1216 ();
 b15zdnd00an1n01x5 FILLER_100_1220 ();
 b15zdnd11an1n08x5 FILLER_100_1237 ();
 b15zdnd11an1n04x5 FILLER_100_1267 ();
 b15zdnd00an1n02x5 FILLER_100_1271 ();
 b15zdnd00an1n01x5 FILLER_100_1273 ();
 b15zdnd11an1n04x5 FILLER_100_1284 ();
 b15zdnd00an1n02x5 FILLER_100_1288 ();
 b15zdnd00an1n01x5 FILLER_100_1290 ();
 b15zdnd11an1n32x5 FILLER_100_1298 ();
 b15zdnd00an1n01x5 FILLER_100_1330 ();
 b15zdnd11an1n08x5 FILLER_100_1335 ();
 b15zdnd11an1n04x5 FILLER_100_1343 ();
 b15zdnd11an1n08x5 FILLER_100_1354 ();
 b15zdnd11an1n64x5 FILLER_100_1376 ();
 b15zdnd11an1n08x5 FILLER_100_1440 ();
 b15zdnd00an1n02x5 FILLER_100_1448 ();
 b15zdnd00an1n01x5 FILLER_100_1450 ();
 b15zdnd11an1n64x5 FILLER_100_1458 ();
 b15zdnd11an1n64x5 FILLER_100_1522 ();
 b15zdnd11an1n16x5 FILLER_100_1586 ();
 b15zdnd11an1n08x5 FILLER_100_1602 ();
 b15zdnd11an1n04x5 FILLER_100_1610 ();
 b15zdnd00an1n02x5 FILLER_100_1614 ();
 b15zdnd11an1n16x5 FILLER_100_1621 ();
 b15zdnd11an1n04x5 FILLER_100_1637 ();
 b15zdnd11an1n16x5 FILLER_100_1661 ();
 b15zdnd11an1n08x5 FILLER_100_1686 ();
 b15zdnd00an1n02x5 FILLER_100_1694 ();
 b15zdnd11an1n32x5 FILLER_100_1707 ();
 b15zdnd11an1n16x5 FILLER_100_1739 ();
 b15zdnd11an1n04x5 FILLER_100_1755 ();
 b15zdnd11an1n08x5 FILLER_100_1765 ();
 b15zdnd00an1n01x5 FILLER_100_1773 ();
 b15zdnd11an1n16x5 FILLER_100_1790 ();
 b15zdnd00an1n01x5 FILLER_100_1806 ();
 b15zdnd11an1n16x5 FILLER_100_1813 ();
 b15zdnd11an1n08x5 FILLER_100_1842 ();
 b15zdnd11an1n04x5 FILLER_100_1850 ();
 b15zdnd00an1n02x5 FILLER_100_1854 ();
 b15zdnd11an1n04x5 FILLER_100_1868 ();
 b15zdnd11an1n64x5 FILLER_100_1881 ();
 b15zdnd11an1n32x5 FILLER_100_1945 ();
 b15zdnd11an1n08x5 FILLER_100_1977 ();
 b15zdnd00an1n02x5 FILLER_100_1985 ();
 b15zdnd00an1n01x5 FILLER_100_1987 ();
 b15zdnd11an1n08x5 FILLER_100_2000 ();
 b15zdnd00an1n02x5 FILLER_100_2008 ();
 b15zdnd00an1n01x5 FILLER_100_2010 ();
 b15zdnd11an1n04x5 FILLER_100_2017 ();
 b15zdnd11an1n64x5 FILLER_100_2028 ();
 b15zdnd11an1n16x5 FILLER_100_2097 ();
 b15zdnd11an1n08x5 FILLER_100_2113 ();
 b15zdnd00an1n02x5 FILLER_100_2121 ();
 b15zdnd00an1n01x5 FILLER_100_2123 ();
 b15zdnd11an1n16x5 FILLER_100_2136 ();
 b15zdnd00an1n02x5 FILLER_100_2152 ();
 b15zdnd11an1n16x5 FILLER_100_2162 ();
 b15zdnd00an1n02x5 FILLER_100_2178 ();
 b15zdnd00an1n01x5 FILLER_100_2180 ();
 b15zdnd11an1n04x5 FILLER_100_2186 ();
 b15zdnd11an1n08x5 FILLER_100_2202 ();
 b15zdnd00an1n02x5 FILLER_100_2210 ();
 b15zdnd11an1n32x5 FILLER_100_2218 ();
 b15zdnd11an1n16x5 FILLER_100_2250 ();
 b15zdnd11an1n08x5 FILLER_100_2266 ();
 b15zdnd00an1n02x5 FILLER_100_2274 ();
 b15zdnd11an1n64x5 FILLER_101_0 ();
 b15zdnd11an1n64x5 FILLER_101_64 ();
 b15zdnd11an1n16x5 FILLER_101_128 ();
 b15zdnd11an1n08x5 FILLER_101_144 ();
 b15zdnd11an1n04x5 FILLER_101_152 ();
 b15zdnd00an1n02x5 FILLER_101_156 ();
 b15zdnd00an1n01x5 FILLER_101_158 ();
 b15zdnd11an1n08x5 FILLER_101_175 ();
 b15zdnd11an1n04x5 FILLER_101_183 ();
 b15zdnd00an1n01x5 FILLER_101_187 ();
 b15zdnd11an1n08x5 FILLER_101_194 ();
 b15zdnd00an1n02x5 FILLER_101_202 ();
 b15zdnd11an1n16x5 FILLER_101_212 ();
 b15zdnd11an1n08x5 FILLER_101_228 ();
 b15zdnd11an1n04x5 FILLER_101_236 ();
 b15zdnd00an1n02x5 FILLER_101_240 ();
 b15zdnd11an1n32x5 FILLER_101_249 ();
 b15zdnd11an1n16x5 FILLER_101_281 ();
 b15zdnd11an1n04x5 FILLER_101_297 ();
 b15zdnd00an1n01x5 FILLER_101_301 ();
 b15zdnd11an1n04x5 FILLER_101_318 ();
 b15zdnd00an1n01x5 FILLER_101_322 ();
 b15zdnd11an1n64x5 FILLER_101_333 ();
 b15zdnd11an1n16x5 FILLER_101_397 ();
 b15zdnd11an1n08x5 FILLER_101_413 ();
 b15zdnd00an1n02x5 FILLER_101_421 ();
 b15zdnd11an1n08x5 FILLER_101_428 ();
 b15zdnd11an1n04x5 FILLER_101_445 ();
 b15zdnd11an1n32x5 FILLER_101_454 ();
 b15zdnd11an1n16x5 FILLER_101_486 ();
 b15zdnd11an1n08x5 FILLER_101_512 ();
 b15zdnd00an1n02x5 FILLER_101_520 ();
 b15zdnd00an1n01x5 FILLER_101_522 ();
 b15zdnd11an1n04x5 FILLER_101_540 ();
 b15zdnd11an1n32x5 FILLER_101_558 ();
 b15zdnd11an1n08x5 FILLER_101_590 ();
 b15zdnd11an1n04x5 FILLER_101_598 ();
 b15zdnd11an1n64x5 FILLER_101_623 ();
 b15zdnd11an1n64x5 FILLER_101_687 ();
 b15zdnd11an1n08x5 FILLER_101_751 ();
 b15zdnd11an1n04x5 FILLER_101_759 ();
 b15zdnd00an1n01x5 FILLER_101_763 ();
 b15zdnd11an1n64x5 FILLER_101_783 ();
 b15zdnd00an1n02x5 FILLER_101_847 ();
 b15zdnd11an1n16x5 FILLER_101_858 ();
 b15zdnd11an1n04x5 FILLER_101_874 ();
 b15zdnd11an1n64x5 FILLER_101_884 ();
 b15zdnd11an1n64x5 FILLER_101_948 ();
 b15zdnd11an1n08x5 FILLER_101_1012 ();
 b15zdnd00an1n01x5 FILLER_101_1020 ();
 b15zdnd11an1n04x5 FILLER_101_1030 ();
 b15zdnd11an1n64x5 FILLER_101_1043 ();
 b15zdnd11an1n04x5 FILLER_101_1107 ();
 b15zdnd00an1n02x5 FILLER_101_1111 ();
 b15zdnd00an1n01x5 FILLER_101_1113 ();
 b15zdnd11an1n16x5 FILLER_101_1125 ();
 b15zdnd00an1n02x5 FILLER_101_1141 ();
 b15zdnd00an1n01x5 FILLER_101_1143 ();
 b15zdnd11an1n32x5 FILLER_101_1155 ();
 b15zdnd11an1n16x5 FILLER_101_1187 ();
 b15zdnd11an1n08x5 FILLER_101_1203 ();
 b15zdnd00an1n02x5 FILLER_101_1211 ();
 b15zdnd11an1n16x5 FILLER_101_1237 ();
 b15zdnd11an1n04x5 FILLER_101_1253 ();
 b15zdnd00an1n02x5 FILLER_101_1257 ();
 b15zdnd00an1n01x5 FILLER_101_1259 ();
 b15zdnd11an1n04x5 FILLER_101_1276 ();
 b15zdnd11an1n08x5 FILLER_101_1296 ();
 b15zdnd00an1n02x5 FILLER_101_1304 ();
 b15zdnd00an1n01x5 FILLER_101_1306 ();
 b15zdnd11an1n16x5 FILLER_101_1317 ();
 b15zdnd11an1n04x5 FILLER_101_1333 ();
 b15zdnd00an1n02x5 FILLER_101_1337 ();
 b15zdnd00an1n01x5 FILLER_101_1339 ();
 b15zdnd11an1n32x5 FILLER_101_1345 ();
 b15zdnd00an1n02x5 FILLER_101_1377 ();
 b15zdnd00an1n01x5 FILLER_101_1379 ();
 b15zdnd11an1n08x5 FILLER_101_1386 ();
 b15zdnd00an1n02x5 FILLER_101_1394 ();
 b15zdnd11an1n04x5 FILLER_101_1402 ();
 b15zdnd11an1n08x5 FILLER_101_1413 ();
 b15zdnd00an1n02x5 FILLER_101_1421 ();
 b15zdnd00an1n01x5 FILLER_101_1423 ();
 b15zdnd11an1n04x5 FILLER_101_1431 ();
 b15zdnd00an1n02x5 FILLER_101_1435 ();
 b15zdnd11an1n08x5 FILLER_101_1447 ();
 b15zdnd11an1n04x5 FILLER_101_1455 ();
 b15zdnd00an1n01x5 FILLER_101_1459 ();
 b15zdnd11an1n04x5 FILLER_101_1469 ();
 b15zdnd11an1n08x5 FILLER_101_1479 ();
 b15zdnd00an1n01x5 FILLER_101_1487 ();
 b15zdnd11an1n32x5 FILLER_101_1497 ();
 b15zdnd11an1n16x5 FILLER_101_1529 ();
 b15zdnd11an1n08x5 FILLER_101_1545 ();
 b15zdnd11an1n32x5 FILLER_101_1571 ();
 b15zdnd11an1n16x5 FILLER_101_1623 ();
 b15zdnd00an1n01x5 FILLER_101_1639 ();
 b15zdnd11an1n16x5 FILLER_101_1645 ();
 b15zdnd00an1n02x5 FILLER_101_1661 ();
 b15zdnd00an1n01x5 FILLER_101_1663 ();
 b15zdnd11an1n32x5 FILLER_101_1690 ();
 b15zdnd11an1n16x5 FILLER_101_1722 ();
 b15zdnd11an1n04x5 FILLER_101_1738 ();
 b15zdnd00an1n01x5 FILLER_101_1742 ();
 b15zdnd11an1n08x5 FILLER_101_1751 ();
 b15zdnd11an1n04x5 FILLER_101_1759 ();
 b15zdnd00an1n02x5 FILLER_101_1763 ();
 b15zdnd00an1n01x5 FILLER_101_1765 ();
 b15zdnd11an1n16x5 FILLER_101_1771 ();
 b15zdnd11an1n08x5 FILLER_101_1787 ();
 b15zdnd00an1n02x5 FILLER_101_1795 ();
 b15zdnd00an1n01x5 FILLER_101_1797 ();
 b15zdnd11an1n16x5 FILLER_101_1814 ();
 b15zdnd11an1n08x5 FILLER_101_1830 ();
 b15zdnd11an1n04x5 FILLER_101_1847 ();
 b15zdnd00an1n01x5 FILLER_101_1851 ();
 b15zdnd11an1n04x5 FILLER_101_1857 ();
 b15zdnd11an1n08x5 FILLER_101_1875 ();
 b15zdnd00an1n01x5 FILLER_101_1883 ();
 b15zdnd11an1n32x5 FILLER_101_1891 ();
 b15zdnd00an1n01x5 FILLER_101_1923 ();
 b15zdnd11an1n16x5 FILLER_101_1928 ();
 b15zdnd11an1n04x5 FILLER_101_1944 ();
 b15zdnd00an1n02x5 FILLER_101_1948 ();
 b15zdnd00an1n01x5 FILLER_101_1950 ();
 b15zdnd11an1n32x5 FILLER_101_1963 ();
 b15zdnd11an1n08x5 FILLER_101_1995 ();
 b15zdnd00an1n02x5 FILLER_101_2003 ();
 b15zdnd11an1n04x5 FILLER_101_2010 ();
 b15zdnd11an1n32x5 FILLER_101_2026 ();
 b15zdnd11an1n08x5 FILLER_101_2058 ();
 b15zdnd11an1n04x5 FILLER_101_2066 ();
 b15zdnd00an1n02x5 FILLER_101_2070 ();
 b15zdnd11an1n04x5 FILLER_101_2077 ();
 b15zdnd11an1n08x5 FILLER_101_2087 ();
 b15zdnd11an1n32x5 FILLER_101_2106 ();
 b15zdnd00an1n02x5 FILLER_101_2138 ();
 b15zdnd00an1n01x5 FILLER_101_2140 ();
 b15zdnd11an1n08x5 FILLER_101_2146 ();
 b15zdnd11an1n04x5 FILLER_101_2154 ();
 b15zdnd00an1n02x5 FILLER_101_2158 ();
 b15zdnd00an1n01x5 FILLER_101_2160 ();
 b15zdnd11an1n64x5 FILLER_101_2169 ();
 b15zdnd11an1n32x5 FILLER_101_2233 ();
 b15zdnd11an1n16x5 FILLER_101_2265 ();
 b15zdnd00an1n02x5 FILLER_101_2281 ();
 b15zdnd00an1n01x5 FILLER_101_2283 ();
 b15zdnd11an1n64x5 FILLER_102_8 ();
 b15zdnd11an1n64x5 FILLER_102_72 ();
 b15zdnd11an1n08x5 FILLER_102_136 ();
 b15zdnd11an1n04x5 FILLER_102_144 ();
 b15zdnd00an1n02x5 FILLER_102_148 ();
 b15zdnd00an1n01x5 FILLER_102_150 ();
 b15zdnd11an1n64x5 FILLER_102_160 ();
 b15zdnd11an1n16x5 FILLER_102_224 ();
 b15zdnd11an1n08x5 FILLER_102_240 ();
 b15zdnd11an1n04x5 FILLER_102_248 ();
 b15zdnd00an1n01x5 FILLER_102_252 ();
 b15zdnd11an1n32x5 FILLER_102_267 ();
 b15zdnd11an1n16x5 FILLER_102_299 ();
 b15zdnd11an1n08x5 FILLER_102_315 ();
 b15zdnd11an1n64x5 FILLER_102_329 ();
 b15zdnd11an1n32x5 FILLER_102_393 ();
 b15zdnd00an1n02x5 FILLER_102_425 ();
 b15zdnd00an1n01x5 FILLER_102_427 ();
 b15zdnd11an1n04x5 FILLER_102_438 ();
 b15zdnd11an1n16x5 FILLER_102_451 ();
 b15zdnd11an1n04x5 FILLER_102_467 ();
 b15zdnd00an1n02x5 FILLER_102_471 ();
 b15zdnd00an1n01x5 FILLER_102_473 ();
 b15zdnd11an1n64x5 FILLER_102_490 ();
 b15zdnd00an1n02x5 FILLER_102_554 ();
 b15zdnd00an1n01x5 FILLER_102_556 ();
 b15zdnd11an1n04x5 FILLER_102_572 ();
 b15zdnd11an1n32x5 FILLER_102_589 ();
 b15zdnd11an1n04x5 FILLER_102_621 ();
 b15zdnd00an1n01x5 FILLER_102_625 ();
 b15zdnd11an1n08x5 FILLER_102_631 ();
 b15zdnd00an1n02x5 FILLER_102_639 ();
 b15zdnd11an1n04x5 FILLER_102_653 ();
 b15zdnd11an1n32x5 FILLER_102_677 ();
 b15zdnd11an1n08x5 FILLER_102_709 ();
 b15zdnd00an1n01x5 FILLER_102_717 ();
 b15zdnd11an1n32x5 FILLER_102_726 ();
 b15zdnd11an1n04x5 FILLER_102_758 ();
 b15zdnd00an1n01x5 FILLER_102_762 ();
 b15zdnd11an1n04x5 FILLER_102_771 ();
 b15zdnd00an1n02x5 FILLER_102_775 ();
 b15zdnd11an1n08x5 FILLER_102_783 ();
 b15zdnd11an1n04x5 FILLER_102_791 ();
 b15zdnd00an1n01x5 FILLER_102_795 ();
 b15zdnd11an1n08x5 FILLER_102_802 ();
 b15zdnd11an1n04x5 FILLER_102_810 ();
 b15zdnd00an1n01x5 FILLER_102_814 ();
 b15zdnd11an1n16x5 FILLER_102_829 ();
 b15zdnd11an1n04x5 FILLER_102_845 ();
 b15zdnd00an1n02x5 FILLER_102_849 ();
 b15zdnd11an1n04x5 FILLER_102_856 ();
 b15zdnd11an1n08x5 FILLER_102_868 ();
 b15zdnd00an1n02x5 FILLER_102_876 ();
 b15zdnd11an1n32x5 FILLER_102_890 ();
 b15zdnd11an1n16x5 FILLER_102_922 ();
 b15zdnd11an1n08x5 FILLER_102_938 ();
 b15zdnd11an1n64x5 FILLER_102_966 ();
 b15zdnd11an1n64x5 FILLER_102_1030 ();
 b15zdnd11an1n32x5 FILLER_102_1094 ();
 b15zdnd11an1n08x5 FILLER_102_1126 ();
 b15zdnd11an1n32x5 FILLER_102_1154 ();
 b15zdnd11an1n16x5 FILLER_102_1186 ();
 b15zdnd11an1n08x5 FILLER_102_1202 ();
 b15zdnd11an1n04x5 FILLER_102_1210 ();
 b15zdnd00an1n01x5 FILLER_102_1214 ();
 b15zdnd11an1n64x5 FILLER_102_1228 ();
 b15zdnd11an1n32x5 FILLER_102_1292 ();
 b15zdnd11an1n32x5 FILLER_102_1349 ();
 b15zdnd11an1n16x5 FILLER_102_1381 ();
 b15zdnd11an1n08x5 FILLER_102_1397 ();
 b15zdnd00an1n02x5 FILLER_102_1405 ();
 b15zdnd11an1n32x5 FILLER_102_1413 ();
 b15zdnd11an1n04x5 FILLER_102_1445 ();
 b15zdnd00an1n02x5 FILLER_102_1449 ();
 b15zdnd00an1n01x5 FILLER_102_1451 ();
 b15zdnd11an1n16x5 FILLER_102_1467 ();
 b15zdnd11an1n08x5 FILLER_102_1483 ();
 b15zdnd11an1n04x5 FILLER_102_1491 ();
 b15zdnd00an1n01x5 FILLER_102_1495 ();
 b15zdnd11an1n08x5 FILLER_102_1501 ();
 b15zdnd11an1n04x5 FILLER_102_1509 ();
 b15zdnd00an1n02x5 FILLER_102_1513 ();
 b15zdnd00an1n01x5 FILLER_102_1515 ();
 b15zdnd11an1n04x5 FILLER_102_1531 ();
 b15zdnd11an1n32x5 FILLER_102_1541 ();
 b15zdnd11an1n08x5 FILLER_102_1573 ();
 b15zdnd11an1n08x5 FILLER_102_1591 ();
 b15zdnd11an1n04x5 FILLER_102_1599 ();
 b15zdnd00an1n01x5 FILLER_102_1603 ();
 b15zdnd11an1n64x5 FILLER_102_1635 ();
 b15zdnd11an1n32x5 FILLER_102_1699 ();
 b15zdnd11an1n08x5 FILLER_102_1731 ();
 b15zdnd11an1n04x5 FILLER_102_1739 ();
 b15zdnd11an1n64x5 FILLER_102_1759 ();
 b15zdnd11an1n08x5 FILLER_102_1823 ();
 b15zdnd11an1n04x5 FILLER_102_1831 ();
 b15zdnd11an1n08x5 FILLER_102_1851 ();
 b15zdnd11an1n16x5 FILLER_102_1863 ();
 b15zdnd11an1n08x5 FILLER_102_1879 ();
 b15zdnd11an1n04x5 FILLER_102_1887 ();
 b15zdnd11an1n04x5 FILLER_102_1896 ();
 b15zdnd11an1n16x5 FILLER_102_1905 ();
 b15zdnd11an1n08x5 FILLER_102_1921 ();
 b15zdnd11an1n04x5 FILLER_102_1929 ();
 b15zdnd00an1n02x5 FILLER_102_1933 ();
 b15zdnd00an1n01x5 FILLER_102_1935 ();
 b15zdnd11an1n04x5 FILLER_102_1942 ();
 b15zdnd11an1n04x5 FILLER_102_1953 ();
 b15zdnd11an1n32x5 FILLER_102_1961 ();
 b15zdnd11an1n16x5 FILLER_102_1993 ();
 b15zdnd11an1n08x5 FILLER_102_2009 ();
 b15zdnd11an1n04x5 FILLER_102_2017 ();
 b15zdnd00an1n02x5 FILLER_102_2021 ();
 b15zdnd11an1n64x5 FILLER_102_2033 ();
 b15zdnd11an1n04x5 FILLER_102_2097 ();
 b15zdnd11an1n16x5 FILLER_102_2106 ();
 b15zdnd11an1n08x5 FILLER_102_2122 ();
 b15zdnd00an1n01x5 FILLER_102_2130 ();
 b15zdnd11an1n04x5 FILLER_102_2135 ();
 b15zdnd00an1n02x5 FILLER_102_2152 ();
 b15zdnd11an1n64x5 FILLER_102_2162 ();
 b15zdnd11an1n32x5 FILLER_102_2226 ();
 b15zdnd00an1n02x5 FILLER_102_2258 ();
 b15zdnd11an1n04x5 FILLER_102_2266 ();
 b15zdnd00an1n02x5 FILLER_102_2274 ();
 b15zdnd11an1n64x5 FILLER_103_0 ();
 b15zdnd11an1n64x5 FILLER_103_64 ();
 b15zdnd11an1n64x5 FILLER_103_128 ();
 b15zdnd11an1n32x5 FILLER_103_192 ();
 b15zdnd11an1n16x5 FILLER_103_224 ();
 b15zdnd11an1n04x5 FILLER_103_247 ();
 b15zdnd11an1n64x5 FILLER_103_261 ();
 b15zdnd11an1n64x5 FILLER_103_325 ();
 b15zdnd11an1n64x5 FILLER_103_389 ();
 b15zdnd11an1n64x5 FILLER_103_453 ();
 b15zdnd11an1n16x5 FILLER_103_517 ();
 b15zdnd00an1n02x5 FILLER_103_533 ();
 b15zdnd00an1n01x5 FILLER_103_535 ();
 b15zdnd11an1n04x5 FILLER_103_545 ();
 b15zdnd11an1n08x5 FILLER_103_569 ();
 b15zdnd00an1n01x5 FILLER_103_577 ();
 b15zdnd11an1n32x5 FILLER_103_584 ();
 b15zdnd11an1n08x5 FILLER_103_616 ();
 b15zdnd00an1n02x5 FILLER_103_624 ();
 b15zdnd00an1n01x5 FILLER_103_626 ();
 b15zdnd11an1n08x5 FILLER_103_642 ();
 b15zdnd11an1n04x5 FILLER_103_650 ();
 b15zdnd00an1n01x5 FILLER_103_654 ();
 b15zdnd11an1n16x5 FILLER_103_670 ();
 b15zdnd11an1n04x5 FILLER_103_686 ();
 b15zdnd00an1n01x5 FILLER_103_690 ();
 b15zdnd11an1n64x5 FILLER_103_703 ();
 b15zdnd11an1n08x5 FILLER_103_767 ();
 b15zdnd11an1n04x5 FILLER_103_775 ();
 b15zdnd00an1n01x5 FILLER_103_779 ();
 b15zdnd11an1n64x5 FILLER_103_801 ();
 b15zdnd11an1n32x5 FILLER_103_865 ();
 b15zdnd11an1n08x5 FILLER_103_897 ();
 b15zdnd11an1n04x5 FILLER_103_905 ();
 b15zdnd00an1n02x5 FILLER_103_909 ();
 b15zdnd11an1n04x5 FILLER_103_918 ();
 b15zdnd11an1n32x5 FILLER_103_927 ();
 b15zdnd11an1n16x5 FILLER_103_959 ();
 b15zdnd11an1n08x5 FILLER_103_975 ();
 b15zdnd11an1n04x5 FILLER_103_983 ();
 b15zdnd00an1n02x5 FILLER_103_987 ();
 b15zdnd00an1n01x5 FILLER_103_989 ();
 b15zdnd11an1n64x5 FILLER_103_995 ();
 b15zdnd11an1n64x5 FILLER_103_1059 ();
 b15zdnd11an1n64x5 FILLER_103_1123 ();
 b15zdnd11an1n16x5 FILLER_103_1187 ();
 b15zdnd11an1n08x5 FILLER_103_1203 ();
 b15zdnd11an1n32x5 FILLER_103_1227 ();
 b15zdnd11an1n08x5 FILLER_103_1259 ();
 b15zdnd00an1n01x5 FILLER_103_1267 ();
 b15zdnd11an1n64x5 FILLER_103_1273 ();
 b15zdnd11an1n08x5 FILLER_103_1337 ();
 b15zdnd11an1n04x5 FILLER_103_1345 ();
 b15zdnd00an1n01x5 FILLER_103_1349 ();
 b15zdnd11an1n64x5 FILLER_103_1366 ();
 b15zdnd11an1n64x5 FILLER_103_1430 ();
 b15zdnd00an1n02x5 FILLER_103_1494 ();
 b15zdnd11an1n16x5 FILLER_103_1503 ();
 b15zdnd11an1n08x5 FILLER_103_1519 ();
 b15zdnd11an1n04x5 FILLER_103_1527 ();
 b15zdnd00an1n01x5 FILLER_103_1531 ();
 b15zdnd11an1n16x5 FILLER_103_1546 ();
 b15zdnd11an1n08x5 FILLER_103_1562 ();
 b15zdnd11an1n04x5 FILLER_103_1570 ();
 b15zdnd00an1n01x5 FILLER_103_1574 ();
 b15zdnd11an1n64x5 FILLER_103_1591 ();
 b15zdnd11an1n64x5 FILLER_103_1655 ();
 b15zdnd11an1n16x5 FILLER_103_1719 ();
 b15zdnd11an1n04x5 FILLER_103_1735 ();
 b15zdnd00an1n02x5 FILLER_103_1739 ();
 b15zdnd11an1n64x5 FILLER_103_1751 ();
 b15zdnd11an1n64x5 FILLER_103_1815 ();
 b15zdnd11an1n64x5 FILLER_103_1879 ();
 b15zdnd11an1n32x5 FILLER_103_1943 ();
 b15zdnd11an1n08x5 FILLER_103_1975 ();
 b15zdnd11an1n32x5 FILLER_103_2004 ();
 b15zdnd11an1n16x5 FILLER_103_2036 ();
 b15zdnd00an1n02x5 FILLER_103_2052 ();
 b15zdnd00an1n01x5 FILLER_103_2054 ();
 b15zdnd11an1n16x5 FILLER_103_2061 ();
 b15zdnd00an1n01x5 FILLER_103_2077 ();
 b15zdnd11an1n08x5 FILLER_103_2088 ();
 b15zdnd00an1n02x5 FILLER_103_2096 ();
 b15zdnd11an1n32x5 FILLER_103_2110 ();
 b15zdnd11an1n16x5 FILLER_103_2142 ();
 b15zdnd11an1n08x5 FILLER_103_2158 ();
 b15zdnd11an1n04x5 FILLER_103_2166 ();
 b15zdnd00an1n02x5 FILLER_103_2170 ();
 b15zdnd11an1n64x5 FILLER_103_2176 ();
 b15zdnd11an1n08x5 FILLER_103_2240 ();
 b15zdnd11an1n04x5 FILLER_103_2248 ();
 b15zdnd00an1n01x5 FILLER_103_2252 ();
 b15zdnd11an1n04x5 FILLER_103_2273 ();
 b15zdnd00an1n01x5 FILLER_103_2277 ();
 b15zdnd00an1n02x5 FILLER_103_2282 ();
 b15zdnd11an1n64x5 FILLER_104_8 ();
 b15zdnd11an1n64x5 FILLER_104_72 ();
 b15zdnd11an1n64x5 FILLER_104_136 ();
 b15zdnd11an1n64x5 FILLER_104_200 ();
 b15zdnd11an1n64x5 FILLER_104_264 ();
 b15zdnd11an1n64x5 FILLER_104_328 ();
 b15zdnd11an1n64x5 FILLER_104_392 ();
 b15zdnd11an1n16x5 FILLER_104_456 ();
 b15zdnd11an1n32x5 FILLER_104_493 ();
 b15zdnd11an1n08x5 FILLER_104_525 ();
 b15zdnd00an1n02x5 FILLER_104_533 ();
 b15zdnd11an1n16x5 FILLER_104_540 ();
 b15zdnd11an1n32x5 FILLER_104_569 ();
 b15zdnd11an1n16x5 FILLER_104_601 ();
 b15zdnd00an1n01x5 FILLER_104_617 ();
 b15zdnd11an1n04x5 FILLER_104_638 ();
 b15zdnd11an1n16x5 FILLER_104_662 ();
 b15zdnd00an1n02x5 FILLER_104_678 ();
 b15zdnd11an1n04x5 FILLER_104_701 ();
 b15zdnd00an1n02x5 FILLER_104_705 ();
 b15zdnd00an1n02x5 FILLER_104_716 ();
 b15zdnd11an1n08x5 FILLER_104_726 ();
 b15zdnd11an1n04x5 FILLER_104_748 ();
 b15zdnd11an1n16x5 FILLER_104_759 ();
 b15zdnd11an1n32x5 FILLER_104_780 ();
 b15zdnd11an1n08x5 FILLER_104_812 ();
 b15zdnd11an1n04x5 FILLER_104_820 ();
 b15zdnd00an1n02x5 FILLER_104_824 ();
 b15zdnd00an1n01x5 FILLER_104_826 ();
 b15zdnd11an1n16x5 FILLER_104_840 ();
 b15zdnd11an1n64x5 FILLER_104_861 ();
 b15zdnd00an1n02x5 FILLER_104_925 ();
 b15zdnd00an1n01x5 FILLER_104_927 ();
 b15zdnd11an1n04x5 FILLER_104_954 ();
 b15zdnd11an1n16x5 FILLER_104_967 ();
 b15zdnd11an1n04x5 FILLER_104_983 ();
 b15zdnd00an1n02x5 FILLER_104_987 ();
 b15zdnd00an1n01x5 FILLER_104_989 ();
 b15zdnd11an1n64x5 FILLER_104_999 ();
 b15zdnd11an1n64x5 FILLER_104_1063 ();
 b15zdnd11an1n32x5 FILLER_104_1127 ();
 b15zdnd11an1n16x5 FILLER_104_1159 ();
 b15zdnd00an1n02x5 FILLER_104_1175 ();
 b15zdnd11an1n64x5 FILLER_104_1197 ();
 b15zdnd11an1n08x5 FILLER_104_1261 ();
 b15zdnd00an1n02x5 FILLER_104_1269 ();
 b15zdnd00an1n01x5 FILLER_104_1271 ();
 b15zdnd11an1n16x5 FILLER_104_1278 ();
 b15zdnd11an1n08x5 FILLER_104_1294 ();
 b15zdnd11an1n04x5 FILLER_104_1302 ();
 b15zdnd00an1n01x5 FILLER_104_1306 ();
 b15zdnd11an1n16x5 FILLER_104_1317 ();
 b15zdnd11an1n08x5 FILLER_104_1333 ();
 b15zdnd00an1n01x5 FILLER_104_1341 ();
 b15zdnd11an1n16x5 FILLER_104_1353 ();
 b15zdnd11an1n04x5 FILLER_104_1369 ();
 b15zdnd00an1n02x5 FILLER_104_1373 ();
 b15zdnd00an1n01x5 FILLER_104_1375 ();
 b15zdnd11an1n08x5 FILLER_104_1380 ();
 b15zdnd11an1n04x5 FILLER_104_1388 ();
 b15zdnd00an1n02x5 FILLER_104_1392 ();
 b15zdnd00an1n01x5 FILLER_104_1394 ();
 b15zdnd11an1n32x5 FILLER_104_1400 ();
 b15zdnd11an1n16x5 FILLER_104_1432 ();
 b15zdnd11an1n04x5 FILLER_104_1448 ();
 b15zdnd00an1n02x5 FILLER_104_1452 ();
 b15zdnd00an1n01x5 FILLER_104_1454 ();
 b15zdnd11an1n32x5 FILLER_104_1466 ();
 b15zdnd11an1n08x5 FILLER_104_1510 ();
 b15zdnd00an1n02x5 FILLER_104_1518 ();
 b15zdnd11an1n64x5 FILLER_104_1546 ();
 b15zdnd11an1n64x5 FILLER_104_1610 ();
 b15zdnd11an1n32x5 FILLER_104_1674 ();
 b15zdnd11an1n08x5 FILLER_104_1706 ();
 b15zdnd11an1n04x5 FILLER_104_1714 ();
 b15zdnd00an1n02x5 FILLER_104_1718 ();
 b15zdnd00an1n01x5 FILLER_104_1720 ();
 b15zdnd11an1n16x5 FILLER_104_1747 ();
 b15zdnd00an1n01x5 FILLER_104_1763 ();
 b15zdnd11an1n64x5 FILLER_104_1769 ();
 b15zdnd11an1n16x5 FILLER_104_1833 ();
 b15zdnd00an1n02x5 FILLER_104_1849 ();
 b15zdnd00an1n01x5 FILLER_104_1851 ();
 b15zdnd11an1n64x5 FILLER_104_1858 ();
 b15zdnd11an1n32x5 FILLER_104_1922 ();
 b15zdnd11an1n16x5 FILLER_104_1954 ();
 b15zdnd11an1n08x5 FILLER_104_1970 ();
 b15zdnd00an1n02x5 FILLER_104_1978 ();
 b15zdnd00an1n01x5 FILLER_104_1980 ();
 b15zdnd11an1n16x5 FILLER_104_1992 ();
 b15zdnd11an1n04x5 FILLER_104_2008 ();
 b15zdnd00an1n02x5 FILLER_104_2012 ();
 b15zdnd00an1n01x5 FILLER_104_2014 ();
 b15zdnd11an1n64x5 FILLER_104_2019 ();
 b15zdnd11an1n64x5 FILLER_104_2083 ();
 b15zdnd11an1n04x5 FILLER_104_2147 ();
 b15zdnd00an1n02x5 FILLER_104_2151 ();
 b15zdnd00an1n01x5 FILLER_104_2153 ();
 b15zdnd11an1n04x5 FILLER_104_2162 ();
 b15zdnd00an1n01x5 FILLER_104_2166 ();
 b15zdnd11an1n16x5 FILLER_104_2180 ();
 b15zdnd11an1n04x5 FILLER_104_2196 ();
 b15zdnd00an1n02x5 FILLER_104_2200 ();
 b15zdnd00an1n01x5 FILLER_104_2202 ();
 b15zdnd11an1n32x5 FILLER_104_2219 ();
 b15zdnd11an1n08x5 FILLER_104_2251 ();
 b15zdnd00an1n02x5 FILLER_104_2259 ();
 b15zdnd11an1n08x5 FILLER_104_2266 ();
 b15zdnd00an1n02x5 FILLER_104_2274 ();
 b15zdnd11an1n64x5 FILLER_105_0 ();
 b15zdnd11an1n64x5 FILLER_105_64 ();
 b15zdnd11an1n64x5 FILLER_105_128 ();
 b15zdnd11an1n64x5 FILLER_105_192 ();
 b15zdnd11an1n64x5 FILLER_105_256 ();
 b15zdnd11an1n64x5 FILLER_105_320 ();
 b15zdnd11an1n32x5 FILLER_105_384 ();
 b15zdnd11an1n16x5 FILLER_105_416 ();
 b15zdnd11an1n08x5 FILLER_105_432 ();
 b15zdnd11an1n04x5 FILLER_105_440 ();
 b15zdnd00an1n01x5 FILLER_105_444 ();
 b15zdnd11an1n08x5 FILLER_105_466 ();
 b15zdnd11an1n04x5 FILLER_105_474 ();
 b15zdnd00an1n02x5 FILLER_105_478 ();
 b15zdnd00an1n01x5 FILLER_105_480 ();
 b15zdnd11an1n16x5 FILLER_105_487 ();
 b15zdnd11an1n08x5 FILLER_105_503 ();
 b15zdnd11an1n04x5 FILLER_105_511 ();
 b15zdnd00an1n02x5 FILLER_105_515 ();
 b15zdnd00an1n01x5 FILLER_105_517 ();
 b15zdnd11an1n32x5 FILLER_105_534 ();
 b15zdnd11an1n16x5 FILLER_105_566 ();
 b15zdnd00an1n02x5 FILLER_105_582 ();
 b15zdnd11an1n08x5 FILLER_105_599 ();
 b15zdnd11an1n04x5 FILLER_105_607 ();
 b15zdnd00an1n02x5 FILLER_105_611 ();
 b15zdnd11an1n32x5 FILLER_105_625 ();
 b15zdnd11an1n08x5 FILLER_105_657 ();
 b15zdnd11an1n04x5 FILLER_105_665 ();
 b15zdnd11an1n64x5 FILLER_105_681 ();
 b15zdnd11an1n16x5 FILLER_105_745 ();
 b15zdnd11an1n08x5 FILLER_105_761 ();
 b15zdnd00an1n02x5 FILLER_105_769 ();
 b15zdnd00an1n01x5 FILLER_105_771 ();
 b15zdnd11an1n64x5 FILLER_105_785 ();
 b15zdnd11an1n08x5 FILLER_105_849 ();
 b15zdnd11an1n04x5 FILLER_105_857 ();
 b15zdnd00an1n02x5 FILLER_105_861 ();
 b15zdnd11an1n08x5 FILLER_105_875 ();
 b15zdnd11an1n04x5 FILLER_105_883 ();
 b15zdnd00an1n01x5 FILLER_105_887 ();
 b15zdnd11an1n04x5 FILLER_105_894 ();
 b15zdnd11an1n32x5 FILLER_105_903 ();
 b15zdnd11an1n16x5 FILLER_105_935 ();
 b15zdnd00an1n02x5 FILLER_105_951 ();
 b15zdnd00an1n01x5 FILLER_105_953 ();
 b15zdnd11an1n64x5 FILLER_105_959 ();
 b15zdnd11an1n08x5 FILLER_105_1023 ();
 b15zdnd00an1n02x5 FILLER_105_1031 ();
 b15zdnd11an1n32x5 FILLER_105_1053 ();
 b15zdnd11an1n16x5 FILLER_105_1085 ();
 b15zdnd11an1n04x5 FILLER_105_1101 ();
 b15zdnd11an1n32x5 FILLER_105_1125 ();
 b15zdnd11an1n16x5 FILLER_105_1157 ();
 b15zdnd11an1n08x5 FILLER_105_1173 ();
 b15zdnd00an1n02x5 FILLER_105_1181 ();
 b15zdnd11an1n32x5 FILLER_105_1188 ();
 b15zdnd11an1n08x5 FILLER_105_1220 ();
 b15zdnd00an1n02x5 FILLER_105_1228 ();
 b15zdnd11an1n08x5 FILLER_105_1248 ();
 b15zdnd00an1n01x5 FILLER_105_1256 ();
 b15zdnd11an1n64x5 FILLER_105_1267 ();
 b15zdnd11an1n04x5 FILLER_105_1336 ();
 b15zdnd11an1n16x5 FILLER_105_1353 ();
 b15zdnd11an1n04x5 FILLER_105_1369 ();
 b15zdnd00an1n02x5 FILLER_105_1373 ();
 b15zdnd11an1n32x5 FILLER_105_1390 ();
 b15zdnd11an1n08x5 FILLER_105_1422 ();
 b15zdnd11an1n04x5 FILLER_105_1430 ();
 b15zdnd00an1n02x5 FILLER_105_1434 ();
 b15zdnd11an1n08x5 FILLER_105_1441 ();
 b15zdnd11an1n04x5 FILLER_105_1449 ();
 b15zdnd00an1n02x5 FILLER_105_1453 ();
 b15zdnd00an1n01x5 FILLER_105_1455 ();
 b15zdnd11an1n64x5 FILLER_105_1460 ();
 b15zdnd11an1n04x5 FILLER_105_1524 ();
 b15zdnd00an1n02x5 FILLER_105_1528 ();
 b15zdnd11an1n08x5 FILLER_105_1542 ();
 b15zdnd11an1n04x5 FILLER_105_1550 ();
 b15zdnd00an1n02x5 FILLER_105_1554 ();
 b15zdnd00an1n01x5 FILLER_105_1556 ();
 b15zdnd11an1n04x5 FILLER_105_1580 ();
 b15zdnd00an1n01x5 FILLER_105_1584 ();
 b15zdnd11an1n64x5 FILLER_105_1593 ();
 b15zdnd11an1n64x5 FILLER_105_1657 ();
 b15zdnd11an1n32x5 FILLER_105_1721 ();
 b15zdnd11an1n04x5 FILLER_105_1760 ();
 b15zdnd11an1n04x5 FILLER_105_1771 ();
 b15zdnd00an1n02x5 FILLER_105_1775 ();
 b15zdnd11an1n16x5 FILLER_105_1783 ();
 b15zdnd11an1n08x5 FILLER_105_1799 ();
 b15zdnd11an1n04x5 FILLER_105_1813 ();
 b15zdnd00an1n01x5 FILLER_105_1817 ();
 b15zdnd11an1n64x5 FILLER_105_1826 ();
 b15zdnd11an1n16x5 FILLER_105_1890 ();
 b15zdnd11an1n08x5 FILLER_105_1906 ();
 b15zdnd11an1n04x5 FILLER_105_1914 ();
 b15zdnd00an1n01x5 FILLER_105_1918 ();
 b15zdnd11an1n16x5 FILLER_105_1926 ();
 b15zdnd11an1n04x5 FILLER_105_1942 ();
 b15zdnd00an1n01x5 FILLER_105_1946 ();
 b15zdnd11an1n04x5 FILLER_105_1954 ();
 b15zdnd11an1n08x5 FILLER_105_1970 ();
 b15zdnd11an1n04x5 FILLER_105_1978 ();
 b15zdnd00an1n02x5 FILLER_105_1982 ();
 b15zdnd00an1n01x5 FILLER_105_1984 ();
 b15zdnd11an1n16x5 FILLER_105_2002 ();
 b15zdnd11an1n32x5 FILLER_105_2023 ();
 b15zdnd11an1n08x5 FILLER_105_2055 ();
 b15zdnd11an1n04x5 FILLER_105_2063 ();
 b15zdnd00an1n02x5 FILLER_105_2067 ();
 b15zdnd11an1n64x5 FILLER_105_2083 ();
 b15zdnd11an1n04x5 FILLER_105_2147 ();
 b15zdnd00an1n02x5 FILLER_105_2151 ();
 b15zdnd00an1n01x5 FILLER_105_2153 ();
 b15zdnd11an1n04x5 FILLER_105_2167 ();
 b15zdnd11an1n04x5 FILLER_105_2184 ();
 b15zdnd11an1n32x5 FILLER_105_2192 ();
 b15zdnd11an1n08x5 FILLER_105_2224 ();
 b15zdnd00an1n01x5 FILLER_105_2232 ();
 b15zdnd11an1n16x5 FILLER_105_2237 ();
 b15zdnd11an1n08x5 FILLER_105_2253 ();
 b15zdnd11an1n04x5 FILLER_105_2261 ();
 b15zdnd00an1n02x5 FILLER_105_2265 ();
 b15zdnd11an1n08x5 FILLER_105_2271 ();
 b15zdnd11an1n04x5 FILLER_105_2279 ();
 b15zdnd00an1n01x5 FILLER_105_2283 ();
 b15zdnd11an1n64x5 FILLER_106_8 ();
 b15zdnd11an1n64x5 FILLER_106_72 ();
 b15zdnd11an1n64x5 FILLER_106_136 ();
 b15zdnd11an1n64x5 FILLER_106_200 ();
 b15zdnd11an1n64x5 FILLER_106_264 ();
 b15zdnd11an1n64x5 FILLER_106_328 ();
 b15zdnd11an1n32x5 FILLER_106_392 ();
 b15zdnd11an1n08x5 FILLER_106_424 ();
 b15zdnd00an1n02x5 FILLER_106_432 ();
 b15zdnd00an1n01x5 FILLER_106_434 ();
 b15zdnd11an1n16x5 FILLER_106_439 ();
 b15zdnd00an1n01x5 FILLER_106_455 ();
 b15zdnd11an1n04x5 FILLER_106_468 ();
 b15zdnd11an1n04x5 FILLER_106_481 ();
 b15zdnd00an1n02x5 FILLER_106_485 ();
 b15zdnd00an1n01x5 FILLER_106_487 ();
 b15zdnd11an1n16x5 FILLER_106_493 ();
 b15zdnd11an1n08x5 FILLER_106_509 ();
 b15zdnd00an1n02x5 FILLER_106_517 ();
 b15zdnd11an1n64x5 FILLER_106_529 ();
 b15zdnd11an1n04x5 FILLER_106_593 ();
 b15zdnd11an1n64x5 FILLER_106_618 ();
 b15zdnd11an1n32x5 FILLER_106_682 ();
 b15zdnd11an1n04x5 FILLER_106_714 ();
 b15zdnd00an1n02x5 FILLER_106_726 ();
 b15zdnd11an1n04x5 FILLER_106_742 ();
 b15zdnd11an1n04x5 FILLER_106_752 ();
 b15zdnd11an1n32x5 FILLER_106_769 ();
 b15zdnd11an1n16x5 FILLER_106_801 ();
 b15zdnd11an1n08x5 FILLER_106_817 ();
 b15zdnd11an1n04x5 FILLER_106_825 ();
 b15zdnd00an1n02x5 FILLER_106_829 ();
 b15zdnd00an1n01x5 FILLER_106_831 ();
 b15zdnd11an1n32x5 FILLER_106_842 ();
 b15zdnd11an1n16x5 FILLER_106_874 ();
 b15zdnd00an1n02x5 FILLER_106_890 ();
 b15zdnd00an1n01x5 FILLER_106_892 ();
 b15zdnd11an1n64x5 FILLER_106_906 ();
 b15zdnd11an1n32x5 FILLER_106_970 ();
 b15zdnd11an1n08x5 FILLER_106_1002 ();
 b15zdnd11an1n04x5 FILLER_106_1010 ();
 b15zdnd00an1n02x5 FILLER_106_1014 ();
 b15zdnd11an1n64x5 FILLER_106_1042 ();
 b15zdnd11an1n64x5 FILLER_106_1106 ();
 b15zdnd11an1n32x5 FILLER_106_1170 ();
 b15zdnd11an1n16x5 FILLER_106_1202 ();
 b15zdnd00an1n02x5 FILLER_106_1218 ();
 b15zdnd11an1n04x5 FILLER_106_1236 ();
 b15zdnd11an1n64x5 FILLER_106_1256 ();
 b15zdnd11an1n08x5 FILLER_106_1320 ();
 b15zdnd00an1n02x5 FILLER_106_1328 ();
 b15zdnd00an1n01x5 FILLER_106_1330 ();
 b15zdnd11an1n08x5 FILLER_106_1338 ();
 b15zdnd00an1n01x5 FILLER_106_1346 ();
 b15zdnd11an1n16x5 FILLER_106_1353 ();
 b15zdnd11an1n08x5 FILLER_106_1369 ();
 b15zdnd11an1n04x5 FILLER_106_1377 ();
 b15zdnd00an1n02x5 FILLER_106_1381 ();
 b15zdnd11an1n04x5 FILLER_106_1400 ();
 b15zdnd11an1n16x5 FILLER_106_1411 ();
 b15zdnd11an1n08x5 FILLER_106_1427 ();
 b15zdnd11an1n04x5 FILLER_106_1435 ();
 b15zdnd11an1n16x5 FILLER_106_1447 ();
 b15zdnd11an1n08x5 FILLER_106_1463 ();
 b15zdnd00an1n02x5 FILLER_106_1471 ();
 b15zdnd11an1n08x5 FILLER_106_1479 ();
 b15zdnd11an1n04x5 FILLER_106_1487 ();
 b15zdnd00an1n02x5 FILLER_106_1491 ();
 b15zdnd11an1n16x5 FILLER_106_1499 ();
 b15zdnd11an1n08x5 FILLER_106_1515 ();
 b15zdnd11an1n16x5 FILLER_106_1533 ();
 b15zdnd11an1n08x5 FILLER_106_1549 ();
 b15zdnd11an1n08x5 FILLER_106_1566 ();
 b15zdnd11an1n04x5 FILLER_106_1574 ();
 b15zdnd00an1n01x5 FILLER_106_1578 ();
 b15zdnd11an1n08x5 FILLER_106_1600 ();
 b15zdnd11an1n04x5 FILLER_106_1608 ();
 b15zdnd00an1n02x5 FILLER_106_1612 ();
 b15zdnd00an1n01x5 FILLER_106_1614 ();
 b15zdnd11an1n08x5 FILLER_106_1631 ();
 b15zdnd11an1n04x5 FILLER_106_1639 ();
 b15zdnd00an1n02x5 FILLER_106_1643 ();
 b15zdnd11an1n16x5 FILLER_106_1661 ();
 b15zdnd00an1n01x5 FILLER_106_1677 ();
 b15zdnd11an1n64x5 FILLER_106_1698 ();
 b15zdnd11an1n16x5 FILLER_106_1762 ();
 b15zdnd11an1n32x5 FILLER_106_1788 ();
 b15zdnd11an1n16x5 FILLER_106_1820 ();
 b15zdnd11an1n04x5 FILLER_106_1836 ();
 b15zdnd11an1n08x5 FILLER_106_1850 ();
 b15zdnd11an1n04x5 FILLER_106_1858 ();
 b15zdnd00an1n02x5 FILLER_106_1862 ();
 b15zdnd11an1n32x5 FILLER_106_1880 ();
 b15zdnd11an1n64x5 FILLER_106_1917 ();
 b15zdnd00an1n02x5 FILLER_106_1981 ();
 b15zdnd00an1n01x5 FILLER_106_1983 ();
 b15zdnd11an1n16x5 FILLER_106_1991 ();
 b15zdnd11an1n08x5 FILLER_106_2007 ();
 b15zdnd11an1n04x5 FILLER_106_2015 ();
 b15zdnd11an1n04x5 FILLER_106_2024 ();
 b15zdnd11an1n32x5 FILLER_106_2036 ();
 b15zdnd11an1n04x5 FILLER_106_2068 ();
 b15zdnd11an1n08x5 FILLER_106_2078 ();
 b15zdnd00an1n02x5 FILLER_106_2086 ();
 b15zdnd00an1n01x5 FILLER_106_2088 ();
 b15zdnd11an1n04x5 FILLER_106_2095 ();
 b15zdnd11an1n32x5 FILLER_106_2108 ();
 b15zdnd11an1n08x5 FILLER_106_2140 ();
 b15zdnd11an1n04x5 FILLER_106_2148 ();
 b15zdnd00an1n02x5 FILLER_106_2152 ();
 b15zdnd00an1n02x5 FILLER_106_2162 ();
 b15zdnd11an1n64x5 FILLER_106_2168 ();
 b15zdnd11an1n16x5 FILLER_106_2232 ();
 b15zdnd11an1n08x5 FILLER_106_2248 ();
 b15zdnd11an1n04x5 FILLER_106_2256 ();
 b15zdnd00an1n02x5 FILLER_106_2260 ();
 b15zdnd11an1n04x5 FILLER_106_2266 ();
 b15zdnd00an1n02x5 FILLER_106_2274 ();
 b15zdnd11an1n64x5 FILLER_107_0 ();
 b15zdnd11an1n64x5 FILLER_107_64 ();
 b15zdnd11an1n64x5 FILLER_107_128 ();
 b15zdnd11an1n64x5 FILLER_107_192 ();
 b15zdnd11an1n64x5 FILLER_107_256 ();
 b15zdnd11an1n64x5 FILLER_107_320 ();
 b15zdnd11an1n32x5 FILLER_107_384 ();
 b15zdnd11an1n08x5 FILLER_107_416 ();
 b15zdnd11an1n04x5 FILLER_107_424 ();
 b15zdnd11an1n04x5 FILLER_107_434 ();
 b15zdnd11an1n64x5 FILLER_107_444 ();
 b15zdnd11an1n04x5 FILLER_107_508 ();
 b15zdnd00an1n02x5 FILLER_107_512 ();
 b15zdnd11an1n04x5 FILLER_107_529 ();
 b15zdnd11an1n32x5 FILLER_107_539 ();
 b15zdnd11an1n16x5 FILLER_107_571 ();
 b15zdnd11an1n08x5 FILLER_107_587 ();
 b15zdnd11an1n04x5 FILLER_107_595 ();
 b15zdnd00an1n02x5 FILLER_107_599 ();
 b15zdnd11an1n64x5 FILLER_107_605 ();
 b15zdnd11an1n64x5 FILLER_107_669 ();
 b15zdnd11an1n64x5 FILLER_107_733 ();
 b15zdnd11an1n16x5 FILLER_107_797 ();
 b15zdnd00an1n01x5 FILLER_107_813 ();
 b15zdnd11an1n08x5 FILLER_107_820 ();
 b15zdnd11an1n04x5 FILLER_107_828 ();
 b15zdnd00an1n02x5 FILLER_107_832 ();
 b15zdnd11an1n08x5 FILLER_107_846 ();
 b15zdnd00an1n02x5 FILLER_107_854 ();
 b15zdnd11an1n16x5 FILLER_107_874 ();
 b15zdnd11an1n08x5 FILLER_107_890 ();
 b15zdnd11an1n04x5 FILLER_107_898 ();
 b15zdnd00an1n02x5 FILLER_107_902 ();
 b15zdnd00an1n01x5 FILLER_107_904 ();
 b15zdnd11an1n64x5 FILLER_107_931 ();
 b15zdnd11an1n08x5 FILLER_107_999 ();
 b15zdnd11an1n04x5 FILLER_107_1007 ();
 b15zdnd00an1n01x5 FILLER_107_1011 ();
 b15zdnd11an1n64x5 FILLER_107_1021 ();
 b15zdnd11an1n08x5 FILLER_107_1085 ();
 b15zdnd11an1n04x5 FILLER_107_1093 ();
 b15zdnd00an1n02x5 FILLER_107_1097 ();
 b15zdnd11an1n64x5 FILLER_107_1130 ();
 b15zdnd11an1n16x5 FILLER_107_1194 ();
 b15zdnd00an1n02x5 FILLER_107_1210 ();
 b15zdnd11an1n32x5 FILLER_107_1222 ();
 b15zdnd11an1n16x5 FILLER_107_1254 ();
 b15zdnd11an1n08x5 FILLER_107_1270 ();
 b15zdnd11an1n04x5 FILLER_107_1278 ();
 b15zdnd00an1n01x5 FILLER_107_1282 ();
 b15zdnd11an1n08x5 FILLER_107_1298 ();
 b15zdnd11an1n04x5 FILLER_107_1306 ();
 b15zdnd00an1n01x5 FILLER_107_1310 ();
 b15zdnd11an1n04x5 FILLER_107_1315 ();
 b15zdnd11an1n64x5 FILLER_107_1325 ();
 b15zdnd11an1n08x5 FILLER_107_1389 ();
 b15zdnd00an1n02x5 FILLER_107_1397 ();
 b15zdnd00an1n01x5 FILLER_107_1399 ();
 b15zdnd11an1n32x5 FILLER_107_1408 ();
 b15zdnd00an1n01x5 FILLER_107_1440 ();
 b15zdnd11an1n04x5 FILLER_107_1451 ();
 b15zdnd11an1n32x5 FILLER_107_1461 ();
 b15zdnd11an1n08x5 FILLER_107_1493 ();
 b15zdnd11an1n64x5 FILLER_107_1508 ();
 b15zdnd11an1n32x5 FILLER_107_1572 ();
 b15zdnd11an1n16x5 FILLER_107_1604 ();
 b15zdnd00an1n02x5 FILLER_107_1620 ();
 b15zdnd00an1n01x5 FILLER_107_1622 ();
 b15zdnd11an1n64x5 FILLER_107_1644 ();
 b15zdnd11an1n32x5 FILLER_107_1708 ();
 b15zdnd00an1n01x5 FILLER_107_1740 ();
 b15zdnd11an1n04x5 FILLER_107_1748 ();
 b15zdnd11an1n32x5 FILLER_107_1757 ();
 b15zdnd11an1n16x5 FILLER_107_1789 ();
 b15zdnd11an1n08x5 FILLER_107_1805 ();
 b15zdnd11an1n04x5 FILLER_107_1813 ();
 b15zdnd00an1n02x5 FILLER_107_1817 ();
 b15zdnd11an1n16x5 FILLER_107_1824 ();
 b15zdnd11an1n04x5 FILLER_107_1840 ();
 b15zdnd11an1n08x5 FILLER_107_1850 ();
 b15zdnd00an1n01x5 FILLER_107_1858 ();
 b15zdnd11an1n04x5 FILLER_107_1866 ();
 b15zdnd00an1n01x5 FILLER_107_1870 ();
 b15zdnd11an1n16x5 FILLER_107_1879 ();
 b15zdnd11an1n08x5 FILLER_107_1895 ();
 b15zdnd11an1n04x5 FILLER_107_1908 ();
 b15zdnd11an1n04x5 FILLER_107_1917 ();
 b15zdnd11an1n64x5 FILLER_107_1927 ();
 b15zdnd11an1n04x5 FILLER_107_1991 ();
 b15zdnd00an1n01x5 FILLER_107_1995 ();
 b15zdnd11an1n32x5 FILLER_107_2001 ();
 b15zdnd11an1n16x5 FILLER_107_2033 ();
 b15zdnd00an1n02x5 FILLER_107_2049 ();
 b15zdnd11an1n04x5 FILLER_107_2067 ();
 b15zdnd00an1n02x5 FILLER_107_2071 ();
 b15zdnd11an1n04x5 FILLER_107_2083 ();
 b15zdnd00an1n02x5 FILLER_107_2087 ();
 b15zdnd00an1n01x5 FILLER_107_2089 ();
 b15zdnd11an1n04x5 FILLER_107_2101 ();
 b15zdnd00an1n02x5 FILLER_107_2105 ();
 b15zdnd00an1n01x5 FILLER_107_2107 ();
 b15zdnd11an1n04x5 FILLER_107_2113 ();
 b15zdnd11an1n04x5 FILLER_107_2123 ();
 b15zdnd00an1n01x5 FILLER_107_2127 ();
 b15zdnd11an1n32x5 FILLER_107_2133 ();
 b15zdnd11an1n04x5 FILLER_107_2165 ();
 b15zdnd00an1n02x5 FILLER_107_2169 ();
 b15zdnd11an1n32x5 FILLER_107_2183 ();
 b15zdnd11an1n16x5 FILLER_107_2215 ();
 b15zdnd11an1n08x5 FILLER_107_2231 ();
 b15zdnd11an1n04x5 FILLER_107_2239 ();
 b15zdnd00an1n02x5 FILLER_107_2243 ();
 b15zdnd00an1n01x5 FILLER_107_2245 ();
 b15zdnd11an1n16x5 FILLER_107_2250 ();
 b15zdnd11an1n08x5 FILLER_107_2266 ();
 b15zdnd11an1n04x5 FILLER_107_2274 ();
 b15zdnd00an1n02x5 FILLER_107_2282 ();
 b15zdnd11an1n64x5 FILLER_108_8 ();
 b15zdnd11an1n64x5 FILLER_108_72 ();
 b15zdnd11an1n64x5 FILLER_108_136 ();
 b15zdnd11an1n64x5 FILLER_108_200 ();
 b15zdnd11an1n64x5 FILLER_108_264 ();
 b15zdnd11an1n64x5 FILLER_108_328 ();
 b15zdnd11an1n32x5 FILLER_108_392 ();
 b15zdnd11an1n08x5 FILLER_108_424 ();
 b15zdnd00an1n02x5 FILLER_108_432 ();
 b15zdnd00an1n01x5 FILLER_108_434 ();
 b15zdnd11an1n32x5 FILLER_108_441 ();
 b15zdnd11an1n16x5 FILLER_108_473 ();
 b15zdnd11an1n08x5 FILLER_108_489 ();
 b15zdnd11an1n04x5 FILLER_108_497 ();
 b15zdnd11an1n32x5 FILLER_108_511 ();
 b15zdnd11an1n16x5 FILLER_108_543 ();
 b15zdnd00an1n01x5 FILLER_108_559 ();
 b15zdnd11an1n64x5 FILLER_108_567 ();
 b15zdnd11an1n08x5 FILLER_108_631 ();
 b15zdnd11an1n16x5 FILLER_108_645 ();
 b15zdnd11an1n08x5 FILLER_108_661 ();
 b15zdnd11an1n04x5 FILLER_108_669 ();
 b15zdnd00an1n01x5 FILLER_108_673 ();
 b15zdnd11an1n16x5 FILLER_108_680 ();
 b15zdnd11an1n04x5 FILLER_108_696 ();
 b15zdnd00an1n02x5 FILLER_108_700 ();
 b15zdnd00an1n01x5 FILLER_108_702 ();
 b15zdnd00an1n02x5 FILLER_108_716 ();
 b15zdnd11an1n32x5 FILLER_108_726 ();
 b15zdnd00an1n01x5 FILLER_108_758 ();
 b15zdnd11an1n04x5 FILLER_108_765 ();
 b15zdnd11an1n16x5 FILLER_108_776 ();
 b15zdnd11an1n08x5 FILLER_108_792 ();
 b15zdnd00an1n01x5 FILLER_108_800 ();
 b15zdnd11an1n16x5 FILLER_108_814 ();
 b15zdnd11an1n04x5 FILLER_108_830 ();
 b15zdnd00an1n02x5 FILLER_108_834 ();
 b15zdnd00an1n01x5 FILLER_108_836 ();
 b15zdnd11an1n08x5 FILLER_108_847 ();
 b15zdnd11an1n32x5 FILLER_108_871 ();
 b15zdnd11an1n04x5 FILLER_108_903 ();
 b15zdnd00an1n02x5 FILLER_108_907 ();
 b15zdnd00an1n01x5 FILLER_108_909 ();
 b15zdnd11an1n64x5 FILLER_108_914 ();
 b15zdnd11an1n64x5 FILLER_108_978 ();
 b15zdnd11an1n64x5 FILLER_108_1042 ();
 b15zdnd11an1n32x5 FILLER_108_1106 ();
 b15zdnd11an1n08x5 FILLER_108_1138 ();
 b15zdnd11an1n32x5 FILLER_108_1166 ();
 b15zdnd11an1n04x5 FILLER_108_1198 ();
 b15zdnd00an1n02x5 FILLER_108_1202 ();
 b15zdnd00an1n01x5 FILLER_108_1204 ();
 b15zdnd11an1n32x5 FILLER_108_1212 ();
 b15zdnd11an1n04x5 FILLER_108_1244 ();
 b15zdnd11an1n08x5 FILLER_108_1257 ();
 b15zdnd11an1n04x5 FILLER_108_1265 ();
 b15zdnd11an1n04x5 FILLER_108_1273 ();
 b15zdnd11an1n04x5 FILLER_108_1282 ();
 b15zdnd11an1n64x5 FILLER_108_1318 ();
 b15zdnd11an1n16x5 FILLER_108_1382 ();
 b15zdnd11an1n08x5 FILLER_108_1398 ();
 b15zdnd11an1n64x5 FILLER_108_1412 ();
 b15zdnd00an1n01x5 FILLER_108_1476 ();
 b15zdnd11an1n64x5 FILLER_108_1486 ();
 b15zdnd11an1n64x5 FILLER_108_1550 ();
 b15zdnd11an1n08x5 FILLER_108_1614 ();
 b15zdnd00an1n02x5 FILLER_108_1622 ();
 b15zdnd00an1n01x5 FILLER_108_1624 ();
 b15zdnd11an1n08x5 FILLER_108_1629 ();
 b15zdnd11an1n04x5 FILLER_108_1637 ();
 b15zdnd11an1n04x5 FILLER_108_1673 ();
 b15zdnd00an1n01x5 FILLER_108_1677 ();
 b15zdnd11an1n32x5 FILLER_108_1687 ();
 b15zdnd11an1n16x5 FILLER_108_1719 ();
 b15zdnd11an1n04x5 FILLER_108_1735 ();
 b15zdnd11an1n32x5 FILLER_108_1749 ();
 b15zdnd11an1n08x5 FILLER_108_1781 ();
 b15zdnd11an1n16x5 FILLER_108_1794 ();
 b15zdnd00an1n02x5 FILLER_108_1810 ();
 b15zdnd00an1n01x5 FILLER_108_1812 ();
 b15zdnd11an1n32x5 FILLER_108_1822 ();
 b15zdnd11an1n04x5 FILLER_108_1854 ();
 b15zdnd00an1n02x5 FILLER_108_1858 ();
 b15zdnd00an1n01x5 FILLER_108_1860 ();
 b15zdnd11an1n64x5 FILLER_108_1866 ();
 b15zdnd11an1n04x5 FILLER_108_1930 ();
 b15zdnd11an1n16x5 FILLER_108_1941 ();
 b15zdnd11an1n08x5 FILLER_108_1957 ();
 b15zdnd11an1n04x5 FILLER_108_1965 ();
 b15zdnd00an1n02x5 FILLER_108_1969 ();
 b15zdnd00an1n01x5 FILLER_108_1971 ();
 b15zdnd11an1n08x5 FILLER_108_1982 ();
 b15zdnd00an1n02x5 FILLER_108_1990 ();
 b15zdnd00an1n01x5 FILLER_108_1992 ();
 b15zdnd11an1n64x5 FILLER_108_2002 ();
 b15zdnd11an1n32x5 FILLER_108_2066 ();
 b15zdnd11an1n16x5 FILLER_108_2098 ();
 b15zdnd11an1n04x5 FILLER_108_2114 ();
 b15zdnd00an1n02x5 FILLER_108_2118 ();
 b15zdnd00an1n01x5 FILLER_108_2120 ();
 b15zdnd11an1n04x5 FILLER_108_2130 ();
 b15zdnd11an1n08x5 FILLER_108_2142 ();
 b15zdnd11an1n04x5 FILLER_108_2150 ();
 b15zdnd11an1n16x5 FILLER_108_2162 ();
 b15zdnd11an1n08x5 FILLER_108_2178 ();
 b15zdnd00an1n02x5 FILLER_108_2186 ();
 b15zdnd11an1n16x5 FILLER_108_2209 ();
 b15zdnd11an1n08x5 FILLER_108_2225 ();
 b15zdnd00an1n02x5 FILLER_108_2233 ();
 b15zdnd00an1n01x5 FILLER_108_2235 ();
 b15zdnd11an1n32x5 FILLER_108_2241 ();
 b15zdnd00an1n02x5 FILLER_108_2273 ();
 b15zdnd00an1n01x5 FILLER_108_2275 ();
 b15zdnd11an1n64x5 FILLER_109_0 ();
 b15zdnd11an1n64x5 FILLER_109_64 ();
 b15zdnd11an1n64x5 FILLER_109_128 ();
 b15zdnd11an1n64x5 FILLER_109_192 ();
 b15zdnd11an1n64x5 FILLER_109_256 ();
 b15zdnd11an1n64x5 FILLER_109_320 ();
 b15zdnd11an1n64x5 FILLER_109_384 ();
 b15zdnd11an1n64x5 FILLER_109_448 ();
 b15zdnd11an1n16x5 FILLER_109_512 ();
 b15zdnd11an1n04x5 FILLER_109_528 ();
 b15zdnd00an1n01x5 FILLER_109_532 ();
 b15zdnd11an1n08x5 FILLER_109_537 ();
 b15zdnd11an1n04x5 FILLER_109_545 ();
 b15zdnd00an1n01x5 FILLER_109_549 ();
 b15zdnd11an1n64x5 FILLER_109_558 ();
 b15zdnd11an1n16x5 FILLER_109_622 ();
 b15zdnd11an1n08x5 FILLER_109_638 ();
 b15zdnd11an1n04x5 FILLER_109_646 ();
 b15zdnd11an1n16x5 FILLER_109_674 ();
 b15zdnd11an1n04x5 FILLER_109_690 ();
 b15zdnd11an1n64x5 FILLER_109_710 ();
 b15zdnd11an1n32x5 FILLER_109_774 ();
 b15zdnd11an1n08x5 FILLER_109_806 ();
 b15zdnd00an1n02x5 FILLER_109_814 ();
 b15zdnd11an1n32x5 FILLER_109_848 ();
 b15zdnd11an1n32x5 FILLER_109_894 ();
 b15zdnd11an1n16x5 FILLER_109_926 ();
 b15zdnd11an1n04x5 FILLER_109_942 ();
 b15zdnd11an1n64x5 FILLER_109_966 ();
 b15zdnd11an1n32x5 FILLER_109_1030 ();
 b15zdnd00an1n02x5 FILLER_109_1062 ();
 b15zdnd00an1n01x5 FILLER_109_1064 ();
 b15zdnd11an1n16x5 FILLER_109_1077 ();
 b15zdnd11an1n32x5 FILLER_109_1097 ();
 b15zdnd11an1n08x5 FILLER_109_1129 ();
 b15zdnd11an1n04x5 FILLER_109_1162 ();
 b15zdnd11an1n04x5 FILLER_109_1197 ();
 b15zdnd11an1n04x5 FILLER_109_1222 ();
 b15zdnd11an1n16x5 FILLER_109_1236 ();
 b15zdnd11an1n08x5 FILLER_109_1252 ();
 b15zdnd00an1n02x5 FILLER_109_1260 ();
 b15zdnd00an1n01x5 FILLER_109_1262 ();
 b15zdnd11an1n04x5 FILLER_109_1268 ();
 b15zdnd11an1n32x5 FILLER_109_1283 ();
 b15zdnd11an1n16x5 FILLER_109_1315 ();
 b15zdnd11an1n08x5 FILLER_109_1331 ();
 b15zdnd00an1n01x5 FILLER_109_1339 ();
 b15zdnd11an1n32x5 FILLER_109_1348 ();
 b15zdnd00an1n01x5 FILLER_109_1380 ();
 b15zdnd11an1n04x5 FILLER_109_1395 ();
 b15zdnd11an1n64x5 FILLER_109_1409 ();
 b15zdnd00an1n01x5 FILLER_109_1473 ();
 b15zdnd11an1n64x5 FILLER_109_1482 ();
 b15zdnd11an1n16x5 FILLER_109_1546 ();
 b15zdnd00an1n02x5 FILLER_109_1562 ();
 b15zdnd00an1n01x5 FILLER_109_1564 ();
 b15zdnd11an1n04x5 FILLER_109_1570 ();
 b15zdnd11an1n08x5 FILLER_109_1581 ();
 b15zdnd00an1n01x5 FILLER_109_1589 ();
 b15zdnd11an1n64x5 FILLER_109_1594 ();
 b15zdnd11an1n08x5 FILLER_109_1658 ();
 b15zdnd11an1n04x5 FILLER_109_1666 ();
 b15zdnd00an1n02x5 FILLER_109_1670 ();
 b15zdnd00an1n01x5 FILLER_109_1672 ();
 b15zdnd11an1n64x5 FILLER_109_1685 ();
 b15zdnd11an1n32x5 FILLER_109_1749 ();
 b15zdnd00an1n02x5 FILLER_109_1781 ();
 b15zdnd11an1n64x5 FILLER_109_1790 ();
 b15zdnd11an1n16x5 FILLER_109_1854 ();
 b15zdnd11an1n08x5 FILLER_109_1870 ();
 b15zdnd11an1n16x5 FILLER_109_1897 ();
 b15zdnd11an1n08x5 FILLER_109_1913 ();
 b15zdnd00an1n02x5 FILLER_109_1921 ();
 b15zdnd11an1n16x5 FILLER_109_1931 ();
 b15zdnd00an1n02x5 FILLER_109_1947 ();
 b15zdnd00an1n01x5 FILLER_109_1949 ();
 b15zdnd11an1n32x5 FILLER_109_1970 ();
 b15zdnd11an1n16x5 FILLER_109_2002 ();
 b15zdnd11an1n08x5 FILLER_109_2018 ();
 b15zdnd11an1n04x5 FILLER_109_2026 ();
 b15zdnd00an1n02x5 FILLER_109_2030 ();
 b15zdnd11an1n64x5 FILLER_109_2049 ();
 b15zdnd11an1n04x5 FILLER_109_2113 ();
 b15zdnd00an1n02x5 FILLER_109_2117 ();
 b15zdnd11an1n32x5 FILLER_109_2129 ();
 b15zdnd11an1n08x5 FILLER_109_2161 ();
 b15zdnd11an1n04x5 FILLER_109_2169 ();
 b15zdnd00an1n01x5 FILLER_109_2173 ();
 b15zdnd11an1n04x5 FILLER_109_2184 ();
 b15zdnd11an1n04x5 FILLER_109_2192 ();
 b15zdnd11an1n04x5 FILLER_109_2207 ();
 b15zdnd11an1n08x5 FILLER_109_2215 ();
 b15zdnd11an1n04x5 FILLER_109_2223 ();
 b15zdnd00an1n02x5 FILLER_109_2227 ();
 b15zdnd11an1n32x5 FILLER_109_2249 ();
 b15zdnd00an1n02x5 FILLER_109_2281 ();
 b15zdnd00an1n01x5 FILLER_109_2283 ();
 b15zdnd11an1n64x5 FILLER_110_8 ();
 b15zdnd11an1n64x5 FILLER_110_72 ();
 b15zdnd11an1n64x5 FILLER_110_136 ();
 b15zdnd11an1n64x5 FILLER_110_200 ();
 b15zdnd11an1n64x5 FILLER_110_264 ();
 b15zdnd11an1n64x5 FILLER_110_328 ();
 b15zdnd11an1n16x5 FILLER_110_392 ();
 b15zdnd11an1n08x5 FILLER_110_408 ();
 b15zdnd11an1n04x5 FILLER_110_416 ();
 b15zdnd00an1n02x5 FILLER_110_420 ();
 b15zdnd00an1n01x5 FILLER_110_422 ();
 b15zdnd11an1n32x5 FILLER_110_431 ();
 b15zdnd11an1n64x5 FILLER_110_474 ();
 b15zdnd11an1n16x5 FILLER_110_546 ();
 b15zdnd11an1n04x5 FILLER_110_566 ();
 b15zdnd11an1n04x5 FILLER_110_580 ();
 b15zdnd11an1n08x5 FILLER_110_589 ();
 b15zdnd11an1n04x5 FILLER_110_597 ();
 b15zdnd11an1n32x5 FILLER_110_613 ();
 b15zdnd00an1n01x5 FILLER_110_645 ();
 b15zdnd11an1n04x5 FILLER_110_667 ();
 b15zdnd11an1n04x5 FILLER_110_675 ();
 b15zdnd00an1n02x5 FILLER_110_679 ();
 b15zdnd00an1n01x5 FILLER_110_681 ();
 b15zdnd11an1n08x5 FILLER_110_687 ();
 b15zdnd00an1n01x5 FILLER_110_695 ();
 b15zdnd11an1n08x5 FILLER_110_709 ();
 b15zdnd00an1n01x5 FILLER_110_717 ();
 b15zdnd11an1n16x5 FILLER_110_726 ();
 b15zdnd11an1n08x5 FILLER_110_742 ();
 b15zdnd00an1n02x5 FILLER_110_750 ();
 b15zdnd00an1n01x5 FILLER_110_752 ();
 b15zdnd11an1n08x5 FILLER_110_759 ();
 b15zdnd11an1n04x5 FILLER_110_767 ();
 b15zdnd00an1n02x5 FILLER_110_771 ();
 b15zdnd11an1n32x5 FILLER_110_778 ();
 b15zdnd11an1n16x5 FILLER_110_810 ();
 b15zdnd11an1n08x5 FILLER_110_826 ();
 b15zdnd11an1n04x5 FILLER_110_834 ();
 b15zdnd00an1n01x5 FILLER_110_838 ();
 b15zdnd11an1n08x5 FILLER_110_853 ();
 b15zdnd00an1n01x5 FILLER_110_861 ();
 b15zdnd11an1n16x5 FILLER_110_876 ();
 b15zdnd11an1n08x5 FILLER_110_892 ();
 b15zdnd00an1n01x5 FILLER_110_900 ();
 b15zdnd11an1n64x5 FILLER_110_909 ();
 b15zdnd11an1n04x5 FILLER_110_973 ();
 b15zdnd00an1n02x5 FILLER_110_977 ();
 b15zdnd11an1n32x5 FILLER_110_999 ();
 b15zdnd11an1n16x5 FILLER_110_1031 ();
 b15zdnd11an1n08x5 FILLER_110_1047 ();
 b15zdnd11an1n04x5 FILLER_110_1055 ();
 b15zdnd00an1n02x5 FILLER_110_1059 ();
 b15zdnd00an1n01x5 FILLER_110_1061 ();
 b15zdnd11an1n08x5 FILLER_110_1072 ();
 b15zdnd11an1n64x5 FILLER_110_1085 ();
 b15zdnd11an1n32x5 FILLER_110_1149 ();
 b15zdnd11an1n16x5 FILLER_110_1181 ();
 b15zdnd11an1n04x5 FILLER_110_1197 ();
 b15zdnd11an1n08x5 FILLER_110_1211 ();
 b15zdnd11an1n04x5 FILLER_110_1219 ();
 b15zdnd00an1n02x5 FILLER_110_1223 ();
 b15zdnd00an1n01x5 FILLER_110_1225 ();
 b15zdnd11an1n04x5 FILLER_110_1242 ();
 b15zdnd11an1n64x5 FILLER_110_1259 ();
 b15zdnd11an1n08x5 FILLER_110_1323 ();
 b15zdnd11an1n04x5 FILLER_110_1331 ();
 b15zdnd00an1n02x5 FILLER_110_1335 ();
 b15zdnd00an1n01x5 FILLER_110_1337 ();
 b15zdnd11an1n32x5 FILLER_110_1351 ();
 b15zdnd11an1n16x5 FILLER_110_1383 ();
 b15zdnd11an1n08x5 FILLER_110_1405 ();
 b15zdnd11an1n04x5 FILLER_110_1413 ();
 b15zdnd00an1n02x5 FILLER_110_1417 ();
 b15zdnd11an1n64x5 FILLER_110_1425 ();
 b15zdnd11an1n16x5 FILLER_110_1489 ();
 b15zdnd11an1n08x5 FILLER_110_1505 ();
 b15zdnd11an1n04x5 FILLER_110_1513 ();
 b15zdnd00an1n01x5 FILLER_110_1517 ();
 b15zdnd11an1n16x5 FILLER_110_1539 ();
 b15zdnd11an1n08x5 FILLER_110_1555 ();
 b15zdnd00an1n02x5 FILLER_110_1563 ();
 b15zdnd11an1n04x5 FILLER_110_1585 ();
 b15zdnd11an1n04x5 FILLER_110_1595 ();
 b15zdnd11an1n08x5 FILLER_110_1603 ();
 b15zdnd00an1n01x5 FILLER_110_1611 ();
 b15zdnd11an1n64x5 FILLER_110_1617 ();
 b15zdnd11an1n32x5 FILLER_110_1681 ();
 b15zdnd11an1n16x5 FILLER_110_1713 ();
 b15zdnd00an1n02x5 FILLER_110_1729 ();
 b15zdnd00an1n01x5 FILLER_110_1731 ();
 b15zdnd11an1n04x5 FILLER_110_1739 ();
 b15zdnd11an1n08x5 FILLER_110_1749 ();
 b15zdnd11an1n04x5 FILLER_110_1757 ();
 b15zdnd11an1n64x5 FILLER_110_1766 ();
 b15zdnd11an1n16x5 FILLER_110_1830 ();
 b15zdnd11an1n08x5 FILLER_110_1846 ();
 b15zdnd00an1n02x5 FILLER_110_1854 ();
 b15zdnd00an1n01x5 FILLER_110_1856 ();
 b15zdnd11an1n32x5 FILLER_110_1867 ();
 b15zdnd11an1n16x5 FILLER_110_1899 ();
 b15zdnd11an1n04x5 FILLER_110_1915 ();
 b15zdnd00an1n01x5 FILLER_110_1919 ();
 b15zdnd11an1n64x5 FILLER_110_1927 ();
 b15zdnd11an1n64x5 FILLER_110_1991 ();
 b15zdnd11an1n16x5 FILLER_110_2055 ();
 b15zdnd11an1n04x5 FILLER_110_2071 ();
 b15zdnd00an1n01x5 FILLER_110_2075 ();
 b15zdnd11an1n16x5 FILLER_110_2082 ();
 b15zdnd11an1n08x5 FILLER_110_2098 ();
 b15zdnd11an1n04x5 FILLER_110_2106 ();
 b15zdnd00an1n02x5 FILLER_110_2110 ();
 b15zdnd00an1n01x5 FILLER_110_2112 ();
 b15zdnd11an1n08x5 FILLER_110_2139 ();
 b15zdnd11an1n04x5 FILLER_110_2147 ();
 b15zdnd00an1n02x5 FILLER_110_2151 ();
 b15zdnd00an1n01x5 FILLER_110_2153 ();
 b15zdnd11an1n08x5 FILLER_110_2162 ();
 b15zdnd00an1n02x5 FILLER_110_2170 ();
 b15zdnd11an1n32x5 FILLER_110_2188 ();
 b15zdnd11an1n16x5 FILLER_110_2220 ();
 b15zdnd11an1n04x5 FILLER_110_2236 ();
 b15zdnd11an1n32x5 FILLER_110_2244 ();
 b15zdnd11an1n64x5 FILLER_111_0 ();
 b15zdnd11an1n64x5 FILLER_111_64 ();
 b15zdnd11an1n64x5 FILLER_111_128 ();
 b15zdnd11an1n64x5 FILLER_111_192 ();
 b15zdnd11an1n64x5 FILLER_111_256 ();
 b15zdnd11an1n64x5 FILLER_111_320 ();
 b15zdnd11an1n32x5 FILLER_111_384 ();
 b15zdnd11an1n08x5 FILLER_111_416 ();
 b15zdnd11an1n04x5 FILLER_111_424 ();
 b15zdnd00an1n02x5 FILLER_111_428 ();
 b15zdnd00an1n01x5 FILLER_111_430 ();
 b15zdnd11an1n04x5 FILLER_111_457 ();
 b15zdnd11an1n04x5 FILLER_111_481 ();
 b15zdnd11an1n08x5 FILLER_111_511 ();
 b15zdnd11an1n04x5 FILLER_111_519 ();
 b15zdnd11an1n16x5 FILLER_111_536 ();
 b15zdnd11an1n08x5 FILLER_111_552 ();
 b15zdnd11an1n16x5 FILLER_111_568 ();
 b15zdnd11an1n04x5 FILLER_111_584 ();
 b15zdnd00an1n01x5 FILLER_111_588 ();
 b15zdnd11an1n16x5 FILLER_111_595 ();
 b15zdnd11an1n16x5 FILLER_111_616 ();
 b15zdnd11an1n08x5 FILLER_111_632 ();
 b15zdnd11an1n04x5 FILLER_111_640 ();
 b15zdnd00an1n01x5 FILLER_111_644 ();
 b15zdnd11an1n32x5 FILLER_111_657 ();
 b15zdnd11an1n16x5 FILLER_111_689 ();
 b15zdnd00an1n02x5 FILLER_111_705 ();
 b15zdnd00an1n01x5 FILLER_111_707 ();
 b15zdnd11an1n04x5 FILLER_111_712 ();
 b15zdnd11an1n04x5 FILLER_111_722 ();
 b15zdnd11an1n16x5 FILLER_111_732 ();
 b15zdnd11an1n08x5 FILLER_111_748 ();
 b15zdnd00an1n01x5 FILLER_111_756 ();
 b15zdnd11an1n04x5 FILLER_111_766 ();
 b15zdnd00an1n02x5 FILLER_111_770 ();
 b15zdnd00an1n01x5 FILLER_111_772 ();
 b15zdnd11an1n08x5 FILLER_111_781 ();
 b15zdnd00an1n01x5 FILLER_111_789 ();
 b15zdnd11an1n04x5 FILLER_111_795 ();
 b15zdnd11an1n04x5 FILLER_111_803 ();
 b15zdnd11an1n16x5 FILLER_111_817 ();
 b15zdnd00an1n02x5 FILLER_111_833 ();
 b15zdnd00an1n01x5 FILLER_111_835 ();
 b15zdnd11an1n16x5 FILLER_111_847 ();
 b15zdnd00an1n02x5 FILLER_111_863 ();
 b15zdnd11an1n16x5 FILLER_111_877 ();
 b15zdnd00an1n02x5 FILLER_111_893 ();
 b15zdnd00an1n01x5 FILLER_111_895 ();
 b15zdnd11an1n64x5 FILLER_111_903 ();
 b15zdnd11an1n64x5 FILLER_111_967 ();
 b15zdnd11an1n32x5 FILLER_111_1031 ();
 b15zdnd11an1n08x5 FILLER_111_1068 ();
 b15zdnd00an1n01x5 FILLER_111_1076 ();
 b15zdnd11an1n32x5 FILLER_111_1097 ();
 b15zdnd11an1n08x5 FILLER_111_1129 ();
 b15zdnd00an1n02x5 FILLER_111_1137 ();
 b15zdnd11an1n64x5 FILLER_111_1143 ();
 b15zdnd00an1n01x5 FILLER_111_1207 ();
 b15zdnd11an1n64x5 FILLER_111_1218 ();
 b15zdnd11an1n16x5 FILLER_111_1282 ();
 b15zdnd11an1n08x5 FILLER_111_1298 ();
 b15zdnd00an1n02x5 FILLER_111_1306 ();
 b15zdnd00an1n01x5 FILLER_111_1308 ();
 b15zdnd11an1n16x5 FILLER_111_1316 ();
 b15zdnd00an1n01x5 FILLER_111_1332 ();
 b15zdnd11an1n16x5 FILLER_111_1353 ();
 b15zdnd11an1n08x5 FILLER_111_1369 ();
 b15zdnd00an1n01x5 FILLER_111_1377 ();
 b15zdnd11an1n08x5 FILLER_111_1383 ();
 b15zdnd11an1n04x5 FILLER_111_1391 ();
 b15zdnd00an1n01x5 FILLER_111_1395 ();
 b15zdnd11an1n32x5 FILLER_111_1401 ();
 b15zdnd11an1n08x5 FILLER_111_1433 ();
 b15zdnd11an1n04x5 FILLER_111_1441 ();
 b15zdnd00an1n01x5 FILLER_111_1445 ();
 b15zdnd11an1n04x5 FILLER_111_1458 ();
 b15zdnd00an1n02x5 FILLER_111_1462 ();
 b15zdnd11an1n04x5 FILLER_111_1489 ();
 b15zdnd00an1n01x5 FILLER_111_1493 ();
 b15zdnd11an1n04x5 FILLER_111_1504 ();
 b15zdnd11an1n32x5 FILLER_111_1513 ();
 b15zdnd11an1n04x5 FILLER_111_1545 ();
 b15zdnd11an1n32x5 FILLER_111_1556 ();
 b15zdnd11an1n16x5 FILLER_111_1588 ();
 b15zdnd11an1n08x5 FILLER_111_1604 ();
 b15zdnd00an1n02x5 FILLER_111_1612 ();
 b15zdnd11an1n64x5 FILLER_111_1619 ();
 b15zdnd11an1n64x5 FILLER_111_1683 ();
 b15zdnd11an1n08x5 FILLER_111_1747 ();
 b15zdnd11an1n04x5 FILLER_111_1755 ();
 b15zdnd00an1n02x5 FILLER_111_1759 ();
 b15zdnd11an1n32x5 FILLER_111_1767 ();
 b15zdnd00an1n02x5 FILLER_111_1799 ();
 b15zdnd00an1n01x5 FILLER_111_1801 ();
 b15zdnd11an1n04x5 FILLER_111_1817 ();
 b15zdnd11an1n04x5 FILLER_111_1827 ();
 b15zdnd11an1n08x5 FILLER_111_1837 ();
 b15zdnd11an1n04x5 FILLER_111_1845 ();
 b15zdnd00an1n02x5 FILLER_111_1849 ();
 b15zdnd00an1n01x5 FILLER_111_1851 ();
 b15zdnd11an1n64x5 FILLER_111_1876 ();
 b15zdnd11an1n32x5 FILLER_111_1940 ();
 b15zdnd11an1n16x5 FILLER_111_1972 ();
 b15zdnd11an1n04x5 FILLER_111_1988 ();
 b15zdnd00an1n01x5 FILLER_111_1992 ();
 b15zdnd11an1n08x5 FILLER_111_2001 ();
 b15zdnd11an1n04x5 FILLER_111_2009 ();
 b15zdnd00an1n02x5 FILLER_111_2013 ();
 b15zdnd00an1n01x5 FILLER_111_2015 ();
 b15zdnd11an1n16x5 FILLER_111_2022 ();
 b15zdnd11an1n04x5 FILLER_111_2038 ();
 b15zdnd00an1n02x5 FILLER_111_2042 ();
 b15zdnd00an1n01x5 FILLER_111_2044 ();
 b15zdnd11an1n04x5 FILLER_111_2061 ();
 b15zdnd11an1n04x5 FILLER_111_2070 ();
 b15zdnd00an1n01x5 FILLER_111_2074 ();
 b15zdnd11an1n16x5 FILLER_111_2087 ();
 b15zdnd00an1n02x5 FILLER_111_2103 ();
 b15zdnd11an1n32x5 FILLER_111_2110 ();
 b15zdnd00an1n02x5 FILLER_111_2142 ();
 b15zdnd00an1n01x5 FILLER_111_2144 ();
 b15zdnd11an1n64x5 FILLER_111_2157 ();
 b15zdnd11an1n32x5 FILLER_111_2221 ();
 b15zdnd00an1n01x5 FILLER_111_2253 ();
 b15zdnd11an1n16x5 FILLER_111_2258 ();
 b15zdnd11an1n08x5 FILLER_111_2274 ();
 b15zdnd00an1n02x5 FILLER_111_2282 ();
 b15zdnd11an1n64x5 FILLER_112_8 ();
 b15zdnd11an1n64x5 FILLER_112_72 ();
 b15zdnd11an1n64x5 FILLER_112_136 ();
 b15zdnd11an1n64x5 FILLER_112_200 ();
 b15zdnd11an1n64x5 FILLER_112_264 ();
 b15zdnd11an1n64x5 FILLER_112_328 ();
 b15zdnd11an1n32x5 FILLER_112_392 ();
 b15zdnd11an1n08x5 FILLER_112_424 ();
 b15zdnd11an1n16x5 FILLER_112_447 ();
 b15zdnd11an1n04x5 FILLER_112_463 ();
 b15zdnd00an1n01x5 FILLER_112_467 ();
 b15zdnd11an1n16x5 FILLER_112_481 ();
 b15zdnd11an1n08x5 FILLER_112_504 ();
 b15zdnd00an1n02x5 FILLER_112_512 ();
 b15zdnd00an1n01x5 FILLER_112_514 ();
 b15zdnd11an1n04x5 FILLER_112_525 ();
 b15zdnd11an1n32x5 FILLER_112_535 ();
 b15zdnd11an1n16x5 FILLER_112_567 ();
 b15zdnd00an1n02x5 FILLER_112_583 ();
 b15zdnd00an1n01x5 FILLER_112_585 ();
 b15zdnd11an1n16x5 FILLER_112_592 ();
 b15zdnd00an1n02x5 FILLER_112_608 ();
 b15zdnd00an1n01x5 FILLER_112_610 ();
 b15zdnd11an1n64x5 FILLER_112_616 ();
 b15zdnd11an1n08x5 FILLER_112_680 ();
 b15zdnd00an1n02x5 FILLER_112_688 ();
 b15zdnd00an1n02x5 FILLER_112_716 ();
 b15zdnd11an1n32x5 FILLER_112_726 ();
 b15zdnd11an1n08x5 FILLER_112_758 ();
 b15zdnd11an1n04x5 FILLER_112_766 ();
 b15zdnd00an1n01x5 FILLER_112_770 ();
 b15zdnd11an1n16x5 FILLER_112_783 ();
 b15zdnd11an1n08x5 FILLER_112_799 ();
 b15zdnd00an1n02x5 FILLER_112_807 ();
 b15zdnd00an1n01x5 FILLER_112_809 ();
 b15zdnd11an1n08x5 FILLER_112_836 ();
 b15zdnd11an1n64x5 FILLER_112_849 ();
 b15zdnd11an1n04x5 FILLER_112_913 ();
 b15zdnd11an1n04x5 FILLER_112_930 ();
 b15zdnd11an1n04x5 FILLER_112_939 ();
 b15zdnd11an1n64x5 FILLER_112_955 ();
 b15zdnd11an1n16x5 FILLER_112_1019 ();
 b15zdnd11an1n32x5 FILLER_112_1055 ();
 b15zdnd00an1n02x5 FILLER_112_1087 ();
 b15zdnd11an1n16x5 FILLER_112_1092 ();
 b15zdnd11an1n08x5 FILLER_112_1108 ();
 b15zdnd11an1n04x5 FILLER_112_1116 ();
 b15zdnd00an1n02x5 FILLER_112_1120 ();
 b15zdnd00an1n01x5 FILLER_112_1122 ();
 b15zdnd11an1n64x5 FILLER_112_1128 ();
 b15zdnd11an1n08x5 FILLER_112_1192 ();
 b15zdnd11an1n04x5 FILLER_112_1200 ();
 b15zdnd00an1n02x5 FILLER_112_1204 ();
 b15zdnd00an1n01x5 FILLER_112_1206 ();
 b15zdnd11an1n16x5 FILLER_112_1222 ();
 b15zdnd11an1n08x5 FILLER_112_1238 ();
 b15zdnd00an1n01x5 FILLER_112_1246 ();
 b15zdnd11an1n16x5 FILLER_112_1256 ();
 b15zdnd11an1n08x5 FILLER_112_1272 ();
 b15zdnd11an1n04x5 FILLER_112_1280 ();
 b15zdnd00an1n02x5 FILLER_112_1284 ();
 b15zdnd00an1n01x5 FILLER_112_1286 ();
 b15zdnd11an1n04x5 FILLER_112_1293 ();
 b15zdnd11an1n16x5 FILLER_112_1310 ();
 b15zdnd11an1n32x5 FILLER_112_1344 ();
 b15zdnd11an1n04x5 FILLER_112_1376 ();
 b15zdnd11an1n64x5 FILLER_112_1385 ();
 b15zdnd00an1n02x5 FILLER_112_1449 ();
 b15zdnd00an1n01x5 FILLER_112_1451 ();
 b15zdnd11an1n04x5 FILLER_112_1468 ();
 b15zdnd00an1n02x5 FILLER_112_1472 ();
 b15zdnd00an1n01x5 FILLER_112_1474 ();
 b15zdnd11an1n16x5 FILLER_112_1479 ();
 b15zdnd11an1n04x5 FILLER_112_1495 ();
 b15zdnd11an1n32x5 FILLER_112_1520 ();
 b15zdnd00an1n01x5 FILLER_112_1552 ();
 b15zdnd11an1n16x5 FILLER_112_1558 ();
 b15zdnd00an1n02x5 FILLER_112_1574 ();
 b15zdnd11an1n04x5 FILLER_112_1588 ();
 b15zdnd00an1n01x5 FILLER_112_1592 ();
 b15zdnd11an1n64x5 FILLER_112_1598 ();
 b15zdnd11an1n64x5 FILLER_112_1662 ();
 b15zdnd11an1n08x5 FILLER_112_1726 ();
 b15zdnd00an1n01x5 FILLER_112_1734 ();
 b15zdnd11an1n32x5 FILLER_112_1741 ();
 b15zdnd11an1n04x5 FILLER_112_1773 ();
 b15zdnd00an1n02x5 FILLER_112_1777 ();
 b15zdnd00an1n01x5 FILLER_112_1779 ();
 b15zdnd11an1n04x5 FILLER_112_1787 ();
 b15zdnd11an1n16x5 FILLER_112_1796 ();
 b15zdnd11an1n04x5 FILLER_112_1812 ();
 b15zdnd00an1n01x5 FILLER_112_1816 ();
 b15zdnd11an1n04x5 FILLER_112_1823 ();
 b15zdnd11an1n16x5 FILLER_112_1833 ();
 b15zdnd11an1n08x5 FILLER_112_1849 ();
 b15zdnd11an1n04x5 FILLER_112_1857 ();
 b15zdnd00an1n02x5 FILLER_112_1861 ();
 b15zdnd11an1n16x5 FILLER_112_1874 ();
 b15zdnd11an1n04x5 FILLER_112_1890 ();
 b15zdnd00an1n01x5 FILLER_112_1894 ();
 b15zdnd11an1n16x5 FILLER_112_1907 ();
 b15zdnd11an1n04x5 FILLER_112_1923 ();
 b15zdnd11an1n04x5 FILLER_112_1931 ();
 b15zdnd00an1n02x5 FILLER_112_1935 ();
 b15zdnd11an1n08x5 FILLER_112_1946 ();
 b15zdnd11an1n04x5 FILLER_112_1954 ();
 b15zdnd00an1n02x5 FILLER_112_1958 ();
 b15zdnd00an1n01x5 FILLER_112_1960 ();
 b15zdnd11an1n32x5 FILLER_112_1967 ();
 b15zdnd11an1n08x5 FILLER_112_1999 ();
 b15zdnd00an1n02x5 FILLER_112_2007 ();
 b15zdnd11an1n32x5 FILLER_112_2040 ();
 b15zdnd11an1n16x5 FILLER_112_2072 ();
 b15zdnd00an1n01x5 FILLER_112_2088 ();
 b15zdnd11an1n04x5 FILLER_112_2095 ();
 b15zdnd00an1n01x5 FILLER_112_2099 ();
 b15zdnd11an1n04x5 FILLER_112_2115 ();
 b15zdnd11an1n08x5 FILLER_112_2139 ();
 b15zdnd11an1n04x5 FILLER_112_2147 ();
 b15zdnd00an1n02x5 FILLER_112_2151 ();
 b15zdnd00an1n01x5 FILLER_112_2153 ();
 b15zdnd11an1n04x5 FILLER_112_2162 ();
 b15zdnd00an1n02x5 FILLER_112_2166 ();
 b15zdnd11an1n64x5 FILLER_112_2180 ();
 b15zdnd11an1n08x5 FILLER_112_2244 ();
 b15zdnd11an1n08x5 FILLER_112_2261 ();
 b15zdnd11an1n04x5 FILLER_112_2269 ();
 b15zdnd00an1n02x5 FILLER_112_2273 ();
 b15zdnd00an1n01x5 FILLER_112_2275 ();
 b15zdnd11an1n64x5 FILLER_113_0 ();
 b15zdnd11an1n64x5 FILLER_113_64 ();
 b15zdnd11an1n16x5 FILLER_113_128 ();
 b15zdnd11an1n08x5 FILLER_113_144 ();
 b15zdnd11an1n04x5 FILLER_113_152 ();
 b15zdnd00an1n01x5 FILLER_113_156 ();
 b15zdnd11an1n64x5 FILLER_113_166 ();
 b15zdnd11an1n16x5 FILLER_113_230 ();
 b15zdnd11an1n04x5 FILLER_113_246 ();
 b15zdnd00an1n01x5 FILLER_113_250 ();
 b15zdnd11an1n16x5 FILLER_113_267 ();
 b15zdnd11an1n08x5 FILLER_113_283 ();
 b15zdnd00an1n02x5 FILLER_113_291 ();
 b15zdnd00an1n01x5 FILLER_113_293 ();
 b15zdnd11an1n64x5 FILLER_113_298 ();
 b15zdnd11an1n64x5 FILLER_113_362 ();
 b15zdnd11an1n32x5 FILLER_113_426 ();
 b15zdnd11an1n04x5 FILLER_113_458 ();
 b15zdnd00an1n01x5 FILLER_113_462 ();
 b15zdnd11an1n32x5 FILLER_113_470 ();
 b15zdnd00an1n02x5 FILLER_113_502 ();
 b15zdnd11an1n08x5 FILLER_113_512 ();
 b15zdnd11an1n04x5 FILLER_113_520 ();
 b15zdnd00an1n01x5 FILLER_113_524 ();
 b15zdnd11an1n64x5 FILLER_113_530 ();
 b15zdnd11an1n16x5 FILLER_113_594 ();
 b15zdnd11an1n08x5 FILLER_113_610 ();
 b15zdnd00an1n01x5 FILLER_113_618 ();
 b15zdnd11an1n64x5 FILLER_113_635 ();
 b15zdnd11an1n32x5 FILLER_113_699 ();
 b15zdnd11an1n16x5 FILLER_113_731 ();
 b15zdnd00an1n02x5 FILLER_113_747 ();
 b15zdnd00an1n01x5 FILLER_113_749 ();
 b15zdnd11an1n08x5 FILLER_113_754 ();
 b15zdnd00an1n02x5 FILLER_113_762 ();
 b15zdnd00an1n01x5 FILLER_113_764 ();
 b15zdnd11an1n32x5 FILLER_113_777 ();
 b15zdnd11an1n04x5 FILLER_113_809 ();
 b15zdnd00an1n02x5 FILLER_113_813 ();
 b15zdnd11an1n64x5 FILLER_113_825 ();
 b15zdnd11an1n64x5 FILLER_113_889 ();
 b15zdnd11an1n64x5 FILLER_113_953 ();
 b15zdnd11an1n08x5 FILLER_113_1017 ();
 b15zdnd00an1n02x5 FILLER_113_1025 ();
 b15zdnd00an1n01x5 FILLER_113_1027 ();
 b15zdnd11an1n64x5 FILLER_113_1054 ();
 b15zdnd11an1n04x5 FILLER_113_1118 ();
 b15zdnd00an1n02x5 FILLER_113_1122 ();
 b15zdnd11an1n32x5 FILLER_113_1144 ();
 b15zdnd11an1n16x5 FILLER_113_1176 ();
 b15zdnd11an1n04x5 FILLER_113_1192 ();
 b15zdnd11an1n32x5 FILLER_113_1209 ();
 b15zdnd11an1n08x5 FILLER_113_1241 ();
 b15zdnd11an1n04x5 FILLER_113_1249 ();
 b15zdnd00an1n01x5 FILLER_113_1253 ();
 b15zdnd11an1n16x5 FILLER_113_1261 ();
 b15zdnd11an1n08x5 FILLER_113_1277 ();
 b15zdnd11an1n04x5 FILLER_113_1285 ();
 b15zdnd11an1n04x5 FILLER_113_1295 ();
 b15zdnd11an1n16x5 FILLER_113_1307 ();
 b15zdnd11an1n08x5 FILLER_113_1323 ();
 b15zdnd00an1n01x5 FILLER_113_1331 ();
 b15zdnd11an1n64x5 FILLER_113_1341 ();
 b15zdnd11an1n08x5 FILLER_113_1405 ();
 b15zdnd11an1n04x5 FILLER_113_1413 ();
 b15zdnd00an1n01x5 FILLER_113_1417 ();
 b15zdnd11an1n08x5 FILLER_113_1431 ();
 b15zdnd11an1n04x5 FILLER_113_1439 ();
 b15zdnd00an1n01x5 FILLER_113_1443 ();
 b15zdnd11an1n04x5 FILLER_113_1459 ();
 b15zdnd11an1n04x5 FILLER_113_1469 ();
 b15zdnd11an1n16x5 FILLER_113_1488 ();
 b15zdnd11an1n04x5 FILLER_113_1520 ();
 b15zdnd11an1n64x5 FILLER_113_1540 ();
 b15zdnd11an1n08x5 FILLER_113_1604 ();
 b15zdnd11an1n16x5 FILLER_113_1628 ();
 b15zdnd11an1n08x5 FILLER_113_1644 ();
 b15zdnd11an1n64x5 FILLER_113_1656 ();
 b15zdnd11an1n64x5 FILLER_113_1720 ();
 b15zdnd11an1n04x5 FILLER_113_1784 ();
 b15zdnd00an1n02x5 FILLER_113_1788 ();
 b15zdnd11an1n04x5 FILLER_113_1799 ();
 b15zdnd11an1n64x5 FILLER_113_1812 ();
 b15zdnd11an1n16x5 FILLER_113_1876 ();
 b15zdnd11an1n04x5 FILLER_113_1892 ();
 b15zdnd00an1n02x5 FILLER_113_1896 ();
 b15zdnd00an1n01x5 FILLER_113_1898 ();
 b15zdnd11an1n16x5 FILLER_113_1912 ();
 b15zdnd11an1n08x5 FILLER_113_1928 ();
 b15zdnd00an1n02x5 FILLER_113_1936 ();
 b15zdnd11an1n04x5 FILLER_113_1951 ();
 b15zdnd00an1n02x5 FILLER_113_1955 ();
 b15zdnd00an1n01x5 FILLER_113_1957 ();
 b15zdnd11an1n16x5 FILLER_113_1968 ();
 b15zdnd00an1n01x5 FILLER_113_1984 ();
 b15zdnd11an1n04x5 FILLER_113_1989 ();
 b15zdnd11an1n32x5 FILLER_113_2005 ();
 b15zdnd11an1n08x5 FILLER_113_2037 ();
 b15zdnd11an1n32x5 FILLER_113_2050 ();
 b15zdnd00an1n02x5 FILLER_113_2082 ();
 b15zdnd11an1n64x5 FILLER_113_2094 ();
 b15zdnd00an1n01x5 FILLER_113_2158 ();
 b15zdnd11an1n04x5 FILLER_113_2179 ();
 b15zdnd11an1n16x5 FILLER_113_2207 ();
 b15zdnd00an1n02x5 FILLER_113_2223 ();
 b15zdnd00an1n01x5 FILLER_113_2225 ();
 b15zdnd11an1n04x5 FILLER_113_2246 ();
 b15zdnd00an1n02x5 FILLER_113_2282 ();
 b15zdnd11an1n64x5 FILLER_114_8 ();
 b15zdnd11an1n08x5 FILLER_114_72 ();
 b15zdnd11an1n16x5 FILLER_114_87 ();
 b15zdnd11an1n08x5 FILLER_114_103 ();
 b15zdnd11an1n04x5 FILLER_114_125 ();
 b15zdnd00an1n02x5 FILLER_114_129 ();
 b15zdnd11an1n08x5 FILLER_114_149 ();
 b15zdnd11an1n04x5 FILLER_114_157 ();
 b15zdnd11an1n16x5 FILLER_114_173 ();
 b15zdnd11an1n04x5 FILLER_114_189 ();
 b15zdnd00an1n01x5 FILLER_114_193 ();
 b15zdnd11an1n16x5 FILLER_114_204 ();
 b15zdnd11an1n08x5 FILLER_114_220 ();
 b15zdnd00an1n02x5 FILLER_114_228 ();
 b15zdnd00an1n01x5 FILLER_114_230 ();
 b15zdnd11an1n04x5 FILLER_114_237 ();
 b15zdnd00an1n01x5 FILLER_114_241 ();
 b15zdnd11an1n04x5 FILLER_114_247 ();
 b15zdnd11an1n04x5 FILLER_114_267 ();
 b15zdnd11an1n64x5 FILLER_114_278 ();
 b15zdnd11an1n64x5 FILLER_114_342 ();
 b15zdnd11an1n64x5 FILLER_114_406 ();
 b15zdnd11an1n32x5 FILLER_114_470 ();
 b15zdnd11an1n16x5 FILLER_114_502 ();
 b15zdnd11an1n08x5 FILLER_114_518 ();
 b15zdnd11an1n04x5 FILLER_114_526 ();
 b15zdnd11an1n16x5 FILLER_114_540 ();
 b15zdnd00an1n02x5 FILLER_114_556 ();
 b15zdnd00an1n01x5 FILLER_114_558 ();
 b15zdnd11an1n32x5 FILLER_114_570 ();
 b15zdnd11an1n16x5 FILLER_114_602 ();
 b15zdnd00an1n01x5 FILLER_114_618 ();
 b15zdnd11an1n32x5 FILLER_114_628 ();
 b15zdnd11an1n16x5 FILLER_114_660 ();
 b15zdnd11an1n08x5 FILLER_114_676 ();
 b15zdnd00an1n02x5 FILLER_114_684 ();
 b15zdnd00an1n01x5 FILLER_114_686 ();
 b15zdnd11an1n04x5 FILLER_114_691 ();
 b15zdnd11an1n08x5 FILLER_114_705 ();
 b15zdnd11an1n04x5 FILLER_114_713 ();
 b15zdnd00an1n01x5 FILLER_114_717 ();
 b15zdnd11an1n04x5 FILLER_114_726 ();
 b15zdnd00an1n02x5 FILLER_114_730 ();
 b15zdnd11an1n64x5 FILLER_114_742 ();
 b15zdnd11an1n32x5 FILLER_114_806 ();
 b15zdnd11an1n04x5 FILLER_114_838 ();
 b15zdnd11an1n16x5 FILLER_114_867 ();
 b15zdnd11an1n08x5 FILLER_114_883 ();
 b15zdnd11an1n04x5 FILLER_114_891 ();
 b15zdnd00an1n01x5 FILLER_114_895 ();
 b15zdnd11an1n08x5 FILLER_114_905 ();
 b15zdnd00an1n01x5 FILLER_114_913 ();
 b15zdnd11an1n32x5 FILLER_114_924 ();
 b15zdnd11an1n16x5 FILLER_114_956 ();
 b15zdnd11an1n08x5 FILLER_114_972 ();
 b15zdnd00an1n01x5 FILLER_114_980 ();
 b15zdnd11an1n32x5 FILLER_114_1001 ();
 b15zdnd11an1n16x5 FILLER_114_1033 ();
 b15zdnd11an1n08x5 FILLER_114_1049 ();
 b15zdnd11an1n04x5 FILLER_114_1057 ();
 b15zdnd00an1n02x5 FILLER_114_1061 ();
 b15zdnd00an1n01x5 FILLER_114_1063 ();
 b15zdnd11an1n64x5 FILLER_114_1095 ();
 b15zdnd11an1n08x5 FILLER_114_1159 ();
 b15zdnd11an1n04x5 FILLER_114_1167 ();
 b15zdnd00an1n01x5 FILLER_114_1171 ();
 b15zdnd11an1n32x5 FILLER_114_1183 ();
 b15zdnd11an1n04x5 FILLER_114_1215 ();
 b15zdnd11an1n04x5 FILLER_114_1226 ();
 b15zdnd11an1n16x5 FILLER_114_1239 ();
 b15zdnd11an1n04x5 FILLER_114_1255 ();
 b15zdnd00an1n02x5 FILLER_114_1259 ();
 b15zdnd00an1n01x5 FILLER_114_1261 ();
 b15zdnd11an1n04x5 FILLER_114_1283 ();
 b15zdnd00an1n02x5 FILLER_114_1287 ();
 b15zdnd00an1n01x5 FILLER_114_1289 ();
 b15zdnd11an1n64x5 FILLER_114_1299 ();
 b15zdnd11an1n08x5 FILLER_114_1363 ();
 b15zdnd11an1n04x5 FILLER_114_1371 ();
 b15zdnd00an1n02x5 FILLER_114_1375 ();
 b15zdnd11an1n04x5 FILLER_114_1389 ();
 b15zdnd11an1n16x5 FILLER_114_1399 ();
 b15zdnd11an1n08x5 FILLER_114_1415 ();
 b15zdnd11an1n64x5 FILLER_114_1433 ();
 b15zdnd11an1n16x5 FILLER_114_1497 ();
 b15zdnd11an1n08x5 FILLER_114_1513 ();
 b15zdnd11an1n04x5 FILLER_114_1521 ();
 b15zdnd00an1n02x5 FILLER_114_1525 ();
 b15zdnd11an1n16x5 FILLER_114_1532 ();
 b15zdnd00an1n02x5 FILLER_114_1548 ();
 b15zdnd11an1n64x5 FILLER_114_1555 ();
 b15zdnd11an1n08x5 FILLER_114_1619 ();
 b15zdnd00an1n02x5 FILLER_114_1627 ();
 b15zdnd11an1n16x5 FILLER_114_1649 ();
 b15zdnd11an1n08x5 FILLER_114_1665 ();
 b15zdnd11an1n64x5 FILLER_114_1693 ();
 b15zdnd11an1n32x5 FILLER_114_1757 ();
 b15zdnd11an1n16x5 FILLER_114_1789 ();
 b15zdnd11an1n64x5 FILLER_114_1810 ();
 b15zdnd11an1n64x5 FILLER_114_1874 ();
 b15zdnd11an1n16x5 FILLER_114_1938 ();
 b15zdnd11an1n16x5 FILLER_114_1968 ();
 b15zdnd00an1n02x5 FILLER_114_1984 ();
 b15zdnd00an1n01x5 FILLER_114_1986 ();
 b15zdnd11an1n16x5 FILLER_114_1996 ();
 b15zdnd00an1n02x5 FILLER_114_2012 ();
 b15zdnd11an1n64x5 FILLER_114_2024 ();
 b15zdnd11an1n64x5 FILLER_114_2088 ();
 b15zdnd00an1n02x5 FILLER_114_2152 ();
 b15zdnd11an1n64x5 FILLER_114_2162 ();
 b15zdnd00an1n02x5 FILLER_114_2226 ();
 b15zdnd00an1n01x5 FILLER_114_2228 ();
 b15zdnd11an1n08x5 FILLER_114_2249 ();
 b15zdnd11an1n04x5 FILLER_114_2257 ();
 b15zdnd11an1n08x5 FILLER_114_2265 ();
 b15zdnd00an1n02x5 FILLER_114_2273 ();
 b15zdnd00an1n01x5 FILLER_114_2275 ();
 b15zdnd11an1n32x5 FILLER_115_0 ();
 b15zdnd11an1n16x5 FILLER_115_32 ();
 b15zdnd11an1n08x5 FILLER_115_48 ();
 b15zdnd11an1n04x5 FILLER_115_63 ();
 b15zdnd11an1n08x5 FILLER_115_74 ();
 b15zdnd00an1n01x5 FILLER_115_82 ();
 b15zdnd11an1n04x5 FILLER_115_91 ();
 b15zdnd00an1n02x5 FILLER_115_95 ();
 b15zdnd00an1n01x5 FILLER_115_97 ();
 b15zdnd11an1n08x5 FILLER_115_114 ();
 b15zdnd00an1n02x5 FILLER_115_122 ();
 b15zdnd11an1n16x5 FILLER_115_144 ();
 b15zdnd11an1n04x5 FILLER_115_160 ();
 b15zdnd00an1n01x5 FILLER_115_164 ();
 b15zdnd11an1n08x5 FILLER_115_169 ();
 b15zdnd11an1n04x5 FILLER_115_177 ();
 b15zdnd11an1n08x5 FILLER_115_192 ();
 b15zdnd11an1n04x5 FILLER_115_205 ();
 b15zdnd11an1n08x5 FILLER_115_223 ();
 b15zdnd00an1n01x5 FILLER_115_231 ();
 b15zdnd11an1n04x5 FILLER_115_236 ();
 b15zdnd11an1n08x5 FILLER_115_250 ();
 b15zdnd11an1n04x5 FILLER_115_258 ();
 b15zdnd00an1n02x5 FILLER_115_262 ();
 b15zdnd00an1n01x5 FILLER_115_264 ();
 b15zdnd11an1n16x5 FILLER_115_291 ();
 b15zdnd11an1n08x5 FILLER_115_307 ();
 b15zdnd00an1n02x5 FILLER_115_315 ();
 b15zdnd11an1n08x5 FILLER_115_334 ();
 b15zdnd11an1n64x5 FILLER_115_354 ();
 b15zdnd11an1n64x5 FILLER_115_418 ();
 b15zdnd11an1n64x5 FILLER_115_482 ();
 b15zdnd11an1n32x5 FILLER_115_546 ();
 b15zdnd11an1n16x5 FILLER_115_578 ();
 b15zdnd00an1n02x5 FILLER_115_594 ();
 b15zdnd00an1n01x5 FILLER_115_596 ();
 b15zdnd11an1n04x5 FILLER_115_603 ();
 b15zdnd11an1n32x5 FILLER_115_612 ();
 b15zdnd00an1n02x5 FILLER_115_644 ();
 b15zdnd00an1n01x5 FILLER_115_646 ();
 b15zdnd11an1n04x5 FILLER_115_655 ();
 b15zdnd11an1n16x5 FILLER_115_663 ();
 b15zdnd00an1n02x5 FILLER_115_679 ();
 b15zdnd00an1n01x5 FILLER_115_681 ();
 b15zdnd11an1n16x5 FILLER_115_694 ();
 b15zdnd11an1n08x5 FILLER_115_710 ();
 b15zdnd11an1n04x5 FILLER_115_718 ();
 b15zdnd00an1n01x5 FILLER_115_722 ();
 b15zdnd11an1n64x5 FILLER_115_739 ();
 b15zdnd11an1n32x5 FILLER_115_803 ();
 b15zdnd11an1n08x5 FILLER_115_835 ();
 b15zdnd11an1n04x5 FILLER_115_843 ();
 b15zdnd00an1n02x5 FILLER_115_847 ();
 b15zdnd00an1n01x5 FILLER_115_849 ();
 b15zdnd11an1n16x5 FILLER_115_860 ();
 b15zdnd11an1n04x5 FILLER_115_876 ();
 b15zdnd00an1n02x5 FILLER_115_880 ();
 b15zdnd00an1n01x5 FILLER_115_882 ();
 b15zdnd11an1n04x5 FILLER_115_888 ();
 b15zdnd11an1n08x5 FILLER_115_898 ();
 b15zdnd00an1n01x5 FILLER_115_906 ();
 b15zdnd11an1n04x5 FILLER_115_921 ();
 b15zdnd11an1n64x5 FILLER_115_932 ();
 b15zdnd11an1n16x5 FILLER_115_996 ();
 b15zdnd11an1n08x5 FILLER_115_1012 ();
 b15zdnd11an1n04x5 FILLER_115_1040 ();
 b15zdnd11an1n04x5 FILLER_115_1054 ();
 b15zdnd00an1n01x5 FILLER_115_1058 ();
 b15zdnd11an1n64x5 FILLER_115_1063 ();
 b15zdnd11an1n64x5 FILLER_115_1127 ();
 b15zdnd11an1n08x5 FILLER_115_1191 ();
 b15zdnd00an1n01x5 FILLER_115_1199 ();
 b15zdnd11an1n32x5 FILLER_115_1218 ();
 b15zdnd11an1n16x5 FILLER_115_1250 ();
 b15zdnd00an1n01x5 FILLER_115_1266 ();
 b15zdnd11an1n08x5 FILLER_115_1271 ();
 b15zdnd11an1n04x5 FILLER_115_1279 ();
 b15zdnd00an1n02x5 FILLER_115_1283 ();
 b15zdnd11an1n32x5 FILLER_115_1291 ();
 b15zdnd11an1n04x5 FILLER_115_1323 ();
 b15zdnd00an1n02x5 FILLER_115_1327 ();
 b15zdnd00an1n01x5 FILLER_115_1329 ();
 b15zdnd11an1n64x5 FILLER_115_1336 ();
 b15zdnd11an1n16x5 FILLER_115_1400 ();
 b15zdnd00an1n02x5 FILLER_115_1416 ();
 b15zdnd00an1n01x5 FILLER_115_1418 ();
 b15zdnd11an1n64x5 FILLER_115_1434 ();
 b15zdnd11an1n32x5 FILLER_115_1498 ();
 b15zdnd11an1n08x5 FILLER_115_1530 ();
 b15zdnd00an1n02x5 FILLER_115_1538 ();
 b15zdnd00an1n01x5 FILLER_115_1540 ();
 b15zdnd11an1n32x5 FILLER_115_1564 ();
 b15zdnd11an1n08x5 FILLER_115_1596 ();
 b15zdnd11an1n08x5 FILLER_115_1624 ();
 b15zdnd11an1n64x5 FILLER_115_1656 ();
 b15zdnd11an1n16x5 FILLER_115_1720 ();
 b15zdnd11an1n08x5 FILLER_115_1736 ();
 b15zdnd00an1n01x5 FILLER_115_1744 ();
 b15zdnd11an1n04x5 FILLER_115_1752 ();
 b15zdnd11an1n04x5 FILLER_115_1761 ();
 b15zdnd00an1n02x5 FILLER_115_1765 ();
 b15zdnd11an1n04x5 FILLER_115_1774 ();
 b15zdnd11an1n64x5 FILLER_115_1783 ();
 b15zdnd11an1n08x5 FILLER_115_1847 ();
 b15zdnd11an1n04x5 FILLER_115_1855 ();
 b15zdnd00an1n02x5 FILLER_115_1859 ();
 b15zdnd11an1n64x5 FILLER_115_1869 ();
 b15zdnd11an1n32x5 FILLER_115_1933 ();
 b15zdnd11an1n16x5 FILLER_115_1965 ();
 b15zdnd11an1n08x5 FILLER_115_1981 ();
 b15zdnd11an1n04x5 FILLER_115_1989 ();
 b15zdnd00an1n02x5 FILLER_115_1993 ();
 b15zdnd00an1n01x5 FILLER_115_1995 ();
 b15zdnd11an1n64x5 FILLER_115_2013 ();
 b15zdnd11an1n64x5 FILLER_115_2077 ();
 b15zdnd11an1n04x5 FILLER_115_2141 ();
 b15zdnd11an1n04x5 FILLER_115_2151 ();
 b15zdnd11an1n08x5 FILLER_115_2167 ();
 b15zdnd11an1n04x5 FILLER_115_2175 ();
 b15zdnd11an1n64x5 FILLER_115_2195 ();
 b15zdnd11an1n16x5 FILLER_115_2259 ();
 b15zdnd11an1n08x5 FILLER_115_2275 ();
 b15zdnd00an1n01x5 FILLER_115_2283 ();
 b15zdnd11an1n16x5 FILLER_116_8 ();
 b15zdnd11an1n08x5 FILLER_116_24 ();
 b15zdnd00an1n02x5 FILLER_116_32 ();
 b15zdnd00an1n01x5 FILLER_116_34 ();
 b15zdnd11an1n04x5 FILLER_116_66 ();
 b15zdnd11an1n32x5 FILLER_116_77 ();
 b15zdnd11an1n04x5 FILLER_116_109 ();
 b15zdnd00an1n02x5 FILLER_116_113 ();
 b15zdnd11an1n08x5 FILLER_116_121 ();
 b15zdnd00an1n02x5 FILLER_116_129 ();
 b15zdnd00an1n01x5 FILLER_116_131 ();
 b15zdnd11an1n04x5 FILLER_116_144 ();
 b15zdnd11an1n64x5 FILLER_116_158 ();
 b15zdnd11an1n32x5 FILLER_116_222 ();
 b15zdnd11an1n16x5 FILLER_116_254 ();
 b15zdnd00an1n02x5 FILLER_116_270 ();
 b15zdnd00an1n01x5 FILLER_116_272 ();
 b15zdnd11an1n08x5 FILLER_116_285 ();
 b15zdnd11an1n04x5 FILLER_116_293 ();
 b15zdnd00an1n01x5 FILLER_116_297 ();
 b15zdnd11an1n08x5 FILLER_116_310 ();
 b15zdnd11an1n04x5 FILLER_116_318 ();
 b15zdnd00an1n02x5 FILLER_116_322 ();
 b15zdnd11an1n04x5 FILLER_116_336 ();
 b15zdnd11an1n64x5 FILLER_116_363 ();
 b15zdnd11an1n08x5 FILLER_116_427 ();
 b15zdnd00an1n02x5 FILLER_116_435 ();
 b15zdnd11an1n16x5 FILLER_116_447 ();
 b15zdnd11an1n04x5 FILLER_116_463 ();
 b15zdnd11an1n16x5 FILLER_116_480 ();
 b15zdnd11an1n08x5 FILLER_116_496 ();
 b15zdnd11an1n04x5 FILLER_116_509 ();
 b15zdnd00an1n01x5 FILLER_116_513 ();
 b15zdnd11an1n08x5 FILLER_116_524 ();
 b15zdnd00an1n01x5 FILLER_116_532 ();
 b15zdnd11an1n16x5 FILLER_116_539 ();
 b15zdnd11an1n04x5 FILLER_116_555 ();
 b15zdnd00an1n02x5 FILLER_116_559 ();
 b15zdnd00an1n01x5 FILLER_116_561 ();
 b15zdnd11an1n04x5 FILLER_116_568 ();
 b15zdnd11an1n16x5 FILLER_116_585 ();
 b15zdnd00an1n02x5 FILLER_116_601 ();
 b15zdnd00an1n01x5 FILLER_116_603 ();
 b15zdnd11an1n16x5 FILLER_116_624 ();
 b15zdnd00an1n02x5 FILLER_116_640 ();
 b15zdnd00an1n01x5 FILLER_116_642 ();
 b15zdnd11an1n08x5 FILLER_116_673 ();
 b15zdnd11an1n04x5 FILLER_116_681 ();
 b15zdnd11an1n16x5 FILLER_116_700 ();
 b15zdnd00an1n02x5 FILLER_116_716 ();
 b15zdnd00an1n02x5 FILLER_116_726 ();
 b15zdnd11an1n08x5 FILLER_116_760 ();
 b15zdnd11an1n04x5 FILLER_116_768 ();
 b15zdnd11an1n16x5 FILLER_116_780 ();
 b15zdnd11an1n16x5 FILLER_116_822 ();
 b15zdnd00an1n01x5 FILLER_116_838 ();
 b15zdnd11an1n08x5 FILLER_116_865 ();
 b15zdnd00an1n02x5 FILLER_116_873 ();
 b15zdnd00an1n01x5 FILLER_116_875 ();
 b15zdnd11an1n64x5 FILLER_116_902 ();
 b15zdnd11an1n32x5 FILLER_116_966 ();
 b15zdnd00an1n02x5 FILLER_116_998 ();
 b15zdnd11an1n16x5 FILLER_116_1020 ();
 b15zdnd00an1n02x5 FILLER_116_1036 ();
 b15zdnd11an1n64x5 FILLER_116_1049 ();
 b15zdnd11an1n32x5 FILLER_116_1113 ();
 b15zdnd11an1n16x5 FILLER_116_1145 ();
 b15zdnd00an1n02x5 FILLER_116_1161 ();
 b15zdnd11an1n32x5 FILLER_116_1183 ();
 b15zdnd11an1n16x5 FILLER_116_1215 ();
 b15zdnd11an1n04x5 FILLER_116_1231 ();
 b15zdnd00an1n01x5 FILLER_116_1235 ();
 b15zdnd11an1n16x5 FILLER_116_1249 ();
 b15zdnd11an1n04x5 FILLER_116_1265 ();
 b15zdnd00an1n02x5 FILLER_116_1269 ();
 b15zdnd11an1n64x5 FILLER_116_1281 ();
 b15zdnd11an1n16x5 FILLER_116_1345 ();
 b15zdnd11an1n04x5 FILLER_116_1361 ();
 b15zdnd00an1n02x5 FILLER_116_1365 ();
 b15zdnd00an1n01x5 FILLER_116_1367 ();
 b15zdnd11an1n08x5 FILLER_116_1372 ();
 b15zdnd11an1n08x5 FILLER_116_1385 ();
 b15zdnd11an1n64x5 FILLER_116_1407 ();
 b15zdnd11an1n32x5 FILLER_116_1471 ();
 b15zdnd11an1n16x5 FILLER_116_1503 ();
 b15zdnd11an1n08x5 FILLER_116_1519 ();
 b15zdnd11an1n04x5 FILLER_116_1527 ();
 b15zdnd00an1n02x5 FILLER_116_1531 ();
 b15zdnd00an1n01x5 FILLER_116_1533 ();
 b15zdnd11an1n16x5 FILLER_116_1546 ();
 b15zdnd11an1n04x5 FILLER_116_1568 ();
 b15zdnd11an1n08x5 FILLER_116_1577 ();
 b15zdnd00an1n01x5 FILLER_116_1585 ();
 b15zdnd11an1n04x5 FILLER_116_1596 ();
 b15zdnd00an1n02x5 FILLER_116_1600 ();
 b15zdnd00an1n01x5 FILLER_116_1602 ();
 b15zdnd11an1n04x5 FILLER_116_1609 ();
 b15zdnd11an1n16x5 FILLER_116_1618 ();
 b15zdnd00an1n02x5 FILLER_116_1634 ();
 b15zdnd11an1n64x5 FILLER_116_1648 ();
 b15zdnd11an1n32x5 FILLER_116_1712 ();
 b15zdnd11an1n16x5 FILLER_116_1744 ();
 b15zdnd11an1n04x5 FILLER_116_1760 ();
 b15zdnd00an1n01x5 FILLER_116_1764 ();
 b15zdnd11an1n08x5 FILLER_116_1771 ();
 b15zdnd11an1n04x5 FILLER_116_1779 ();
 b15zdnd00an1n01x5 FILLER_116_1783 ();
 b15zdnd11an1n16x5 FILLER_116_1791 ();
 b15zdnd11an1n08x5 FILLER_116_1807 ();
 b15zdnd11an1n04x5 FILLER_116_1815 ();
 b15zdnd00an1n02x5 FILLER_116_1819 ();
 b15zdnd00an1n01x5 FILLER_116_1821 ();
 b15zdnd11an1n16x5 FILLER_116_1832 ();
 b15zdnd11an1n04x5 FILLER_116_1848 ();
 b15zdnd00an1n02x5 FILLER_116_1852 ();
 b15zdnd00an1n01x5 FILLER_116_1854 ();
 b15zdnd11an1n32x5 FILLER_116_1860 ();
 b15zdnd00an1n02x5 FILLER_116_1892 ();
 b15zdnd00an1n01x5 FILLER_116_1894 ();
 b15zdnd11an1n04x5 FILLER_116_1902 ();
 b15zdnd11an1n16x5 FILLER_116_1912 ();
 b15zdnd11an1n04x5 FILLER_116_1928 ();
 b15zdnd11an1n32x5 FILLER_116_1941 ();
 b15zdnd11an1n16x5 FILLER_116_1973 ();
 b15zdnd11an1n32x5 FILLER_116_1993 ();
 b15zdnd11an1n16x5 FILLER_116_2025 ();
 b15zdnd11an1n04x5 FILLER_116_2041 ();
 b15zdnd00an1n02x5 FILLER_116_2045 ();
 b15zdnd11an1n08x5 FILLER_116_2056 ();
 b15zdnd11an1n08x5 FILLER_116_2069 ();
 b15zdnd00an1n02x5 FILLER_116_2077 ();
 b15zdnd00an1n01x5 FILLER_116_2079 ();
 b15zdnd11an1n16x5 FILLER_116_2092 ();
 b15zdnd11an1n08x5 FILLER_116_2108 ();
 b15zdnd11an1n16x5 FILLER_116_2130 ();
 b15zdnd11an1n08x5 FILLER_116_2146 ();
 b15zdnd11an1n64x5 FILLER_116_2162 ();
 b15zdnd11an1n32x5 FILLER_116_2226 ();
 b15zdnd11an1n08x5 FILLER_116_2263 ();
 b15zdnd11an1n04x5 FILLER_116_2271 ();
 b15zdnd00an1n01x5 FILLER_116_2275 ();
 b15zdnd11an1n32x5 FILLER_117_0 ();
 b15zdnd11an1n04x5 FILLER_117_32 ();
 b15zdnd11an1n04x5 FILLER_117_54 ();
 b15zdnd11an1n32x5 FILLER_117_80 ();
 b15zdnd11an1n16x5 FILLER_117_112 ();
 b15zdnd11an1n08x5 FILLER_117_128 ();
 b15zdnd00an1n01x5 FILLER_117_136 ();
 b15zdnd11an1n64x5 FILLER_117_156 ();
 b15zdnd11an1n32x5 FILLER_117_220 ();
 b15zdnd11an1n08x5 FILLER_117_252 ();
 b15zdnd11an1n04x5 FILLER_117_260 ();
 b15zdnd11an1n64x5 FILLER_117_278 ();
 b15zdnd11an1n64x5 FILLER_117_342 ();
 b15zdnd11an1n16x5 FILLER_117_406 ();
 b15zdnd00an1n02x5 FILLER_117_422 ();
 b15zdnd00an1n01x5 FILLER_117_424 ();
 b15zdnd11an1n04x5 FILLER_117_432 ();
 b15zdnd11an1n16x5 FILLER_117_450 ();
 b15zdnd11an1n04x5 FILLER_117_466 ();
 b15zdnd11an1n16x5 FILLER_117_474 ();
 b15zdnd11an1n04x5 FILLER_117_490 ();
 b15zdnd11an1n16x5 FILLER_117_506 ();
 b15zdnd11an1n16x5 FILLER_117_538 ();
 b15zdnd00an1n02x5 FILLER_117_554 ();
 b15zdnd00an1n01x5 FILLER_117_556 ();
 b15zdnd11an1n64x5 FILLER_117_568 ();
 b15zdnd11an1n16x5 FILLER_117_632 ();
 b15zdnd11an1n08x5 FILLER_117_648 ();
 b15zdnd11an1n04x5 FILLER_117_656 ();
 b15zdnd00an1n02x5 FILLER_117_660 ();
 b15zdnd11an1n32x5 FILLER_117_666 ();
 b15zdnd11an1n16x5 FILLER_117_698 ();
 b15zdnd11an1n08x5 FILLER_117_714 ();
 b15zdnd11an1n04x5 FILLER_117_722 ();
 b15zdnd00an1n02x5 FILLER_117_726 ();
 b15zdnd00an1n01x5 FILLER_117_728 ();
 b15zdnd11an1n16x5 FILLER_117_738 ();
 b15zdnd11an1n08x5 FILLER_117_754 ();
 b15zdnd11an1n04x5 FILLER_117_762 ();
 b15zdnd00an1n01x5 FILLER_117_766 ();
 b15zdnd11an1n04x5 FILLER_117_783 ();
 b15zdnd11an1n08x5 FILLER_117_793 ();
 b15zdnd11an1n04x5 FILLER_117_806 ();
 b15zdnd11an1n04x5 FILLER_117_815 ();
 b15zdnd00an1n01x5 FILLER_117_819 ();
 b15zdnd11an1n16x5 FILLER_117_828 ();
 b15zdnd11an1n08x5 FILLER_117_844 ();
 b15zdnd11an1n04x5 FILLER_117_852 ();
 b15zdnd11an1n32x5 FILLER_117_868 ();
 b15zdnd11an1n16x5 FILLER_117_906 ();
 b15zdnd11an1n64x5 FILLER_117_948 ();
 b15zdnd11an1n08x5 FILLER_117_1012 ();
 b15zdnd11an1n04x5 FILLER_117_1020 ();
 b15zdnd11an1n64x5 FILLER_117_1044 ();
 b15zdnd11an1n16x5 FILLER_117_1108 ();
 b15zdnd11an1n08x5 FILLER_117_1124 ();
 b15zdnd00an1n01x5 FILLER_117_1132 ();
 b15zdnd11an1n32x5 FILLER_117_1137 ();
 b15zdnd11an1n16x5 FILLER_117_1169 ();
 b15zdnd11an1n08x5 FILLER_117_1185 ();
 b15zdnd11an1n32x5 FILLER_117_1205 ();
 b15zdnd11an1n08x5 FILLER_117_1237 ();
 b15zdnd11an1n04x5 FILLER_117_1252 ();
 b15zdnd11an1n64x5 FILLER_117_1263 ();
 b15zdnd11an1n08x5 FILLER_117_1327 ();
 b15zdnd11an1n04x5 FILLER_117_1335 ();
 b15zdnd00an1n02x5 FILLER_117_1339 ();
 b15zdnd11an1n64x5 FILLER_117_1348 ();
 b15zdnd11an1n16x5 FILLER_117_1412 ();
 b15zdnd11an1n08x5 FILLER_117_1428 ();
 b15zdnd11an1n04x5 FILLER_117_1436 ();
 b15zdnd00an1n01x5 FILLER_117_1440 ();
 b15zdnd11an1n08x5 FILLER_117_1447 ();
 b15zdnd00an1n02x5 FILLER_117_1455 ();
 b15zdnd00an1n01x5 FILLER_117_1457 ();
 b15zdnd11an1n32x5 FILLER_117_1468 ();
 b15zdnd11an1n16x5 FILLER_117_1500 ();
 b15zdnd11an1n08x5 FILLER_117_1516 ();
 b15zdnd11an1n04x5 FILLER_117_1524 ();
 b15zdnd11an1n16x5 FILLER_117_1533 ();
 b15zdnd11an1n08x5 FILLER_117_1549 ();
 b15zdnd11an1n04x5 FILLER_117_1557 ();
 b15zdnd00an1n01x5 FILLER_117_1561 ();
 b15zdnd11an1n04x5 FILLER_117_1588 ();
 b15zdnd11an1n64x5 FILLER_117_1597 ();
 b15zdnd11an1n64x5 FILLER_117_1661 ();
 b15zdnd11an1n16x5 FILLER_117_1725 ();
 b15zdnd11an1n04x5 FILLER_117_1741 ();
 b15zdnd00an1n01x5 FILLER_117_1745 ();
 b15zdnd11an1n16x5 FILLER_117_1777 ();
 b15zdnd11an1n08x5 FILLER_117_1793 ();
 b15zdnd11an1n04x5 FILLER_117_1801 ();
 b15zdnd00an1n01x5 FILLER_117_1805 ();
 b15zdnd11an1n32x5 FILLER_117_1810 ();
 b15zdnd11an1n04x5 FILLER_117_1842 ();
 b15zdnd00an1n01x5 FILLER_117_1846 ();
 b15zdnd11an1n04x5 FILLER_117_1851 ();
 b15zdnd11an1n64x5 FILLER_117_1864 ();
 b15zdnd11an1n64x5 FILLER_117_1928 ();
 b15zdnd11an1n64x5 FILLER_117_1992 ();
 b15zdnd11an1n04x5 FILLER_117_2056 ();
 b15zdnd00an1n02x5 FILLER_117_2060 ();
 b15zdnd00an1n01x5 FILLER_117_2062 ();
 b15zdnd11an1n08x5 FILLER_117_2072 ();
 b15zdnd11an1n04x5 FILLER_117_2080 ();
 b15zdnd00an1n01x5 FILLER_117_2084 ();
 b15zdnd11an1n32x5 FILLER_117_2097 ();
 b15zdnd00an1n01x5 FILLER_117_2129 ();
 b15zdnd11an1n04x5 FILLER_117_2142 ();
 b15zdnd11an1n08x5 FILLER_117_2161 ();
 b15zdnd11an1n04x5 FILLER_117_2169 ();
 b15zdnd00an1n02x5 FILLER_117_2173 ();
 b15zdnd00an1n01x5 FILLER_117_2175 ();
 b15zdnd11an1n08x5 FILLER_117_2185 ();
 b15zdnd11an1n04x5 FILLER_117_2193 ();
 b15zdnd00an1n02x5 FILLER_117_2197 ();
 b15zdnd11an1n32x5 FILLER_117_2217 ();
 b15zdnd11an1n04x5 FILLER_117_2249 ();
 b15zdnd11an1n04x5 FILLER_117_2273 ();
 b15zdnd00an1n02x5 FILLER_117_2281 ();
 b15zdnd00an1n01x5 FILLER_117_2283 ();
 b15zdnd11an1n64x5 FILLER_118_8 ();
 b15zdnd11an1n64x5 FILLER_118_72 ();
 b15zdnd11an1n32x5 FILLER_118_136 ();
 b15zdnd11an1n16x5 FILLER_118_168 ();
 b15zdnd11an1n08x5 FILLER_118_190 ();
 b15zdnd11an1n04x5 FILLER_118_207 ();
 b15zdnd11an1n04x5 FILLER_118_217 ();
 b15zdnd11an1n64x5 FILLER_118_228 ();
 b15zdnd11an1n64x5 FILLER_118_292 ();
 b15zdnd11an1n64x5 FILLER_118_356 ();
 b15zdnd11an1n16x5 FILLER_118_420 ();
 b15zdnd11an1n08x5 FILLER_118_436 ();
 b15zdnd11an1n04x5 FILLER_118_444 ();
 b15zdnd00an1n02x5 FILLER_118_448 ();
 b15zdnd11an1n04x5 FILLER_118_457 ();
 b15zdnd11an1n32x5 FILLER_118_473 ();
 b15zdnd11an1n16x5 FILLER_118_505 ();
 b15zdnd11an1n04x5 FILLER_118_521 ();
 b15zdnd00an1n02x5 FILLER_118_525 ();
 b15zdnd11an1n16x5 FILLER_118_532 ();
 b15zdnd00an1n02x5 FILLER_118_548 ();
 b15zdnd00an1n01x5 FILLER_118_550 ();
 b15zdnd11an1n16x5 FILLER_118_559 ();
 b15zdnd11an1n08x5 FILLER_118_575 ();
 b15zdnd11an1n04x5 FILLER_118_583 ();
 b15zdnd00an1n01x5 FILLER_118_587 ();
 b15zdnd11an1n16x5 FILLER_118_593 ();
 b15zdnd11an1n08x5 FILLER_118_609 ();
 b15zdnd00an1n01x5 FILLER_118_617 ();
 b15zdnd11an1n16x5 FILLER_118_629 ();
 b15zdnd11an1n08x5 FILLER_118_645 ();
 b15zdnd11an1n04x5 FILLER_118_653 ();
 b15zdnd00an1n02x5 FILLER_118_657 ();
 b15zdnd00an1n01x5 FILLER_118_659 ();
 b15zdnd11an1n04x5 FILLER_118_666 ();
 b15zdnd11an1n08x5 FILLER_118_680 ();
 b15zdnd11an1n04x5 FILLER_118_688 ();
 b15zdnd00an1n02x5 FILLER_118_692 ();
 b15zdnd00an1n01x5 FILLER_118_694 ();
 b15zdnd11an1n16x5 FILLER_118_701 ();
 b15zdnd00an1n01x5 FILLER_118_717 ();
 b15zdnd11an1n16x5 FILLER_118_726 ();
 b15zdnd11an1n08x5 FILLER_118_748 ();
 b15zdnd00an1n02x5 FILLER_118_756 ();
 b15zdnd11an1n32x5 FILLER_118_763 ();
 b15zdnd11an1n16x5 FILLER_118_795 ();
 b15zdnd00an1n02x5 FILLER_118_811 ();
 b15zdnd00an1n01x5 FILLER_118_813 ();
 b15zdnd11an1n04x5 FILLER_118_820 ();
 b15zdnd00an1n02x5 FILLER_118_824 ();
 b15zdnd11an1n32x5 FILLER_118_831 ();
 b15zdnd11an1n16x5 FILLER_118_863 ();
 b15zdnd11an1n08x5 FILLER_118_879 ();
 b15zdnd11an1n04x5 FILLER_118_887 ();
 b15zdnd11an1n04x5 FILLER_118_897 ();
 b15zdnd11an1n64x5 FILLER_118_912 ();
 b15zdnd11an1n64x5 FILLER_118_976 ();
 b15zdnd11an1n64x5 FILLER_118_1040 ();
 b15zdnd11an1n64x5 FILLER_118_1104 ();
 b15zdnd11an1n32x5 FILLER_118_1168 ();
 b15zdnd11an1n04x5 FILLER_118_1200 ();
 b15zdnd00an1n02x5 FILLER_118_1204 ();
 b15zdnd11an1n08x5 FILLER_118_1212 ();
 b15zdnd11an1n32x5 FILLER_118_1230 ();
 b15zdnd11an1n16x5 FILLER_118_1262 ();
 b15zdnd11an1n08x5 FILLER_118_1278 ();
 b15zdnd00an1n02x5 FILLER_118_1286 ();
 b15zdnd00an1n01x5 FILLER_118_1288 ();
 b15zdnd11an1n04x5 FILLER_118_1304 ();
 b15zdnd11an1n16x5 FILLER_118_1323 ();
 b15zdnd11an1n04x5 FILLER_118_1339 ();
 b15zdnd00an1n01x5 FILLER_118_1343 ();
 b15zdnd11an1n64x5 FILLER_118_1351 ();
 b15zdnd00an1n01x5 FILLER_118_1415 ();
 b15zdnd11an1n08x5 FILLER_118_1427 ();
 b15zdnd11an1n04x5 FILLER_118_1435 ();
 b15zdnd00an1n01x5 FILLER_118_1439 ();
 b15zdnd11an1n08x5 FILLER_118_1449 ();
 b15zdnd11an1n04x5 FILLER_118_1457 ();
 b15zdnd00an1n01x5 FILLER_118_1461 ();
 b15zdnd11an1n16x5 FILLER_118_1476 ();
 b15zdnd00an1n01x5 FILLER_118_1492 ();
 b15zdnd11an1n16x5 FILLER_118_1500 ();
 b15zdnd11an1n08x5 FILLER_118_1516 ();
 b15zdnd11an1n04x5 FILLER_118_1530 ();
 b15zdnd11an1n32x5 FILLER_118_1541 ();
 b15zdnd11an1n08x5 FILLER_118_1573 ();
 b15zdnd11an1n04x5 FILLER_118_1591 ();
 b15zdnd00an1n02x5 FILLER_118_1595 ();
 b15zdnd11an1n08x5 FILLER_118_1603 ();
 b15zdnd11an1n04x5 FILLER_118_1611 ();
 b15zdnd00an1n02x5 FILLER_118_1615 ();
 b15zdnd11an1n32x5 FILLER_118_1621 ();
 b15zdnd11an1n16x5 FILLER_118_1653 ();
 b15zdnd11an1n08x5 FILLER_118_1669 ();
 b15zdnd11an1n04x5 FILLER_118_1677 ();
 b15zdnd00an1n02x5 FILLER_118_1681 ();
 b15zdnd11an1n64x5 FILLER_118_1703 ();
 b15zdnd11an1n32x5 FILLER_118_1767 ();
 b15zdnd11an1n16x5 FILLER_118_1816 ();
 b15zdnd11an1n08x5 FILLER_118_1832 ();
 b15zdnd00an1n02x5 FILLER_118_1840 ();
 b15zdnd11an1n08x5 FILLER_118_1846 ();
 b15zdnd11an1n32x5 FILLER_118_1863 ();
 b15zdnd11an1n08x5 FILLER_118_1895 ();
 b15zdnd11an1n04x5 FILLER_118_1903 ();
 b15zdnd11an1n32x5 FILLER_118_1915 ();
 b15zdnd11an1n08x5 FILLER_118_1947 ();
 b15zdnd00an1n02x5 FILLER_118_1955 ();
 b15zdnd11an1n04x5 FILLER_118_1961 ();
 b15zdnd00an1n02x5 FILLER_118_1965 ();
 b15zdnd00an1n01x5 FILLER_118_1967 ();
 b15zdnd11an1n04x5 FILLER_118_1977 ();
 b15zdnd11an1n16x5 FILLER_118_1985 ();
 b15zdnd11an1n08x5 FILLER_118_2001 ();
 b15zdnd00an1n01x5 FILLER_118_2009 ();
 b15zdnd11an1n04x5 FILLER_118_2021 ();
 b15zdnd11an1n04x5 FILLER_118_2034 ();
 b15zdnd11an1n04x5 FILLER_118_2043 ();
 b15zdnd11an1n04x5 FILLER_118_2052 ();
 b15zdnd00an1n02x5 FILLER_118_2056 ();
 b15zdnd00an1n01x5 FILLER_118_2058 ();
 b15zdnd11an1n04x5 FILLER_118_2074 ();
 b15zdnd11an1n16x5 FILLER_118_2084 ();
 b15zdnd00an1n01x5 FILLER_118_2100 ();
 b15zdnd11an1n04x5 FILLER_118_2111 ();
 b15zdnd11an1n16x5 FILLER_118_2129 ();
 b15zdnd11an1n08x5 FILLER_118_2145 ();
 b15zdnd00an1n01x5 FILLER_118_2153 ();
 b15zdnd00an1n02x5 FILLER_118_2162 ();
 b15zdnd11an1n64x5 FILLER_118_2172 ();
 b15zdnd11an1n16x5 FILLER_118_2236 ();
 b15zdnd11an1n04x5 FILLER_118_2252 ();
 b15zdnd00an1n01x5 FILLER_118_2256 ();
 b15zdnd11an1n16x5 FILLER_118_2260 ();
 b15zdnd11an1n64x5 FILLER_119_0 ();
 b15zdnd00an1n02x5 FILLER_119_64 ();
 b15zdnd00an1n01x5 FILLER_119_66 ();
 b15zdnd11an1n64x5 FILLER_119_74 ();
 b15zdnd11an1n08x5 FILLER_119_138 ();
 b15zdnd00an1n02x5 FILLER_119_146 ();
 b15zdnd11an1n04x5 FILLER_119_155 ();
 b15zdnd11an1n04x5 FILLER_119_167 ();
 b15zdnd00an1n01x5 FILLER_119_171 ();
 b15zdnd11an1n04x5 FILLER_119_188 ();
 b15zdnd11an1n32x5 FILLER_119_208 ();
 b15zdnd11an1n08x5 FILLER_119_240 ();
 b15zdnd00an1n01x5 FILLER_119_248 ();
 b15zdnd11an1n04x5 FILLER_119_254 ();
 b15zdnd11an1n04x5 FILLER_119_266 ();
 b15zdnd11an1n32x5 FILLER_119_276 ();
 b15zdnd00an1n01x5 FILLER_119_308 ();
 b15zdnd11an1n04x5 FILLER_119_325 ();
 b15zdnd11an1n16x5 FILLER_119_336 ();
 b15zdnd00an1n02x5 FILLER_119_352 ();
 b15zdnd11an1n04x5 FILLER_119_362 ();
 b15zdnd11an1n32x5 FILLER_119_386 ();
 b15zdnd11an1n16x5 FILLER_119_418 ();
 b15zdnd11an1n04x5 FILLER_119_434 ();
 b15zdnd00an1n02x5 FILLER_119_438 ();
 b15zdnd11an1n64x5 FILLER_119_453 ();
 b15zdnd11an1n32x5 FILLER_119_517 ();
 b15zdnd11an1n04x5 FILLER_119_549 ();
 b15zdnd11an1n32x5 FILLER_119_557 ();
 b15zdnd11an1n16x5 FILLER_119_589 ();
 b15zdnd00an1n02x5 FILLER_119_605 ();
 b15zdnd00an1n01x5 FILLER_119_607 ();
 b15zdnd11an1n08x5 FILLER_119_613 ();
 b15zdnd11an1n32x5 FILLER_119_634 ();
 b15zdnd11an1n16x5 FILLER_119_666 ();
 b15zdnd11an1n08x5 FILLER_119_682 ();
 b15zdnd11an1n04x5 FILLER_119_690 ();
 b15zdnd11an1n32x5 FILLER_119_700 ();
 b15zdnd00an1n02x5 FILLER_119_732 ();
 b15zdnd00an1n01x5 FILLER_119_734 ();
 b15zdnd11an1n64x5 FILLER_119_748 ();
 b15zdnd11an1n04x5 FILLER_119_812 ();
 b15zdnd00an1n02x5 FILLER_119_816 ();
 b15zdnd11an1n04x5 FILLER_119_828 ();
 b15zdnd00an1n02x5 FILLER_119_832 ();
 b15zdnd11an1n08x5 FILLER_119_838 ();
 b15zdnd11an1n04x5 FILLER_119_846 ();
 b15zdnd00an1n01x5 FILLER_119_850 ();
 b15zdnd11an1n64x5 FILLER_119_858 ();
 b15zdnd11an1n64x5 FILLER_119_922 ();
 b15zdnd11an1n64x5 FILLER_119_986 ();
 b15zdnd11an1n08x5 FILLER_119_1050 ();
 b15zdnd11an1n04x5 FILLER_119_1058 ();
 b15zdnd00an1n02x5 FILLER_119_1062 ();
 b15zdnd00an1n01x5 FILLER_119_1064 ();
 b15zdnd11an1n64x5 FILLER_119_1085 ();
 b15zdnd11an1n32x5 FILLER_119_1149 ();
 b15zdnd11an1n16x5 FILLER_119_1181 ();
 b15zdnd11an1n04x5 FILLER_119_1197 ();
 b15zdnd00an1n01x5 FILLER_119_1201 ();
 b15zdnd11an1n08x5 FILLER_119_1209 ();
 b15zdnd11an1n04x5 FILLER_119_1217 ();
 b15zdnd00an1n02x5 FILLER_119_1221 ();
 b15zdnd11an1n04x5 FILLER_119_1229 ();
 b15zdnd00an1n02x5 FILLER_119_1233 ();
 b15zdnd11an1n16x5 FILLER_119_1245 ();
 b15zdnd11an1n08x5 FILLER_119_1261 ();
 b15zdnd11an1n04x5 FILLER_119_1269 ();
 b15zdnd00an1n02x5 FILLER_119_1273 ();
 b15zdnd00an1n01x5 FILLER_119_1275 ();
 b15zdnd11an1n04x5 FILLER_119_1283 ();
 b15zdnd11an1n04x5 FILLER_119_1307 ();
 b15zdnd11an1n04x5 FILLER_119_1315 ();
 b15zdnd11an1n04x5 FILLER_119_1326 ();
 b15zdnd00an1n01x5 FILLER_119_1330 ();
 b15zdnd11an1n16x5 FILLER_119_1343 ();
 b15zdnd11an1n04x5 FILLER_119_1359 ();
 b15zdnd00an1n02x5 FILLER_119_1363 ();
 b15zdnd11an1n04x5 FILLER_119_1371 ();
 b15zdnd11an1n04x5 FILLER_119_1380 ();
 b15zdnd00an1n01x5 FILLER_119_1384 ();
 b15zdnd11an1n08x5 FILLER_119_1390 ();
 b15zdnd00an1n01x5 FILLER_119_1398 ();
 b15zdnd11an1n32x5 FILLER_119_1403 ();
 b15zdnd11an1n16x5 FILLER_119_1435 ();
 b15zdnd11an1n08x5 FILLER_119_1451 ();
 b15zdnd00an1n02x5 FILLER_119_1459 ();
 b15zdnd11an1n16x5 FILLER_119_1466 ();
 b15zdnd00an1n02x5 FILLER_119_1482 ();
 b15zdnd11an1n04x5 FILLER_119_1489 ();
 b15zdnd11an1n16x5 FILLER_119_1505 ();
 b15zdnd11an1n08x5 FILLER_119_1521 ();
 b15zdnd00an1n01x5 FILLER_119_1529 ();
 b15zdnd11an1n64x5 FILLER_119_1535 ();
 b15zdnd11an1n16x5 FILLER_119_1599 ();
 b15zdnd00an1n01x5 FILLER_119_1615 ();
 b15zdnd11an1n08x5 FILLER_119_1622 ();
 b15zdnd11an1n16x5 FILLER_119_1656 ();
 b15zdnd11an1n08x5 FILLER_119_1672 ();
 b15zdnd00an1n02x5 FILLER_119_1680 ();
 b15zdnd00an1n01x5 FILLER_119_1682 ();
 b15zdnd11an1n08x5 FILLER_119_1688 ();
 b15zdnd11an1n04x5 FILLER_119_1696 ();
 b15zdnd11an1n32x5 FILLER_119_1703 ();
 b15zdnd11an1n16x5 FILLER_119_1735 ();
 b15zdnd11an1n08x5 FILLER_119_1751 ();
 b15zdnd00an1n02x5 FILLER_119_1759 ();
 b15zdnd00an1n01x5 FILLER_119_1761 ();
 b15zdnd11an1n08x5 FILLER_119_1772 ();
 b15zdnd11an1n04x5 FILLER_119_1780 ();
 b15zdnd00an1n02x5 FILLER_119_1784 ();
 b15zdnd11an1n04x5 FILLER_119_1790 ();
 b15zdnd00an1n02x5 FILLER_119_1794 ();
 b15zdnd11an1n04x5 FILLER_119_1805 ();
 b15zdnd11an1n04x5 FILLER_119_1832 ();
 b15zdnd11an1n08x5 FILLER_119_1846 ();
 b15zdnd11an1n04x5 FILLER_119_1854 ();
 b15zdnd00an1n02x5 FILLER_119_1858 ();
 b15zdnd00an1n01x5 FILLER_119_1860 ();
 b15zdnd11an1n16x5 FILLER_119_1865 ();
 b15zdnd11an1n08x5 FILLER_119_1881 ();
 b15zdnd11an1n04x5 FILLER_119_1889 ();
 b15zdnd00an1n02x5 FILLER_119_1893 ();
 b15zdnd00an1n01x5 FILLER_119_1895 ();
 b15zdnd11an1n04x5 FILLER_119_1901 ();
 b15zdnd11an1n04x5 FILLER_119_1910 ();
 b15zdnd00an1n02x5 FILLER_119_1914 ();
 b15zdnd11an1n04x5 FILLER_119_1922 ();
 b15zdnd11an1n16x5 FILLER_119_1930 ();
 b15zdnd11an1n08x5 FILLER_119_1946 ();
 b15zdnd00an1n01x5 FILLER_119_1954 ();
 b15zdnd11an1n16x5 FILLER_119_1962 ();
 b15zdnd11an1n04x5 FILLER_119_1996 ();
 b15zdnd00an1n02x5 FILLER_119_2000 ();
 b15zdnd00an1n01x5 FILLER_119_2002 ();
 b15zdnd11an1n64x5 FILLER_119_2019 ();
 b15zdnd00an1n02x5 FILLER_119_2083 ();
 b15zdnd00an1n01x5 FILLER_119_2085 ();
 b15zdnd11an1n08x5 FILLER_119_2092 ();
 b15zdnd11an1n04x5 FILLER_119_2126 ();
 b15zdnd11an1n32x5 FILLER_119_2136 ();
 b15zdnd11an1n04x5 FILLER_119_2168 ();
 b15zdnd00an1n02x5 FILLER_119_2172 ();
 b15zdnd00an1n01x5 FILLER_119_2174 ();
 b15zdnd11an1n64x5 FILLER_119_2198 ();
 b15zdnd11an1n16x5 FILLER_119_2262 ();
 b15zdnd11an1n04x5 FILLER_119_2278 ();
 b15zdnd00an1n02x5 FILLER_119_2282 ();
 b15zdnd11an1n16x5 FILLER_120_8 ();
 b15zdnd11an1n08x5 FILLER_120_24 ();
 b15zdnd11an1n04x5 FILLER_120_32 ();
 b15zdnd00an1n02x5 FILLER_120_36 ();
 b15zdnd11an1n04x5 FILLER_120_54 ();
 b15zdnd11an1n32x5 FILLER_120_70 ();
 b15zdnd11an1n08x5 FILLER_120_102 ();
 b15zdnd00an1n01x5 FILLER_120_110 ();
 b15zdnd11an1n32x5 FILLER_120_118 ();
 b15zdnd11an1n16x5 FILLER_120_150 ();
 b15zdnd11an1n08x5 FILLER_120_166 ();
 b15zdnd11an1n04x5 FILLER_120_174 ();
 b15zdnd00an1n01x5 FILLER_120_178 ();
 b15zdnd11an1n04x5 FILLER_120_192 ();
 b15zdnd11an1n16x5 FILLER_120_205 ();
 b15zdnd00an1n02x5 FILLER_120_221 ();
 b15zdnd00an1n01x5 FILLER_120_223 ();
 b15zdnd11an1n16x5 FILLER_120_236 ();
 b15zdnd11an1n04x5 FILLER_120_252 ();
 b15zdnd00an1n01x5 FILLER_120_256 ();
 b15zdnd11an1n16x5 FILLER_120_262 ();
 b15zdnd00an1n02x5 FILLER_120_278 ();
 b15zdnd11an1n32x5 FILLER_120_298 ();
 b15zdnd00an1n01x5 FILLER_120_330 ();
 b15zdnd11an1n64x5 FILLER_120_340 ();
 b15zdnd11an1n16x5 FILLER_120_404 ();
 b15zdnd11an1n08x5 FILLER_120_420 ();
 b15zdnd00an1n01x5 FILLER_120_428 ();
 b15zdnd11an1n16x5 FILLER_120_438 ();
 b15zdnd11an1n04x5 FILLER_120_463 ();
 b15zdnd00an1n02x5 FILLER_120_467 ();
 b15zdnd11an1n04x5 FILLER_120_475 ();
 b15zdnd11an1n04x5 FILLER_120_486 ();
 b15zdnd00an1n02x5 FILLER_120_490 ();
 b15zdnd11an1n32x5 FILLER_120_498 ();
 b15zdnd11an1n08x5 FILLER_120_530 ();
 b15zdnd11an1n04x5 FILLER_120_538 ();
 b15zdnd00an1n02x5 FILLER_120_542 ();
 b15zdnd11an1n16x5 FILLER_120_567 ();
 b15zdnd11an1n08x5 FILLER_120_583 ();
 b15zdnd11an1n04x5 FILLER_120_591 ();
 b15zdnd11an1n08x5 FILLER_120_616 ();
 b15zdnd11an1n04x5 FILLER_120_624 ();
 b15zdnd11an1n16x5 FILLER_120_632 ();
 b15zdnd00an1n02x5 FILLER_120_648 ();
 b15zdnd11an1n32x5 FILLER_120_657 ();
 b15zdnd11an1n16x5 FILLER_120_689 ();
 b15zdnd11an1n08x5 FILLER_120_705 ();
 b15zdnd11an1n04x5 FILLER_120_713 ();
 b15zdnd00an1n01x5 FILLER_120_717 ();
 b15zdnd11an1n04x5 FILLER_120_726 ();
 b15zdnd11an1n64x5 FILLER_120_751 ();
 b15zdnd00an1n02x5 FILLER_120_815 ();
 b15zdnd11an1n32x5 FILLER_120_829 ();
 b15zdnd11an1n32x5 FILLER_120_882 ();
 b15zdnd11an1n16x5 FILLER_120_914 ();
 b15zdnd11an1n04x5 FILLER_120_930 ();
 b15zdnd00an1n02x5 FILLER_120_934 ();
 b15zdnd00an1n01x5 FILLER_120_936 ();
 b15zdnd11an1n64x5 FILLER_120_957 ();
 b15zdnd11an1n32x5 FILLER_120_1021 ();
 b15zdnd11an1n08x5 FILLER_120_1053 ();
 b15zdnd00an1n02x5 FILLER_120_1061 ();
 b15zdnd11an1n64x5 FILLER_120_1074 ();
 b15zdnd11an1n32x5 FILLER_120_1138 ();
 b15zdnd11an1n04x5 FILLER_120_1170 ();
 b15zdnd11an1n32x5 FILLER_120_1205 ();
 b15zdnd11an1n16x5 FILLER_120_1237 ();
 b15zdnd11an1n08x5 FILLER_120_1253 ();
 b15zdnd11an1n04x5 FILLER_120_1261 ();
 b15zdnd00an1n01x5 FILLER_120_1265 ();
 b15zdnd11an1n04x5 FILLER_120_1270 ();
 b15zdnd11an1n04x5 FILLER_120_1281 ();
 b15zdnd00an1n01x5 FILLER_120_1285 ();
 b15zdnd11an1n32x5 FILLER_120_1294 ();
 b15zdnd11an1n08x5 FILLER_120_1326 ();
 b15zdnd00an1n01x5 FILLER_120_1334 ();
 b15zdnd11an1n08x5 FILLER_120_1348 ();
 b15zdnd11an1n04x5 FILLER_120_1356 ();
 b15zdnd00an1n01x5 FILLER_120_1360 ();
 b15zdnd11an1n16x5 FILLER_120_1373 ();
 b15zdnd11an1n04x5 FILLER_120_1389 ();
 b15zdnd00an1n02x5 FILLER_120_1393 ();
 b15zdnd00an1n01x5 FILLER_120_1395 ();
 b15zdnd11an1n64x5 FILLER_120_1402 ();
 b15zdnd11an1n16x5 FILLER_120_1466 ();
 b15zdnd11an1n08x5 FILLER_120_1482 ();
 b15zdnd00an1n02x5 FILLER_120_1490 ();
 b15zdnd00an1n01x5 FILLER_120_1492 ();
 b15zdnd11an1n08x5 FILLER_120_1511 ();
 b15zdnd00an1n02x5 FILLER_120_1519 ();
 b15zdnd00an1n01x5 FILLER_120_1521 ();
 b15zdnd11an1n32x5 FILLER_120_1527 ();
 b15zdnd11an1n16x5 FILLER_120_1559 ();
 b15zdnd11an1n08x5 FILLER_120_1575 ();
 b15zdnd11an1n04x5 FILLER_120_1583 ();
 b15zdnd00an1n02x5 FILLER_120_1587 ();
 b15zdnd00an1n01x5 FILLER_120_1589 ();
 b15zdnd11an1n16x5 FILLER_120_1596 ();
 b15zdnd11an1n08x5 FILLER_120_1612 ();
 b15zdnd00an1n02x5 FILLER_120_1620 ();
 b15zdnd00an1n01x5 FILLER_120_1622 ();
 b15zdnd11an1n04x5 FILLER_120_1631 ();
 b15zdnd11an1n64x5 FILLER_120_1651 ();
 b15zdnd11an1n16x5 FILLER_120_1715 ();
 b15zdnd11an1n08x5 FILLER_120_1731 ();
 b15zdnd11an1n08x5 FILLER_120_1757 ();
 b15zdnd11an1n04x5 FILLER_120_1765 ();
 b15zdnd00an1n01x5 FILLER_120_1769 ();
 b15zdnd11an1n04x5 FILLER_120_1784 ();
 b15zdnd11an1n64x5 FILLER_120_1793 ();
 b15zdnd11an1n08x5 FILLER_120_1857 ();
 b15zdnd00an1n02x5 FILLER_120_1865 ();
 b15zdnd11an1n16x5 FILLER_120_1883 ();
 b15zdnd11an1n08x5 FILLER_120_1899 ();
 b15zdnd00an1n01x5 FILLER_120_1907 ();
 b15zdnd11an1n16x5 FILLER_120_1912 ();
 b15zdnd11an1n04x5 FILLER_120_1928 ();
 b15zdnd00an1n02x5 FILLER_120_1932 ();
 b15zdnd11an1n08x5 FILLER_120_1942 ();
 b15zdnd11an1n04x5 FILLER_120_1950 ();
 b15zdnd00an1n02x5 FILLER_120_1954 ();
 b15zdnd00an1n01x5 FILLER_120_1956 ();
 b15zdnd11an1n64x5 FILLER_120_1961 ();
 b15zdnd11an1n64x5 FILLER_120_2025 ();
 b15zdnd11an1n64x5 FILLER_120_2089 ();
 b15zdnd00an1n01x5 FILLER_120_2153 ();
 b15zdnd11an1n16x5 FILLER_120_2162 ();
 b15zdnd00an1n02x5 FILLER_120_2178 ();
 b15zdnd00an1n01x5 FILLER_120_2180 ();
 b15zdnd11an1n16x5 FILLER_120_2197 ();
 b15zdnd11an1n08x5 FILLER_120_2213 ();
 b15zdnd11an1n04x5 FILLER_120_2221 ();
 b15zdnd00an1n02x5 FILLER_120_2225 ();
 b15zdnd00an1n01x5 FILLER_120_2227 ();
 b15zdnd11an1n32x5 FILLER_120_2233 ();
 b15zdnd11an1n08x5 FILLER_120_2265 ();
 b15zdnd00an1n02x5 FILLER_120_2273 ();
 b15zdnd00an1n01x5 FILLER_120_2275 ();
 b15zdnd11an1n32x5 FILLER_121_0 ();
 b15zdnd11an1n08x5 FILLER_121_32 ();
 b15zdnd11an1n04x5 FILLER_121_40 ();
 b15zdnd00an1n02x5 FILLER_121_44 ();
 b15zdnd00an1n01x5 FILLER_121_46 ();
 b15zdnd11an1n08x5 FILLER_121_65 ();
 b15zdnd11an1n04x5 FILLER_121_73 ();
 b15zdnd00an1n01x5 FILLER_121_77 ();
 b15zdnd11an1n04x5 FILLER_121_96 ();
 b15zdnd11an1n04x5 FILLER_121_105 ();
 b15zdnd11an1n04x5 FILLER_121_116 ();
 b15zdnd11an1n16x5 FILLER_121_125 ();
 b15zdnd11an1n08x5 FILLER_121_141 ();
 b15zdnd00an1n02x5 FILLER_121_149 ();
 b15zdnd00an1n01x5 FILLER_121_151 ();
 b15zdnd11an1n32x5 FILLER_121_175 ();
 b15zdnd11an1n16x5 FILLER_121_207 ();
 b15zdnd11an1n04x5 FILLER_121_223 ();
 b15zdnd11an1n64x5 FILLER_121_232 ();
 b15zdnd11an1n32x5 FILLER_121_296 ();
 b15zdnd11an1n04x5 FILLER_121_328 ();
 b15zdnd00an1n02x5 FILLER_121_332 ();
 b15zdnd00an1n01x5 FILLER_121_334 ();
 b15zdnd11an1n64x5 FILLER_121_344 ();
 b15zdnd11an1n16x5 FILLER_121_408 ();
 b15zdnd11an1n04x5 FILLER_121_424 ();
 b15zdnd00an1n02x5 FILLER_121_428 ();
 b15zdnd00an1n01x5 FILLER_121_430 ();
 b15zdnd11an1n16x5 FILLER_121_443 ();
 b15zdnd11an1n08x5 FILLER_121_459 ();
 b15zdnd11an1n16x5 FILLER_121_499 ();
 b15zdnd11an1n08x5 FILLER_121_515 ();
 b15zdnd11an1n16x5 FILLER_121_539 ();
 b15zdnd11an1n08x5 FILLER_121_555 ();
 b15zdnd11an1n04x5 FILLER_121_563 ();
 b15zdnd00an1n02x5 FILLER_121_567 ();
 b15zdnd11an1n64x5 FILLER_121_574 ();
 b15zdnd11an1n16x5 FILLER_121_638 ();
 b15zdnd11an1n04x5 FILLER_121_654 ();
 b15zdnd11an1n16x5 FILLER_121_664 ();
 b15zdnd11an1n08x5 FILLER_121_680 ();
 b15zdnd11an1n04x5 FILLER_121_688 ();
 b15zdnd00an1n02x5 FILLER_121_692 ();
 b15zdnd11an1n08x5 FILLER_121_709 ();
 b15zdnd00an1n02x5 FILLER_121_717 ();
 b15zdnd00an1n01x5 FILLER_121_719 ();
 b15zdnd11an1n04x5 FILLER_121_726 ();
 b15zdnd11an1n32x5 FILLER_121_734 ();
 b15zdnd11an1n08x5 FILLER_121_766 ();
 b15zdnd00an1n01x5 FILLER_121_774 ();
 b15zdnd11an1n16x5 FILLER_121_779 ();
 b15zdnd11an1n08x5 FILLER_121_795 ();
 b15zdnd11an1n04x5 FILLER_121_803 ();
 b15zdnd00an1n02x5 FILLER_121_807 ();
 b15zdnd11an1n16x5 FILLER_121_817 ();
 b15zdnd11an1n08x5 FILLER_121_833 ();
 b15zdnd11an1n04x5 FILLER_121_841 ();
 b15zdnd00an1n02x5 FILLER_121_845 ();
 b15zdnd11an1n64x5 FILLER_121_853 ();
 b15zdnd11an1n32x5 FILLER_121_917 ();
 b15zdnd11an1n08x5 FILLER_121_949 ();
 b15zdnd00an1n02x5 FILLER_121_957 ();
 b15zdnd00an1n01x5 FILLER_121_959 ();
 b15zdnd11an1n04x5 FILLER_121_980 ();
 b15zdnd11an1n16x5 FILLER_121_1009 ();
 b15zdnd11an1n04x5 FILLER_121_1025 ();
 b15zdnd00an1n02x5 FILLER_121_1029 ();
 b15zdnd11an1n16x5 FILLER_121_1051 ();
 b15zdnd11an1n04x5 FILLER_121_1067 ();
 b15zdnd00an1n02x5 FILLER_121_1071 ();
 b15zdnd00an1n01x5 FILLER_121_1073 ();
 b15zdnd11an1n08x5 FILLER_121_1094 ();
 b15zdnd11an1n04x5 FILLER_121_1102 ();
 b15zdnd00an1n01x5 FILLER_121_1106 ();
 b15zdnd11an1n04x5 FILLER_121_1127 ();
 b15zdnd11an1n64x5 FILLER_121_1136 ();
 b15zdnd11an1n64x5 FILLER_121_1200 ();
 b15zdnd11an1n64x5 FILLER_121_1271 ();
 b15zdnd11an1n32x5 FILLER_121_1335 ();
 b15zdnd11an1n16x5 FILLER_121_1367 ();
 b15zdnd11an1n08x5 FILLER_121_1383 ();
 b15zdnd00an1n01x5 FILLER_121_1391 ();
 b15zdnd11an1n04x5 FILLER_121_1408 ();
 b15zdnd11an1n64x5 FILLER_121_1422 ();
 b15zdnd11an1n32x5 FILLER_121_1486 ();
 b15zdnd11an1n16x5 FILLER_121_1518 ();
 b15zdnd11an1n08x5 FILLER_121_1534 ();
 b15zdnd11an1n04x5 FILLER_121_1542 ();
 b15zdnd11an1n64x5 FILLER_121_1551 ();
 b15zdnd11an1n08x5 FILLER_121_1615 ();
 b15zdnd00an1n02x5 FILLER_121_1623 ();
 b15zdnd00an1n01x5 FILLER_121_1625 ();
 b15zdnd11an1n64x5 FILLER_121_1632 ();
 b15zdnd11an1n64x5 FILLER_121_1696 ();
 b15zdnd00an1n01x5 FILLER_121_1760 ();
 b15zdnd11an1n04x5 FILLER_121_1781 ();
 b15zdnd00an1n02x5 FILLER_121_1785 ();
 b15zdnd00an1n01x5 FILLER_121_1787 ();
 b15zdnd11an1n64x5 FILLER_121_1795 ();
 b15zdnd11an1n32x5 FILLER_121_1859 ();
 b15zdnd11an1n08x5 FILLER_121_1891 ();
 b15zdnd11an1n04x5 FILLER_121_1899 ();
 b15zdnd11an1n64x5 FILLER_121_1913 ();
 b15zdnd11an1n64x5 FILLER_121_1977 ();
 b15zdnd11an1n04x5 FILLER_121_2041 ();
 b15zdnd00an1n01x5 FILLER_121_2045 ();
 b15zdnd11an1n08x5 FILLER_121_2053 ();
 b15zdnd11an1n04x5 FILLER_121_2061 ();
 b15zdnd00an1n01x5 FILLER_121_2065 ();
 b15zdnd11an1n64x5 FILLER_121_2073 ();
 b15zdnd11an1n04x5 FILLER_121_2137 ();
 b15zdnd00an1n02x5 FILLER_121_2141 ();
 b15zdnd11an1n04x5 FILLER_121_2164 ();
 b15zdnd11an1n16x5 FILLER_121_2200 ();
 b15zdnd11an1n04x5 FILLER_121_2216 ();
 b15zdnd00an1n02x5 FILLER_121_2220 ();
 b15zdnd11an1n32x5 FILLER_121_2242 ();
 b15zdnd11an1n08x5 FILLER_121_2274 ();
 b15zdnd00an1n02x5 FILLER_121_2282 ();
 b15zdnd11an1n64x5 FILLER_122_8 ();
 b15zdnd11an1n64x5 FILLER_122_72 ();
 b15zdnd11an1n08x5 FILLER_122_136 ();
 b15zdnd00an1n02x5 FILLER_122_144 ();
 b15zdnd00an1n01x5 FILLER_122_146 ();
 b15zdnd11an1n64x5 FILLER_122_153 ();
 b15zdnd11an1n08x5 FILLER_122_217 ();
 b15zdnd00an1n02x5 FILLER_122_225 ();
 b15zdnd11an1n32x5 FILLER_122_235 ();
 b15zdnd11an1n04x5 FILLER_122_267 ();
 b15zdnd00an1n02x5 FILLER_122_271 ();
 b15zdnd11an1n04x5 FILLER_122_280 ();
 b15zdnd11an1n32x5 FILLER_122_288 ();
 b15zdnd11an1n64x5 FILLER_122_344 ();
 b15zdnd11an1n32x5 FILLER_122_408 ();
 b15zdnd11an1n08x5 FILLER_122_440 ();
 b15zdnd11an1n04x5 FILLER_122_448 ();
 b15zdnd11an1n32x5 FILLER_122_460 ();
 b15zdnd11an1n16x5 FILLER_122_492 ();
 b15zdnd00an1n02x5 FILLER_122_508 ();
 b15zdnd11an1n08x5 FILLER_122_514 ();
 b15zdnd11an1n04x5 FILLER_122_522 ();
 b15zdnd11an1n16x5 FILLER_122_530 ();
 b15zdnd00an1n02x5 FILLER_122_546 ();
 b15zdnd11an1n04x5 FILLER_122_556 ();
 b15zdnd11an1n16x5 FILLER_122_572 ();
 b15zdnd11an1n04x5 FILLER_122_588 ();
 b15zdnd00an1n01x5 FILLER_122_592 ();
 b15zdnd11an1n32x5 FILLER_122_605 ();
 b15zdnd11an1n16x5 FILLER_122_637 ();
 b15zdnd11an1n04x5 FILLER_122_653 ();
 b15zdnd00an1n02x5 FILLER_122_657 ();
 b15zdnd00an1n01x5 FILLER_122_659 ();
 b15zdnd11an1n08x5 FILLER_122_677 ();
 b15zdnd00an1n02x5 FILLER_122_685 ();
 b15zdnd00an1n01x5 FILLER_122_687 ();
 b15zdnd11an1n16x5 FILLER_122_697 ();
 b15zdnd11an1n04x5 FILLER_122_713 ();
 b15zdnd00an1n01x5 FILLER_122_717 ();
 b15zdnd11an1n32x5 FILLER_122_726 ();
 b15zdnd11an1n08x5 FILLER_122_758 ();
 b15zdnd00an1n01x5 FILLER_122_766 ();
 b15zdnd11an1n04x5 FILLER_122_772 ();
 b15zdnd11an1n08x5 FILLER_122_789 ();
 b15zdnd11an1n64x5 FILLER_122_809 ();
 b15zdnd11an1n16x5 FILLER_122_873 ();
 b15zdnd11an1n08x5 FILLER_122_889 ();
 b15zdnd00an1n02x5 FILLER_122_897 ();
 b15zdnd00an1n01x5 FILLER_122_899 ();
 b15zdnd11an1n32x5 FILLER_122_910 ();
 b15zdnd11an1n04x5 FILLER_122_942 ();
 b15zdnd00an1n02x5 FILLER_122_946 ();
 b15zdnd00an1n01x5 FILLER_122_948 ();
 b15zdnd11an1n04x5 FILLER_122_975 ();
 b15zdnd11an1n64x5 FILLER_122_1019 ();
 b15zdnd11an1n08x5 FILLER_122_1083 ();
 b15zdnd11an1n04x5 FILLER_122_1091 ();
 b15zdnd00an1n02x5 FILLER_122_1095 ();
 b15zdnd00an1n01x5 FILLER_122_1097 ();
 b15zdnd11an1n04x5 FILLER_122_1118 ();
 b15zdnd11an1n16x5 FILLER_122_1142 ();
 b15zdnd00an1n02x5 FILLER_122_1158 ();
 b15zdnd00an1n01x5 FILLER_122_1160 ();
 b15zdnd11an1n16x5 FILLER_122_1192 ();
 b15zdnd11an1n08x5 FILLER_122_1208 ();
 b15zdnd11an1n04x5 FILLER_122_1216 ();
 b15zdnd11an1n32x5 FILLER_122_1241 ();
 b15zdnd00an1n02x5 FILLER_122_1273 ();
 b15zdnd11an1n64x5 FILLER_122_1281 ();
 b15zdnd11an1n64x5 FILLER_122_1345 ();
 b15zdnd11an1n64x5 FILLER_122_1409 ();
 b15zdnd11an1n32x5 FILLER_122_1473 ();
 b15zdnd11an1n08x5 FILLER_122_1505 ();
 b15zdnd00an1n01x5 FILLER_122_1513 ();
 b15zdnd11an1n32x5 FILLER_122_1527 ();
 b15zdnd00an1n02x5 FILLER_122_1559 ();
 b15zdnd00an1n01x5 FILLER_122_1561 ();
 b15zdnd11an1n04x5 FILLER_122_1567 ();
 b15zdnd11an1n32x5 FILLER_122_1584 ();
 b15zdnd11an1n04x5 FILLER_122_1616 ();
 b15zdnd11an1n64x5 FILLER_122_1625 ();
 b15zdnd11an1n04x5 FILLER_122_1689 ();
 b15zdnd00an1n01x5 FILLER_122_1693 ();
 b15zdnd11an1n64x5 FILLER_122_1703 ();
 b15zdnd11an1n32x5 FILLER_122_1767 ();
 b15zdnd11an1n16x5 FILLER_122_1799 ();
 b15zdnd11an1n04x5 FILLER_122_1815 ();
 b15zdnd00an1n02x5 FILLER_122_1819 ();
 b15zdnd11an1n64x5 FILLER_122_1852 ();
 b15zdnd11an1n08x5 FILLER_122_1916 ();
 b15zdnd11an1n04x5 FILLER_122_1924 ();
 b15zdnd11an1n32x5 FILLER_122_1937 ();
 b15zdnd11an1n08x5 FILLER_122_1969 ();
 b15zdnd00an1n01x5 FILLER_122_1977 ();
 b15zdnd11an1n32x5 FILLER_122_2004 ();
 b15zdnd11an1n16x5 FILLER_122_2036 ();
 b15zdnd11an1n04x5 FILLER_122_2052 ();
 b15zdnd00an1n02x5 FILLER_122_2056 ();
 b15zdnd11an1n04x5 FILLER_122_2076 ();
 b15zdnd11an1n64x5 FILLER_122_2084 ();
 b15zdnd11an1n04x5 FILLER_122_2148 ();
 b15zdnd00an1n02x5 FILLER_122_2152 ();
 b15zdnd11an1n64x5 FILLER_122_2162 ();
 b15zdnd11an1n08x5 FILLER_122_2226 ();
 b15zdnd11an1n04x5 FILLER_122_2234 ();
 b15zdnd00an1n02x5 FILLER_122_2238 ();
 b15zdnd11an1n16x5 FILLER_122_2243 ();
 b15zdnd00an1n02x5 FILLER_122_2259 ();
 b15zdnd11an1n08x5 FILLER_122_2265 ();
 b15zdnd00an1n02x5 FILLER_122_2273 ();
 b15zdnd00an1n01x5 FILLER_122_2275 ();
 b15zdnd11an1n64x5 FILLER_123_0 ();
 b15zdnd11an1n64x5 FILLER_123_64 ();
 b15zdnd11an1n16x5 FILLER_123_128 ();
 b15zdnd11an1n08x5 FILLER_123_144 ();
 b15zdnd11an1n04x5 FILLER_123_152 ();
 b15zdnd00an1n01x5 FILLER_123_156 ();
 b15zdnd11an1n16x5 FILLER_123_166 ();
 b15zdnd11an1n04x5 FILLER_123_182 ();
 b15zdnd00an1n02x5 FILLER_123_186 ();
 b15zdnd11an1n64x5 FILLER_123_192 ();
 b15zdnd11an1n08x5 FILLER_123_256 ();
 b15zdnd11an1n04x5 FILLER_123_264 ();
 b15zdnd00an1n02x5 FILLER_123_268 ();
 b15zdnd11an1n08x5 FILLER_123_275 ();
 b15zdnd11an1n64x5 FILLER_123_288 ();
 b15zdnd11an1n64x5 FILLER_123_352 ();
 b15zdnd11an1n16x5 FILLER_123_416 ();
 b15zdnd11an1n08x5 FILLER_123_432 ();
 b15zdnd00an1n01x5 FILLER_123_440 ();
 b15zdnd11an1n16x5 FILLER_123_450 ();
 b15zdnd00an1n02x5 FILLER_123_466 ();
 b15zdnd11an1n04x5 FILLER_123_484 ();
 b15zdnd11an1n04x5 FILLER_123_500 ();
 b15zdnd11an1n64x5 FILLER_123_514 ();
 b15zdnd11an1n08x5 FILLER_123_578 ();
 b15zdnd11an1n04x5 FILLER_123_586 ();
 b15zdnd11an1n16x5 FILLER_123_596 ();
 b15zdnd11an1n08x5 FILLER_123_612 ();
 b15zdnd11an1n04x5 FILLER_123_620 ();
 b15zdnd00an1n01x5 FILLER_123_624 ();
 b15zdnd11an1n04x5 FILLER_123_642 ();
 b15zdnd11an1n64x5 FILLER_123_653 ();
 b15zdnd11an1n16x5 FILLER_123_717 ();
 b15zdnd11an1n08x5 FILLER_123_733 ();
 b15zdnd11an1n04x5 FILLER_123_741 ();
 b15zdnd00an1n02x5 FILLER_123_745 ();
 b15zdnd00an1n01x5 FILLER_123_747 ();
 b15zdnd11an1n32x5 FILLER_123_757 ();
 b15zdnd11an1n08x5 FILLER_123_789 ();
 b15zdnd11an1n16x5 FILLER_123_802 ();
 b15zdnd11an1n08x5 FILLER_123_818 ();
 b15zdnd00an1n02x5 FILLER_123_826 ();
 b15zdnd00an1n01x5 FILLER_123_828 ();
 b15zdnd11an1n08x5 FILLER_123_835 ();
 b15zdnd00an1n02x5 FILLER_123_843 ();
 b15zdnd00an1n01x5 FILLER_123_845 ();
 b15zdnd11an1n04x5 FILLER_123_852 ();
 b15zdnd00an1n01x5 FILLER_123_856 ();
 b15zdnd11an1n04x5 FILLER_123_877 ();
 b15zdnd00an1n02x5 FILLER_123_881 ();
 b15zdnd11an1n04x5 FILLER_123_899 ();
 b15zdnd00an1n01x5 FILLER_123_903 ();
 b15zdnd11an1n64x5 FILLER_123_912 ();
 b15zdnd11an1n32x5 FILLER_123_976 ();
 b15zdnd00an1n02x5 FILLER_123_1008 ();
 b15zdnd11an1n64x5 FILLER_123_1028 ();
 b15zdnd11an1n64x5 FILLER_123_1092 ();
 b15zdnd11an1n32x5 FILLER_123_1156 ();
 b15zdnd11an1n16x5 FILLER_123_1188 ();
 b15zdnd11an1n08x5 FILLER_123_1204 ();
 b15zdnd00an1n02x5 FILLER_123_1212 ();
 b15zdnd11an1n64x5 FILLER_123_1221 ();
 b15zdnd11an1n08x5 FILLER_123_1285 ();
 b15zdnd00an1n01x5 FILLER_123_1293 ();
 b15zdnd11an1n32x5 FILLER_123_1300 ();
 b15zdnd11an1n16x5 FILLER_123_1332 ();
 b15zdnd00an1n02x5 FILLER_123_1348 ();
 b15zdnd11an1n64x5 FILLER_123_1355 ();
 b15zdnd11an1n08x5 FILLER_123_1419 ();
 b15zdnd11an1n04x5 FILLER_123_1427 ();
 b15zdnd11an1n08x5 FILLER_123_1441 ();
 b15zdnd11an1n04x5 FILLER_123_1449 ();
 b15zdnd00an1n02x5 FILLER_123_1453 ();
 b15zdnd11an1n64x5 FILLER_123_1462 ();
 b15zdnd11an1n32x5 FILLER_123_1526 ();
 b15zdnd11an1n16x5 FILLER_123_1558 ();
 b15zdnd00an1n01x5 FILLER_123_1574 ();
 b15zdnd11an1n04x5 FILLER_123_1579 ();
 b15zdnd00an1n01x5 FILLER_123_1583 ();
 b15zdnd11an1n04x5 FILLER_123_1590 ();
 b15zdnd00an1n02x5 FILLER_123_1594 ();
 b15zdnd11an1n04x5 FILLER_123_1614 ();
 b15zdnd00an1n02x5 FILLER_123_1618 ();
 b15zdnd11an1n04x5 FILLER_123_1626 ();
 b15zdnd00an1n02x5 FILLER_123_1630 ();
 b15zdnd00an1n01x5 FILLER_123_1632 ();
 b15zdnd11an1n32x5 FILLER_123_1639 ();
 b15zdnd11an1n16x5 FILLER_123_1671 ();
 b15zdnd11an1n04x5 FILLER_123_1687 ();
 b15zdnd00an1n02x5 FILLER_123_1691 ();
 b15zdnd00an1n01x5 FILLER_123_1693 ();
 b15zdnd11an1n64x5 FILLER_123_1705 ();
 b15zdnd00an1n02x5 FILLER_123_1769 ();
 b15zdnd11an1n16x5 FILLER_123_1785 ();
 b15zdnd00an1n02x5 FILLER_123_1801 ();
 b15zdnd00an1n01x5 FILLER_123_1803 ();
 b15zdnd11an1n08x5 FILLER_123_1809 ();
 b15zdnd00an1n01x5 FILLER_123_1817 ();
 b15zdnd11an1n04x5 FILLER_123_1827 ();
 b15zdnd11an1n08x5 FILLER_123_1847 ();
 b15zdnd00an1n02x5 FILLER_123_1855 ();
 b15zdnd11an1n04x5 FILLER_123_1862 ();
 b15zdnd11an1n04x5 FILLER_123_1873 ();
 b15zdnd11an1n16x5 FILLER_123_1889 ();
 b15zdnd11an1n08x5 FILLER_123_1905 ();
 b15zdnd11an1n04x5 FILLER_123_1913 ();
 b15zdnd00an1n02x5 FILLER_123_1917 ();
 b15zdnd00an1n01x5 FILLER_123_1919 ();
 b15zdnd11an1n08x5 FILLER_123_1936 ();
 b15zdnd11an1n04x5 FILLER_123_1944 ();
 b15zdnd00an1n01x5 FILLER_123_1948 ();
 b15zdnd11an1n32x5 FILLER_123_1975 ();
 b15zdnd11an1n32x5 FILLER_123_2018 ();
 b15zdnd11an1n16x5 FILLER_123_2050 ();
 b15zdnd11an1n08x5 FILLER_123_2066 ();
 b15zdnd11an1n04x5 FILLER_123_2074 ();
 b15zdnd00an1n02x5 FILLER_123_2078 ();
 b15zdnd00an1n01x5 FILLER_123_2080 ();
 b15zdnd11an1n04x5 FILLER_123_2090 ();
 b15zdnd11an1n16x5 FILLER_123_2106 ();
 b15zdnd11an1n04x5 FILLER_123_2122 ();
 b15zdnd11an1n08x5 FILLER_123_2130 ();
 b15zdnd11an1n04x5 FILLER_123_2138 ();
 b15zdnd11an1n64x5 FILLER_123_2162 ();
 b15zdnd11an1n16x5 FILLER_123_2226 ();
 b15zdnd11an1n04x5 FILLER_123_2242 ();
 b15zdnd00an1n01x5 FILLER_123_2246 ();
 b15zdnd11an1n16x5 FILLER_123_2267 ();
 b15zdnd00an1n01x5 FILLER_123_2283 ();
 b15zdnd11an1n32x5 FILLER_124_8 ();
 b15zdnd00an1n02x5 FILLER_124_40 ();
 b15zdnd00an1n01x5 FILLER_124_42 ();
 b15zdnd11an1n04x5 FILLER_124_61 ();
 b15zdnd11an1n16x5 FILLER_124_73 ();
 b15zdnd11an1n08x5 FILLER_124_89 ();
 b15zdnd11an1n04x5 FILLER_124_97 ();
 b15zdnd00an1n02x5 FILLER_124_101 ();
 b15zdnd11an1n04x5 FILLER_124_115 ();
 b15zdnd11an1n32x5 FILLER_124_131 ();
 b15zdnd11an1n08x5 FILLER_124_171 ();
 b15zdnd11an1n04x5 FILLER_124_179 ();
 b15zdnd00an1n02x5 FILLER_124_183 ();
 b15zdnd11an1n32x5 FILLER_124_190 ();
 b15zdnd11an1n04x5 FILLER_124_222 ();
 b15zdnd00an1n02x5 FILLER_124_226 ();
 b15zdnd11an1n32x5 FILLER_124_234 ();
 b15zdnd11an1n16x5 FILLER_124_266 ();
 b15zdnd11an1n08x5 FILLER_124_282 ();
 b15zdnd11an1n04x5 FILLER_124_290 ();
 b15zdnd11an1n04x5 FILLER_124_314 ();
 b15zdnd11an1n08x5 FILLER_124_331 ();
 b15zdnd11an1n04x5 FILLER_124_339 ();
 b15zdnd00an1n02x5 FILLER_124_343 ();
 b15zdnd00an1n01x5 FILLER_124_345 ();
 b15zdnd11an1n04x5 FILLER_124_358 ();
 b15zdnd00an1n02x5 FILLER_124_362 ();
 b15zdnd11an1n64x5 FILLER_124_372 ();
 b15zdnd11an1n64x5 FILLER_124_462 ();
 b15zdnd11an1n64x5 FILLER_124_526 ();
 b15zdnd11an1n32x5 FILLER_124_590 ();
 b15zdnd00an1n02x5 FILLER_124_622 ();
 b15zdnd00an1n01x5 FILLER_124_624 ();
 b15zdnd11an1n16x5 FILLER_124_638 ();
 b15zdnd11an1n08x5 FILLER_124_654 ();
 b15zdnd11an1n32x5 FILLER_124_667 ();
 b15zdnd11an1n16x5 FILLER_124_699 ();
 b15zdnd00an1n02x5 FILLER_124_715 ();
 b15zdnd00an1n01x5 FILLER_124_717 ();
 b15zdnd11an1n16x5 FILLER_124_726 ();
 b15zdnd11an1n04x5 FILLER_124_742 ();
 b15zdnd00an1n01x5 FILLER_124_746 ();
 b15zdnd11an1n32x5 FILLER_124_759 ();
 b15zdnd11an1n04x5 FILLER_124_791 ();
 b15zdnd00an1n02x5 FILLER_124_795 ();
 b15zdnd00an1n01x5 FILLER_124_797 ();
 b15zdnd11an1n32x5 FILLER_124_818 ();
 b15zdnd11an1n08x5 FILLER_124_850 ();
 b15zdnd11an1n04x5 FILLER_124_858 ();
 b15zdnd00an1n02x5 FILLER_124_862 ();
 b15zdnd11an1n04x5 FILLER_124_880 ();
 b15zdnd11an1n64x5 FILLER_124_904 ();
 b15zdnd11an1n16x5 FILLER_124_968 ();
 b15zdnd00an1n01x5 FILLER_124_984 ();
 b15zdnd11an1n64x5 FILLER_124_994 ();
 b15zdnd11an1n32x5 FILLER_124_1058 ();
 b15zdnd11an1n16x5 FILLER_124_1090 ();
 b15zdnd11an1n04x5 FILLER_124_1115 ();
 b15zdnd11an1n64x5 FILLER_124_1145 ();
 b15zdnd11an1n64x5 FILLER_124_1209 ();
 b15zdnd00an1n02x5 FILLER_124_1273 ();
 b15zdnd11an1n04x5 FILLER_124_1288 ();
 b15zdnd11an1n04x5 FILLER_124_1299 ();
 b15zdnd11an1n04x5 FILLER_124_1307 ();
 b15zdnd11an1n16x5 FILLER_124_1316 ();
 b15zdnd11an1n04x5 FILLER_124_1332 ();
 b15zdnd11an1n08x5 FILLER_124_1342 ();
 b15zdnd00an1n01x5 FILLER_124_1350 ();
 b15zdnd11an1n16x5 FILLER_124_1361 ();
 b15zdnd11an1n04x5 FILLER_124_1377 ();
 b15zdnd00an1n02x5 FILLER_124_1381 ();
 b15zdnd00an1n01x5 FILLER_124_1383 ();
 b15zdnd11an1n04x5 FILLER_124_1390 ();
 b15zdnd11an1n08x5 FILLER_124_1400 ();
 b15zdnd00an1n01x5 FILLER_124_1408 ();
 b15zdnd11an1n04x5 FILLER_124_1423 ();
 b15zdnd11an1n08x5 FILLER_124_1443 ();
 b15zdnd11an1n04x5 FILLER_124_1451 ();
 b15zdnd00an1n02x5 FILLER_124_1455 ();
 b15zdnd00an1n01x5 FILLER_124_1457 ();
 b15zdnd11an1n04x5 FILLER_124_1464 ();
 b15zdnd11an1n08x5 FILLER_124_1481 ();
 b15zdnd11an1n04x5 FILLER_124_1489 ();
 b15zdnd00an1n01x5 FILLER_124_1493 ();
 b15zdnd11an1n16x5 FILLER_124_1499 ();
 b15zdnd11an1n08x5 FILLER_124_1522 ();
 b15zdnd00an1n02x5 FILLER_124_1530 ();
 b15zdnd11an1n64x5 FILLER_124_1537 ();
 b15zdnd11an1n16x5 FILLER_124_1601 ();
 b15zdnd11an1n08x5 FILLER_124_1617 ();
 b15zdnd00an1n01x5 FILLER_124_1625 ();
 b15zdnd11an1n04x5 FILLER_124_1640 ();
 b15zdnd11an1n64x5 FILLER_124_1656 ();
 b15zdnd11an1n16x5 FILLER_124_1720 ();
 b15zdnd11an1n08x5 FILLER_124_1736 ();
 b15zdnd11an1n04x5 FILLER_124_1744 ();
 b15zdnd00an1n01x5 FILLER_124_1748 ();
 b15zdnd11an1n16x5 FILLER_124_1780 ();
 b15zdnd11an1n04x5 FILLER_124_1796 ();
 b15zdnd00an1n02x5 FILLER_124_1800 ();
 b15zdnd11an1n64x5 FILLER_124_1806 ();
 b15zdnd11an1n04x5 FILLER_124_1870 ();
 b15zdnd00an1n02x5 FILLER_124_1874 ();
 b15zdnd00an1n01x5 FILLER_124_1876 ();
 b15zdnd11an1n04x5 FILLER_124_1889 ();
 b15zdnd00an1n02x5 FILLER_124_1893 ();
 b15zdnd00an1n01x5 FILLER_124_1895 ();
 b15zdnd11an1n04x5 FILLER_124_1908 ();
 b15zdnd11an1n16x5 FILLER_124_1921 ();
 b15zdnd11an1n08x5 FILLER_124_1937 ();
 b15zdnd11an1n04x5 FILLER_124_1945 ();
 b15zdnd00an1n02x5 FILLER_124_1949 ();
 b15zdnd00an1n01x5 FILLER_124_1951 ();
 b15zdnd11an1n04x5 FILLER_124_1962 ();
 b15zdnd11an1n04x5 FILLER_124_1971 ();
 b15zdnd11an1n16x5 FILLER_124_1982 ();
 b15zdnd11an1n04x5 FILLER_124_1998 ();
 b15zdnd00an1n02x5 FILLER_124_2002 ();
 b15zdnd00an1n01x5 FILLER_124_2004 ();
 b15zdnd11an1n04x5 FILLER_124_2012 ();
 b15zdnd11an1n08x5 FILLER_124_2023 ();
 b15zdnd11an1n04x5 FILLER_124_2031 ();
 b15zdnd00an1n02x5 FILLER_124_2035 ();
 b15zdnd11an1n04x5 FILLER_124_2051 ();
 b15zdnd11an1n16x5 FILLER_124_2064 ();
 b15zdnd00an1n02x5 FILLER_124_2080 ();
 b15zdnd00an1n01x5 FILLER_124_2082 ();
 b15zdnd11an1n16x5 FILLER_124_2099 ();
 b15zdnd11an1n04x5 FILLER_124_2115 ();
 b15zdnd00an1n01x5 FILLER_124_2119 ();
 b15zdnd11an1n04x5 FILLER_124_2150 ();
 b15zdnd00an1n02x5 FILLER_124_2162 ();
 b15zdnd00an1n01x5 FILLER_124_2164 ();
 b15zdnd11an1n64x5 FILLER_124_2177 ();
 b15zdnd11an1n32x5 FILLER_124_2241 ();
 b15zdnd00an1n02x5 FILLER_124_2273 ();
 b15zdnd00an1n01x5 FILLER_124_2275 ();
 b15zdnd11an1n32x5 FILLER_125_0 ();
 b15zdnd11an1n16x5 FILLER_125_32 ();
 b15zdnd11an1n08x5 FILLER_125_48 ();
 b15zdnd00an1n01x5 FILLER_125_56 ();
 b15zdnd11an1n16x5 FILLER_125_89 ();
 b15zdnd00an1n02x5 FILLER_125_105 ();
 b15zdnd11an1n04x5 FILLER_125_114 ();
 b15zdnd11an1n32x5 FILLER_125_139 ();
 b15zdnd11an1n08x5 FILLER_125_171 ();
 b15zdnd11an1n04x5 FILLER_125_179 ();
 b15zdnd00an1n02x5 FILLER_125_183 ();
 b15zdnd11an1n16x5 FILLER_125_192 ();
 b15zdnd11an1n08x5 FILLER_125_208 ();
 b15zdnd11an1n04x5 FILLER_125_216 ();
 b15zdnd00an1n02x5 FILLER_125_220 ();
 b15zdnd00an1n01x5 FILLER_125_222 ();
 b15zdnd11an1n32x5 FILLER_125_230 ();
 b15zdnd00an1n02x5 FILLER_125_262 ();
 b15zdnd11an1n32x5 FILLER_125_272 ();
 b15zdnd00an1n02x5 FILLER_125_304 ();
 b15zdnd00an1n01x5 FILLER_125_306 ();
 b15zdnd11an1n04x5 FILLER_125_327 ();
 b15zdnd00an1n02x5 FILLER_125_331 ();
 b15zdnd00an1n01x5 FILLER_125_333 ();
 b15zdnd11an1n04x5 FILLER_125_351 ();
 b15zdnd11an1n64x5 FILLER_125_365 ();
 b15zdnd11an1n64x5 FILLER_125_429 ();
 b15zdnd11an1n08x5 FILLER_125_493 ();
 b15zdnd00an1n02x5 FILLER_125_501 ();
 b15zdnd11an1n16x5 FILLER_125_506 ();
 b15zdnd11an1n08x5 FILLER_125_522 ();
 b15zdnd11an1n04x5 FILLER_125_530 ();
 b15zdnd00an1n02x5 FILLER_125_534 ();
 b15zdnd11an1n32x5 FILLER_125_546 ();
 b15zdnd11an1n08x5 FILLER_125_578 ();
 b15zdnd00an1n02x5 FILLER_125_586 ();
 b15zdnd11an1n32x5 FILLER_125_592 ();
 b15zdnd00an1n02x5 FILLER_125_624 ();
 b15zdnd11an1n16x5 FILLER_125_639 ();
 b15zdnd11an1n04x5 FILLER_125_655 ();
 b15zdnd11an1n16x5 FILLER_125_674 ();
 b15zdnd00an1n01x5 FILLER_125_690 ();
 b15zdnd11an1n64x5 FILLER_125_696 ();
 b15zdnd11an1n16x5 FILLER_125_760 ();
 b15zdnd11an1n04x5 FILLER_125_776 ();
 b15zdnd00an1n02x5 FILLER_125_780 ();
 b15zdnd00an1n01x5 FILLER_125_782 ();
 b15zdnd11an1n08x5 FILLER_125_795 ();
 b15zdnd11an1n04x5 FILLER_125_803 ();
 b15zdnd00an1n02x5 FILLER_125_807 ();
 b15zdnd00an1n01x5 FILLER_125_809 ();
 b15zdnd11an1n08x5 FILLER_125_819 ();
 b15zdnd00an1n01x5 FILLER_125_827 ();
 b15zdnd11an1n04x5 FILLER_125_837 ();
 b15zdnd11an1n04x5 FILLER_125_846 ();
 b15zdnd00an1n02x5 FILLER_125_850 ();
 b15zdnd11an1n04x5 FILLER_125_872 ();
 b15zdnd11an1n08x5 FILLER_125_894 ();
 b15zdnd00an1n02x5 FILLER_125_902 ();
 b15zdnd00an1n01x5 FILLER_125_904 ();
 b15zdnd11an1n04x5 FILLER_125_931 ();
 b15zdnd11an1n16x5 FILLER_125_955 ();
 b15zdnd11an1n08x5 FILLER_125_971 ();
 b15zdnd00an1n02x5 FILLER_125_979 ();
 b15zdnd00an1n01x5 FILLER_125_981 ();
 b15zdnd11an1n64x5 FILLER_125_991 ();
 b15zdnd11an1n32x5 FILLER_125_1055 ();
 b15zdnd11an1n08x5 FILLER_125_1087 ();
 b15zdnd00an1n02x5 FILLER_125_1095 ();
 b15zdnd11an1n04x5 FILLER_125_1103 ();
 b15zdnd11an1n64x5 FILLER_125_1112 ();
 b15zdnd11an1n16x5 FILLER_125_1176 ();
 b15zdnd11an1n04x5 FILLER_125_1192 ();
 b15zdnd00an1n02x5 FILLER_125_1196 ();
 b15zdnd00an1n01x5 FILLER_125_1198 ();
 b15zdnd11an1n08x5 FILLER_125_1218 ();
 b15zdnd00an1n02x5 FILLER_125_1226 ();
 b15zdnd11an1n32x5 FILLER_125_1233 ();
 b15zdnd11an1n04x5 FILLER_125_1265 ();
 b15zdnd00an1n02x5 FILLER_125_1269 ();
 b15zdnd00an1n01x5 FILLER_125_1271 ();
 b15zdnd11an1n08x5 FILLER_125_1278 ();
 b15zdnd11an1n04x5 FILLER_125_1286 ();
 b15zdnd00an1n01x5 FILLER_125_1290 ();
 b15zdnd11an1n64x5 FILLER_125_1304 ();
 b15zdnd11an1n16x5 FILLER_125_1368 ();
 b15zdnd11an1n08x5 FILLER_125_1384 ();
 b15zdnd11an1n04x5 FILLER_125_1392 ();
 b15zdnd11an1n16x5 FILLER_125_1402 ();
 b15zdnd11an1n08x5 FILLER_125_1418 ();
 b15zdnd00an1n02x5 FILLER_125_1426 ();
 b15zdnd11an1n08x5 FILLER_125_1438 ();
 b15zdnd11an1n04x5 FILLER_125_1446 ();
 b15zdnd00an1n02x5 FILLER_125_1450 ();
 b15zdnd11an1n04x5 FILLER_125_1459 ();
 b15zdnd11an1n32x5 FILLER_125_1467 ();
 b15zdnd11an1n08x5 FILLER_125_1499 ();
 b15zdnd11an1n04x5 FILLER_125_1507 ();
 b15zdnd00an1n01x5 FILLER_125_1511 ();
 b15zdnd11an1n08x5 FILLER_125_1518 ();
 b15zdnd11an1n04x5 FILLER_125_1526 ();
 b15zdnd00an1n01x5 FILLER_125_1530 ();
 b15zdnd11an1n64x5 FILLER_125_1551 ();
 b15zdnd11an1n04x5 FILLER_125_1615 ();
 b15zdnd00an1n01x5 FILLER_125_1619 ();
 b15zdnd11an1n32x5 FILLER_125_1629 ();
 b15zdnd11an1n16x5 FILLER_125_1661 ();
 b15zdnd11an1n08x5 FILLER_125_1677 ();
 b15zdnd00an1n02x5 FILLER_125_1685 ();
 b15zdnd11an1n64x5 FILLER_125_1707 ();
 b15zdnd11an1n16x5 FILLER_125_1771 ();
 b15zdnd11an1n08x5 FILLER_125_1787 ();
 b15zdnd11an1n04x5 FILLER_125_1795 ();
 b15zdnd00an1n02x5 FILLER_125_1799 ();
 b15zdnd00an1n01x5 FILLER_125_1801 ();
 b15zdnd11an1n32x5 FILLER_125_1820 ();
 b15zdnd11an1n08x5 FILLER_125_1852 ();
 b15zdnd11an1n64x5 FILLER_125_1872 ();
 b15zdnd11an1n16x5 FILLER_125_1936 ();
 b15zdnd11an1n08x5 FILLER_125_1952 ();
 b15zdnd00an1n02x5 FILLER_125_1960 ();
 b15zdnd11an1n04x5 FILLER_125_1967 ();
 b15zdnd00an1n02x5 FILLER_125_1971 ();
 b15zdnd11an1n04x5 FILLER_125_1982 ();
 b15zdnd00an1n02x5 FILLER_125_1986 ();
 b15zdnd00an1n01x5 FILLER_125_1988 ();
 b15zdnd11an1n04x5 FILLER_125_1996 ();
 b15zdnd00an1n02x5 FILLER_125_2000 ();
 b15zdnd00an1n01x5 FILLER_125_2002 ();
 b15zdnd11an1n32x5 FILLER_125_2017 ();
 b15zdnd11an1n08x5 FILLER_125_2049 ();
 b15zdnd11an1n04x5 FILLER_125_2083 ();
 b15zdnd11an1n32x5 FILLER_125_2097 ();
 b15zdnd00an1n01x5 FILLER_125_2129 ();
 b15zdnd11an1n08x5 FILLER_125_2145 ();
 b15zdnd11an1n04x5 FILLER_125_2153 ();
 b15zdnd00an1n02x5 FILLER_125_2157 ();
 b15zdnd11an1n16x5 FILLER_125_2170 ();
 b15zdnd11an1n08x5 FILLER_125_2186 ();
 b15zdnd11an1n64x5 FILLER_125_2210 ();
 b15zdnd11an1n04x5 FILLER_125_2274 ();
 b15zdnd00an1n02x5 FILLER_125_2282 ();
 b15zdnd11an1n16x5 FILLER_126_8 ();
 b15zdnd11an1n08x5 FILLER_126_24 ();
 b15zdnd11an1n04x5 FILLER_126_32 ();
 b15zdnd00an1n02x5 FILLER_126_36 ();
 b15zdnd11an1n32x5 FILLER_126_54 ();
 b15zdnd11an1n16x5 FILLER_126_86 ();
 b15zdnd00an1n02x5 FILLER_126_102 ();
 b15zdnd11an1n16x5 FILLER_126_109 ();
 b15zdnd11an1n04x5 FILLER_126_125 ();
 b15zdnd00an1n01x5 FILLER_126_129 ();
 b15zdnd11an1n32x5 FILLER_126_137 ();
 b15zdnd11an1n16x5 FILLER_126_169 ();
 b15zdnd11an1n04x5 FILLER_126_185 ();
 b15zdnd00an1n02x5 FILLER_126_189 ();
 b15zdnd00an1n01x5 FILLER_126_191 ();
 b15zdnd11an1n16x5 FILLER_126_204 ();
 b15zdnd11an1n04x5 FILLER_126_220 ();
 b15zdnd11an1n04x5 FILLER_126_234 ();
 b15zdnd00an1n01x5 FILLER_126_238 ();
 b15zdnd11an1n08x5 FILLER_126_244 ();
 b15zdnd00an1n01x5 FILLER_126_252 ();
 b15zdnd11an1n04x5 FILLER_126_271 ();
 b15zdnd11an1n32x5 FILLER_126_280 ();
 b15zdnd11an1n04x5 FILLER_126_312 ();
 b15zdnd00an1n02x5 FILLER_126_316 ();
 b15zdnd11an1n04x5 FILLER_126_325 ();
 b15zdnd00an1n02x5 FILLER_126_329 ();
 b15zdnd11an1n08x5 FILLER_126_337 ();
 b15zdnd11an1n04x5 FILLER_126_345 ();
 b15zdnd00an1n02x5 FILLER_126_349 ();
 b15zdnd00an1n01x5 FILLER_126_351 ();
 b15zdnd11an1n04x5 FILLER_126_357 ();
 b15zdnd11an1n64x5 FILLER_126_369 ();
 b15zdnd11an1n16x5 FILLER_126_433 ();
 b15zdnd11an1n08x5 FILLER_126_449 ();
 b15zdnd00an1n02x5 FILLER_126_457 ();
 b15zdnd11an1n16x5 FILLER_126_472 ();
 b15zdnd00an1n02x5 FILLER_126_488 ();
 b15zdnd00an1n01x5 FILLER_126_490 ();
 b15zdnd11an1n04x5 FILLER_126_497 ();
 b15zdnd11an1n16x5 FILLER_126_515 ();
 b15zdnd00an1n02x5 FILLER_126_531 ();
 b15zdnd00an1n01x5 FILLER_126_533 ();
 b15zdnd11an1n08x5 FILLER_126_541 ();
 b15zdnd11an1n04x5 FILLER_126_549 ();
 b15zdnd11an1n08x5 FILLER_126_573 ();
 b15zdnd11an1n32x5 FILLER_126_602 ();
 b15zdnd11an1n16x5 FILLER_126_634 ();
 b15zdnd11an1n08x5 FILLER_126_650 ();
 b15zdnd00an1n01x5 FILLER_126_658 ();
 b15zdnd11an1n16x5 FILLER_126_664 ();
 b15zdnd00an1n01x5 FILLER_126_680 ();
 b15zdnd11an1n16x5 FILLER_126_697 ();
 b15zdnd11an1n04x5 FILLER_126_713 ();
 b15zdnd00an1n01x5 FILLER_126_717 ();
 b15zdnd00an1n02x5 FILLER_126_726 ();
 b15zdnd11an1n32x5 FILLER_126_733 ();
 b15zdnd11an1n16x5 FILLER_126_765 ();
 b15zdnd00an1n02x5 FILLER_126_781 ();
 b15zdnd00an1n01x5 FILLER_126_783 ();
 b15zdnd11an1n08x5 FILLER_126_793 ();
 b15zdnd11an1n04x5 FILLER_126_801 ();
 b15zdnd00an1n02x5 FILLER_126_805 ();
 b15zdnd00an1n01x5 FILLER_126_807 ();
 b15zdnd11an1n08x5 FILLER_126_824 ();
 b15zdnd11an1n04x5 FILLER_126_832 ();
 b15zdnd00an1n02x5 FILLER_126_836 ();
 b15zdnd00an1n01x5 FILLER_126_838 ();
 b15zdnd11an1n16x5 FILLER_126_845 ();
 b15zdnd11an1n08x5 FILLER_126_861 ();
 b15zdnd11an1n04x5 FILLER_126_869 ();
 b15zdnd11an1n32x5 FILLER_126_878 ();
 b15zdnd11an1n16x5 FILLER_126_910 ();
 b15zdnd11an1n08x5 FILLER_126_926 ();
 b15zdnd11an1n08x5 FILLER_126_939 ();
 b15zdnd11an1n04x5 FILLER_126_947 ();
 b15zdnd00an1n02x5 FILLER_126_951 ();
 b15zdnd11an1n08x5 FILLER_126_956 ();
 b15zdnd11an1n04x5 FILLER_126_964 ();
 b15zdnd00an1n01x5 FILLER_126_968 ();
 b15zdnd11an1n16x5 FILLER_126_980 ();
 b15zdnd11an1n04x5 FILLER_126_996 ();
 b15zdnd00an1n02x5 FILLER_126_1000 ();
 b15zdnd11an1n04x5 FILLER_126_1033 ();
 b15zdnd11an1n32x5 FILLER_126_1060 ();
 b15zdnd00an1n02x5 FILLER_126_1092 ();
 b15zdnd11an1n16x5 FILLER_126_1114 ();
 b15zdnd00an1n02x5 FILLER_126_1130 ();
 b15zdnd11an1n16x5 FILLER_126_1153 ();
 b15zdnd11an1n04x5 FILLER_126_1169 ();
 b15zdnd00an1n01x5 FILLER_126_1173 ();
 b15zdnd11an1n04x5 FILLER_126_1205 ();
 b15zdnd11an1n04x5 FILLER_126_1215 ();
 b15zdnd11an1n64x5 FILLER_126_1231 ();
 b15zdnd11an1n64x5 FILLER_126_1295 ();
 b15zdnd11an1n16x5 FILLER_126_1359 ();
 b15zdnd00an1n02x5 FILLER_126_1375 ();
 b15zdnd00an1n01x5 FILLER_126_1377 ();
 b15zdnd11an1n16x5 FILLER_126_1382 ();
 b15zdnd00an1n02x5 FILLER_126_1398 ();
 b15zdnd11an1n32x5 FILLER_126_1404 ();
 b15zdnd11an1n08x5 FILLER_126_1436 ();
 b15zdnd11an1n04x5 FILLER_126_1444 ();
 b15zdnd00an1n02x5 FILLER_126_1448 ();
 b15zdnd00an1n01x5 FILLER_126_1450 ();
 b15zdnd11an1n32x5 FILLER_126_1455 ();
 b15zdnd11an1n16x5 FILLER_126_1487 ();
 b15zdnd11an1n08x5 FILLER_126_1503 ();
 b15zdnd11an1n04x5 FILLER_126_1511 ();
 b15zdnd00an1n01x5 FILLER_126_1515 ();
 b15zdnd11an1n08x5 FILLER_126_1526 ();
 b15zdnd11an1n32x5 FILLER_126_1538 ();
 b15zdnd11an1n08x5 FILLER_126_1570 ();
 b15zdnd00an1n01x5 FILLER_126_1578 ();
 b15zdnd11an1n64x5 FILLER_126_1590 ();
 b15zdnd11an1n64x5 FILLER_126_1654 ();
 b15zdnd11an1n32x5 FILLER_126_1718 ();
 b15zdnd11an1n16x5 FILLER_126_1750 ();
 b15zdnd11an1n08x5 FILLER_126_1766 ();
 b15zdnd00an1n01x5 FILLER_126_1774 ();
 b15zdnd11an1n64x5 FILLER_126_1786 ();
 b15zdnd11an1n64x5 FILLER_126_1850 ();
 b15zdnd11an1n64x5 FILLER_126_1914 ();
 b15zdnd11an1n32x5 FILLER_126_1978 ();
 b15zdnd11an1n16x5 FILLER_126_2010 ();
 b15zdnd00an1n01x5 FILLER_126_2026 ();
 b15zdnd11an1n04x5 FILLER_126_2053 ();
 b15zdnd11an1n64x5 FILLER_126_2062 ();
 b15zdnd11an1n16x5 FILLER_126_2126 ();
 b15zdnd11an1n08x5 FILLER_126_2142 ();
 b15zdnd11an1n04x5 FILLER_126_2150 ();
 b15zdnd11an1n16x5 FILLER_126_2162 ();
 b15zdnd11an1n08x5 FILLER_126_2178 ();
 b15zdnd00an1n02x5 FILLER_126_2186 ();
 b15zdnd00an1n01x5 FILLER_126_2188 ();
 b15zdnd11an1n32x5 FILLER_126_2215 ();
 b15zdnd11an1n04x5 FILLER_126_2247 ();
 b15zdnd00an1n02x5 FILLER_126_2251 ();
 b15zdnd11an1n16x5 FILLER_126_2258 ();
 b15zdnd00an1n02x5 FILLER_126_2274 ();
 b15zdnd11an1n64x5 FILLER_127_0 ();
 b15zdnd11an1n32x5 FILLER_127_64 ();
 b15zdnd11an1n08x5 FILLER_127_96 ();
 b15zdnd00an1n02x5 FILLER_127_104 ();
 b15zdnd00an1n01x5 FILLER_127_106 ();
 b15zdnd11an1n16x5 FILLER_127_113 ();
 b15zdnd11an1n08x5 FILLER_127_129 ();
 b15zdnd00an1n01x5 FILLER_127_137 ();
 b15zdnd11an1n04x5 FILLER_127_145 ();
 b15zdnd11an1n08x5 FILLER_127_167 ();
 b15zdnd11an1n04x5 FILLER_127_175 ();
 b15zdnd00an1n02x5 FILLER_127_179 ();
 b15zdnd11an1n04x5 FILLER_127_186 ();
 b15zdnd11an1n08x5 FILLER_127_196 ();
 b15zdnd11an1n04x5 FILLER_127_204 ();
 b15zdnd11an1n64x5 FILLER_127_220 ();
 b15zdnd11an1n16x5 FILLER_127_284 ();
 b15zdnd11an1n04x5 FILLER_127_300 ();
 b15zdnd00an1n02x5 FILLER_127_304 ();
 b15zdnd00an1n01x5 FILLER_127_306 ();
 b15zdnd11an1n32x5 FILLER_127_327 ();
 b15zdnd00an1n02x5 FILLER_127_359 ();
 b15zdnd00an1n01x5 FILLER_127_361 ();
 b15zdnd11an1n64x5 FILLER_127_370 ();
 b15zdnd11an1n16x5 FILLER_127_434 ();
 b15zdnd11an1n04x5 FILLER_127_466 ();
 b15zdnd11an1n04x5 FILLER_127_491 ();
 b15zdnd11an1n16x5 FILLER_127_507 ();
 b15zdnd00an1n01x5 FILLER_127_523 ();
 b15zdnd11an1n08x5 FILLER_127_540 ();
 b15zdnd11an1n04x5 FILLER_127_548 ();
 b15zdnd11an1n04x5 FILLER_127_556 ();
 b15zdnd11an1n32x5 FILLER_127_573 ();
 b15zdnd00an1n02x5 FILLER_127_605 ();
 b15zdnd11an1n16x5 FILLER_127_625 ();
 b15zdnd11an1n08x5 FILLER_127_641 ();
 b15zdnd00an1n01x5 FILLER_127_649 ();
 b15zdnd11an1n32x5 FILLER_127_656 ();
 b15zdnd11an1n16x5 FILLER_127_688 ();
 b15zdnd11an1n08x5 FILLER_127_704 ();
 b15zdnd00an1n01x5 FILLER_127_712 ();
 b15zdnd11an1n04x5 FILLER_127_720 ();
 b15zdnd11an1n04x5 FILLER_127_734 ();
 b15zdnd11an1n04x5 FILLER_127_745 ();
 b15zdnd11an1n04x5 FILLER_127_754 ();
 b15zdnd11an1n16x5 FILLER_127_778 ();
 b15zdnd00an1n01x5 FILLER_127_794 ();
 b15zdnd11an1n32x5 FILLER_127_807 ();
 b15zdnd11an1n08x5 FILLER_127_839 ();
 b15zdnd11an1n04x5 FILLER_127_847 ();
 b15zdnd00an1n01x5 FILLER_127_851 ();
 b15zdnd11an1n04x5 FILLER_127_870 ();
 b15zdnd00an1n01x5 FILLER_127_874 ();
 b15zdnd11an1n04x5 FILLER_127_901 ();
 b15zdnd11an1n04x5 FILLER_127_931 ();
 b15zdnd11an1n64x5 FILLER_127_939 ();
 b15zdnd11an1n64x5 FILLER_127_1003 ();
 b15zdnd11an1n64x5 FILLER_127_1067 ();
 b15zdnd11an1n32x5 FILLER_127_1131 ();
 b15zdnd00an1n01x5 FILLER_127_1163 ();
 b15zdnd11an1n32x5 FILLER_127_1175 ();
 b15zdnd11an1n16x5 FILLER_127_1207 ();
 b15zdnd11an1n32x5 FILLER_127_1227 ();
 b15zdnd11an1n04x5 FILLER_127_1259 ();
 b15zdnd00an1n02x5 FILLER_127_1263 ();
 b15zdnd11an1n04x5 FILLER_127_1270 ();
 b15zdnd11an1n64x5 FILLER_127_1280 ();
 b15zdnd00an1n02x5 FILLER_127_1344 ();
 b15zdnd11an1n16x5 FILLER_127_1361 ();
 b15zdnd11an1n04x5 FILLER_127_1377 ();
 b15zdnd00an1n02x5 FILLER_127_1381 ();
 b15zdnd11an1n04x5 FILLER_127_1393 ();
 b15zdnd11an1n16x5 FILLER_127_1402 ();
 b15zdnd11an1n08x5 FILLER_127_1418 ();
 b15zdnd00an1n02x5 FILLER_127_1426 ();
 b15zdnd11an1n08x5 FILLER_127_1434 ();
 b15zdnd11an1n04x5 FILLER_127_1442 ();
 b15zdnd00an1n02x5 FILLER_127_1446 ();
 b15zdnd11an1n32x5 FILLER_127_1456 ();
 b15zdnd11an1n16x5 FILLER_127_1488 ();
 b15zdnd11an1n08x5 FILLER_127_1504 ();
 b15zdnd00an1n01x5 FILLER_127_1512 ();
 b15zdnd11an1n08x5 FILLER_127_1527 ();
 b15zdnd11an1n32x5 FILLER_127_1540 ();
 b15zdnd11an1n08x5 FILLER_127_1572 ();
 b15zdnd00an1n02x5 FILLER_127_1580 ();
 b15zdnd00an1n01x5 FILLER_127_1582 ();
 b15zdnd11an1n64x5 FILLER_127_1587 ();
 b15zdnd11an1n32x5 FILLER_127_1651 ();
 b15zdnd11an1n16x5 FILLER_127_1683 ();
 b15zdnd11an1n04x5 FILLER_127_1699 ();
 b15zdnd00an1n02x5 FILLER_127_1703 ();
 b15zdnd11an1n32x5 FILLER_127_1716 ();
 b15zdnd11an1n04x5 FILLER_127_1748 ();
 b15zdnd00an1n02x5 FILLER_127_1752 ();
 b15zdnd11an1n04x5 FILLER_127_1786 ();
 b15zdnd11an1n04x5 FILLER_127_1798 ();
 b15zdnd11an1n32x5 FILLER_127_1818 ();
 b15zdnd11an1n16x5 FILLER_127_1850 ();
 b15zdnd11an1n04x5 FILLER_127_1872 ();
 b15zdnd11an1n16x5 FILLER_127_1881 ();
 b15zdnd00an1n01x5 FILLER_127_1897 ();
 b15zdnd11an1n16x5 FILLER_127_1911 ();
 b15zdnd11an1n08x5 FILLER_127_1927 ();
 b15zdnd11an1n08x5 FILLER_127_1940 ();
 b15zdnd11an1n04x5 FILLER_127_1948 ();
 b15zdnd11an1n64x5 FILLER_127_1956 ();
 b15zdnd11an1n32x5 FILLER_127_2020 ();
 b15zdnd11an1n16x5 FILLER_127_2052 ();
 b15zdnd11an1n08x5 FILLER_127_2068 ();
 b15zdnd11an1n04x5 FILLER_127_2076 ();
 b15zdnd00an1n01x5 FILLER_127_2080 ();
 b15zdnd11an1n32x5 FILLER_127_2095 ();
 b15zdnd11an1n16x5 FILLER_127_2127 ();
 b15zdnd11an1n08x5 FILLER_127_2143 ();
 b15zdnd11an1n04x5 FILLER_127_2151 ();
 b15zdnd00an1n02x5 FILLER_127_2155 ();
 b15zdnd00an1n01x5 FILLER_127_2157 ();
 b15zdnd11an1n04x5 FILLER_127_2189 ();
 b15zdnd11an1n32x5 FILLER_127_2216 ();
 b15zdnd00an1n02x5 FILLER_127_2248 ();
 b15zdnd00an1n01x5 FILLER_127_2250 ();
 b15zdnd11an1n08x5 FILLER_127_2271 ();
 b15zdnd11an1n04x5 FILLER_127_2279 ();
 b15zdnd00an1n01x5 FILLER_127_2283 ();
 b15zdnd11an1n16x5 FILLER_128_8 ();
 b15zdnd11an1n08x5 FILLER_128_24 ();
 b15zdnd11an1n04x5 FILLER_128_32 ();
 b15zdnd00an1n02x5 FILLER_128_36 ();
 b15zdnd00an1n01x5 FILLER_128_38 ();
 b15zdnd11an1n16x5 FILLER_128_57 ();
 b15zdnd11an1n04x5 FILLER_128_73 ();
 b15zdnd00an1n02x5 FILLER_128_77 ();
 b15zdnd11an1n16x5 FILLER_128_91 ();
 b15zdnd11an1n04x5 FILLER_128_107 ();
 b15zdnd00an1n02x5 FILLER_128_111 ();
 b15zdnd00an1n01x5 FILLER_128_113 ();
 b15zdnd11an1n32x5 FILLER_128_118 ();
 b15zdnd00an1n01x5 FILLER_128_150 ();
 b15zdnd11an1n04x5 FILLER_128_156 ();
 b15zdnd00an1n02x5 FILLER_128_160 ();
 b15zdnd00an1n01x5 FILLER_128_162 ();
 b15zdnd11an1n04x5 FILLER_128_175 ();
 b15zdnd11an1n64x5 FILLER_128_186 ();
 b15zdnd00an1n02x5 FILLER_128_250 ();
 b15zdnd11an1n16x5 FILLER_128_256 ();
 b15zdnd11an1n08x5 FILLER_128_272 ();
 b15zdnd00an1n02x5 FILLER_128_280 ();
 b15zdnd00an1n01x5 FILLER_128_282 ();
 b15zdnd11an1n04x5 FILLER_128_290 ();
 b15zdnd11an1n04x5 FILLER_128_306 ();
 b15zdnd11an1n64x5 FILLER_128_323 ();
 b15zdnd11an1n64x5 FILLER_128_387 ();
 b15zdnd11an1n16x5 FILLER_128_451 ();
 b15zdnd11an1n04x5 FILLER_128_467 ();
 b15zdnd00an1n02x5 FILLER_128_471 ();
 b15zdnd11an1n04x5 FILLER_128_494 ();
 b15zdnd11an1n16x5 FILLER_128_514 ();
 b15zdnd11an1n08x5 FILLER_128_540 ();
 b15zdnd11an1n04x5 FILLER_128_548 ();
 b15zdnd11an1n16x5 FILLER_128_558 ();
 b15zdnd11an1n08x5 FILLER_128_574 ();
 b15zdnd11an1n04x5 FILLER_128_582 ();
 b15zdnd00an1n02x5 FILLER_128_586 ();
 b15zdnd00an1n01x5 FILLER_128_588 ();
 b15zdnd11an1n08x5 FILLER_128_602 ();
 b15zdnd11an1n04x5 FILLER_128_610 ();
 b15zdnd00an1n02x5 FILLER_128_614 ();
 b15zdnd00an1n01x5 FILLER_128_616 ();
 b15zdnd11an1n16x5 FILLER_128_630 ();
 b15zdnd11an1n08x5 FILLER_128_646 ();
 b15zdnd11an1n04x5 FILLER_128_654 ();
 b15zdnd11an1n16x5 FILLER_128_662 ();
 b15zdnd11an1n08x5 FILLER_128_678 ();
 b15zdnd11an1n04x5 FILLER_128_686 ();
 b15zdnd00an1n01x5 FILLER_128_690 ();
 b15zdnd11an1n08x5 FILLER_128_705 ();
 b15zdnd11an1n04x5 FILLER_128_713 ();
 b15zdnd00an1n01x5 FILLER_128_717 ();
 b15zdnd11an1n16x5 FILLER_128_726 ();
 b15zdnd11an1n08x5 FILLER_128_742 ();
 b15zdnd00an1n01x5 FILLER_128_750 ();
 b15zdnd11an1n08x5 FILLER_128_764 ();
 b15zdnd11an1n04x5 FILLER_128_772 ();
 b15zdnd00an1n02x5 FILLER_128_776 ();
 b15zdnd00an1n01x5 FILLER_128_778 ();
 b15zdnd11an1n32x5 FILLER_128_795 ();
 b15zdnd11an1n64x5 FILLER_128_850 ();
 b15zdnd11an1n32x5 FILLER_128_914 ();
 b15zdnd11an1n16x5 FILLER_128_946 ();
 b15zdnd11an1n08x5 FILLER_128_962 ();
 b15zdnd00an1n02x5 FILLER_128_970 ();
 b15zdnd00an1n01x5 FILLER_128_972 ();
 b15zdnd11an1n32x5 FILLER_128_982 ();
 b15zdnd11an1n16x5 FILLER_128_1014 ();
 b15zdnd11an1n04x5 FILLER_128_1030 ();
 b15zdnd00an1n02x5 FILLER_128_1034 ();
 b15zdnd00an1n01x5 FILLER_128_1036 ();
 b15zdnd11an1n64x5 FILLER_128_1046 ();
 b15zdnd11an1n32x5 FILLER_128_1110 ();
 b15zdnd11an1n08x5 FILLER_128_1142 ();
 b15zdnd11an1n04x5 FILLER_128_1150 ();
 b15zdnd11an1n16x5 FILLER_128_1174 ();
 b15zdnd11an1n08x5 FILLER_128_1190 ();
 b15zdnd00an1n02x5 FILLER_128_1198 ();
 b15zdnd00an1n01x5 FILLER_128_1200 ();
 b15zdnd11an1n04x5 FILLER_128_1206 ();
 b15zdnd11an1n32x5 FILLER_128_1217 ();
 b15zdnd11an1n16x5 FILLER_128_1249 ();
 b15zdnd11an1n04x5 FILLER_128_1265 ();
 b15zdnd00an1n02x5 FILLER_128_1269 ();
 b15zdnd11an1n64x5 FILLER_128_1277 ();
 b15zdnd11an1n64x5 FILLER_128_1341 ();
 b15zdnd11an1n64x5 FILLER_128_1405 ();
 b15zdnd11an1n32x5 FILLER_128_1469 ();
 b15zdnd11an1n08x5 FILLER_128_1501 ();
 b15zdnd11an1n04x5 FILLER_128_1509 ();
 b15zdnd11an1n32x5 FILLER_128_1518 ();
 b15zdnd11an1n04x5 FILLER_128_1550 ();
 b15zdnd11an1n32x5 FILLER_128_1563 ();
 b15zdnd11an1n08x5 FILLER_128_1595 ();
 b15zdnd11an1n04x5 FILLER_128_1603 ();
 b15zdnd11an1n04x5 FILLER_128_1620 ();
 b15zdnd11an1n64x5 FILLER_128_1634 ();
 b15zdnd11an1n08x5 FILLER_128_1698 ();
 b15zdnd00an1n02x5 FILLER_128_1706 ();
 b15zdnd00an1n01x5 FILLER_128_1708 ();
 b15zdnd11an1n16x5 FILLER_128_1718 ();
 b15zdnd11an1n08x5 FILLER_128_1734 ();
 b15zdnd11an1n04x5 FILLER_128_1742 ();
 b15zdnd00an1n02x5 FILLER_128_1746 ();
 b15zdnd00an1n01x5 FILLER_128_1748 ();
 b15zdnd11an1n04x5 FILLER_128_1767 ();
 b15zdnd00an1n02x5 FILLER_128_1771 ();
 b15zdnd00an1n01x5 FILLER_128_1773 ();
 b15zdnd11an1n08x5 FILLER_128_1795 ();
 b15zdnd11an1n04x5 FILLER_128_1803 ();
 b15zdnd00an1n02x5 FILLER_128_1807 ();
 b15zdnd00an1n01x5 FILLER_128_1809 ();
 b15zdnd11an1n04x5 FILLER_128_1816 ();
 b15zdnd11an1n32x5 FILLER_128_1826 ();
 b15zdnd11an1n04x5 FILLER_128_1858 ();
 b15zdnd00an1n02x5 FILLER_128_1862 ();
 b15zdnd11an1n08x5 FILLER_128_1871 ();
 b15zdnd11an1n16x5 FILLER_128_1884 ();
 b15zdnd11an1n04x5 FILLER_128_1900 ();
 b15zdnd00an1n02x5 FILLER_128_1904 ();
 b15zdnd11an1n16x5 FILLER_128_1920 ();
 b15zdnd11an1n04x5 FILLER_128_1936 ();
 b15zdnd11an1n08x5 FILLER_128_1950 ();
 b15zdnd00an1n01x5 FILLER_128_1958 ();
 b15zdnd11an1n32x5 FILLER_128_1970 ();
 b15zdnd11an1n04x5 FILLER_128_2002 ();
 b15zdnd00an1n02x5 FILLER_128_2006 ();
 b15zdnd00an1n01x5 FILLER_128_2008 ();
 b15zdnd11an1n16x5 FILLER_128_2014 ();
 b15zdnd11an1n04x5 FILLER_128_2030 ();
 b15zdnd00an1n02x5 FILLER_128_2034 ();
 b15zdnd00an1n01x5 FILLER_128_2036 ();
 b15zdnd11an1n16x5 FILLER_128_2041 ();
 b15zdnd00an1n01x5 FILLER_128_2057 ();
 b15zdnd11an1n08x5 FILLER_128_2072 ();
 b15zdnd11an1n04x5 FILLER_128_2080 ();
 b15zdnd11an1n04x5 FILLER_128_2091 ();
 b15zdnd11an1n04x5 FILLER_128_2111 ();
 b15zdnd11an1n16x5 FILLER_128_2135 ();
 b15zdnd00an1n02x5 FILLER_128_2151 ();
 b15zdnd00an1n01x5 FILLER_128_2153 ();
 b15zdnd11an1n64x5 FILLER_128_2162 ();
 b15zdnd11an1n32x5 FILLER_128_2226 ();
 b15zdnd00an1n01x5 FILLER_128_2258 ();
 b15zdnd11an1n08x5 FILLER_128_2263 ();
 b15zdnd11an1n04x5 FILLER_128_2271 ();
 b15zdnd00an1n01x5 FILLER_128_2275 ();
 b15zdnd11an1n32x5 FILLER_129_0 ();
 b15zdnd00an1n02x5 FILLER_129_32 ();
 b15zdnd11an1n08x5 FILLER_129_39 ();
 b15zdnd11an1n04x5 FILLER_129_47 ();
 b15zdnd00an1n02x5 FILLER_129_51 ();
 b15zdnd00an1n01x5 FILLER_129_53 ();
 b15zdnd11an1n08x5 FILLER_129_61 ();
 b15zdnd00an1n02x5 FILLER_129_69 ();
 b15zdnd11an1n64x5 FILLER_129_81 ();
 b15zdnd11an1n04x5 FILLER_129_145 ();
 b15zdnd00an1n02x5 FILLER_129_149 ();
 b15zdnd00an1n01x5 FILLER_129_151 ();
 b15zdnd11an1n32x5 FILLER_129_165 ();
 b15zdnd11an1n16x5 FILLER_129_197 ();
 b15zdnd00an1n02x5 FILLER_129_213 ();
 b15zdnd11an1n16x5 FILLER_129_226 ();
 b15zdnd11an1n08x5 FILLER_129_242 ();
 b15zdnd00an1n01x5 FILLER_129_250 ();
 b15zdnd11an1n16x5 FILLER_129_258 ();
 b15zdnd11an1n04x5 FILLER_129_284 ();
 b15zdnd11an1n04x5 FILLER_129_304 ();
 b15zdnd00an1n02x5 FILLER_129_308 ();
 b15zdnd11an1n08x5 FILLER_129_314 ();
 b15zdnd00an1n02x5 FILLER_129_322 ();
 b15zdnd11an1n04x5 FILLER_129_341 ();
 b15zdnd11an1n32x5 FILLER_129_363 ();
 b15zdnd11an1n16x5 FILLER_129_395 ();
 b15zdnd11an1n08x5 FILLER_129_411 ();
 b15zdnd11an1n04x5 FILLER_129_419 ();
 b15zdnd00an1n01x5 FILLER_129_423 ();
 b15zdnd11an1n08x5 FILLER_129_429 ();
 b15zdnd11an1n04x5 FILLER_129_437 ();
 b15zdnd00an1n02x5 FILLER_129_441 ();
 b15zdnd00an1n01x5 FILLER_129_443 ();
 b15zdnd11an1n64x5 FILLER_129_451 ();
 b15zdnd11an1n64x5 FILLER_129_515 ();
 b15zdnd11an1n32x5 FILLER_129_579 ();
 b15zdnd00an1n01x5 FILLER_129_611 ();
 b15zdnd11an1n32x5 FILLER_129_619 ();
 b15zdnd11an1n08x5 FILLER_129_651 ();
 b15zdnd11an1n64x5 FILLER_129_669 ();
 b15zdnd11an1n16x5 FILLER_129_733 ();
 b15zdnd11an1n08x5 FILLER_129_749 ();
 b15zdnd11an1n64x5 FILLER_129_767 ();
 b15zdnd11an1n16x5 FILLER_129_831 ();
 b15zdnd11an1n32x5 FILLER_129_873 ();
 b15zdnd11an1n04x5 FILLER_129_905 ();
 b15zdnd11an1n64x5 FILLER_129_929 ();
 b15zdnd11an1n64x5 FILLER_129_993 ();
 b15zdnd11an1n64x5 FILLER_129_1057 ();
 b15zdnd11an1n64x5 FILLER_129_1121 ();
 b15zdnd11an1n08x5 FILLER_129_1185 ();
 b15zdnd00an1n01x5 FILLER_129_1193 ();
 b15zdnd11an1n08x5 FILLER_129_1201 ();
 b15zdnd00an1n02x5 FILLER_129_1209 ();
 b15zdnd11an1n32x5 FILLER_129_1218 ();
 b15zdnd11an1n04x5 FILLER_129_1250 ();
 b15zdnd00an1n02x5 FILLER_129_1254 ();
 b15zdnd00an1n01x5 FILLER_129_1256 ();
 b15zdnd11an1n04x5 FILLER_129_1262 ();
 b15zdnd11an1n08x5 FILLER_129_1281 ();
 b15zdnd00an1n02x5 FILLER_129_1289 ();
 b15zdnd00an1n01x5 FILLER_129_1291 ();
 b15zdnd11an1n04x5 FILLER_129_1301 ();
 b15zdnd11an1n04x5 FILLER_129_1317 ();
 b15zdnd11an1n16x5 FILLER_129_1325 ();
 b15zdnd11an1n08x5 FILLER_129_1341 ();
 b15zdnd11an1n64x5 FILLER_129_1355 ();
 b15zdnd11an1n64x5 FILLER_129_1419 ();
 b15zdnd11an1n04x5 FILLER_129_1483 ();
 b15zdnd00an1n02x5 FILLER_129_1487 ();
 b15zdnd11an1n16x5 FILLER_129_1510 ();
 b15zdnd11an1n08x5 FILLER_129_1526 ();
 b15zdnd00an1n02x5 FILLER_129_1534 ();
 b15zdnd11an1n04x5 FILLER_129_1541 ();
 b15zdnd11an1n32x5 FILLER_129_1559 ();
 b15zdnd00an1n01x5 FILLER_129_1591 ();
 b15zdnd11an1n04x5 FILLER_129_1596 ();
 b15zdnd00an1n02x5 FILLER_129_1600 ();
 b15zdnd00an1n01x5 FILLER_129_1602 ();
 b15zdnd11an1n64x5 FILLER_129_1619 ();
 b15zdnd11an1n32x5 FILLER_129_1683 ();
 b15zdnd11an1n04x5 FILLER_129_1715 ();
 b15zdnd00an1n02x5 FILLER_129_1719 ();
 b15zdnd00an1n01x5 FILLER_129_1721 ();
 b15zdnd11an1n32x5 FILLER_129_1742 ();
 b15zdnd11an1n16x5 FILLER_129_1774 ();
 b15zdnd00an1n02x5 FILLER_129_1790 ();
 b15zdnd00an1n01x5 FILLER_129_1792 ();
 b15zdnd11an1n08x5 FILLER_129_1825 ();
 b15zdnd11an1n64x5 FILLER_129_1845 ();
 b15zdnd11an1n64x5 FILLER_129_1909 ();
 b15zdnd11an1n04x5 FILLER_129_1973 ();
 b15zdnd00an1n01x5 FILLER_129_1977 ();
 b15zdnd11an1n04x5 FILLER_129_1984 ();
 b15zdnd11an1n08x5 FILLER_129_1994 ();
 b15zdnd11an1n04x5 FILLER_129_2002 ();
 b15zdnd11an1n04x5 FILLER_129_2013 ();
 b15zdnd11an1n16x5 FILLER_129_2023 ();
 b15zdnd11an1n08x5 FILLER_129_2039 ();
 b15zdnd11an1n08x5 FILLER_129_2055 ();
 b15zdnd00an1n02x5 FILLER_129_2063 ();
 b15zdnd00an1n01x5 FILLER_129_2065 ();
 b15zdnd11an1n04x5 FILLER_129_2092 ();
 b15zdnd11an1n16x5 FILLER_129_2106 ();
 b15zdnd11an1n08x5 FILLER_129_2122 ();
 b15zdnd00an1n01x5 FILLER_129_2130 ();
 b15zdnd11an1n08x5 FILLER_129_2143 ();
 b15zdnd00an1n01x5 FILLER_129_2151 ();
 b15zdnd11an1n04x5 FILLER_129_2166 ();
 b15zdnd00an1n01x5 FILLER_129_2170 ();
 b15zdnd11an1n04x5 FILLER_129_2176 ();
 b15zdnd11an1n04x5 FILLER_129_2189 ();
 b15zdnd11an1n64x5 FILLER_129_2213 ();
 b15zdnd11an1n04x5 FILLER_129_2277 ();
 b15zdnd00an1n02x5 FILLER_129_2281 ();
 b15zdnd00an1n01x5 FILLER_129_2283 ();
 b15zdnd11an1n32x5 FILLER_130_8 ();
 b15zdnd11an1n16x5 FILLER_130_40 ();
 b15zdnd11an1n08x5 FILLER_130_56 ();
 b15zdnd00an1n02x5 FILLER_130_64 ();
 b15zdnd11an1n32x5 FILLER_130_70 ();
 b15zdnd00an1n02x5 FILLER_130_102 ();
 b15zdnd00an1n01x5 FILLER_130_104 ();
 b15zdnd11an1n04x5 FILLER_130_116 ();
 b15zdnd11an1n16x5 FILLER_130_136 ();
 b15zdnd00an1n02x5 FILLER_130_152 ();
 b15zdnd00an1n01x5 FILLER_130_154 ();
 b15zdnd11an1n16x5 FILLER_130_160 ();
 b15zdnd11an1n32x5 FILLER_130_183 ();
 b15zdnd00an1n02x5 FILLER_130_215 ();
 b15zdnd11an1n64x5 FILLER_130_229 ();
 b15zdnd11an1n64x5 FILLER_130_293 ();
 b15zdnd11an1n04x5 FILLER_130_357 ();
 b15zdnd11an1n32x5 FILLER_130_374 ();
 b15zdnd11an1n16x5 FILLER_130_406 ();
 b15zdnd11an1n08x5 FILLER_130_422 ();
 b15zdnd11an1n04x5 FILLER_130_430 ();
 b15zdnd00an1n01x5 FILLER_130_434 ();
 b15zdnd11an1n08x5 FILLER_130_440 ();
 b15zdnd11an1n64x5 FILLER_130_454 ();
 b15zdnd11an1n64x5 FILLER_130_518 ();
 b15zdnd11an1n32x5 FILLER_130_582 ();
 b15zdnd11an1n04x5 FILLER_130_614 ();
 b15zdnd11an1n64x5 FILLER_130_626 ();
 b15zdnd11an1n16x5 FILLER_130_690 ();
 b15zdnd11an1n08x5 FILLER_130_706 ();
 b15zdnd11an1n04x5 FILLER_130_714 ();
 b15zdnd00an1n02x5 FILLER_130_726 ();
 b15zdnd11an1n32x5 FILLER_130_735 ();
 b15zdnd11an1n16x5 FILLER_130_767 ();
 b15zdnd11an1n08x5 FILLER_130_783 ();
 b15zdnd00an1n02x5 FILLER_130_791 ();
 b15zdnd00an1n01x5 FILLER_130_793 ();
 b15zdnd11an1n16x5 FILLER_130_802 ();
 b15zdnd11an1n08x5 FILLER_130_818 ();
 b15zdnd11an1n04x5 FILLER_130_826 ();
 b15zdnd00an1n01x5 FILLER_130_830 ();
 b15zdnd11an1n64x5 FILLER_130_838 ();
 b15zdnd11an1n04x5 FILLER_130_902 ();
 b15zdnd00an1n01x5 FILLER_130_906 ();
 b15zdnd11an1n64x5 FILLER_130_927 ();
 b15zdnd11an1n08x5 FILLER_130_991 ();
 b15zdnd00an1n02x5 FILLER_130_999 ();
 b15zdnd11an1n64x5 FILLER_130_1033 ();
 b15zdnd11an1n04x5 FILLER_130_1097 ();
 b15zdnd00an1n02x5 FILLER_130_1101 ();
 b15zdnd00an1n01x5 FILLER_130_1103 ();
 b15zdnd11an1n64x5 FILLER_130_1125 ();
 b15zdnd11an1n08x5 FILLER_130_1189 ();
 b15zdnd11an1n04x5 FILLER_130_1197 ();
 b15zdnd11an1n04x5 FILLER_130_1206 ();
 b15zdnd11an1n32x5 FILLER_130_1216 ();
 b15zdnd11an1n16x5 FILLER_130_1248 ();
 b15zdnd11an1n08x5 FILLER_130_1264 ();
 b15zdnd00an1n02x5 FILLER_130_1272 ();
 b15zdnd11an1n16x5 FILLER_130_1281 ();
 b15zdnd11an1n08x5 FILLER_130_1297 ();
 b15zdnd00an1n02x5 FILLER_130_1305 ();
 b15zdnd11an1n08x5 FILLER_130_1313 ();
 b15zdnd00an1n01x5 FILLER_130_1321 ();
 b15zdnd11an1n08x5 FILLER_130_1329 ();
 b15zdnd00an1n01x5 FILLER_130_1337 ();
 b15zdnd11an1n04x5 FILLER_130_1350 ();
 b15zdnd11an1n08x5 FILLER_130_1358 ();
 b15zdnd11an1n04x5 FILLER_130_1366 ();
 b15zdnd11an1n08x5 FILLER_130_1374 ();
 b15zdnd11an1n04x5 FILLER_130_1382 ();
 b15zdnd00an1n02x5 FILLER_130_1386 ();
 b15zdnd11an1n16x5 FILLER_130_1394 ();
 b15zdnd11an1n08x5 FILLER_130_1410 ();
 b15zdnd00an1n02x5 FILLER_130_1418 ();
 b15zdnd00an1n01x5 FILLER_130_1420 ();
 b15zdnd11an1n04x5 FILLER_130_1432 ();
 b15zdnd11an1n32x5 FILLER_130_1442 ();
 b15zdnd11an1n16x5 FILLER_130_1474 ();
 b15zdnd11an1n04x5 FILLER_130_1490 ();
 b15zdnd00an1n01x5 FILLER_130_1494 ();
 b15zdnd11an1n32x5 FILLER_130_1507 ();
 b15zdnd11an1n16x5 FILLER_130_1539 ();
 b15zdnd11an1n04x5 FILLER_130_1555 ();
 b15zdnd11an1n32x5 FILLER_130_1564 ();
 b15zdnd11an1n16x5 FILLER_130_1596 ();
 b15zdnd00an1n02x5 FILLER_130_1612 ();
 b15zdnd11an1n08x5 FILLER_130_1618 ();
 b15zdnd11an1n04x5 FILLER_130_1626 ();
 b15zdnd11an1n64x5 FILLER_130_1637 ();
 b15zdnd11an1n64x5 FILLER_130_1701 ();
 b15zdnd11an1n16x5 FILLER_130_1765 ();
 b15zdnd11an1n04x5 FILLER_130_1781 ();
 b15zdnd11an1n04x5 FILLER_130_1811 ();
 b15zdnd00an1n01x5 FILLER_130_1815 ();
 b15zdnd11an1n04x5 FILLER_130_1820 ();
 b15zdnd00an1n02x5 FILLER_130_1824 ();
 b15zdnd11an1n04x5 FILLER_130_1831 ();
 b15zdnd11an1n32x5 FILLER_130_1839 ();
 b15zdnd11an1n08x5 FILLER_130_1871 ();
 b15zdnd00an1n02x5 FILLER_130_1879 ();
 b15zdnd11an1n04x5 FILLER_130_1913 ();
 b15zdnd00an1n01x5 FILLER_130_1917 ();
 b15zdnd11an1n04x5 FILLER_130_1923 ();
 b15zdnd11an1n04x5 FILLER_130_1933 ();
 b15zdnd11an1n04x5 FILLER_130_1957 ();
 b15zdnd11an1n16x5 FILLER_130_1982 ();
 b15zdnd11an1n04x5 FILLER_130_1998 ();
 b15zdnd11an1n04x5 FILLER_130_2007 ();
 b15zdnd11an1n04x5 FILLER_130_2021 ();
 b15zdnd11an1n16x5 FILLER_130_2031 ();
 b15zdnd11an1n08x5 FILLER_130_2047 ();
 b15zdnd00an1n02x5 FILLER_130_2055 ();
 b15zdnd11an1n04x5 FILLER_130_2064 ();
 b15zdnd00an1n02x5 FILLER_130_2068 ();
 b15zdnd00an1n01x5 FILLER_130_2070 ();
 b15zdnd11an1n08x5 FILLER_130_2078 ();
 b15zdnd00an1n01x5 FILLER_130_2086 ();
 b15zdnd11an1n04x5 FILLER_130_2113 ();
 b15zdnd11an1n16x5 FILLER_130_2138 ();
 b15zdnd00an1n02x5 FILLER_130_2162 ();
 b15zdnd11an1n64x5 FILLER_130_2184 ();
 b15zdnd11an1n04x5 FILLER_130_2248 ();
 b15zdnd00an1n02x5 FILLER_130_2252 ();
 b15zdnd00an1n02x5 FILLER_130_2274 ();
 b15zdnd11an1n16x5 FILLER_131_0 ();
 b15zdnd11an1n08x5 FILLER_131_16 ();
 b15zdnd11an1n04x5 FILLER_131_24 ();
 b15zdnd00an1n02x5 FILLER_131_28 ();
 b15zdnd11an1n04x5 FILLER_131_39 ();
 b15zdnd11an1n16x5 FILLER_131_48 ();
 b15zdnd11an1n04x5 FILLER_131_64 ();
 b15zdnd11an1n64x5 FILLER_131_75 ();
 b15zdnd11an1n32x5 FILLER_131_139 ();
 b15zdnd00an1n02x5 FILLER_131_171 ();
 b15zdnd00an1n01x5 FILLER_131_173 ();
 b15zdnd11an1n08x5 FILLER_131_187 ();
 b15zdnd11an1n04x5 FILLER_131_195 ();
 b15zdnd00an1n01x5 FILLER_131_199 ();
 b15zdnd11an1n32x5 FILLER_131_205 ();
 b15zdnd11an1n16x5 FILLER_131_237 ();
 b15zdnd11an1n08x5 FILLER_131_253 ();
 b15zdnd00an1n02x5 FILLER_131_261 ();
 b15zdnd00an1n01x5 FILLER_131_263 ();
 b15zdnd11an1n64x5 FILLER_131_269 ();
 b15zdnd11an1n64x5 FILLER_131_333 ();
 b15zdnd11an1n64x5 FILLER_131_397 ();
 b15zdnd11an1n08x5 FILLER_131_461 ();
 b15zdnd11an1n04x5 FILLER_131_485 ();
 b15zdnd11an1n32x5 FILLER_131_495 ();
 b15zdnd11an1n16x5 FILLER_131_527 ();
 b15zdnd00an1n02x5 FILLER_131_543 ();
 b15zdnd00an1n01x5 FILLER_131_545 ();
 b15zdnd11an1n08x5 FILLER_131_558 ();
 b15zdnd00an1n02x5 FILLER_131_566 ();
 b15zdnd00an1n01x5 FILLER_131_568 ();
 b15zdnd11an1n16x5 FILLER_131_587 ();
 b15zdnd11an1n04x5 FILLER_131_603 ();
 b15zdnd00an1n02x5 FILLER_131_607 ();
 b15zdnd11an1n64x5 FILLER_131_618 ();
 b15zdnd11an1n16x5 FILLER_131_682 ();
 b15zdnd00an1n02x5 FILLER_131_698 ();
 b15zdnd11an1n04x5 FILLER_131_714 ();
 b15zdnd11an1n64x5 FILLER_131_730 ();
 b15zdnd00an1n01x5 FILLER_131_794 ();
 b15zdnd11an1n04x5 FILLER_131_802 ();
 b15zdnd11an1n04x5 FILLER_131_819 ();
 b15zdnd00an1n01x5 FILLER_131_823 ();
 b15zdnd11an1n04x5 FILLER_131_838 ();
 b15zdnd00an1n01x5 FILLER_131_842 ();
 b15zdnd11an1n04x5 FILLER_131_865 ();
 b15zdnd11an1n64x5 FILLER_131_879 ();
 b15zdnd11an1n16x5 FILLER_131_943 ();
 b15zdnd11an1n08x5 FILLER_131_959 ();
 b15zdnd11an1n04x5 FILLER_131_967 ();
 b15zdnd00an1n02x5 FILLER_131_971 ();
 b15zdnd00an1n01x5 FILLER_131_973 ();
 b15zdnd11an1n64x5 FILLER_131_994 ();
 b15zdnd11an1n32x5 FILLER_131_1058 ();
 b15zdnd00an1n02x5 FILLER_131_1090 ();
 b15zdnd11an1n32x5 FILLER_131_1104 ();
 b15zdnd11an1n16x5 FILLER_131_1136 ();
 b15zdnd11an1n08x5 FILLER_131_1152 ();
 b15zdnd11an1n04x5 FILLER_131_1160 ();
 b15zdnd00an1n02x5 FILLER_131_1164 ();
 b15zdnd11an1n64x5 FILLER_131_1191 ();
 b15zdnd11an1n08x5 FILLER_131_1255 ();
 b15zdnd00an1n02x5 FILLER_131_1263 ();
 b15zdnd11an1n16x5 FILLER_131_1272 ();
 b15zdnd11an1n08x5 FILLER_131_1288 ();
 b15zdnd11an1n04x5 FILLER_131_1296 ();
 b15zdnd00an1n02x5 FILLER_131_1300 ();
 b15zdnd00an1n01x5 FILLER_131_1302 ();
 b15zdnd11an1n64x5 FILLER_131_1316 ();
 b15zdnd11an1n08x5 FILLER_131_1380 ();
 b15zdnd00an1n01x5 FILLER_131_1388 ();
 b15zdnd11an1n04x5 FILLER_131_1393 ();
 b15zdnd00an1n02x5 FILLER_131_1397 ();
 b15zdnd11an1n04x5 FILLER_131_1425 ();
 b15zdnd11an1n32x5 FILLER_131_1436 ();
 b15zdnd11an1n16x5 FILLER_131_1468 ();
 b15zdnd11an1n04x5 FILLER_131_1484 ();
 b15zdnd00an1n02x5 FILLER_131_1488 ();
 b15zdnd00an1n01x5 FILLER_131_1490 ();
 b15zdnd11an1n32x5 FILLER_131_1499 ();
 b15zdnd11an1n16x5 FILLER_131_1531 ();
 b15zdnd11an1n08x5 FILLER_131_1547 ();
 b15zdnd00an1n02x5 FILLER_131_1555 ();
 b15zdnd11an1n64x5 FILLER_131_1563 ();
 b15zdnd11an1n08x5 FILLER_131_1627 ();
 b15zdnd00an1n02x5 FILLER_131_1635 ();
 b15zdnd11an1n64x5 FILLER_131_1649 ();
 b15zdnd11an1n64x5 FILLER_131_1713 ();
 b15zdnd11an1n64x5 FILLER_131_1777 ();
 b15zdnd11an1n32x5 FILLER_131_1841 ();
 b15zdnd11an1n04x5 FILLER_131_1899 ();
 b15zdnd11an1n08x5 FILLER_131_1907 ();
 b15zdnd00an1n02x5 FILLER_131_1915 ();
 b15zdnd11an1n16x5 FILLER_131_1922 ();
 b15zdnd11an1n04x5 FILLER_131_1938 ();
 b15zdnd00an1n02x5 FILLER_131_1942 ();
 b15zdnd00an1n01x5 FILLER_131_1944 ();
 b15zdnd11an1n16x5 FILLER_131_1971 ();
 b15zdnd11an1n08x5 FILLER_131_1987 ();
 b15zdnd11an1n04x5 FILLER_131_1995 ();
 b15zdnd00an1n01x5 FILLER_131_1999 ();
 b15zdnd11an1n08x5 FILLER_131_2020 ();
 b15zdnd00an1n02x5 FILLER_131_2028 ();
 b15zdnd11an1n32x5 FILLER_131_2056 ();
 b15zdnd11an1n16x5 FILLER_131_2088 ();
 b15zdnd00an1n02x5 FILLER_131_2104 ();
 b15zdnd00an1n01x5 FILLER_131_2106 ();
 b15zdnd11an1n04x5 FILLER_131_2133 ();
 b15zdnd11an1n64x5 FILLER_131_2142 ();
 b15zdnd11an1n16x5 FILLER_131_2206 ();
 b15zdnd11an1n04x5 FILLER_131_2222 ();
 b15zdnd00an1n01x5 FILLER_131_2226 ();
 b15zdnd11an1n08x5 FILLER_131_2233 ();
 b15zdnd11an1n04x5 FILLER_131_2241 ();
 b15zdnd00an1n02x5 FILLER_131_2245 ();
 b15zdnd11an1n32x5 FILLER_131_2251 ();
 b15zdnd00an1n01x5 FILLER_131_2283 ();
 b15zdnd11an1n32x5 FILLER_132_8 ();
 b15zdnd00an1n02x5 FILLER_132_40 ();
 b15zdnd00an1n01x5 FILLER_132_42 ();
 b15zdnd11an1n04x5 FILLER_132_59 ();
 b15zdnd11an1n32x5 FILLER_132_73 ();
 b15zdnd11an1n16x5 FILLER_132_105 ();
 b15zdnd11an1n08x5 FILLER_132_121 ();
 b15zdnd11an1n04x5 FILLER_132_129 ();
 b15zdnd00an1n02x5 FILLER_132_133 ();
 b15zdnd11an1n32x5 FILLER_132_147 ();
 b15zdnd11an1n16x5 FILLER_132_179 ();
 b15zdnd11an1n04x5 FILLER_132_195 ();
 b15zdnd00an1n02x5 FILLER_132_199 ();
 b15zdnd11an1n16x5 FILLER_132_206 ();
 b15zdnd11an1n04x5 FILLER_132_222 ();
 b15zdnd11an1n08x5 FILLER_132_240 ();
 b15zdnd11an1n04x5 FILLER_132_248 ();
 b15zdnd00an1n01x5 FILLER_132_252 ();
 b15zdnd11an1n04x5 FILLER_132_258 ();
 b15zdnd11an1n32x5 FILLER_132_277 ();
 b15zdnd11an1n16x5 FILLER_132_309 ();
 b15zdnd11an1n08x5 FILLER_132_325 ();
 b15zdnd11an1n04x5 FILLER_132_333 ();
 b15zdnd00an1n01x5 FILLER_132_337 ();
 b15zdnd11an1n64x5 FILLER_132_352 ();
 b15zdnd11an1n32x5 FILLER_132_416 ();
 b15zdnd11an1n16x5 FILLER_132_448 ();
 b15zdnd11an1n08x5 FILLER_132_482 ();
 b15zdnd00an1n02x5 FILLER_132_490 ();
 b15zdnd11an1n32x5 FILLER_132_500 ();
 b15zdnd00an1n02x5 FILLER_132_532 ();
 b15zdnd00an1n01x5 FILLER_132_534 ();
 b15zdnd11an1n04x5 FILLER_132_547 ();
 b15zdnd00an1n02x5 FILLER_132_551 ();
 b15zdnd11an1n16x5 FILLER_132_578 ();
 b15zdnd11an1n04x5 FILLER_132_594 ();
 b15zdnd00an1n01x5 FILLER_132_598 ();
 b15zdnd11an1n16x5 FILLER_132_609 ();
 b15zdnd11an1n04x5 FILLER_132_625 ();
 b15zdnd00an1n02x5 FILLER_132_629 ();
 b15zdnd00an1n01x5 FILLER_132_631 ();
 b15zdnd11an1n16x5 FILLER_132_640 ();
 b15zdnd00an1n02x5 FILLER_132_656 ();
 b15zdnd11an1n32x5 FILLER_132_664 ();
 b15zdnd11an1n08x5 FILLER_132_696 ();
 b15zdnd00an1n02x5 FILLER_132_704 ();
 b15zdnd11an1n04x5 FILLER_132_712 ();
 b15zdnd00an1n02x5 FILLER_132_716 ();
 b15zdnd11an1n16x5 FILLER_132_726 ();
 b15zdnd11an1n32x5 FILLER_132_747 ();
 b15zdnd11an1n16x5 FILLER_132_779 ();
 b15zdnd11an1n08x5 FILLER_132_795 ();
 b15zdnd11an1n04x5 FILLER_132_815 ();
 b15zdnd11an1n04x5 FILLER_132_839 ();
 b15zdnd00an1n02x5 FILLER_132_843 ();
 b15zdnd00an1n01x5 FILLER_132_845 ();
 b15zdnd11an1n08x5 FILLER_132_866 ();
 b15zdnd00an1n02x5 FILLER_132_874 ();
 b15zdnd00an1n01x5 FILLER_132_876 ();
 b15zdnd11an1n04x5 FILLER_132_883 ();
 b15zdnd11an1n16x5 FILLER_132_896 ();
 b15zdnd00an1n02x5 FILLER_132_912 ();
 b15zdnd00an1n01x5 FILLER_132_914 ();
 b15zdnd11an1n16x5 FILLER_132_920 ();
 b15zdnd11an1n08x5 FILLER_132_936 ();
 b15zdnd00an1n02x5 FILLER_132_944 ();
 b15zdnd00an1n01x5 FILLER_132_946 ();
 b15zdnd11an1n04x5 FILLER_132_967 ();
 b15zdnd11an1n64x5 FILLER_132_980 ();
 b15zdnd11an1n32x5 FILLER_132_1044 ();
 b15zdnd11an1n16x5 FILLER_132_1076 ();
 b15zdnd11an1n04x5 FILLER_132_1101 ();
 b15zdnd00an1n01x5 FILLER_132_1105 ();
 b15zdnd11an1n64x5 FILLER_132_1137 ();
 b15zdnd11an1n16x5 FILLER_132_1201 ();
 b15zdnd11an1n08x5 FILLER_132_1217 ();
 b15zdnd00an1n01x5 FILLER_132_1225 ();
 b15zdnd11an1n32x5 FILLER_132_1232 ();
 b15zdnd11an1n04x5 FILLER_132_1264 ();
 b15zdnd11an1n64x5 FILLER_132_1273 ();
 b15zdnd11an1n08x5 FILLER_132_1358 ();
 b15zdnd00an1n02x5 FILLER_132_1366 ();
 b15zdnd00an1n01x5 FILLER_132_1368 ();
 b15zdnd11an1n08x5 FILLER_132_1377 ();
 b15zdnd00an1n01x5 FILLER_132_1385 ();
 b15zdnd11an1n16x5 FILLER_132_1397 ();
 b15zdnd11an1n04x5 FILLER_132_1420 ();
 b15zdnd11an1n32x5 FILLER_132_1429 ();
 b15zdnd00an1n02x5 FILLER_132_1461 ();
 b15zdnd00an1n01x5 FILLER_132_1463 ();
 b15zdnd11an1n16x5 FILLER_132_1476 ();
 b15zdnd11an1n08x5 FILLER_132_1492 ();
 b15zdnd00an1n02x5 FILLER_132_1500 ();
 b15zdnd11an1n08x5 FILLER_132_1512 ();
 b15zdnd11an1n16x5 FILLER_132_1531 ();
 b15zdnd11an1n08x5 FILLER_132_1547 ();
 b15zdnd11an1n16x5 FILLER_132_1561 ();
 b15zdnd11an1n08x5 FILLER_132_1586 ();
 b15zdnd11an1n04x5 FILLER_132_1594 ();
 b15zdnd11an1n16x5 FILLER_132_1615 ();
 b15zdnd11an1n08x5 FILLER_132_1631 ();
 b15zdnd11an1n64x5 FILLER_132_1645 ();
 b15zdnd11an1n64x5 FILLER_132_1709 ();
 b15zdnd11an1n64x5 FILLER_132_1773 ();
 b15zdnd11an1n32x5 FILLER_132_1837 ();
 b15zdnd00an1n02x5 FILLER_132_1869 ();
 b15zdnd11an1n32x5 FILLER_132_1889 ();
 b15zdnd11an1n04x5 FILLER_132_1921 ();
 b15zdnd00an1n01x5 FILLER_132_1925 ();
 b15zdnd11an1n64x5 FILLER_132_1932 ();
 b15zdnd11an1n08x5 FILLER_132_1996 ();
 b15zdnd11an1n04x5 FILLER_132_2004 ();
 b15zdnd00an1n01x5 FILLER_132_2008 ();
 b15zdnd11an1n64x5 FILLER_132_2035 ();
 b15zdnd11an1n32x5 FILLER_132_2099 ();
 b15zdnd11an1n16x5 FILLER_132_2131 ();
 b15zdnd11an1n04x5 FILLER_132_2147 ();
 b15zdnd00an1n02x5 FILLER_132_2151 ();
 b15zdnd00an1n01x5 FILLER_132_2153 ();
 b15zdnd11an1n32x5 FILLER_132_2162 ();
 b15zdnd11an1n16x5 FILLER_132_2194 ();
 b15zdnd11an1n08x5 FILLER_132_2210 ();
 b15zdnd00an1n02x5 FILLER_132_2218 ();
 b15zdnd11an1n32x5 FILLER_132_2240 ();
 b15zdnd11an1n04x5 FILLER_132_2272 ();
 b15zdnd11an1n32x5 FILLER_133_0 ();
 b15zdnd11an1n16x5 FILLER_133_32 ();
 b15zdnd11an1n08x5 FILLER_133_54 ();
 b15zdnd11an1n04x5 FILLER_133_62 ();
 b15zdnd00an1n02x5 FILLER_133_66 ();
 b15zdnd00an1n01x5 FILLER_133_68 ();
 b15zdnd11an1n04x5 FILLER_133_76 ();
 b15zdnd00an1n01x5 FILLER_133_80 ();
 b15zdnd11an1n16x5 FILLER_133_96 ();
 b15zdnd11an1n04x5 FILLER_133_124 ();
 b15zdnd11an1n16x5 FILLER_133_134 ();
 b15zdnd00an1n01x5 FILLER_133_150 ();
 b15zdnd11an1n08x5 FILLER_133_167 ();
 b15zdnd11an1n08x5 FILLER_133_186 ();
 b15zdnd11an1n04x5 FILLER_133_194 ();
 b15zdnd00an1n02x5 FILLER_133_198 ();
 b15zdnd00an1n01x5 FILLER_133_200 ();
 b15zdnd11an1n32x5 FILLER_133_216 ();
 b15zdnd11an1n16x5 FILLER_133_248 ();
 b15zdnd11an1n08x5 FILLER_133_264 ();
 b15zdnd11an1n04x5 FILLER_133_272 ();
 b15zdnd00an1n02x5 FILLER_133_276 ();
 b15zdnd11an1n32x5 FILLER_133_284 ();
 b15zdnd00an1n01x5 FILLER_133_316 ();
 b15zdnd11an1n32x5 FILLER_133_327 ();
 b15zdnd11an1n32x5 FILLER_133_391 ();
 b15zdnd11an1n16x5 FILLER_133_423 ();
 b15zdnd00an1n01x5 FILLER_133_439 ();
 b15zdnd11an1n16x5 FILLER_133_463 ();
 b15zdnd11an1n08x5 FILLER_133_479 ();
 b15zdnd00an1n02x5 FILLER_133_487 ();
 b15zdnd00an1n01x5 FILLER_133_489 ();
 b15zdnd11an1n32x5 FILLER_133_498 ();
 b15zdnd11an1n16x5 FILLER_133_530 ();
 b15zdnd11an1n04x5 FILLER_133_546 ();
 b15zdnd00an1n01x5 FILLER_133_550 ();
 b15zdnd11an1n32x5 FILLER_133_564 ();
 b15zdnd11an1n04x5 FILLER_133_596 ();
 b15zdnd00an1n02x5 FILLER_133_600 ();
 b15zdnd11an1n08x5 FILLER_133_610 ();
 b15zdnd11an1n04x5 FILLER_133_618 ();
 b15zdnd00an1n02x5 FILLER_133_622 ();
 b15zdnd11an1n64x5 FILLER_133_631 ();
 b15zdnd11an1n64x5 FILLER_133_695 ();
 b15zdnd11an1n04x5 FILLER_133_759 ();
 b15zdnd00an1n02x5 FILLER_133_763 ();
 b15zdnd11an1n04x5 FILLER_133_782 ();
 b15zdnd11an1n64x5 FILLER_133_798 ();
 b15zdnd11an1n32x5 FILLER_133_862 ();
 b15zdnd11an1n16x5 FILLER_133_894 ();
 b15zdnd11an1n64x5 FILLER_133_919 ();
 b15zdnd11an1n32x5 FILLER_133_983 ();
 b15zdnd11an1n16x5 FILLER_133_1015 ();
 b15zdnd11an1n08x5 FILLER_133_1031 ();
 b15zdnd11an1n04x5 FILLER_133_1039 ();
 b15zdnd00an1n01x5 FILLER_133_1043 ();
 b15zdnd11an1n64x5 FILLER_133_1064 ();
 b15zdnd11an1n32x5 FILLER_133_1128 ();
 b15zdnd00an1n02x5 FILLER_133_1160 ();
 b15zdnd11an1n08x5 FILLER_133_1188 ();
 b15zdnd11an1n04x5 FILLER_133_1196 ();
 b15zdnd00an1n02x5 FILLER_133_1200 ();
 b15zdnd00an1n01x5 FILLER_133_1202 ();
 b15zdnd11an1n08x5 FILLER_133_1212 ();
 b15zdnd11an1n04x5 FILLER_133_1220 ();
 b15zdnd00an1n02x5 FILLER_133_1224 ();
 b15zdnd00an1n01x5 FILLER_133_1226 ();
 b15zdnd11an1n04x5 FILLER_133_1238 ();
 b15zdnd11an1n16x5 FILLER_133_1249 ();
 b15zdnd11an1n08x5 FILLER_133_1265 ();
 b15zdnd00an1n01x5 FILLER_133_1273 ();
 b15zdnd11an1n32x5 FILLER_133_1285 ();
 b15zdnd11an1n16x5 FILLER_133_1317 ();
 b15zdnd11an1n08x5 FILLER_133_1333 ();
 b15zdnd00an1n02x5 FILLER_133_1341 ();
 b15zdnd11an1n08x5 FILLER_133_1358 ();
 b15zdnd00an1n01x5 FILLER_133_1366 ();
 b15zdnd11an1n64x5 FILLER_133_1377 ();
 b15zdnd11an1n08x5 FILLER_133_1441 ();
 b15zdnd00an1n02x5 FILLER_133_1449 ();
 b15zdnd00an1n01x5 FILLER_133_1451 ();
 b15zdnd11an1n08x5 FILLER_133_1458 ();
 b15zdnd00an1n01x5 FILLER_133_1466 ();
 b15zdnd11an1n32x5 FILLER_133_1476 ();
 b15zdnd11an1n04x5 FILLER_133_1508 ();
 b15zdnd00an1n01x5 FILLER_133_1512 ();
 b15zdnd11an1n04x5 FILLER_133_1517 ();
 b15zdnd11an1n32x5 FILLER_133_1528 ();
 b15zdnd11an1n08x5 FILLER_133_1560 ();
 b15zdnd00an1n02x5 FILLER_133_1568 ();
 b15zdnd00an1n01x5 FILLER_133_1570 ();
 b15zdnd11an1n04x5 FILLER_133_1576 ();
 b15zdnd11an1n04x5 FILLER_133_1584 ();
 b15zdnd11an1n08x5 FILLER_133_1595 ();
 b15zdnd11an1n04x5 FILLER_133_1603 ();
 b15zdnd00an1n02x5 FILLER_133_1607 ();
 b15zdnd11an1n08x5 FILLER_133_1613 ();
 b15zdnd11an1n04x5 FILLER_133_1621 ();
 b15zdnd00an1n01x5 FILLER_133_1625 ();
 b15zdnd11an1n32x5 FILLER_133_1631 ();
 b15zdnd11an1n16x5 FILLER_133_1663 ();
 b15zdnd11an1n04x5 FILLER_133_1679 ();
 b15zdnd00an1n02x5 FILLER_133_1683 ();
 b15zdnd11an1n32x5 FILLER_133_1705 ();
 b15zdnd00an1n01x5 FILLER_133_1737 ();
 b15zdnd11an1n16x5 FILLER_133_1747 ();
 b15zdnd11an1n08x5 FILLER_133_1783 ();
 b15zdnd11an1n64x5 FILLER_133_1800 ();
 b15zdnd11an1n08x5 FILLER_133_1864 ();
 b15zdnd11an1n64x5 FILLER_133_1898 ();
 b15zdnd11an1n64x5 FILLER_133_1962 ();
 b15zdnd11an1n64x5 FILLER_133_2026 ();
 b15zdnd11an1n32x5 FILLER_133_2090 ();
 b15zdnd11an1n16x5 FILLER_133_2122 ();
 b15zdnd11an1n08x5 FILLER_133_2138 ();
 b15zdnd11an1n04x5 FILLER_133_2146 ();
 b15zdnd00an1n02x5 FILLER_133_2150 ();
 b15zdnd00an1n01x5 FILLER_133_2152 ();
 b15zdnd11an1n32x5 FILLER_133_2173 ();
 b15zdnd11an1n16x5 FILLER_133_2205 ();
 b15zdnd11an1n08x5 FILLER_133_2221 ();
 b15zdnd11an1n32x5 FILLER_133_2234 ();
 b15zdnd11an1n16x5 FILLER_133_2266 ();
 b15zdnd00an1n02x5 FILLER_133_2282 ();
 b15zdnd11an1n32x5 FILLER_134_8 ();
 b15zdnd11an1n04x5 FILLER_134_40 ();
 b15zdnd00an1n01x5 FILLER_134_44 ();
 b15zdnd11an1n04x5 FILLER_134_65 ();
 b15zdnd11an1n16x5 FILLER_134_73 ();
 b15zdnd11an1n08x5 FILLER_134_89 ();
 b15zdnd11an1n04x5 FILLER_134_97 ();
 b15zdnd11an1n16x5 FILLER_134_108 ();
 b15zdnd11an1n08x5 FILLER_134_124 ();
 b15zdnd11an1n16x5 FILLER_134_137 ();
 b15zdnd11an1n08x5 FILLER_134_153 ();
 b15zdnd11an1n04x5 FILLER_134_161 ();
 b15zdnd11an1n04x5 FILLER_134_171 ();
 b15zdnd11an1n64x5 FILLER_134_181 ();
 b15zdnd11an1n16x5 FILLER_134_245 ();
 b15zdnd11an1n08x5 FILLER_134_261 ();
 b15zdnd11an1n04x5 FILLER_134_269 ();
 b15zdnd00an1n01x5 FILLER_134_273 ();
 b15zdnd11an1n08x5 FILLER_134_279 ();
 b15zdnd11an1n04x5 FILLER_134_287 ();
 b15zdnd00an1n01x5 FILLER_134_291 ();
 b15zdnd11an1n04x5 FILLER_134_305 ();
 b15zdnd00an1n02x5 FILLER_134_309 ();
 b15zdnd11an1n32x5 FILLER_134_326 ();
 b15zdnd11an1n08x5 FILLER_134_358 ();
 b15zdnd00an1n02x5 FILLER_134_366 ();
 b15zdnd00an1n01x5 FILLER_134_368 ();
 b15zdnd11an1n08x5 FILLER_134_375 ();
 b15zdnd00an1n01x5 FILLER_134_383 ();
 b15zdnd11an1n64x5 FILLER_134_391 ();
 b15zdnd11an1n64x5 FILLER_134_455 ();
 b15zdnd11an1n64x5 FILLER_134_519 ();
 b15zdnd11an1n32x5 FILLER_134_583 ();
 b15zdnd11an1n08x5 FILLER_134_615 ();
 b15zdnd00an1n01x5 FILLER_134_623 ();
 b15zdnd11an1n08x5 FILLER_134_637 ();
 b15zdnd00an1n02x5 FILLER_134_645 ();
 b15zdnd11an1n16x5 FILLER_134_664 ();
 b15zdnd11an1n08x5 FILLER_134_680 ();
 b15zdnd00an1n02x5 FILLER_134_688 ();
 b15zdnd00an1n01x5 FILLER_134_690 ();
 b15zdnd11an1n08x5 FILLER_134_704 ();
 b15zdnd11an1n04x5 FILLER_134_712 ();
 b15zdnd00an1n02x5 FILLER_134_716 ();
 b15zdnd11an1n08x5 FILLER_134_726 ();
 b15zdnd00an1n02x5 FILLER_134_734 ();
 b15zdnd11an1n08x5 FILLER_134_740 ();
 b15zdnd11an1n04x5 FILLER_134_756 ();
 b15zdnd11an1n16x5 FILLER_134_769 ();
 b15zdnd00an1n02x5 FILLER_134_785 ();
 b15zdnd11an1n64x5 FILLER_134_805 ();
 b15zdnd11an1n32x5 FILLER_134_869 ();
 b15zdnd11an1n16x5 FILLER_134_901 ();
 b15zdnd11an1n04x5 FILLER_134_917 ();
 b15zdnd00an1n01x5 FILLER_134_921 ();
 b15zdnd11an1n64x5 FILLER_134_932 ();
 b15zdnd11an1n16x5 FILLER_134_996 ();
 b15zdnd11an1n04x5 FILLER_134_1012 ();
 b15zdnd11an1n32x5 FILLER_134_1034 ();
 b15zdnd11an1n04x5 FILLER_134_1066 ();
 b15zdnd00an1n01x5 FILLER_134_1070 ();
 b15zdnd11an1n64x5 FILLER_134_1086 ();
 b15zdnd11an1n64x5 FILLER_134_1150 ();
 b15zdnd11an1n32x5 FILLER_134_1214 ();
 b15zdnd11an1n04x5 FILLER_134_1246 ();
 b15zdnd11an1n64x5 FILLER_134_1254 ();
 b15zdnd11an1n64x5 FILLER_134_1318 ();
 b15zdnd11an1n64x5 FILLER_134_1382 ();
 b15zdnd11an1n16x5 FILLER_134_1446 ();
 b15zdnd00an1n01x5 FILLER_134_1462 ();
 b15zdnd11an1n32x5 FILLER_134_1469 ();
 b15zdnd11an1n08x5 FILLER_134_1501 ();
 b15zdnd11an1n04x5 FILLER_134_1509 ();
 b15zdnd00an1n02x5 FILLER_134_1513 ();
 b15zdnd11an1n64x5 FILLER_134_1522 ();
 b15zdnd11an1n08x5 FILLER_134_1586 ();
 b15zdnd11an1n04x5 FILLER_134_1594 ();
 b15zdnd00an1n02x5 FILLER_134_1598 ();
 b15zdnd11an1n04x5 FILLER_134_1618 ();
 b15zdnd11an1n64x5 FILLER_134_1634 ();
 b15zdnd11an1n32x5 FILLER_134_1698 ();
 b15zdnd11an1n08x5 FILLER_134_1730 ();
 b15zdnd11an1n04x5 FILLER_134_1738 ();
 b15zdnd00an1n02x5 FILLER_134_1742 ();
 b15zdnd11an1n08x5 FILLER_134_1753 ();
 b15zdnd00an1n02x5 FILLER_134_1761 ();
 b15zdnd00an1n01x5 FILLER_134_1763 ();
 b15zdnd11an1n08x5 FILLER_134_1782 ();
 b15zdnd00an1n02x5 FILLER_134_1790 ();
 b15zdnd00an1n01x5 FILLER_134_1792 ();
 b15zdnd11an1n16x5 FILLER_134_1804 ();
 b15zdnd11an1n04x5 FILLER_134_1820 ();
 b15zdnd00an1n01x5 FILLER_134_1824 ();
 b15zdnd11an1n04x5 FILLER_134_1835 ();
 b15zdnd11an1n64x5 FILLER_134_1850 ();
 b15zdnd11an1n64x5 FILLER_134_1914 ();
 b15zdnd11an1n32x5 FILLER_134_1978 ();
 b15zdnd11an1n16x5 FILLER_134_2010 ();
 b15zdnd00an1n02x5 FILLER_134_2026 ();
 b15zdnd00an1n01x5 FILLER_134_2028 ();
 b15zdnd11an1n32x5 FILLER_134_2046 ();
 b15zdnd11an1n16x5 FILLER_134_2078 ();
 b15zdnd00an1n01x5 FILLER_134_2094 ();
 b15zdnd11an1n32x5 FILLER_134_2121 ();
 b15zdnd00an1n01x5 FILLER_134_2153 ();
 b15zdnd00an1n02x5 FILLER_134_2162 ();
 b15zdnd00an1n01x5 FILLER_134_2164 ();
 b15zdnd11an1n16x5 FILLER_134_2169 ();
 b15zdnd00an1n01x5 FILLER_134_2185 ();
 b15zdnd11an1n64x5 FILLER_134_2206 ();
 b15zdnd11an1n04x5 FILLER_134_2270 ();
 b15zdnd00an1n02x5 FILLER_134_2274 ();
 b15zdnd11an1n64x5 FILLER_135_0 ();
 b15zdnd11an1n16x5 FILLER_135_64 ();
 b15zdnd11an1n08x5 FILLER_135_80 ();
 b15zdnd11an1n04x5 FILLER_135_88 ();
 b15zdnd11an1n32x5 FILLER_135_98 ();
 b15zdnd11an1n04x5 FILLER_135_130 ();
 b15zdnd00an1n02x5 FILLER_135_134 ();
 b15zdnd11an1n16x5 FILLER_135_142 ();
 b15zdnd11an1n08x5 FILLER_135_158 ();
 b15zdnd11an1n32x5 FILLER_135_177 ();
 b15zdnd00an1n02x5 FILLER_135_209 ();
 b15zdnd11an1n32x5 FILLER_135_220 ();
 b15zdnd11an1n08x5 FILLER_135_252 ();
 b15zdnd11an1n04x5 FILLER_135_260 ();
 b15zdnd11an1n08x5 FILLER_135_271 ();
 b15zdnd00an1n02x5 FILLER_135_279 ();
 b15zdnd11an1n04x5 FILLER_135_297 ();
 b15zdnd00an1n01x5 FILLER_135_301 ();
 b15zdnd11an1n08x5 FILLER_135_307 ();
 b15zdnd11an1n04x5 FILLER_135_315 ();
 b15zdnd00an1n01x5 FILLER_135_319 ();
 b15zdnd11an1n16x5 FILLER_135_325 ();
 b15zdnd11an1n04x5 FILLER_135_341 ();
 b15zdnd00an1n02x5 FILLER_135_345 ();
 b15zdnd00an1n01x5 FILLER_135_347 ();
 b15zdnd11an1n08x5 FILLER_135_364 ();
 b15zdnd00an1n01x5 FILLER_135_372 ();
 b15zdnd11an1n64x5 FILLER_135_380 ();
 b15zdnd11an1n16x5 FILLER_135_444 ();
 b15zdnd00an1n02x5 FILLER_135_460 ();
 b15zdnd11an1n64x5 FILLER_135_478 ();
 b15zdnd11an1n64x5 FILLER_135_542 ();
 b15zdnd11an1n08x5 FILLER_135_606 ();
 b15zdnd11an1n04x5 FILLER_135_614 ();
 b15zdnd00an1n01x5 FILLER_135_618 ();
 b15zdnd11an1n08x5 FILLER_135_625 ();
 b15zdnd00an1n02x5 FILLER_135_633 ();
 b15zdnd00an1n01x5 FILLER_135_635 ();
 b15zdnd11an1n04x5 FILLER_135_640 ();
 b15zdnd00an1n02x5 FILLER_135_644 ();
 b15zdnd11an1n04x5 FILLER_135_652 ();
 b15zdnd11an1n16x5 FILLER_135_666 ();
 b15zdnd11an1n08x5 FILLER_135_698 ();
 b15zdnd11an1n04x5 FILLER_135_706 ();
 b15zdnd00an1n02x5 FILLER_135_710 ();
 b15zdnd11an1n08x5 FILLER_135_721 ();
 b15zdnd11an1n04x5 FILLER_135_729 ();
 b15zdnd00an1n02x5 FILLER_135_733 ();
 b15zdnd11an1n04x5 FILLER_135_745 ();
 b15zdnd00an1n02x5 FILLER_135_749 ();
 b15zdnd11an1n16x5 FILLER_135_760 ();
 b15zdnd00an1n01x5 FILLER_135_776 ();
 b15zdnd11an1n64x5 FILLER_135_795 ();
 b15zdnd11an1n08x5 FILLER_135_859 ();
 b15zdnd11an1n04x5 FILLER_135_867 ();
 b15zdnd11an1n16x5 FILLER_135_891 ();
 b15zdnd11an1n08x5 FILLER_135_907 ();
 b15zdnd11an1n04x5 FILLER_135_915 ();
 b15zdnd11an1n32x5 FILLER_135_930 ();
 b15zdnd11an1n04x5 FILLER_135_962 ();
 b15zdnd11an1n04x5 FILLER_135_987 ();
 b15zdnd11an1n16x5 FILLER_135_1016 ();
 b15zdnd11an1n04x5 FILLER_135_1032 ();
 b15zdnd00an1n01x5 FILLER_135_1036 ();
 b15zdnd11an1n16x5 FILLER_135_1047 ();
 b15zdnd11an1n08x5 FILLER_135_1063 ();
 b15zdnd11an1n04x5 FILLER_135_1071 ();
 b15zdnd00an1n01x5 FILLER_135_1075 ();
 b15zdnd11an1n04x5 FILLER_135_1085 ();
 b15zdnd11an1n64x5 FILLER_135_1098 ();
 b15zdnd11an1n32x5 FILLER_135_1162 ();
 b15zdnd11an1n16x5 FILLER_135_1194 ();
 b15zdnd00an1n02x5 FILLER_135_1210 ();
 b15zdnd11an1n32x5 FILLER_135_1216 ();
 b15zdnd11an1n08x5 FILLER_135_1248 ();
 b15zdnd00an1n02x5 FILLER_135_1256 ();
 b15zdnd00an1n01x5 FILLER_135_1258 ();
 b15zdnd11an1n32x5 FILLER_135_1264 ();
 b15zdnd11an1n08x5 FILLER_135_1296 ();
 b15zdnd00an1n02x5 FILLER_135_1304 ();
 b15zdnd11an1n04x5 FILLER_135_1315 ();
 b15zdnd00an1n01x5 FILLER_135_1319 ();
 b15zdnd11an1n32x5 FILLER_135_1334 ();
 b15zdnd00an1n02x5 FILLER_135_1366 ();
 b15zdnd11an1n32x5 FILLER_135_1374 ();
 b15zdnd11an1n08x5 FILLER_135_1406 ();
 b15zdnd11an1n04x5 FILLER_135_1414 ();
 b15zdnd00an1n02x5 FILLER_135_1418 ();
 b15zdnd11an1n32x5 FILLER_135_1426 ();
 b15zdnd11an1n16x5 FILLER_135_1458 ();
 b15zdnd11an1n08x5 FILLER_135_1474 ();
 b15zdnd00an1n02x5 FILLER_135_1482 ();
 b15zdnd11an1n16x5 FILLER_135_1489 ();
 b15zdnd11an1n08x5 FILLER_135_1505 ();
 b15zdnd11an1n32x5 FILLER_135_1519 ();
 b15zdnd11an1n32x5 FILLER_135_1563 ();
 b15zdnd11an1n16x5 FILLER_135_1595 ();
 b15zdnd11an1n08x5 FILLER_135_1611 ();
 b15zdnd11an1n04x5 FILLER_135_1619 ();
 b15zdnd00an1n02x5 FILLER_135_1623 ();
 b15zdnd11an1n64x5 FILLER_135_1630 ();
 b15zdnd11an1n16x5 FILLER_135_1703 ();
 b15zdnd11an1n08x5 FILLER_135_1719 ();
 b15zdnd11an1n04x5 FILLER_135_1727 ();
 b15zdnd00an1n02x5 FILLER_135_1731 ();
 b15zdnd00an1n01x5 FILLER_135_1733 ();
 b15zdnd11an1n32x5 FILLER_135_1743 ();
 b15zdnd11an1n16x5 FILLER_135_1775 ();
 b15zdnd11an1n08x5 FILLER_135_1791 ();
 b15zdnd11an1n04x5 FILLER_135_1799 ();
 b15zdnd00an1n01x5 FILLER_135_1803 ();
 b15zdnd11an1n04x5 FILLER_135_1821 ();
 b15zdnd11an1n32x5 FILLER_135_1835 ();
 b15zdnd11an1n08x5 FILLER_135_1867 ();
 b15zdnd11an1n04x5 FILLER_135_1875 ();
 b15zdnd00an1n01x5 FILLER_135_1879 ();
 b15zdnd11an1n32x5 FILLER_135_1911 ();
 b15zdnd11an1n16x5 FILLER_135_1943 ();
 b15zdnd11an1n04x5 FILLER_135_1959 ();
 b15zdnd00an1n02x5 FILLER_135_1963 ();
 b15zdnd11an1n32x5 FILLER_135_1985 ();
 b15zdnd11an1n16x5 FILLER_135_2017 ();
 b15zdnd11an1n08x5 FILLER_135_2033 ();
 b15zdnd00an1n02x5 FILLER_135_2041 ();
 b15zdnd00an1n01x5 FILLER_135_2043 ();
 b15zdnd11an1n64x5 FILLER_135_2064 ();
 b15zdnd11an1n32x5 FILLER_135_2128 ();
 b15zdnd11an1n04x5 FILLER_135_2160 ();
 b15zdnd00an1n01x5 FILLER_135_2164 ();
 b15zdnd11an1n64x5 FILLER_135_2170 ();
 b15zdnd11an1n08x5 FILLER_135_2234 ();
 b15zdnd00an1n02x5 FILLER_135_2242 ();
 b15zdnd00an1n01x5 FILLER_135_2244 ();
 b15zdnd11an1n32x5 FILLER_135_2249 ();
 b15zdnd00an1n02x5 FILLER_135_2281 ();
 b15zdnd00an1n01x5 FILLER_135_2283 ();
 b15zdnd11an1n64x5 FILLER_136_8 ();
 b15zdnd11an1n64x5 FILLER_136_72 ();
 b15zdnd11an1n64x5 FILLER_136_136 ();
 b15zdnd11an1n08x5 FILLER_136_200 ();
 b15zdnd11an1n04x5 FILLER_136_208 ();
 b15zdnd11an1n64x5 FILLER_136_227 ();
 b15zdnd11an1n08x5 FILLER_136_291 ();
 b15zdnd00an1n02x5 FILLER_136_299 ();
 b15zdnd11an1n64x5 FILLER_136_310 ();
 b15zdnd11an1n64x5 FILLER_136_374 ();
 b15zdnd11an1n64x5 FILLER_136_438 ();
 b15zdnd11an1n64x5 FILLER_136_502 ();
 b15zdnd11an1n64x5 FILLER_136_566 ();
 b15zdnd11an1n32x5 FILLER_136_630 ();
 b15zdnd11an1n08x5 FILLER_136_662 ();
 b15zdnd00an1n02x5 FILLER_136_670 ();
 b15zdnd00an1n01x5 FILLER_136_672 ();
 b15zdnd11an1n32x5 FILLER_136_686 ();
 b15zdnd11an1n64x5 FILLER_136_726 ();
 b15zdnd11an1n32x5 FILLER_136_790 ();
 b15zdnd00an1n02x5 FILLER_136_822 ();
 b15zdnd11an1n16x5 FILLER_136_844 ();
 b15zdnd11an1n08x5 FILLER_136_860 ();
 b15zdnd11an1n04x5 FILLER_136_868 ();
 b15zdnd00an1n02x5 FILLER_136_872 ();
 b15zdnd00an1n01x5 FILLER_136_874 ();
 b15zdnd11an1n04x5 FILLER_136_884 ();
 b15zdnd11an1n64x5 FILLER_136_893 ();
 b15zdnd11an1n16x5 FILLER_136_957 ();
 b15zdnd11an1n04x5 FILLER_136_973 ();
 b15zdnd00an1n02x5 FILLER_136_977 ();
 b15zdnd00an1n01x5 FILLER_136_979 ();
 b15zdnd11an1n64x5 FILLER_136_990 ();
 b15zdnd11an1n32x5 FILLER_136_1054 ();
 b15zdnd11an1n08x5 FILLER_136_1086 ();
 b15zdnd11an1n64x5 FILLER_136_1103 ();
 b15zdnd11an1n32x5 FILLER_136_1167 ();
 b15zdnd11an1n04x5 FILLER_136_1199 ();
 b15zdnd00an1n02x5 FILLER_136_1203 ();
 b15zdnd00an1n01x5 FILLER_136_1205 ();
 b15zdnd11an1n32x5 FILLER_136_1212 ();
 b15zdnd11an1n16x5 FILLER_136_1244 ();
 b15zdnd11an1n04x5 FILLER_136_1260 ();
 b15zdnd00an1n02x5 FILLER_136_1264 ();
 b15zdnd00an1n01x5 FILLER_136_1266 ();
 b15zdnd11an1n08x5 FILLER_136_1275 ();
 b15zdnd00an1n01x5 FILLER_136_1283 ();
 b15zdnd11an1n04x5 FILLER_136_1296 ();
 b15zdnd11an1n04x5 FILLER_136_1321 ();
 b15zdnd11an1n04x5 FILLER_136_1329 ();
 b15zdnd11an1n16x5 FILLER_136_1345 ();
 b15zdnd11an1n04x5 FILLER_136_1361 ();
 b15zdnd00an1n01x5 FILLER_136_1365 ();
 b15zdnd11an1n32x5 FILLER_136_1379 ();
 b15zdnd11an1n08x5 FILLER_136_1411 ();
 b15zdnd00an1n02x5 FILLER_136_1419 ();
 b15zdnd00an1n01x5 FILLER_136_1421 ();
 b15zdnd11an1n64x5 FILLER_136_1442 ();
 b15zdnd11an1n32x5 FILLER_136_1506 ();
 b15zdnd11an1n08x5 FILLER_136_1538 ();
 b15zdnd11an1n32x5 FILLER_136_1558 ();
 b15zdnd11an1n64x5 FILLER_136_1595 ();
 b15zdnd11an1n64x5 FILLER_136_1659 ();
 b15zdnd11an1n64x5 FILLER_136_1723 ();
 b15zdnd11an1n64x5 FILLER_136_1787 ();
 b15zdnd11an1n32x5 FILLER_136_1851 ();
 b15zdnd11an1n16x5 FILLER_136_1883 ();
 b15zdnd11an1n32x5 FILLER_136_1919 ();
 b15zdnd11an1n16x5 FILLER_136_1951 ();
 b15zdnd00an1n02x5 FILLER_136_1967 ();
 b15zdnd11an1n04x5 FILLER_136_1995 ();
 b15zdnd11an1n16x5 FILLER_136_2019 ();
 b15zdnd11an1n04x5 FILLER_136_2035 ();
 b15zdnd11an1n32x5 FILLER_136_2057 ();
 b15zdnd11an1n16x5 FILLER_136_2089 ();
 b15zdnd11an1n08x5 FILLER_136_2105 ();
 b15zdnd00an1n01x5 FILLER_136_2113 ();
 b15zdnd11an1n16x5 FILLER_136_2134 ();
 b15zdnd11an1n04x5 FILLER_136_2150 ();
 b15zdnd11an1n64x5 FILLER_136_2162 ();
 b15zdnd11an1n16x5 FILLER_136_2226 ();
 b15zdnd11an1n08x5 FILLER_136_2242 ();
 b15zdnd11an1n04x5 FILLER_136_2250 ();
 b15zdnd00an1n02x5 FILLER_136_2274 ();
 b15zdnd11an1n64x5 FILLER_137_0 ();
 b15zdnd11an1n64x5 FILLER_137_64 ();
 b15zdnd11an1n64x5 FILLER_137_128 ();
 b15zdnd11an1n08x5 FILLER_137_192 ();
 b15zdnd11an1n04x5 FILLER_137_200 ();
 b15zdnd00an1n02x5 FILLER_137_204 ();
 b15zdnd11an1n04x5 FILLER_137_222 ();
 b15zdnd11an1n16x5 FILLER_137_239 ();
 b15zdnd11an1n04x5 FILLER_137_255 ();
 b15zdnd00an1n02x5 FILLER_137_259 ();
 b15zdnd00an1n01x5 FILLER_137_261 ();
 b15zdnd11an1n16x5 FILLER_137_269 ();
 b15zdnd00an1n02x5 FILLER_137_285 ();
 b15zdnd00an1n01x5 FILLER_137_287 ();
 b15zdnd11an1n04x5 FILLER_137_298 ();
 b15zdnd11an1n16x5 FILLER_137_312 ();
 b15zdnd00an1n02x5 FILLER_137_328 ();
 b15zdnd00an1n01x5 FILLER_137_330 ();
 b15zdnd11an1n04x5 FILLER_137_347 ();
 b15zdnd11an1n64x5 FILLER_137_383 ();
 b15zdnd11an1n64x5 FILLER_137_447 ();
 b15zdnd11an1n64x5 FILLER_137_511 ();
 b15zdnd11an1n64x5 FILLER_137_575 ();
 b15zdnd11an1n32x5 FILLER_137_639 ();
 b15zdnd11an1n16x5 FILLER_137_671 ();
 b15zdnd11an1n64x5 FILLER_137_694 ();
 b15zdnd11an1n64x5 FILLER_137_758 ();
 b15zdnd11an1n08x5 FILLER_137_822 ();
 b15zdnd11an1n64x5 FILLER_137_835 ();
 b15zdnd11an1n64x5 FILLER_137_899 ();
 b15zdnd11an1n08x5 FILLER_137_963 ();
 b15zdnd11an1n04x5 FILLER_137_971 ();
 b15zdnd00an1n01x5 FILLER_137_975 ();
 b15zdnd11an1n64x5 FILLER_137_991 ();
 b15zdnd11an1n08x5 FILLER_137_1055 ();
 b15zdnd11an1n04x5 FILLER_137_1081 ();
 b15zdnd00an1n02x5 FILLER_137_1085 ();
 b15zdnd11an1n64x5 FILLER_137_1096 ();
 b15zdnd11an1n32x5 FILLER_137_1160 ();
 b15zdnd11an1n08x5 FILLER_137_1192 ();
 b15zdnd11an1n04x5 FILLER_137_1200 ();
 b15zdnd11an1n32x5 FILLER_137_1209 ();
 b15zdnd11an1n16x5 FILLER_137_1241 ();
 b15zdnd11an1n08x5 FILLER_137_1257 ();
 b15zdnd00an1n02x5 FILLER_137_1265 ();
 b15zdnd00an1n01x5 FILLER_137_1267 ();
 b15zdnd11an1n08x5 FILLER_137_1275 ();
 b15zdnd00an1n01x5 FILLER_137_1283 ();
 b15zdnd11an1n64x5 FILLER_137_1289 ();
 b15zdnd11an1n64x5 FILLER_137_1353 ();
 b15zdnd00an1n01x5 FILLER_137_1417 ();
 b15zdnd11an1n04x5 FILLER_137_1427 ();
 b15zdnd00an1n02x5 FILLER_137_1431 ();
 b15zdnd00an1n01x5 FILLER_137_1433 ();
 b15zdnd11an1n32x5 FILLER_137_1444 ();
 b15zdnd11an1n16x5 FILLER_137_1476 ();
 b15zdnd11an1n08x5 FILLER_137_1492 ();
 b15zdnd11an1n04x5 FILLER_137_1505 ();
 b15zdnd11an1n16x5 FILLER_137_1519 ();
 b15zdnd11an1n04x5 FILLER_137_1535 ();
 b15zdnd00an1n02x5 FILLER_137_1539 ();
 b15zdnd11an1n32x5 FILLER_137_1550 ();
 b15zdnd11an1n08x5 FILLER_137_1582 ();
 b15zdnd11an1n04x5 FILLER_137_1590 ();
 b15zdnd00an1n02x5 FILLER_137_1594 ();
 b15zdnd11an1n16x5 FILLER_137_1601 ();
 b15zdnd11an1n08x5 FILLER_137_1617 ();
 b15zdnd11an1n04x5 FILLER_137_1651 ();
 b15zdnd11an1n08x5 FILLER_137_1675 ();
 b15zdnd00an1n02x5 FILLER_137_1683 ();
 b15zdnd00an1n01x5 FILLER_137_1685 ();
 b15zdnd11an1n04x5 FILLER_137_1706 ();
 b15zdnd11an1n16x5 FILLER_137_1719 ();
 b15zdnd00an1n01x5 FILLER_137_1735 ();
 b15zdnd11an1n64x5 FILLER_137_1767 ();
 b15zdnd11an1n32x5 FILLER_137_1831 ();
 b15zdnd11an1n16x5 FILLER_137_1863 ();
 b15zdnd11an1n08x5 FILLER_137_1879 ();
 b15zdnd11an1n04x5 FILLER_137_1887 ();
 b15zdnd00an1n02x5 FILLER_137_1891 ();
 b15zdnd00an1n01x5 FILLER_137_1893 ();
 b15zdnd11an1n16x5 FILLER_137_1903 ();
 b15zdnd11an1n04x5 FILLER_137_1919 ();
 b15zdnd00an1n01x5 FILLER_137_1923 ();
 b15zdnd11an1n16x5 FILLER_137_1936 ();
 b15zdnd11an1n08x5 FILLER_137_1952 ();
 b15zdnd11an1n04x5 FILLER_137_1960 ();
 b15zdnd11an1n32x5 FILLER_137_1973 ();
 b15zdnd11an1n08x5 FILLER_137_2005 ();
 b15zdnd11an1n04x5 FILLER_137_2039 ();
 b15zdnd11an1n32x5 FILLER_137_2052 ();
 b15zdnd11an1n16x5 FILLER_137_2084 ();
 b15zdnd11an1n04x5 FILLER_137_2100 ();
 b15zdnd11an1n64x5 FILLER_137_2113 ();
 b15zdnd00an1n02x5 FILLER_137_2177 ();
 b15zdnd00an1n01x5 FILLER_137_2179 ();
 b15zdnd11an1n16x5 FILLER_137_2184 ();
 b15zdnd11an1n08x5 FILLER_137_2200 ();
 b15zdnd11an1n04x5 FILLER_137_2208 ();
 b15zdnd00an1n02x5 FILLER_137_2212 ();
 b15zdnd11an1n32x5 FILLER_137_2234 ();
 b15zdnd11an1n04x5 FILLER_137_2266 ();
 b15zdnd11an1n04x5 FILLER_137_2274 ();
 b15zdnd00an1n02x5 FILLER_137_2282 ();
 b15zdnd11an1n32x5 FILLER_138_8 ();
 b15zdnd11an1n08x5 FILLER_138_40 ();
 b15zdnd00an1n02x5 FILLER_138_48 ();
 b15zdnd11an1n04x5 FILLER_138_62 ();
 b15zdnd11an1n32x5 FILLER_138_70 ();
 b15zdnd11an1n16x5 FILLER_138_102 ();
 b15zdnd11an1n04x5 FILLER_138_118 ();
 b15zdnd11an1n04x5 FILLER_138_127 ();
 b15zdnd11an1n32x5 FILLER_138_135 ();
 b15zdnd11an1n08x5 FILLER_138_167 ();
 b15zdnd11an1n64x5 FILLER_138_182 ();
 b15zdnd11an1n16x5 FILLER_138_246 ();
 b15zdnd11an1n04x5 FILLER_138_268 ();
 b15zdnd11an1n64x5 FILLER_138_276 ();
 b15zdnd11an1n32x5 FILLER_138_340 ();
 b15zdnd00an1n02x5 FILLER_138_372 ();
 b15zdnd00an1n01x5 FILLER_138_374 ();
 b15zdnd11an1n64x5 FILLER_138_387 ();
 b15zdnd11an1n08x5 FILLER_138_451 ();
 b15zdnd00an1n02x5 FILLER_138_459 ();
 b15zdnd00an1n01x5 FILLER_138_461 ();
 b15zdnd11an1n08x5 FILLER_138_478 ();
 b15zdnd11an1n04x5 FILLER_138_486 ();
 b15zdnd11an1n04x5 FILLER_138_498 ();
 b15zdnd00an1n01x5 FILLER_138_502 ();
 b15zdnd11an1n16x5 FILLER_138_515 ();
 b15zdnd11an1n04x5 FILLER_138_531 ();
 b15zdnd11an1n04x5 FILLER_138_541 ();
 b15zdnd00an1n02x5 FILLER_138_545 ();
 b15zdnd00an1n01x5 FILLER_138_547 ();
 b15zdnd11an1n04x5 FILLER_138_552 ();
 b15zdnd00an1n02x5 FILLER_138_556 ();
 b15zdnd11an1n16x5 FILLER_138_564 ();
 b15zdnd11an1n08x5 FILLER_138_580 ();
 b15zdnd11an1n04x5 FILLER_138_588 ();
 b15zdnd00an1n02x5 FILLER_138_592 ();
 b15zdnd00an1n01x5 FILLER_138_594 ();
 b15zdnd11an1n64x5 FILLER_138_602 ();
 b15zdnd11an1n32x5 FILLER_138_666 ();
 b15zdnd11an1n16x5 FILLER_138_698 ();
 b15zdnd11an1n04x5 FILLER_138_714 ();
 b15zdnd11an1n16x5 FILLER_138_726 ();
 b15zdnd11an1n04x5 FILLER_138_742 ();
 b15zdnd00an1n01x5 FILLER_138_746 ();
 b15zdnd11an1n32x5 FILLER_138_767 ();
 b15zdnd11an1n16x5 FILLER_138_799 ();
 b15zdnd11an1n08x5 FILLER_138_815 ();
 b15zdnd11an1n04x5 FILLER_138_823 ();
 b15zdnd00an1n02x5 FILLER_138_827 ();
 b15zdnd00an1n01x5 FILLER_138_829 ();
 b15zdnd11an1n32x5 FILLER_138_839 ();
 b15zdnd11an1n16x5 FILLER_138_871 ();
 b15zdnd11an1n08x5 FILLER_138_887 ();
 b15zdnd11an1n64x5 FILLER_138_904 ();
 b15zdnd00an1n02x5 FILLER_138_968 ();
 b15zdnd11an1n64x5 FILLER_138_979 ();
 b15zdnd11an1n32x5 FILLER_138_1043 ();
 b15zdnd11an1n08x5 FILLER_138_1075 ();
 b15zdnd00an1n01x5 FILLER_138_1083 ();
 b15zdnd11an1n64x5 FILLER_138_1095 ();
 b15zdnd11an1n32x5 FILLER_138_1159 ();
 b15zdnd11an1n08x5 FILLER_138_1191 ();
 b15zdnd11an1n04x5 FILLER_138_1199 ();
 b15zdnd11an1n04x5 FILLER_138_1215 ();
 b15zdnd11an1n08x5 FILLER_138_1226 ();
 b15zdnd00an1n01x5 FILLER_138_1234 ();
 b15zdnd11an1n64x5 FILLER_138_1241 ();
 b15zdnd11an1n64x5 FILLER_138_1305 ();
 b15zdnd11an1n16x5 FILLER_138_1369 ();
 b15zdnd11an1n04x5 FILLER_138_1385 ();
 b15zdnd00an1n01x5 FILLER_138_1389 ();
 b15zdnd11an1n64x5 FILLER_138_1401 ();
 b15zdnd00an1n02x5 FILLER_138_1465 ();
 b15zdnd00an1n01x5 FILLER_138_1467 ();
 b15zdnd11an1n16x5 FILLER_138_1474 ();
 b15zdnd11an1n08x5 FILLER_138_1490 ();
 b15zdnd11an1n08x5 FILLER_138_1508 ();
 b15zdnd11an1n04x5 FILLER_138_1516 ();
 b15zdnd00an1n02x5 FILLER_138_1520 ();
 b15zdnd00an1n01x5 FILLER_138_1522 ();
 b15zdnd11an1n16x5 FILLER_138_1529 ();
 b15zdnd11an1n04x5 FILLER_138_1545 ();
 b15zdnd00an1n02x5 FILLER_138_1549 ();
 b15zdnd00an1n01x5 FILLER_138_1551 ();
 b15zdnd11an1n32x5 FILLER_138_1556 ();
 b15zdnd00an1n02x5 FILLER_138_1588 ();
 b15zdnd11an1n08x5 FILLER_138_1597 ();
 b15zdnd11an1n04x5 FILLER_138_1605 ();
 b15zdnd00an1n02x5 FILLER_138_1609 ();
 b15zdnd11an1n04x5 FILLER_138_1619 ();
 b15zdnd11an1n04x5 FILLER_138_1627 ();
 b15zdnd00an1n01x5 FILLER_138_1631 ();
 b15zdnd11an1n08x5 FILLER_138_1638 ();
 b15zdnd11an1n04x5 FILLER_138_1646 ();
 b15zdnd00an1n02x5 FILLER_138_1650 ();
 b15zdnd00an1n01x5 FILLER_138_1652 ();
 b15zdnd11an1n32x5 FILLER_138_1679 ();
 b15zdnd11an1n04x5 FILLER_138_1711 ();
 b15zdnd00an1n02x5 FILLER_138_1715 ();
 b15zdnd00an1n01x5 FILLER_138_1717 ();
 b15zdnd11an1n64x5 FILLER_138_1723 ();
 b15zdnd11an1n64x5 FILLER_138_1787 ();
 b15zdnd11an1n16x5 FILLER_138_1851 ();
 b15zdnd00an1n02x5 FILLER_138_1867 ();
 b15zdnd00an1n01x5 FILLER_138_1869 ();
 b15zdnd11an1n64x5 FILLER_138_1882 ();
 b15zdnd11an1n16x5 FILLER_138_1946 ();
 b15zdnd00an1n01x5 FILLER_138_1962 ();
 b15zdnd11an1n64x5 FILLER_138_1975 ();
 b15zdnd11an1n08x5 FILLER_138_2039 ();
 b15zdnd00an1n01x5 FILLER_138_2047 ();
 b15zdnd11an1n32x5 FILLER_138_2059 ();
 b15zdnd11an1n08x5 FILLER_138_2091 ();
 b15zdnd00an1n01x5 FILLER_138_2099 ();
 b15zdnd11an1n32x5 FILLER_138_2111 ();
 b15zdnd11an1n08x5 FILLER_138_2143 ();
 b15zdnd00an1n02x5 FILLER_138_2151 ();
 b15zdnd00an1n01x5 FILLER_138_2153 ();
 b15zdnd11an1n32x5 FILLER_138_2162 ();
 b15zdnd11an1n08x5 FILLER_138_2194 ();
 b15zdnd00an1n01x5 FILLER_138_2202 ();
 b15zdnd11an1n16x5 FILLER_138_2223 ();
 b15zdnd00an1n02x5 FILLER_138_2239 ();
 b15zdnd11an1n08x5 FILLER_138_2245 ();
 b15zdnd00an1n01x5 FILLER_138_2253 ();
 b15zdnd11an1n16x5 FILLER_138_2258 ();
 b15zdnd00an1n02x5 FILLER_138_2274 ();
 b15zdnd11an1n32x5 FILLER_139_0 ();
 b15zdnd11an1n08x5 FILLER_139_49 ();
 b15zdnd00an1n02x5 FILLER_139_57 ();
 b15zdnd11an1n32x5 FILLER_139_77 ();
 b15zdnd11an1n16x5 FILLER_139_109 ();
 b15zdnd11an1n08x5 FILLER_139_125 ();
 b15zdnd00an1n01x5 FILLER_139_133 ();
 b15zdnd11an1n04x5 FILLER_139_144 ();
 b15zdnd11an1n08x5 FILLER_139_154 ();
 b15zdnd11an1n04x5 FILLER_139_162 ();
 b15zdnd00an1n02x5 FILLER_139_166 ();
 b15zdnd00an1n01x5 FILLER_139_168 ();
 b15zdnd11an1n16x5 FILLER_139_180 ();
 b15zdnd11an1n16x5 FILLER_139_203 ();
 b15zdnd11an1n16x5 FILLER_139_224 ();
 b15zdnd11an1n08x5 FILLER_139_240 ();
 b15zdnd00an1n02x5 FILLER_139_248 ();
 b15zdnd00an1n01x5 FILLER_139_250 ();
 b15zdnd11an1n16x5 FILLER_139_272 ();
 b15zdnd11an1n08x5 FILLER_139_288 ();
 b15zdnd11an1n04x5 FILLER_139_296 ();
 b15zdnd11an1n08x5 FILLER_139_304 ();
 b15zdnd11an1n04x5 FILLER_139_312 ();
 b15zdnd00an1n02x5 FILLER_139_316 ();
 b15zdnd00an1n01x5 FILLER_139_318 ();
 b15zdnd11an1n64x5 FILLER_139_333 ();
 b15zdnd11an1n16x5 FILLER_139_397 ();
 b15zdnd11an1n08x5 FILLER_139_413 ();
 b15zdnd00an1n01x5 FILLER_139_421 ();
 b15zdnd11an1n04x5 FILLER_139_443 ();
 b15zdnd11an1n08x5 FILLER_139_455 ();
 b15zdnd11an1n04x5 FILLER_139_463 ();
 b15zdnd00an1n02x5 FILLER_139_467 ();
 b15zdnd11an1n08x5 FILLER_139_475 ();
 b15zdnd11an1n04x5 FILLER_139_483 ();
 b15zdnd00an1n01x5 FILLER_139_487 ();
 b15zdnd11an1n08x5 FILLER_139_499 ();
 b15zdnd11an1n04x5 FILLER_139_507 ();
 b15zdnd00an1n02x5 FILLER_139_511 ();
 b15zdnd11an1n08x5 FILLER_139_529 ();
 b15zdnd00an1n02x5 FILLER_139_537 ();
 b15zdnd11an1n04x5 FILLER_139_553 ();
 b15zdnd11an1n16x5 FILLER_139_565 ();
 b15zdnd11an1n08x5 FILLER_139_581 ();
 b15zdnd11an1n04x5 FILLER_139_589 ();
 b15zdnd00an1n01x5 FILLER_139_593 ();
 b15zdnd11an1n04x5 FILLER_139_603 ();
 b15zdnd11an1n64x5 FILLER_139_615 ();
 b15zdnd11an1n64x5 FILLER_139_679 ();
 b15zdnd11an1n04x5 FILLER_139_743 ();
 b15zdnd00an1n02x5 FILLER_139_747 ();
 b15zdnd00an1n01x5 FILLER_139_749 ();
 b15zdnd11an1n32x5 FILLER_139_770 ();
 b15zdnd11an1n04x5 FILLER_139_802 ();
 b15zdnd00an1n01x5 FILLER_139_806 ();
 b15zdnd11an1n64x5 FILLER_139_827 ();
 b15zdnd11an1n64x5 FILLER_139_891 ();
 b15zdnd11an1n04x5 FILLER_139_955 ();
 b15zdnd00an1n01x5 FILLER_139_959 ();
 b15zdnd11an1n64x5 FILLER_139_983 ();
 b15zdnd11an1n64x5 FILLER_139_1047 ();
 b15zdnd11an1n16x5 FILLER_139_1111 ();
 b15zdnd11an1n08x5 FILLER_139_1158 ();
 b15zdnd11an1n04x5 FILLER_139_1166 ();
 b15zdnd00an1n02x5 FILLER_139_1170 ();
 b15zdnd11an1n04x5 FILLER_139_1192 ();
 b15zdnd11an1n04x5 FILLER_139_1214 ();
 b15zdnd11an1n08x5 FILLER_139_1225 ();
 b15zdnd11an1n04x5 FILLER_139_1233 ();
 b15zdnd00an1n01x5 FILLER_139_1237 ();
 b15zdnd11an1n32x5 FILLER_139_1244 ();
 b15zdnd00an1n02x5 FILLER_139_1276 ();
 b15zdnd00an1n01x5 FILLER_139_1278 ();
 b15zdnd11an1n32x5 FILLER_139_1287 ();
 b15zdnd11an1n16x5 FILLER_139_1319 ();
 b15zdnd11an1n04x5 FILLER_139_1335 ();
 b15zdnd11an1n32x5 FILLER_139_1343 ();
 b15zdnd11an1n08x5 FILLER_139_1375 ();
 b15zdnd11an1n04x5 FILLER_139_1383 ();
 b15zdnd00an1n02x5 FILLER_139_1387 ();
 b15zdnd00an1n01x5 FILLER_139_1389 ();
 b15zdnd11an1n32x5 FILLER_139_1396 ();
 b15zdnd00an1n02x5 FILLER_139_1428 ();
 b15zdnd00an1n01x5 FILLER_139_1430 ();
 b15zdnd11an1n08x5 FILLER_139_1446 ();
 b15zdnd11an1n04x5 FILLER_139_1454 ();
 b15zdnd11an1n04x5 FILLER_139_1465 ();
 b15zdnd11an1n16x5 FILLER_139_1477 ();
 b15zdnd11an1n08x5 FILLER_139_1493 ();
 b15zdnd11an1n04x5 FILLER_139_1513 ();
 b15zdnd00an1n02x5 FILLER_139_1517 ();
 b15zdnd00an1n01x5 FILLER_139_1519 ();
 b15zdnd11an1n16x5 FILLER_139_1529 ();
 b15zdnd11an1n08x5 FILLER_139_1545 ();
 b15zdnd00an1n02x5 FILLER_139_1553 ();
 b15zdnd11an1n32x5 FILLER_139_1562 ();
 b15zdnd11an1n08x5 FILLER_139_1594 ();
 b15zdnd11an1n04x5 FILLER_139_1602 ();
 b15zdnd11an1n04x5 FILLER_139_1618 ();
 b15zdnd11an1n32x5 FILLER_139_1634 ();
 b15zdnd11an1n16x5 FILLER_139_1666 ();
 b15zdnd00an1n02x5 FILLER_139_1682 ();
 b15zdnd11an1n04x5 FILLER_139_1715 ();
 b15zdnd11an1n04x5 FILLER_139_1739 ();
 b15zdnd11an1n16x5 FILLER_139_1763 ();
 b15zdnd11an1n08x5 FILLER_139_1779 ();
 b15zdnd11an1n04x5 FILLER_139_1787 ();
 b15zdnd00an1n01x5 FILLER_139_1791 ();
 b15zdnd11an1n64x5 FILLER_139_1804 ();
 b15zdnd11an1n64x5 FILLER_139_1868 ();
 b15zdnd11an1n64x5 FILLER_139_1932 ();
 b15zdnd11an1n64x5 FILLER_139_1996 ();
 b15zdnd11an1n04x5 FILLER_139_2060 ();
 b15zdnd00an1n02x5 FILLER_139_2064 ();
 b15zdnd11an1n64x5 FILLER_139_2086 ();
 b15zdnd11an1n16x5 FILLER_139_2150 ();
 b15zdnd11an1n08x5 FILLER_139_2166 ();
 b15zdnd00an1n02x5 FILLER_139_2174 ();
 b15zdnd11an1n16x5 FILLER_139_2181 ();
 b15zdnd11an1n08x5 FILLER_139_2197 ();
 b15zdnd11an1n04x5 FILLER_139_2210 ();
 b15zdnd11an1n32x5 FILLER_139_2240 ();
 b15zdnd11an1n08x5 FILLER_139_2272 ();
 b15zdnd11an1n04x5 FILLER_139_2280 ();
 b15zdnd11an1n32x5 FILLER_140_8 ();
 b15zdnd11an1n04x5 FILLER_140_40 ();
 b15zdnd00an1n02x5 FILLER_140_44 ();
 b15zdnd00an1n01x5 FILLER_140_46 ();
 b15zdnd11an1n08x5 FILLER_140_51 ();
 b15zdnd11an1n32x5 FILLER_140_77 ();
 b15zdnd00an1n02x5 FILLER_140_109 ();
 b15zdnd00an1n01x5 FILLER_140_111 ();
 b15zdnd11an1n32x5 FILLER_140_124 ();
 b15zdnd11an1n08x5 FILLER_140_156 ();
 b15zdnd00an1n02x5 FILLER_140_164 ();
 b15zdnd11an1n04x5 FILLER_140_173 ();
 b15zdnd11an1n16x5 FILLER_140_184 ();
 b15zdnd11an1n64x5 FILLER_140_207 ();
 b15zdnd11an1n16x5 FILLER_140_271 ();
 b15zdnd11an1n08x5 FILLER_140_287 ();
 b15zdnd00an1n01x5 FILLER_140_295 ();
 b15zdnd11an1n08x5 FILLER_140_305 ();
 b15zdnd00an1n02x5 FILLER_140_313 ();
 b15zdnd00an1n01x5 FILLER_140_315 ();
 b15zdnd11an1n04x5 FILLER_140_325 ();
 b15zdnd00an1n01x5 FILLER_140_329 ();
 b15zdnd11an1n08x5 FILLER_140_342 ();
 b15zdnd00an1n02x5 FILLER_140_350 ();
 b15zdnd00an1n01x5 FILLER_140_352 ();
 b15zdnd11an1n64x5 FILLER_140_373 ();
 b15zdnd11an1n16x5 FILLER_140_437 ();
 b15zdnd11an1n04x5 FILLER_140_453 ();
 b15zdnd00an1n02x5 FILLER_140_457 ();
 b15zdnd00an1n01x5 FILLER_140_459 ();
 b15zdnd11an1n64x5 FILLER_140_466 ();
 b15zdnd11an1n64x5 FILLER_140_530 ();
 b15zdnd11an1n08x5 FILLER_140_594 ();
 b15zdnd11an1n04x5 FILLER_140_617 ();
 b15zdnd11an1n08x5 FILLER_140_624 ();
 b15zdnd00an1n01x5 FILLER_140_632 ();
 b15zdnd11an1n04x5 FILLER_140_640 ();
 b15zdnd11an1n64x5 FILLER_140_648 ();
 b15zdnd11an1n04x5 FILLER_140_712 ();
 b15zdnd00an1n02x5 FILLER_140_716 ();
 b15zdnd11an1n16x5 FILLER_140_726 ();
 b15zdnd11an1n04x5 FILLER_140_742 ();
 b15zdnd00an1n02x5 FILLER_140_746 ();
 b15zdnd11an1n64x5 FILLER_140_774 ();
 b15zdnd11an1n32x5 FILLER_140_838 ();
 b15zdnd00an1n02x5 FILLER_140_870 ();
 b15zdnd11an1n04x5 FILLER_140_892 ();
 b15zdnd11an1n64x5 FILLER_140_916 ();
 b15zdnd11an1n16x5 FILLER_140_980 ();
 b15zdnd11an1n08x5 FILLER_140_996 ();
 b15zdnd00an1n02x5 FILLER_140_1004 ();
 b15zdnd11an1n08x5 FILLER_140_1016 ();
 b15zdnd11an1n04x5 FILLER_140_1039 ();
 b15zdnd00an1n02x5 FILLER_140_1043 ();
 b15zdnd11an1n64x5 FILLER_140_1076 ();
 b15zdnd11an1n64x5 FILLER_140_1140 ();
 b15zdnd11an1n64x5 FILLER_140_1204 ();
 b15zdnd11an1n32x5 FILLER_140_1268 ();
 b15zdnd00an1n01x5 FILLER_140_1300 ();
 b15zdnd11an1n16x5 FILLER_140_1306 ();
 b15zdnd00an1n01x5 FILLER_140_1322 ();
 b15zdnd11an1n32x5 FILLER_140_1328 ();
 b15zdnd11an1n16x5 FILLER_140_1360 ();
 b15zdnd00an1n02x5 FILLER_140_1376 ();
 b15zdnd11an1n04x5 FILLER_140_1385 ();
 b15zdnd00an1n02x5 FILLER_140_1389 ();
 b15zdnd11an1n64x5 FILLER_140_1397 ();
 b15zdnd11an1n04x5 FILLER_140_1461 ();
 b15zdnd00an1n01x5 FILLER_140_1465 ();
 b15zdnd11an1n16x5 FILLER_140_1476 ();
 b15zdnd11an1n08x5 FILLER_140_1492 ();
 b15zdnd00an1n01x5 FILLER_140_1500 ();
 b15zdnd11an1n08x5 FILLER_140_1506 ();
 b15zdnd00an1n01x5 FILLER_140_1514 ();
 b15zdnd11an1n32x5 FILLER_140_1523 ();
 b15zdnd11an1n16x5 FILLER_140_1555 ();
 b15zdnd00an1n02x5 FILLER_140_1571 ();
 b15zdnd00an1n01x5 FILLER_140_1573 ();
 b15zdnd11an1n16x5 FILLER_140_1600 ();
 b15zdnd11an1n08x5 FILLER_140_1616 ();
 b15zdnd11an1n04x5 FILLER_140_1624 ();
 b15zdnd00an1n02x5 FILLER_140_1628 ();
 b15zdnd00an1n01x5 FILLER_140_1630 ();
 b15zdnd11an1n64x5 FILLER_140_1635 ();
 b15zdnd11an1n64x5 FILLER_140_1699 ();
 b15zdnd11an1n32x5 FILLER_140_1763 ();
 b15zdnd11an1n08x5 FILLER_140_1795 ();
 b15zdnd11an1n04x5 FILLER_140_1814 ();
 b15zdnd11an1n16x5 FILLER_140_1849 ();
 b15zdnd00an1n02x5 FILLER_140_1865 ();
 b15zdnd00an1n01x5 FILLER_140_1867 ();
 b15zdnd11an1n64x5 FILLER_140_1877 ();
 b15zdnd11an1n64x5 FILLER_140_1941 ();
 b15zdnd11an1n64x5 FILLER_140_2005 ();
 b15zdnd11an1n64x5 FILLER_140_2069 ();
 b15zdnd11an1n16x5 FILLER_140_2133 ();
 b15zdnd11an1n04x5 FILLER_140_2149 ();
 b15zdnd00an1n01x5 FILLER_140_2153 ();
 b15zdnd11an1n08x5 FILLER_140_2162 ();
 b15zdnd11an1n08x5 FILLER_140_2190 ();
 b15zdnd00an1n02x5 FILLER_140_2198 ();
 b15zdnd00an1n01x5 FILLER_140_2200 ();
 b15zdnd11an1n32x5 FILLER_140_2207 ();
 b15zdnd11an1n08x5 FILLER_140_2239 ();
 b15zdnd00an1n01x5 FILLER_140_2247 ();
 b15zdnd11an1n16x5 FILLER_140_2259 ();
 b15zdnd00an1n01x5 FILLER_140_2275 ();
 b15zdnd11an1n32x5 FILLER_141_0 ();
 b15zdnd11an1n16x5 FILLER_141_32 ();
 b15zdnd00an1n02x5 FILLER_141_48 ();
 b15zdnd11an1n04x5 FILLER_141_54 ();
 b15zdnd11an1n04x5 FILLER_141_64 ();
 b15zdnd00an1n02x5 FILLER_141_68 ();
 b15zdnd11an1n08x5 FILLER_141_79 ();
 b15zdnd00an1n01x5 FILLER_141_87 ();
 b15zdnd11an1n08x5 FILLER_141_105 ();
 b15zdnd00an1n02x5 FILLER_141_113 ();
 b15zdnd11an1n08x5 FILLER_141_121 ();
 b15zdnd11an1n64x5 FILLER_141_145 ();
 b15zdnd11an1n64x5 FILLER_141_209 ();
 b15zdnd00an1n02x5 FILLER_141_273 ();
 b15zdnd11an1n16x5 FILLER_141_290 ();
 b15zdnd11an1n08x5 FILLER_141_306 ();
 b15zdnd00an1n02x5 FILLER_141_314 ();
 b15zdnd00an1n01x5 FILLER_141_316 ();
 b15zdnd11an1n16x5 FILLER_141_329 ();
 b15zdnd11an1n08x5 FILLER_141_345 ();
 b15zdnd11an1n04x5 FILLER_141_353 ();
 b15zdnd11an1n64x5 FILLER_141_365 ();
 b15zdnd11an1n16x5 FILLER_141_429 ();
 b15zdnd11an1n08x5 FILLER_141_445 ();
 b15zdnd00an1n01x5 FILLER_141_453 ();
 b15zdnd11an1n04x5 FILLER_141_469 ();
 b15zdnd00an1n02x5 FILLER_141_473 ();
 b15zdnd11an1n32x5 FILLER_141_490 ();
 b15zdnd11an1n16x5 FILLER_141_522 ();
 b15zdnd11an1n08x5 FILLER_141_538 ();
 b15zdnd00an1n01x5 FILLER_141_546 ();
 b15zdnd11an1n32x5 FILLER_141_573 ();
 b15zdnd11an1n16x5 FILLER_141_605 ();
 b15zdnd11an1n08x5 FILLER_141_621 ();
 b15zdnd11an1n04x5 FILLER_141_629 ();
 b15zdnd00an1n02x5 FILLER_141_633 ();
 b15zdnd11an1n08x5 FILLER_141_644 ();
 b15zdnd11an1n04x5 FILLER_141_652 ();
 b15zdnd00an1n02x5 FILLER_141_656 ();
 b15zdnd11an1n04x5 FILLER_141_676 ();
 b15zdnd11an1n64x5 FILLER_141_692 ();
 b15zdnd11an1n64x5 FILLER_141_756 ();
 b15zdnd11an1n64x5 FILLER_141_820 ();
 b15zdnd11an1n16x5 FILLER_141_884 ();
 b15zdnd11an1n08x5 FILLER_141_900 ();
 b15zdnd00an1n02x5 FILLER_141_908 ();
 b15zdnd00an1n01x5 FILLER_141_910 ();
 b15zdnd11an1n64x5 FILLER_141_920 ();
 b15zdnd11an1n16x5 FILLER_141_984 ();
 b15zdnd11an1n08x5 FILLER_141_1000 ();
 b15zdnd00an1n02x5 FILLER_141_1008 ();
 b15zdnd11an1n08x5 FILLER_141_1019 ();
 b15zdnd11an1n04x5 FILLER_141_1027 ();
 b15zdnd11an1n32x5 FILLER_141_1046 ();
 b15zdnd11an1n16x5 FILLER_141_1078 ();
 b15zdnd11an1n08x5 FILLER_141_1094 ();
 b15zdnd11an1n64x5 FILLER_141_1112 ();
 b15zdnd11an1n32x5 FILLER_141_1176 ();
 b15zdnd11an1n04x5 FILLER_141_1208 ();
 b15zdnd00an1n02x5 FILLER_141_1212 ();
 b15zdnd00an1n01x5 FILLER_141_1214 ();
 b15zdnd11an1n04x5 FILLER_141_1226 ();
 b15zdnd11an1n32x5 FILLER_141_1246 ();
 b15zdnd11an1n04x5 FILLER_141_1278 ();
 b15zdnd00an1n02x5 FILLER_141_1282 ();
 b15zdnd00an1n01x5 FILLER_141_1284 ();
 b15zdnd11an1n04x5 FILLER_141_1301 ();
 b15zdnd11an1n08x5 FILLER_141_1321 ();
 b15zdnd00an1n02x5 FILLER_141_1329 ();
 b15zdnd11an1n16x5 FILLER_141_1338 ();
 b15zdnd00an1n01x5 FILLER_141_1354 ();
 b15zdnd11an1n04x5 FILLER_141_1359 ();
 b15zdnd11an1n16x5 FILLER_141_1377 ();
 b15zdnd11an1n08x5 FILLER_141_1393 ();
 b15zdnd11an1n04x5 FILLER_141_1401 ();
 b15zdnd00an1n01x5 FILLER_141_1405 ();
 b15zdnd11an1n16x5 FILLER_141_1418 ();
 b15zdnd11an1n08x5 FILLER_141_1434 ();
 b15zdnd11an1n04x5 FILLER_141_1442 ();
 b15zdnd11an1n64x5 FILLER_141_1458 ();
 b15zdnd11an1n64x5 FILLER_141_1522 ();
 b15zdnd11an1n64x5 FILLER_141_1586 ();
 b15zdnd11an1n08x5 FILLER_141_1650 ();
 b15zdnd00an1n01x5 FILLER_141_1658 ();
 b15zdnd11an1n64x5 FILLER_141_1679 ();
 b15zdnd11an1n64x5 FILLER_141_1743 ();
 b15zdnd11an1n04x5 FILLER_141_1807 ();
 b15zdnd00an1n02x5 FILLER_141_1811 ();
 b15zdnd00an1n01x5 FILLER_141_1813 ();
 b15zdnd11an1n04x5 FILLER_141_1871 ();
 b15zdnd11an1n64x5 FILLER_141_1884 ();
 b15zdnd11an1n32x5 FILLER_141_1948 ();
 b15zdnd11an1n08x5 FILLER_141_1980 ();
 b15zdnd11an1n04x5 FILLER_141_1988 ();
 b15zdnd00an1n01x5 FILLER_141_1992 ();
 b15zdnd11an1n32x5 FILLER_141_2012 ();
 b15zdnd11an1n16x5 FILLER_141_2044 ();
 b15zdnd11an1n04x5 FILLER_141_2060 ();
 b15zdnd00an1n01x5 FILLER_141_2064 ();
 b15zdnd11an1n32x5 FILLER_141_2074 ();
 b15zdnd11an1n16x5 FILLER_141_2106 ();
 b15zdnd00an1n01x5 FILLER_141_2122 ();
 b15zdnd11an1n04x5 FILLER_141_2143 ();
 b15zdnd11an1n32x5 FILLER_141_2152 ();
 b15zdnd11an1n04x5 FILLER_141_2184 ();
 b15zdnd11an1n32x5 FILLER_141_2192 ();
 b15zdnd11an1n08x5 FILLER_141_2224 ();
 b15zdnd00an1n02x5 FILLER_141_2232 ();
 b15zdnd11an1n08x5 FILLER_141_2254 ();
 b15zdnd11an1n04x5 FILLER_141_2266 ();
 b15zdnd11an1n08x5 FILLER_141_2274 ();
 b15zdnd00an1n02x5 FILLER_141_2282 ();
 b15zdnd11an1n64x5 FILLER_142_8 ();
 b15zdnd11an1n32x5 FILLER_142_72 ();
 b15zdnd11an1n08x5 FILLER_142_104 ();
 b15zdnd00an1n02x5 FILLER_142_112 ();
 b15zdnd11an1n32x5 FILLER_142_120 ();
 b15zdnd11an1n08x5 FILLER_142_152 ();
 b15zdnd11an1n04x5 FILLER_142_160 ();
 b15zdnd00an1n02x5 FILLER_142_164 ();
 b15zdnd11an1n64x5 FILLER_142_175 ();
 b15zdnd11an1n64x5 FILLER_142_239 ();
 b15zdnd11an1n16x5 FILLER_142_303 ();
 b15zdnd11an1n04x5 FILLER_142_319 ();
 b15zdnd00an1n02x5 FILLER_142_323 ();
 b15zdnd11an1n16x5 FILLER_142_329 ();
 b15zdnd11an1n04x5 FILLER_142_345 ();
 b15zdnd11an1n64x5 FILLER_142_354 ();
 b15zdnd11an1n08x5 FILLER_142_418 ();
 b15zdnd00an1n01x5 FILLER_142_426 ();
 b15zdnd11an1n08x5 FILLER_142_443 ();
 b15zdnd11an1n04x5 FILLER_142_451 ();
 b15zdnd00an1n02x5 FILLER_142_455 ();
 b15zdnd11an1n08x5 FILLER_142_475 ();
 b15zdnd00an1n01x5 FILLER_142_483 ();
 b15zdnd11an1n04x5 FILLER_142_490 ();
 b15zdnd00an1n02x5 FILLER_142_494 ();
 b15zdnd11an1n64x5 FILLER_142_502 ();
 b15zdnd11an1n08x5 FILLER_142_566 ();
 b15zdnd00an1n01x5 FILLER_142_574 ();
 b15zdnd11an1n64x5 FILLER_142_585 ();
 b15zdnd11an1n04x5 FILLER_142_649 ();
 b15zdnd00an1n01x5 FILLER_142_653 ();
 b15zdnd11an1n32x5 FILLER_142_680 ();
 b15zdnd11an1n04x5 FILLER_142_712 ();
 b15zdnd00an1n02x5 FILLER_142_716 ();
 b15zdnd11an1n04x5 FILLER_142_726 ();
 b15zdnd00an1n01x5 FILLER_142_730 ();
 b15zdnd11an1n08x5 FILLER_142_739 ();
 b15zdnd11an1n04x5 FILLER_142_747 ();
 b15zdnd00an1n02x5 FILLER_142_751 ();
 b15zdnd11an1n08x5 FILLER_142_779 ();
 b15zdnd00an1n02x5 FILLER_142_787 ();
 b15zdnd00an1n01x5 FILLER_142_789 ();
 b15zdnd11an1n64x5 FILLER_142_793 ();
 b15zdnd11an1n08x5 FILLER_142_857 ();
 b15zdnd11an1n04x5 FILLER_142_865 ();
 b15zdnd00an1n01x5 FILLER_142_869 ();
 b15zdnd11an1n32x5 FILLER_142_881 ();
 b15zdnd11an1n08x5 FILLER_142_913 ();
 b15zdnd00an1n02x5 FILLER_142_921 ();
 b15zdnd00an1n01x5 FILLER_142_923 ();
 b15zdnd11an1n16x5 FILLER_142_944 ();
 b15zdnd11an1n04x5 FILLER_142_960 ();
 b15zdnd00an1n02x5 FILLER_142_964 ();
 b15zdnd11an1n64x5 FILLER_142_970 ();
 b15zdnd11an1n64x5 FILLER_142_1034 ();
 b15zdnd11an1n64x5 FILLER_142_1098 ();
 b15zdnd11an1n08x5 FILLER_142_1162 ();
 b15zdnd11an1n04x5 FILLER_142_1170 ();
 b15zdnd11an1n16x5 FILLER_142_1186 ();
 b15zdnd00an1n02x5 FILLER_142_1202 ();
 b15zdnd11an1n04x5 FILLER_142_1210 ();
 b15zdnd11an1n64x5 FILLER_142_1221 ();
 b15zdnd11an1n04x5 FILLER_142_1285 ();
 b15zdnd11an1n08x5 FILLER_142_1294 ();
 b15zdnd11an1n08x5 FILLER_142_1308 ();
 b15zdnd11an1n04x5 FILLER_142_1316 ();
 b15zdnd11an1n04x5 FILLER_142_1329 ();
 b15zdnd11an1n16x5 FILLER_142_1343 ();
 b15zdnd11an1n04x5 FILLER_142_1359 ();
 b15zdnd11an1n08x5 FILLER_142_1372 ();
 b15zdnd00an1n02x5 FILLER_142_1380 ();
 b15zdnd00an1n01x5 FILLER_142_1382 ();
 b15zdnd11an1n16x5 FILLER_142_1399 ();
 b15zdnd11an1n04x5 FILLER_142_1415 ();
 b15zdnd00an1n02x5 FILLER_142_1419 ();
 b15zdnd00an1n01x5 FILLER_142_1421 ();
 b15zdnd11an1n04x5 FILLER_142_1429 ();
 b15zdnd11an1n64x5 FILLER_142_1437 ();
 b15zdnd11an1n08x5 FILLER_142_1501 ();
 b15zdnd11an1n04x5 FILLER_142_1509 ();
 b15zdnd00an1n02x5 FILLER_142_1513 ();
 b15zdnd00an1n01x5 FILLER_142_1515 ();
 b15zdnd11an1n16x5 FILLER_142_1532 ();
 b15zdnd11an1n04x5 FILLER_142_1554 ();
 b15zdnd11an1n32x5 FILLER_142_1565 ();
 b15zdnd11an1n16x5 FILLER_142_1597 ();
 b15zdnd11an1n08x5 FILLER_142_1613 ();
 b15zdnd11an1n16x5 FILLER_142_1641 ();
 b15zdnd11an1n08x5 FILLER_142_1657 ();
 b15zdnd00an1n01x5 FILLER_142_1665 ();
 b15zdnd11an1n04x5 FILLER_142_1671 ();
 b15zdnd11an1n64x5 FILLER_142_1680 ();
 b15zdnd11an1n64x5 FILLER_142_1744 ();
 b15zdnd11an1n08x5 FILLER_142_1808 ();
 b15zdnd00an1n02x5 FILLER_142_1816 ();
 b15zdnd11an1n32x5 FILLER_142_1827 ();
 b15zdnd11an1n16x5 FILLER_142_1859 ();
 b15zdnd11an1n08x5 FILLER_142_1875 ();
 b15zdnd00an1n02x5 FILLER_142_1883 ();
 b15zdnd00an1n01x5 FILLER_142_1885 ();
 b15zdnd11an1n04x5 FILLER_142_1897 ();
 b15zdnd11an1n08x5 FILLER_142_1910 ();
 b15zdnd11an1n04x5 FILLER_142_1918 ();
 b15zdnd11an1n64x5 FILLER_142_1931 ();
 b15zdnd00an1n02x5 FILLER_142_1995 ();
 b15zdnd00an1n01x5 FILLER_142_1997 ();
 b15zdnd11an1n32x5 FILLER_142_2007 ();
 b15zdnd11an1n16x5 FILLER_142_2039 ();
 b15zdnd11an1n08x5 FILLER_142_2055 ();
 b15zdnd11an1n04x5 FILLER_142_2063 ();
 b15zdnd00an1n02x5 FILLER_142_2067 ();
 b15zdnd11an1n32x5 FILLER_142_2081 ();
 b15zdnd00an1n01x5 FILLER_142_2113 ();
 b15zdnd11an1n08x5 FILLER_142_2134 ();
 b15zdnd11an1n04x5 FILLER_142_2148 ();
 b15zdnd00an1n02x5 FILLER_142_2152 ();
 b15zdnd11an1n32x5 FILLER_142_2162 ();
 b15zdnd11an1n16x5 FILLER_142_2194 ();
 b15zdnd11an1n08x5 FILLER_142_2210 ();
 b15zdnd11an1n04x5 FILLER_142_2218 ();
 b15zdnd11an1n04x5 FILLER_142_2242 ();
 b15zdnd11an1n04x5 FILLER_142_2258 ();
 b15zdnd11an1n04x5 FILLER_142_2266 ();
 b15zdnd00an1n02x5 FILLER_142_2274 ();
 b15zdnd11an1n64x5 FILLER_143_0 ();
 b15zdnd11an1n64x5 FILLER_143_64 ();
 b15zdnd11an1n64x5 FILLER_143_128 ();
 b15zdnd11an1n08x5 FILLER_143_192 ();
 b15zdnd11an1n08x5 FILLER_143_204 ();
 b15zdnd11an1n04x5 FILLER_143_212 ();
 b15zdnd00an1n02x5 FILLER_143_216 ();
 b15zdnd11an1n04x5 FILLER_143_224 ();
 b15zdnd11an1n16x5 FILLER_143_242 ();
 b15zdnd11an1n16x5 FILLER_143_267 ();
 b15zdnd00an1n01x5 FILLER_143_283 ();
 b15zdnd11an1n04x5 FILLER_143_296 ();
 b15zdnd11an1n04x5 FILLER_143_321 ();
 b15zdnd11an1n64x5 FILLER_143_335 ();
 b15zdnd11an1n08x5 FILLER_143_399 ();
 b15zdnd11an1n04x5 FILLER_143_407 ();
 b15zdnd00an1n02x5 FILLER_143_411 ();
 b15zdnd11an1n08x5 FILLER_143_419 ();
 b15zdnd00an1n02x5 FILLER_143_427 ();
 b15zdnd11an1n04x5 FILLER_143_445 ();
 b15zdnd11an1n32x5 FILLER_143_475 ();
 b15zdnd11an1n04x5 FILLER_143_507 ();
 b15zdnd00an1n02x5 FILLER_143_511 ();
 b15zdnd11an1n04x5 FILLER_143_517 ();
 b15zdnd00an1n01x5 FILLER_143_521 ();
 b15zdnd11an1n08x5 FILLER_143_525 ();
 b15zdnd11an1n04x5 FILLER_143_533 ();
 b15zdnd11an1n64x5 FILLER_143_542 ();
 b15zdnd11an1n08x5 FILLER_143_606 ();
 b15zdnd11an1n04x5 FILLER_143_619 ();
 b15zdnd11an1n32x5 FILLER_143_635 ();
 b15zdnd00an1n02x5 FILLER_143_667 ();
 b15zdnd11an1n04x5 FILLER_143_685 ();
 b15zdnd11an1n08x5 FILLER_143_715 ();
 b15zdnd00an1n02x5 FILLER_143_723 ();
 b15zdnd11an1n08x5 FILLER_143_730 ();
 b15zdnd11an1n04x5 FILLER_143_738 ();
 b15zdnd11an1n04x5 FILLER_143_768 ();
 b15zdnd11an1n16x5 FILLER_143_792 ();
 b15zdnd11an1n08x5 FILLER_143_808 ();
 b15zdnd11an1n04x5 FILLER_143_816 ();
 b15zdnd00an1n01x5 FILLER_143_820 ();
 b15zdnd11an1n04x5 FILLER_143_841 ();
 b15zdnd11an1n64x5 FILLER_143_850 ();
 b15zdnd11an1n32x5 FILLER_143_914 ();
 b15zdnd11an1n08x5 FILLER_143_946 ();
 b15zdnd11an1n04x5 FILLER_143_954 ();
 b15zdnd00an1n02x5 FILLER_143_958 ();
 b15zdnd00an1n01x5 FILLER_143_960 ();
 b15zdnd11an1n08x5 FILLER_143_966 ();
 b15zdnd11an1n04x5 FILLER_143_974 ();
 b15zdnd00an1n02x5 FILLER_143_978 ();
 b15zdnd11an1n64x5 FILLER_143_989 ();
 b15zdnd11an1n32x5 FILLER_143_1053 ();
 b15zdnd00an1n01x5 FILLER_143_1085 ();
 b15zdnd11an1n16x5 FILLER_143_1107 ();
 b15zdnd00an1n02x5 FILLER_143_1123 ();
 b15zdnd11an1n64x5 FILLER_143_1134 ();
 b15zdnd11an1n08x5 FILLER_143_1198 ();
 b15zdnd11an1n04x5 FILLER_143_1206 ();
 b15zdnd00an1n02x5 FILLER_143_1210 ();
 b15zdnd00an1n01x5 FILLER_143_1212 ();
 b15zdnd11an1n64x5 FILLER_143_1222 ();
 b15zdnd11an1n04x5 FILLER_143_1286 ();
 b15zdnd11an1n32x5 FILLER_143_1299 ();
 b15zdnd11an1n16x5 FILLER_143_1331 ();
 b15zdnd11an1n08x5 FILLER_143_1347 ();
 b15zdnd11an1n04x5 FILLER_143_1355 ();
 b15zdnd00an1n02x5 FILLER_143_1359 ();
 b15zdnd11an1n64x5 FILLER_143_1371 ();
 b15zdnd11an1n64x5 FILLER_143_1435 ();
 b15zdnd11an1n08x5 FILLER_143_1499 ();
 b15zdnd11an1n04x5 FILLER_143_1507 ();
 b15zdnd00an1n02x5 FILLER_143_1511 ();
 b15zdnd11an1n32x5 FILLER_143_1516 ();
 b15zdnd11an1n04x5 FILLER_143_1548 ();
 b15zdnd00an1n01x5 FILLER_143_1552 ();
 b15zdnd11an1n64x5 FILLER_143_1563 ();
 b15zdnd11an1n64x5 FILLER_143_1627 ();
 b15zdnd11an1n16x5 FILLER_143_1691 ();
 b15zdnd11an1n04x5 FILLER_143_1707 ();
 b15zdnd00an1n01x5 FILLER_143_1711 ();
 b15zdnd11an1n64x5 FILLER_143_1732 ();
 b15zdnd11an1n32x5 FILLER_143_1796 ();
 b15zdnd11an1n08x5 FILLER_143_1828 ();
 b15zdnd00an1n01x5 FILLER_143_1836 ();
 b15zdnd11an1n04x5 FILLER_143_1848 ();
 b15zdnd11an1n04x5 FILLER_143_1883 ();
 b15zdnd11an1n04x5 FILLER_143_1902 ();
 b15zdnd11an1n32x5 FILLER_143_1927 ();
 b15zdnd11an1n08x5 FILLER_143_1959 ();
 b15zdnd00an1n02x5 FILLER_143_1967 ();
 b15zdnd11an1n04x5 FILLER_143_1978 ();
 b15zdnd11an1n04x5 FILLER_143_1991 ();
 b15zdnd11an1n16x5 FILLER_143_2006 ();
 b15zdnd11an1n08x5 FILLER_143_2022 ();
 b15zdnd00an1n02x5 FILLER_143_2030 ();
 b15zdnd11an1n64x5 FILLER_143_2044 ();
 b15zdnd11an1n08x5 FILLER_143_2108 ();
 b15zdnd11an1n04x5 FILLER_143_2116 ();
 b15zdnd11an1n04x5 FILLER_143_2125 ();
 b15zdnd11an1n64x5 FILLER_143_2132 ();
 b15zdnd11an1n32x5 FILLER_143_2196 ();
 b15zdnd11an1n16x5 FILLER_143_2228 ();
 b15zdnd11an1n08x5 FILLER_143_2244 ();
 b15zdnd00an1n01x5 FILLER_143_2252 ();
 b15zdnd11an1n04x5 FILLER_143_2257 ();
 b15zdnd11an1n16x5 FILLER_143_2265 ();
 b15zdnd00an1n02x5 FILLER_143_2281 ();
 b15zdnd00an1n01x5 FILLER_143_2283 ();
 b15zdnd11an1n16x5 FILLER_144_8 ();
 b15zdnd11an1n08x5 FILLER_144_24 ();
 b15zdnd11an1n04x5 FILLER_144_32 ();
 b15zdnd00an1n02x5 FILLER_144_36 ();
 b15zdnd11an1n04x5 FILLER_144_44 ();
 b15zdnd00an1n02x5 FILLER_144_48 ();
 b15zdnd11an1n64x5 FILLER_144_54 ();
 b15zdnd11an1n16x5 FILLER_144_130 ();
 b15zdnd11an1n32x5 FILLER_144_153 ();
 b15zdnd11an1n04x5 FILLER_144_185 ();
 b15zdnd11an1n08x5 FILLER_144_204 ();
 b15zdnd11an1n04x5 FILLER_144_212 ();
 b15zdnd00an1n01x5 FILLER_144_216 ();
 b15zdnd11an1n16x5 FILLER_144_224 ();
 b15zdnd11an1n08x5 FILLER_144_240 ();
 b15zdnd11an1n04x5 FILLER_144_248 ();
 b15zdnd00an1n02x5 FILLER_144_252 ();
 b15zdnd11an1n32x5 FILLER_144_263 ();
 b15zdnd11an1n04x5 FILLER_144_295 ();
 b15zdnd00an1n02x5 FILLER_144_299 ();
 b15zdnd11an1n32x5 FILLER_144_313 ();
 b15zdnd00an1n01x5 FILLER_144_345 ();
 b15zdnd11an1n04x5 FILLER_144_354 ();
 b15zdnd11an1n64x5 FILLER_144_364 ();
 b15zdnd11an1n64x5 FILLER_144_428 ();
 b15zdnd11an1n32x5 FILLER_144_492 ();
 b15zdnd11an1n08x5 FILLER_144_524 ();
 b15zdnd11an1n04x5 FILLER_144_532 ();
 b15zdnd00an1n01x5 FILLER_144_536 ();
 b15zdnd11an1n32x5 FILLER_144_542 ();
 b15zdnd11an1n04x5 FILLER_144_574 ();
 b15zdnd11an1n64x5 FILLER_144_581 ();
 b15zdnd11an1n16x5 FILLER_144_645 ();
 b15zdnd11an1n04x5 FILLER_144_661 ();
 b15zdnd11an1n16x5 FILLER_144_685 ();
 b15zdnd11an1n04x5 FILLER_144_701 ();
 b15zdnd00an1n02x5 FILLER_144_716 ();
 b15zdnd11an1n32x5 FILLER_144_726 ();
 b15zdnd11an1n04x5 FILLER_144_758 ();
 b15zdnd00an1n02x5 FILLER_144_762 ();
 b15zdnd11an1n04x5 FILLER_144_768 ();
 b15zdnd11an1n32x5 FILLER_144_777 ();
 b15zdnd11an1n16x5 FILLER_144_809 ();
 b15zdnd11an1n04x5 FILLER_144_825 ();
 b15zdnd00an1n02x5 FILLER_144_829 ();
 b15zdnd11an1n64x5 FILLER_144_840 ();
 b15zdnd11an1n64x5 FILLER_144_904 ();
 b15zdnd11an1n16x5 FILLER_144_968 ();
 b15zdnd11an1n16x5 FILLER_144_1001 ();
 b15zdnd11an1n08x5 FILLER_144_1017 ();
 b15zdnd00an1n02x5 FILLER_144_1025 ();
 b15zdnd11an1n32x5 FILLER_144_1038 ();
 b15zdnd11an1n16x5 FILLER_144_1070 ();
 b15zdnd11an1n08x5 FILLER_144_1086 ();
 b15zdnd11an1n04x5 FILLER_144_1094 ();
 b15zdnd11an1n04x5 FILLER_144_1102 ();
 b15zdnd11an1n16x5 FILLER_144_1111 ();
 b15zdnd00an1n01x5 FILLER_144_1127 ();
 b15zdnd11an1n16x5 FILLER_144_1148 ();
 b15zdnd11an1n08x5 FILLER_144_1164 ();
 b15zdnd00an1n02x5 FILLER_144_1172 ();
 b15zdnd00an1n01x5 FILLER_144_1174 ();
 b15zdnd11an1n16x5 FILLER_144_1206 ();
 b15zdnd00an1n01x5 FILLER_144_1222 ();
 b15zdnd11an1n04x5 FILLER_144_1228 ();
 b15zdnd11an1n16x5 FILLER_144_1255 ();
 b15zdnd11an1n08x5 FILLER_144_1271 ();
 b15zdnd00an1n02x5 FILLER_144_1279 ();
 b15zdnd00an1n01x5 FILLER_144_1281 ();
 b15zdnd11an1n16x5 FILLER_144_1292 ();
 b15zdnd00an1n02x5 FILLER_144_1308 ();
 b15zdnd00an1n01x5 FILLER_144_1310 ();
 b15zdnd11an1n64x5 FILLER_144_1323 ();
 b15zdnd11an1n04x5 FILLER_144_1387 ();
 b15zdnd00an1n02x5 FILLER_144_1391 ();
 b15zdnd11an1n16x5 FILLER_144_1404 ();
 b15zdnd00an1n02x5 FILLER_144_1420 ();
 b15zdnd00an1n01x5 FILLER_144_1422 ();
 b15zdnd11an1n08x5 FILLER_144_1428 ();
 b15zdnd11an1n04x5 FILLER_144_1436 ();
 b15zdnd00an1n02x5 FILLER_144_1440 ();
 b15zdnd00an1n01x5 FILLER_144_1442 ();
 b15zdnd11an1n04x5 FILLER_144_1461 ();
 b15zdnd00an1n01x5 FILLER_144_1465 ();
 b15zdnd11an1n08x5 FILLER_144_1476 ();
 b15zdnd00an1n02x5 FILLER_144_1484 ();
 b15zdnd11an1n04x5 FILLER_144_1497 ();
 b15zdnd11an1n32x5 FILLER_144_1527 ();
 b15zdnd11an1n16x5 FILLER_144_1559 ();
 b15zdnd00an1n01x5 FILLER_144_1575 ();
 b15zdnd11an1n04x5 FILLER_144_1594 ();
 b15zdnd11an1n04x5 FILLER_144_1607 ();
 b15zdnd11an1n08x5 FILLER_144_1616 ();
 b15zdnd11an1n32x5 FILLER_144_1630 ();
 b15zdnd11an1n08x5 FILLER_144_1662 ();
 b15zdnd11an1n04x5 FILLER_144_1670 ();
 b15zdnd11an1n04x5 FILLER_144_1705 ();
 b15zdnd00an1n02x5 FILLER_144_1709 ();
 b15zdnd00an1n01x5 FILLER_144_1711 ();
 b15zdnd11an1n64x5 FILLER_144_1717 ();
 b15zdnd11an1n08x5 FILLER_144_1781 ();
 b15zdnd00an1n02x5 FILLER_144_1789 ();
 b15zdnd11an1n04x5 FILLER_144_1817 ();
 b15zdnd11an1n04x5 FILLER_144_1862 ();
 b15zdnd11an1n32x5 FILLER_144_1875 ();
 b15zdnd00an1n02x5 FILLER_144_1907 ();
 b15zdnd00an1n01x5 FILLER_144_1909 ();
 b15zdnd11an1n32x5 FILLER_144_1941 ();
 b15zdnd00an1n01x5 FILLER_144_1973 ();
 b15zdnd11an1n16x5 FILLER_144_2005 ();
 b15zdnd11an1n08x5 FILLER_144_2021 ();
 b15zdnd11an1n04x5 FILLER_144_2029 ();
 b15zdnd11an1n64x5 FILLER_144_2042 ();
 b15zdnd11an1n32x5 FILLER_144_2106 ();
 b15zdnd11an1n16x5 FILLER_144_2138 ();
 b15zdnd11an1n64x5 FILLER_144_2162 ();
 b15zdnd11an1n16x5 FILLER_144_2226 ();
 b15zdnd11an1n04x5 FILLER_144_2242 ();
 b15zdnd00an1n01x5 FILLER_144_2246 ();
 b15zdnd11an1n04x5 FILLER_144_2258 ();
 b15zdnd11an1n08x5 FILLER_144_2266 ();
 b15zdnd00an1n02x5 FILLER_144_2274 ();
 b15zdnd11an1n32x5 FILLER_145_0 ();
 b15zdnd11an1n08x5 FILLER_145_32 ();
 b15zdnd11an1n16x5 FILLER_145_56 ();
 b15zdnd11an1n04x5 FILLER_145_72 ();
 b15zdnd00an1n02x5 FILLER_145_76 ();
 b15zdnd11an1n04x5 FILLER_145_83 ();
 b15zdnd11an1n08x5 FILLER_145_96 ();
 b15zdnd11an1n04x5 FILLER_145_104 ();
 b15zdnd00an1n02x5 FILLER_145_108 ();
 b15zdnd00an1n01x5 FILLER_145_110 ();
 b15zdnd11an1n16x5 FILLER_145_115 ();
 b15zdnd00an1n02x5 FILLER_145_131 ();
 b15zdnd11an1n04x5 FILLER_145_143 ();
 b15zdnd11an1n16x5 FILLER_145_157 ();
 b15zdnd00an1n01x5 FILLER_145_173 ();
 b15zdnd11an1n04x5 FILLER_145_193 ();
 b15zdnd11an1n08x5 FILLER_145_203 ();
 b15zdnd11an1n16x5 FILLER_145_225 ();
 b15zdnd11an1n04x5 FILLER_145_241 ();
 b15zdnd11an1n16x5 FILLER_145_252 ();
 b15zdnd11an1n08x5 FILLER_145_268 ();
 b15zdnd11an1n04x5 FILLER_145_276 ();
 b15zdnd00an1n02x5 FILLER_145_280 ();
 b15zdnd00an1n01x5 FILLER_145_282 ();
 b15zdnd11an1n32x5 FILLER_145_295 ();
 b15zdnd11an1n16x5 FILLER_145_327 ();
 b15zdnd11an1n08x5 FILLER_145_343 ();
 b15zdnd00an1n02x5 FILLER_145_351 ();
 b15zdnd11an1n04x5 FILLER_145_358 ();
 b15zdnd00an1n01x5 FILLER_145_362 ();
 b15zdnd11an1n64x5 FILLER_145_369 ();
 b15zdnd11an1n64x5 FILLER_145_433 ();
 b15zdnd11an1n04x5 FILLER_145_497 ();
 b15zdnd00an1n02x5 FILLER_145_501 ();
 b15zdnd11an1n32x5 FILLER_145_508 ();
 b15zdnd00an1n02x5 FILLER_145_540 ();
 b15zdnd00an1n01x5 FILLER_145_542 ();
 b15zdnd11an1n04x5 FILLER_145_551 ();
 b15zdnd00an1n01x5 FILLER_145_555 ();
 b15zdnd11an1n04x5 FILLER_145_560 ();
 b15zdnd11an1n04x5 FILLER_145_572 ();
 b15zdnd11an1n04x5 FILLER_145_581 ();
 b15zdnd11an1n32x5 FILLER_145_591 ();
 b15zdnd11an1n08x5 FILLER_145_623 ();
 b15zdnd11an1n04x5 FILLER_145_631 ();
 b15zdnd00an1n01x5 FILLER_145_635 ();
 b15zdnd11an1n04x5 FILLER_145_642 ();
 b15zdnd11an1n64x5 FILLER_145_659 ();
 b15zdnd00an1n02x5 FILLER_145_723 ();
 b15zdnd00an1n01x5 FILLER_145_725 ();
 b15zdnd11an1n64x5 FILLER_145_741 ();
 b15zdnd11an1n64x5 FILLER_145_805 ();
 b15zdnd00an1n02x5 FILLER_145_869 ();
 b15zdnd00an1n01x5 FILLER_145_871 ();
 b15zdnd11an1n16x5 FILLER_145_877 ();
 b15zdnd11an1n32x5 FILLER_145_896 ();
 b15zdnd11an1n16x5 FILLER_145_928 ();
 b15zdnd00an1n02x5 FILLER_145_944 ();
 b15zdnd00an1n01x5 FILLER_145_946 ();
 b15zdnd11an1n64x5 FILLER_145_967 ();
 b15zdnd00an1n01x5 FILLER_145_1031 ();
 b15zdnd11an1n64x5 FILLER_145_1041 ();
 b15zdnd11an1n64x5 FILLER_145_1105 ();
 b15zdnd11an1n32x5 FILLER_145_1169 ();
 b15zdnd11an1n08x5 FILLER_145_1201 ();
 b15zdnd00an1n02x5 FILLER_145_1209 ();
 b15zdnd00an1n01x5 FILLER_145_1211 ();
 b15zdnd11an1n04x5 FILLER_145_1222 ();
 b15zdnd11an1n16x5 FILLER_145_1231 ();
 b15zdnd11an1n32x5 FILLER_145_1252 ();
 b15zdnd11an1n16x5 FILLER_145_1288 ();
 b15zdnd11an1n04x5 FILLER_145_1304 ();
 b15zdnd00an1n02x5 FILLER_145_1308 ();
 b15zdnd00an1n01x5 FILLER_145_1310 ();
 b15zdnd11an1n64x5 FILLER_145_1332 ();
 b15zdnd11an1n32x5 FILLER_145_1396 ();
 b15zdnd11an1n08x5 FILLER_145_1428 ();
 b15zdnd11an1n04x5 FILLER_145_1436 ();
 b15zdnd00an1n01x5 FILLER_145_1440 ();
 b15zdnd11an1n32x5 FILLER_145_1453 ();
 b15zdnd11an1n08x5 FILLER_145_1485 ();
 b15zdnd11an1n04x5 FILLER_145_1493 ();
 b15zdnd00an1n02x5 FILLER_145_1497 ();
 b15zdnd11an1n04x5 FILLER_145_1520 ();
 b15zdnd11an1n04x5 FILLER_145_1529 ();
 b15zdnd11an1n16x5 FILLER_145_1537 ();
 b15zdnd11an1n04x5 FILLER_145_1553 ();
 b15zdnd11an1n08x5 FILLER_145_1563 ();
 b15zdnd11an1n04x5 FILLER_145_1571 ();
 b15zdnd00an1n02x5 FILLER_145_1575 ();
 b15zdnd11an1n32x5 FILLER_145_1600 ();
 b15zdnd11an1n08x5 FILLER_145_1632 ();
 b15zdnd00an1n02x5 FILLER_145_1640 ();
 b15zdnd00an1n01x5 FILLER_145_1642 ();
 b15zdnd11an1n32x5 FILLER_145_1663 ();
 b15zdnd11an1n16x5 FILLER_145_1695 ();
 b15zdnd00an1n02x5 FILLER_145_1711 ();
 b15zdnd00an1n01x5 FILLER_145_1713 ();
 b15zdnd11an1n32x5 FILLER_145_1723 ();
 b15zdnd11an1n16x5 FILLER_145_1755 ();
 b15zdnd11an1n08x5 FILLER_145_1771 ();
 b15zdnd00an1n02x5 FILLER_145_1779 ();
 b15zdnd11an1n64x5 FILLER_145_1799 ();
 b15zdnd00an1n02x5 FILLER_145_1863 ();
 b15zdnd11an1n16x5 FILLER_145_1896 ();
 b15zdnd11an1n04x5 FILLER_145_1912 ();
 b15zdnd11an1n64x5 FILLER_145_1931 ();
 b15zdnd11an1n64x5 FILLER_145_1995 ();
 b15zdnd11an1n64x5 FILLER_145_2059 ();
 b15zdnd11an1n32x5 FILLER_145_2123 ();
 b15zdnd11an1n16x5 FILLER_145_2155 ();
 b15zdnd11an1n08x5 FILLER_145_2171 ();
 b15zdnd00an1n01x5 FILLER_145_2179 ();
 b15zdnd11an1n32x5 FILLER_145_2200 ();
 b15zdnd11an1n08x5 FILLER_145_2232 ();
 b15zdnd00an1n02x5 FILLER_145_2240 ();
 b15zdnd00an1n01x5 FILLER_145_2242 ();
 b15zdnd11an1n16x5 FILLER_145_2263 ();
 b15zdnd11an1n04x5 FILLER_145_2279 ();
 b15zdnd00an1n01x5 FILLER_145_2283 ();
 b15zdnd11an1n16x5 FILLER_146_8 ();
 b15zdnd11an1n08x5 FILLER_146_24 ();
 b15zdnd11an1n04x5 FILLER_146_36 ();
 b15zdnd11an1n04x5 FILLER_146_49 ();
 b15zdnd11an1n32x5 FILLER_146_60 ();
 b15zdnd11an1n32x5 FILLER_146_101 ();
 b15zdnd00an1n01x5 FILLER_146_133 ();
 b15zdnd11an1n04x5 FILLER_146_140 ();
 b15zdnd11an1n16x5 FILLER_146_150 ();
 b15zdnd11an1n08x5 FILLER_146_166 ();
 b15zdnd11an1n04x5 FILLER_146_174 ();
 b15zdnd00an1n02x5 FILLER_146_178 ();
 b15zdnd00an1n01x5 FILLER_146_180 ();
 b15zdnd11an1n32x5 FILLER_146_189 ();
 b15zdnd11an1n16x5 FILLER_146_221 ();
 b15zdnd11an1n04x5 FILLER_146_237 ();
 b15zdnd00an1n02x5 FILLER_146_241 ();
 b15zdnd00an1n01x5 FILLER_146_243 ();
 b15zdnd11an1n64x5 FILLER_146_253 ();
 b15zdnd11an1n16x5 FILLER_146_317 ();
 b15zdnd11an1n04x5 FILLER_146_333 ();
 b15zdnd00an1n01x5 FILLER_146_337 ();
 b15zdnd11an1n04x5 FILLER_146_350 ();
 b15zdnd11an1n64x5 FILLER_146_361 ();
 b15zdnd11an1n16x5 FILLER_146_425 ();
 b15zdnd11an1n04x5 FILLER_146_441 ();
 b15zdnd00an1n02x5 FILLER_146_445 ();
 b15zdnd00an1n01x5 FILLER_146_447 ();
 b15zdnd11an1n04x5 FILLER_146_461 ();
 b15zdnd00an1n01x5 FILLER_146_465 ();
 b15zdnd11an1n16x5 FILLER_146_479 ();
 b15zdnd00an1n02x5 FILLER_146_495 ();
 b15zdnd00an1n01x5 FILLER_146_497 ();
 b15zdnd11an1n32x5 FILLER_146_504 ();
 b15zdnd00an1n02x5 FILLER_146_536 ();
 b15zdnd11an1n16x5 FILLER_146_548 ();
 b15zdnd11an1n08x5 FILLER_146_564 ();
 b15zdnd11an1n04x5 FILLER_146_572 ();
 b15zdnd00an1n02x5 FILLER_146_576 ();
 b15zdnd00an1n01x5 FILLER_146_578 ();
 b15zdnd11an1n16x5 FILLER_146_605 ();
 b15zdnd11an1n08x5 FILLER_146_621 ();
 b15zdnd11an1n04x5 FILLER_146_629 ();
 b15zdnd00an1n02x5 FILLER_146_633 ();
 b15zdnd11an1n16x5 FILLER_146_661 ();
 b15zdnd00an1n01x5 FILLER_146_677 ();
 b15zdnd11an1n16x5 FILLER_146_696 ();
 b15zdnd11an1n04x5 FILLER_146_712 ();
 b15zdnd00an1n02x5 FILLER_146_716 ();
 b15zdnd11an1n16x5 FILLER_146_726 ();
 b15zdnd11an1n08x5 FILLER_146_742 ();
 b15zdnd11an1n64x5 FILLER_146_776 ();
 b15zdnd11an1n32x5 FILLER_146_840 ();
 b15zdnd00an1n02x5 FILLER_146_872 ();
 b15zdnd11an1n08x5 FILLER_146_894 ();
 b15zdnd00an1n02x5 FILLER_146_902 ();
 b15zdnd11an1n32x5 FILLER_146_924 ();
 b15zdnd11an1n16x5 FILLER_146_956 ();
 b15zdnd11an1n08x5 FILLER_146_972 ();
 b15zdnd11an1n04x5 FILLER_146_980 ();
 b15zdnd00an1n01x5 FILLER_146_984 ();
 b15zdnd11an1n16x5 FILLER_146_1004 ();
 b15zdnd11an1n08x5 FILLER_146_1020 ();
 b15zdnd00an1n02x5 FILLER_146_1028 ();
 b15zdnd00an1n01x5 FILLER_146_1030 ();
 b15zdnd11an1n16x5 FILLER_146_1041 ();
 b15zdnd11an1n08x5 FILLER_146_1057 ();
 b15zdnd00an1n02x5 FILLER_146_1065 ();
 b15zdnd11an1n64x5 FILLER_146_1106 ();
 b15zdnd11an1n32x5 FILLER_146_1170 ();
 b15zdnd11an1n16x5 FILLER_146_1202 ();
 b15zdnd11an1n08x5 FILLER_146_1218 ();
 b15zdnd11an1n04x5 FILLER_146_1226 ();
 b15zdnd00an1n02x5 FILLER_146_1230 ();
 b15zdnd11an1n16x5 FILLER_146_1236 ();
 b15zdnd00an1n01x5 FILLER_146_1252 ();
 b15zdnd11an1n16x5 FILLER_146_1269 ();
 b15zdnd00an1n01x5 FILLER_146_1285 ();
 b15zdnd11an1n16x5 FILLER_146_1295 ();
 b15zdnd11an1n04x5 FILLER_146_1311 ();
 b15zdnd00an1n02x5 FILLER_146_1315 ();
 b15zdnd11an1n08x5 FILLER_146_1329 ();
 b15zdnd00an1n01x5 FILLER_146_1337 ();
 b15zdnd11an1n16x5 FILLER_146_1348 ();
 b15zdnd11an1n04x5 FILLER_146_1364 ();
 b15zdnd00an1n02x5 FILLER_146_1368 ();
 b15zdnd00an1n01x5 FILLER_146_1370 ();
 b15zdnd11an1n04x5 FILLER_146_1375 ();
 b15zdnd11an1n04x5 FILLER_146_1385 ();
 b15zdnd11an1n32x5 FILLER_146_1405 ();
 b15zdnd11an1n16x5 FILLER_146_1437 ();
 b15zdnd11an1n16x5 FILLER_146_1458 ();
 b15zdnd11an1n08x5 FILLER_146_1474 ();
 b15zdnd11an1n08x5 FILLER_146_1508 ();
 b15zdnd11an1n04x5 FILLER_146_1516 ();
 b15zdnd00an1n02x5 FILLER_146_1520 ();
 b15zdnd00an1n01x5 FILLER_146_1522 ();
 b15zdnd11an1n16x5 FILLER_146_1529 ();
 b15zdnd11an1n04x5 FILLER_146_1545 ();
 b15zdnd00an1n02x5 FILLER_146_1549 ();
 b15zdnd11an1n64x5 FILLER_146_1569 ();
 b15zdnd11an1n64x5 FILLER_146_1633 ();
 b15zdnd11an1n64x5 FILLER_146_1697 ();
 b15zdnd11an1n32x5 FILLER_146_1761 ();
 b15zdnd11an1n16x5 FILLER_146_1793 ();
 b15zdnd11an1n64x5 FILLER_146_1834 ();
 b15zdnd11an1n32x5 FILLER_146_1898 ();
 b15zdnd11an1n16x5 FILLER_146_1930 ();
 b15zdnd11an1n08x5 FILLER_146_1946 ();
 b15zdnd11an1n04x5 FILLER_146_1954 ();
 b15zdnd11an1n64x5 FILLER_146_1970 ();
 b15zdnd11an1n32x5 FILLER_146_2034 ();
 b15zdnd00an1n02x5 FILLER_146_2066 ();
 b15zdnd00an1n01x5 FILLER_146_2068 ();
 b15zdnd11an1n32x5 FILLER_146_2080 ();
 b15zdnd11an1n08x5 FILLER_146_2112 ();
 b15zdnd00an1n02x5 FILLER_146_2120 ();
 b15zdnd11an1n16x5 FILLER_146_2126 ();
 b15zdnd11an1n08x5 FILLER_146_2142 ();
 b15zdnd11an1n04x5 FILLER_146_2150 ();
 b15zdnd11an1n16x5 FILLER_146_2162 ();
 b15zdnd00an1n02x5 FILLER_146_2178 ();
 b15zdnd11an1n08x5 FILLER_146_2185 ();
 b15zdnd00an1n02x5 FILLER_146_2193 ();
 b15zdnd11an1n16x5 FILLER_146_2215 ();
 b15zdnd11an1n08x5 FILLER_146_2231 ();
 b15zdnd11an1n04x5 FILLER_146_2239 ();
 b15zdnd11an1n04x5 FILLER_146_2249 ();
 b15zdnd11an1n16x5 FILLER_146_2258 ();
 b15zdnd00an1n02x5 FILLER_146_2274 ();
 b15zdnd11an1n32x5 FILLER_147_0 ();
 b15zdnd11an1n08x5 FILLER_147_32 ();
 b15zdnd00an1n01x5 FILLER_147_40 ();
 b15zdnd11an1n32x5 FILLER_147_55 ();
 b15zdnd11an1n08x5 FILLER_147_87 ();
 b15zdnd11an1n04x5 FILLER_147_95 ();
 b15zdnd00an1n01x5 FILLER_147_99 ();
 b15zdnd11an1n64x5 FILLER_147_109 ();
 b15zdnd11an1n16x5 FILLER_147_173 ();
 b15zdnd11an1n32x5 FILLER_147_203 ();
 b15zdnd11an1n16x5 FILLER_147_235 ();
 b15zdnd11an1n08x5 FILLER_147_251 ();
 b15zdnd11an1n04x5 FILLER_147_259 ();
 b15zdnd00an1n02x5 FILLER_147_263 ();
 b15zdnd11an1n04x5 FILLER_147_272 ();
 b15zdnd11an1n08x5 FILLER_147_286 ();
 b15zdnd11an1n04x5 FILLER_147_294 ();
 b15zdnd11an1n08x5 FILLER_147_314 ();
 b15zdnd11an1n04x5 FILLER_147_322 ();
 b15zdnd11an1n04x5 FILLER_147_344 ();
 b15zdnd00an1n01x5 FILLER_147_348 ();
 b15zdnd11an1n64x5 FILLER_147_355 ();
 b15zdnd00an1n01x5 FILLER_147_419 ();
 b15zdnd11an1n04x5 FILLER_147_436 ();
 b15zdnd11an1n04x5 FILLER_147_458 ();
 b15zdnd11an1n04x5 FILLER_147_468 ();
 b15zdnd11an1n08x5 FILLER_147_486 ();
 b15zdnd11an1n04x5 FILLER_147_494 ();
 b15zdnd00an1n02x5 FILLER_147_498 ();
 b15zdnd11an1n64x5 FILLER_147_510 ();
 b15zdnd11an1n08x5 FILLER_147_574 ();
 b15zdnd00an1n02x5 FILLER_147_582 ();
 b15zdnd11an1n08x5 FILLER_147_598 ();
 b15zdnd00an1n02x5 FILLER_147_606 ();
 b15zdnd11an1n04x5 FILLER_147_620 ();
 b15zdnd11an1n04x5 FILLER_147_629 ();
 b15zdnd11an1n16x5 FILLER_147_644 ();
 b15zdnd11an1n08x5 FILLER_147_669 ();
 b15zdnd00an1n02x5 FILLER_147_677 ();
 b15zdnd00an1n01x5 FILLER_147_679 ();
 b15zdnd11an1n16x5 FILLER_147_706 ();
 b15zdnd11an1n04x5 FILLER_147_722 ();
 b15zdnd00an1n02x5 FILLER_147_726 ();
 b15zdnd00an1n01x5 FILLER_147_728 ();
 b15zdnd11an1n04x5 FILLER_147_741 ();
 b15zdnd11an1n32x5 FILLER_147_771 ();
 b15zdnd11an1n64x5 FILLER_147_814 ();
 b15zdnd11an1n16x5 FILLER_147_878 ();
 b15zdnd11an1n08x5 FILLER_147_894 ();
 b15zdnd00an1n01x5 FILLER_147_902 ();
 b15zdnd11an1n16x5 FILLER_147_908 ();
 b15zdnd11an1n16x5 FILLER_147_927 ();
 b15zdnd11an1n08x5 FILLER_147_943 ();
 b15zdnd11an1n04x5 FILLER_147_951 ();
 b15zdnd00an1n02x5 FILLER_147_955 ();
 b15zdnd00an1n01x5 FILLER_147_957 ();
 b15zdnd11an1n08x5 FILLER_147_989 ();
 b15zdnd00an1n02x5 FILLER_147_997 ();
 b15zdnd11an1n64x5 FILLER_147_1030 ();
 b15zdnd11an1n64x5 FILLER_147_1094 ();
 b15zdnd11an1n64x5 FILLER_147_1158 ();
 b15zdnd11an1n64x5 FILLER_147_1222 ();
 b15zdnd11an1n32x5 FILLER_147_1286 ();
 b15zdnd00an1n01x5 FILLER_147_1318 ();
 b15zdnd11an1n64x5 FILLER_147_1343 ();
 b15zdnd11an1n16x5 FILLER_147_1407 ();
 b15zdnd11an1n08x5 FILLER_147_1423 ();
 b15zdnd11an1n04x5 FILLER_147_1431 ();
 b15zdnd00an1n01x5 FILLER_147_1435 ();
 b15zdnd11an1n08x5 FILLER_147_1442 ();
 b15zdnd00an1n01x5 FILLER_147_1450 ();
 b15zdnd11an1n08x5 FILLER_147_1455 ();
 b15zdnd00an1n01x5 FILLER_147_1463 ();
 b15zdnd11an1n32x5 FILLER_147_1468 ();
 b15zdnd11an1n04x5 FILLER_147_1500 ();
 b15zdnd00an1n02x5 FILLER_147_1504 ();
 b15zdnd11an1n16x5 FILLER_147_1511 ();
 b15zdnd11an1n08x5 FILLER_147_1527 ();
 b15zdnd11an1n04x5 FILLER_147_1535 ();
 b15zdnd00an1n02x5 FILLER_147_1539 ();
 b15zdnd00an1n01x5 FILLER_147_1541 ();
 b15zdnd11an1n04x5 FILLER_147_1547 ();
 b15zdnd11an1n32x5 FILLER_147_1567 ();
 b15zdnd11an1n08x5 FILLER_147_1599 ();
 b15zdnd11an1n04x5 FILLER_147_1607 ();
 b15zdnd00an1n01x5 FILLER_147_1611 ();
 b15zdnd11an1n64x5 FILLER_147_1630 ();
 b15zdnd11an1n64x5 FILLER_147_1694 ();
 b15zdnd11an1n16x5 FILLER_147_1758 ();
 b15zdnd11an1n08x5 FILLER_147_1774 ();
 b15zdnd11an1n04x5 FILLER_147_1782 ();
 b15zdnd11an1n64x5 FILLER_147_1827 ();
 b15zdnd11an1n16x5 FILLER_147_1891 ();
 b15zdnd11an1n08x5 FILLER_147_1907 ();
 b15zdnd11an1n04x5 FILLER_147_1915 ();
 b15zdnd00an1n01x5 FILLER_147_1919 ();
 b15zdnd11an1n64x5 FILLER_147_1935 ();
 b15zdnd00an1n02x5 FILLER_147_1999 ();
 b15zdnd11an1n08x5 FILLER_147_2010 ();
 b15zdnd00an1n02x5 FILLER_147_2018 ();
 b15zdnd00an1n01x5 FILLER_147_2020 ();
 b15zdnd11an1n16x5 FILLER_147_2032 ();
 b15zdnd11an1n04x5 FILLER_147_2048 ();
 b15zdnd00an1n02x5 FILLER_147_2052 ();
 b15zdnd00an1n01x5 FILLER_147_2054 ();
 b15zdnd11an1n16x5 FILLER_147_2075 ();
 b15zdnd00an1n02x5 FILLER_147_2091 ();
 b15zdnd11an1n16x5 FILLER_147_2113 ();
 b15zdnd11an1n04x5 FILLER_147_2129 ();
 b15zdnd00an1n01x5 FILLER_147_2133 ();
 b15zdnd11an1n16x5 FILLER_147_2154 ();
 b15zdnd11an1n08x5 FILLER_147_2170 ();
 b15zdnd00an1n01x5 FILLER_147_2178 ();
 b15zdnd11an1n16x5 FILLER_147_2185 ();
 b15zdnd11an1n32x5 FILLER_147_2210 ();
 b15zdnd11an1n16x5 FILLER_147_2242 ();
 b15zdnd11an1n08x5 FILLER_147_2258 ();
 b15zdnd00an1n02x5 FILLER_147_2266 ();
 b15zdnd00an1n01x5 FILLER_147_2268 ();
 b15zdnd11an1n04x5 FILLER_147_2273 ();
 b15zdnd00an1n01x5 FILLER_147_2277 ();
 b15zdnd00an1n02x5 FILLER_147_2282 ();
 b15zdnd11an1n32x5 FILLER_148_8 ();
 b15zdnd11an1n64x5 FILLER_148_58 ();
 b15zdnd11an1n08x5 FILLER_148_122 ();
 b15zdnd11an1n04x5 FILLER_148_130 ();
 b15zdnd00an1n02x5 FILLER_148_134 ();
 b15zdnd11an1n08x5 FILLER_148_144 ();
 b15zdnd00an1n02x5 FILLER_148_152 ();
 b15zdnd00an1n01x5 FILLER_148_154 ();
 b15zdnd11an1n32x5 FILLER_148_159 ();
 b15zdnd11an1n16x5 FILLER_148_191 ();
 b15zdnd11an1n04x5 FILLER_148_207 ();
 b15zdnd11an1n08x5 FILLER_148_219 ();
 b15zdnd11an1n04x5 FILLER_148_227 ();
 b15zdnd00an1n02x5 FILLER_148_231 ();
 b15zdnd00an1n01x5 FILLER_148_233 ();
 b15zdnd11an1n16x5 FILLER_148_244 ();
 b15zdnd11an1n04x5 FILLER_148_260 ();
 b15zdnd00an1n01x5 FILLER_148_264 ();
 b15zdnd11an1n64x5 FILLER_148_274 ();
 b15zdnd11an1n64x5 FILLER_148_338 ();
 b15zdnd11an1n64x5 FILLER_148_402 ();
 b15zdnd11an1n32x5 FILLER_148_466 ();
 b15zdnd00an1n01x5 FILLER_148_498 ();
 b15zdnd11an1n16x5 FILLER_148_521 ();
 b15zdnd11an1n08x5 FILLER_148_537 ();
 b15zdnd11an1n04x5 FILLER_148_545 ();
 b15zdnd00an1n02x5 FILLER_148_549 ();
 b15zdnd11an1n64x5 FILLER_148_561 ();
 b15zdnd11an1n04x5 FILLER_148_625 ();
 b15zdnd00an1n02x5 FILLER_148_629 ();
 b15zdnd00an1n01x5 FILLER_148_631 ();
 b15zdnd11an1n16x5 FILLER_148_642 ();
 b15zdnd11an1n04x5 FILLER_148_658 ();
 b15zdnd00an1n02x5 FILLER_148_662 ();
 b15zdnd00an1n01x5 FILLER_148_664 ();
 b15zdnd11an1n08x5 FILLER_148_670 ();
 b15zdnd11an1n04x5 FILLER_148_678 ();
 b15zdnd00an1n01x5 FILLER_148_682 ();
 b15zdnd11an1n08x5 FILLER_148_695 ();
 b15zdnd11an1n04x5 FILLER_148_703 ();
 b15zdnd00an1n02x5 FILLER_148_707 ();
 b15zdnd00an1n02x5 FILLER_148_716 ();
 b15zdnd11an1n64x5 FILLER_148_726 ();
 b15zdnd11an1n16x5 FILLER_148_790 ();
 b15zdnd11an1n16x5 FILLER_148_826 ();
 b15zdnd11an1n08x5 FILLER_148_842 ();
 b15zdnd00an1n02x5 FILLER_148_850 ();
 b15zdnd11an1n04x5 FILLER_148_857 ();
 b15zdnd11an1n64x5 FILLER_148_865 ();
 b15zdnd11an1n64x5 FILLER_148_929 ();
 b15zdnd11an1n64x5 FILLER_148_993 ();
 b15zdnd11an1n16x5 FILLER_148_1057 ();
 b15zdnd11an1n04x5 FILLER_148_1073 ();
 b15zdnd00an1n02x5 FILLER_148_1077 ();
 b15zdnd11an1n64x5 FILLER_148_1089 ();
 b15zdnd11an1n04x5 FILLER_148_1153 ();
 b15zdnd00an1n02x5 FILLER_148_1157 ();
 b15zdnd11an1n04x5 FILLER_148_1184 ();
 b15zdnd11an1n64x5 FILLER_148_1203 ();
 b15zdnd11an1n32x5 FILLER_148_1267 ();
 b15zdnd11an1n08x5 FILLER_148_1299 ();
 b15zdnd11an1n08x5 FILLER_148_1315 ();
 b15zdnd11an1n04x5 FILLER_148_1323 ();
 b15zdnd00an1n02x5 FILLER_148_1327 ();
 b15zdnd11an1n32x5 FILLER_148_1342 ();
 b15zdnd11an1n16x5 FILLER_148_1374 ();
 b15zdnd11an1n08x5 FILLER_148_1390 ();
 b15zdnd11an1n04x5 FILLER_148_1398 ();
 b15zdnd11an1n04x5 FILLER_148_1408 ();
 b15zdnd11an1n04x5 FILLER_148_1424 ();
 b15zdnd11an1n08x5 FILLER_148_1438 ();
 b15zdnd11an1n04x5 FILLER_148_1446 ();
 b15zdnd00an1n02x5 FILLER_148_1450 ();
 b15zdnd11an1n04x5 FILLER_148_1459 ();
 b15zdnd11an1n16x5 FILLER_148_1470 ();
 b15zdnd11an1n08x5 FILLER_148_1486 ();
 b15zdnd00an1n01x5 FILLER_148_1494 ();
 b15zdnd11an1n08x5 FILLER_148_1507 ();
 b15zdnd11an1n04x5 FILLER_148_1515 ();
 b15zdnd00an1n02x5 FILLER_148_1519 ();
 b15zdnd00an1n01x5 FILLER_148_1521 ();
 b15zdnd11an1n16x5 FILLER_148_1532 ();
 b15zdnd11an1n04x5 FILLER_148_1568 ();
 b15zdnd11an1n64x5 FILLER_148_1588 ();
 b15zdnd11an1n32x5 FILLER_148_1652 ();
 b15zdnd11an1n08x5 FILLER_148_1684 ();
 b15zdnd11an1n04x5 FILLER_148_1692 ();
 b15zdnd00an1n02x5 FILLER_148_1696 ();
 b15zdnd00an1n01x5 FILLER_148_1698 ();
 b15zdnd11an1n64x5 FILLER_148_1730 ();
 b15zdnd11an1n64x5 FILLER_148_1794 ();
 b15zdnd11an1n16x5 FILLER_148_1858 ();
 b15zdnd11an1n08x5 FILLER_148_1889 ();
 b15zdnd11an1n08x5 FILLER_148_1936 ();
 b15zdnd11an1n16x5 FILLER_148_1965 ();
 b15zdnd00an1n02x5 FILLER_148_1981 ();
 b15zdnd11an1n64x5 FILLER_148_2014 ();
 b15zdnd11an1n64x5 FILLER_148_2078 ();
 b15zdnd11an1n08x5 FILLER_148_2142 ();
 b15zdnd11an1n04x5 FILLER_148_2150 ();
 b15zdnd11an1n64x5 FILLER_148_2162 ();
 b15zdnd11an1n16x5 FILLER_148_2226 ();
 b15zdnd11an1n04x5 FILLER_148_2242 ();
 b15zdnd11an1n04x5 FILLER_148_2258 ();
 b15zdnd11an1n04x5 FILLER_148_2266 ();
 b15zdnd00an1n02x5 FILLER_148_2274 ();
 b15zdnd11an1n64x5 FILLER_149_0 ();
 b15zdnd11an1n32x5 FILLER_149_68 ();
 b15zdnd11an1n04x5 FILLER_149_100 ();
 b15zdnd11an1n16x5 FILLER_149_117 ();
 b15zdnd11an1n08x5 FILLER_149_133 ();
 b15zdnd11an1n04x5 FILLER_149_141 ();
 b15zdnd00an1n01x5 FILLER_149_145 ();
 b15zdnd11an1n04x5 FILLER_149_152 ();
 b15zdnd11an1n32x5 FILLER_149_186 ();
 b15zdnd11an1n08x5 FILLER_149_218 ();
 b15zdnd11an1n04x5 FILLER_149_226 ();
 b15zdnd11an1n04x5 FILLER_149_234 ();
 b15zdnd11an1n08x5 FILLER_149_258 ();
 b15zdnd00an1n01x5 FILLER_149_266 ();
 b15zdnd11an1n32x5 FILLER_149_271 ();
 b15zdnd00an1n02x5 FILLER_149_303 ();
 b15zdnd00an1n01x5 FILLER_149_305 ();
 b15zdnd11an1n64x5 FILLER_149_315 ();
 b15zdnd11an1n32x5 FILLER_149_379 ();
 b15zdnd11an1n08x5 FILLER_149_411 ();
 b15zdnd11an1n04x5 FILLER_149_419 ();
 b15zdnd00an1n02x5 FILLER_149_423 ();
 b15zdnd11an1n04x5 FILLER_149_448 ();
 b15zdnd11an1n64x5 FILLER_149_483 ();
 b15zdnd11an1n32x5 FILLER_149_547 ();
 b15zdnd11an1n16x5 FILLER_149_579 ();
 b15zdnd11an1n08x5 FILLER_149_595 ();
 b15zdnd11an1n16x5 FILLER_149_607 ();
 b15zdnd11an1n16x5 FILLER_149_628 ();
 b15zdnd11an1n08x5 FILLER_149_644 ();
 b15zdnd11an1n04x5 FILLER_149_652 ();
 b15zdnd00an1n02x5 FILLER_149_656 ();
 b15zdnd00an1n01x5 FILLER_149_658 ();
 b15zdnd11an1n32x5 FILLER_149_664 ();
 b15zdnd11an1n08x5 FILLER_149_696 ();
 b15zdnd11an1n04x5 FILLER_149_704 ();
 b15zdnd00an1n02x5 FILLER_149_708 ();
 b15zdnd00an1n01x5 FILLER_149_710 ();
 b15zdnd11an1n04x5 FILLER_149_716 ();
 b15zdnd11an1n16x5 FILLER_149_740 ();
 b15zdnd11an1n16x5 FILLER_149_782 ();
 b15zdnd00an1n02x5 FILLER_149_798 ();
 b15zdnd00an1n01x5 FILLER_149_800 ();
 b15zdnd11an1n16x5 FILLER_149_812 ();
 b15zdnd11an1n08x5 FILLER_149_828 ();
 b15zdnd00an1n01x5 FILLER_149_836 ();
 b15zdnd11an1n64x5 FILLER_149_857 ();
 b15zdnd11an1n32x5 FILLER_149_921 ();
 b15zdnd11an1n08x5 FILLER_149_953 ();
 b15zdnd11an1n16x5 FILLER_149_981 ();
 b15zdnd11an1n08x5 FILLER_149_997 ();
 b15zdnd00an1n02x5 FILLER_149_1005 ();
 b15zdnd00an1n01x5 FILLER_149_1007 ();
 b15zdnd11an1n04x5 FILLER_149_1012 ();
 b15zdnd00an1n02x5 FILLER_149_1016 ();
 b15zdnd00an1n01x5 FILLER_149_1018 ();
 b15zdnd11an1n32x5 FILLER_149_1024 ();
 b15zdnd11an1n16x5 FILLER_149_1056 ();
 b15zdnd00an1n01x5 FILLER_149_1072 ();
 b15zdnd11an1n32x5 FILLER_149_1082 ();
 b15zdnd11an1n16x5 FILLER_149_1114 ();
 b15zdnd11an1n08x5 FILLER_149_1130 ();
 b15zdnd11an1n04x5 FILLER_149_1138 ();
 b15zdnd11an1n32x5 FILLER_149_1153 ();
 b15zdnd11an1n04x5 FILLER_149_1185 ();
 b15zdnd11an1n08x5 FILLER_149_1201 ();
 b15zdnd11an1n64x5 FILLER_149_1227 ();
 b15zdnd11an1n04x5 FILLER_149_1291 ();
 b15zdnd00an1n01x5 FILLER_149_1295 ();
 b15zdnd11an1n04x5 FILLER_149_1304 ();
 b15zdnd11an1n04x5 FILLER_149_1320 ();
 b15zdnd00an1n02x5 FILLER_149_1324 ();
 b15zdnd11an1n16x5 FILLER_149_1331 ();
 b15zdnd11an1n08x5 FILLER_149_1347 ();
 b15zdnd11an1n04x5 FILLER_149_1355 ();
 b15zdnd00an1n01x5 FILLER_149_1359 ();
 b15zdnd11an1n16x5 FILLER_149_1366 ();
 b15zdnd11an1n08x5 FILLER_149_1382 ();
 b15zdnd00an1n01x5 FILLER_149_1390 ();
 b15zdnd11an1n32x5 FILLER_149_1398 ();
 b15zdnd11an1n16x5 FILLER_149_1430 ();
 b15zdnd11an1n08x5 FILLER_149_1446 ();
 b15zdnd00an1n02x5 FILLER_149_1454 ();
 b15zdnd11an1n04x5 FILLER_149_1463 ();
 b15zdnd11an1n32x5 FILLER_149_1472 ();
 b15zdnd00an1n02x5 FILLER_149_1504 ();
 b15zdnd11an1n16x5 FILLER_149_1513 ();
 b15zdnd00an1n02x5 FILLER_149_1529 ();
 b15zdnd11an1n64x5 FILLER_149_1557 ();
 b15zdnd00an1n02x5 FILLER_149_1621 ();
 b15zdnd11an1n32x5 FILLER_149_1649 ();
 b15zdnd11an1n16x5 FILLER_149_1681 ();
 b15zdnd00an1n02x5 FILLER_149_1697 ();
 b15zdnd11an1n64x5 FILLER_149_1719 ();
 b15zdnd11an1n32x5 FILLER_149_1783 ();
 b15zdnd11an1n16x5 FILLER_149_1815 ();
 b15zdnd11an1n04x5 FILLER_149_1831 ();
 b15zdnd00an1n01x5 FILLER_149_1835 ();
 b15zdnd11an1n32x5 FILLER_149_1845 ();
 b15zdnd11an1n16x5 FILLER_149_1877 ();
 b15zdnd00an1n02x5 FILLER_149_1893 ();
 b15zdnd00an1n01x5 FILLER_149_1895 ();
 b15zdnd11an1n16x5 FILLER_149_1921 ();
 b15zdnd11an1n08x5 FILLER_149_1937 ();
 b15zdnd11an1n64x5 FILLER_149_1955 ();
 b15zdnd11an1n16x5 FILLER_149_2019 ();
 b15zdnd00an1n01x5 FILLER_149_2035 ();
 b15zdnd11an1n32x5 FILLER_149_2068 ();
 b15zdnd00an1n01x5 FILLER_149_2100 ();
 b15zdnd11an1n64x5 FILLER_149_2112 ();
 b15zdnd11an1n64x5 FILLER_149_2176 ();
 b15zdnd11an1n08x5 FILLER_149_2240 ();
 b15zdnd00an1n01x5 FILLER_149_2248 ();
 b15zdnd11an1n08x5 FILLER_149_2253 ();
 b15zdnd11an1n04x5 FILLER_149_2261 ();
 b15zdnd00an1n01x5 FILLER_149_2265 ();
 b15zdnd11an1n04x5 FILLER_149_2270 ();
 b15zdnd00an1n02x5 FILLER_149_2274 ();
 b15zdnd00an1n01x5 FILLER_149_2276 ();
 b15zdnd00an1n02x5 FILLER_149_2282 ();
 b15zdnd11an1n32x5 FILLER_150_8 ();
 b15zdnd11an1n16x5 FILLER_150_40 ();
 b15zdnd11an1n08x5 FILLER_150_56 ();
 b15zdnd11an1n16x5 FILLER_150_76 ();
 b15zdnd11an1n04x5 FILLER_150_100 ();
 b15zdnd00an1n01x5 FILLER_150_104 ();
 b15zdnd11an1n32x5 FILLER_150_112 ();
 b15zdnd11an1n08x5 FILLER_150_144 ();
 b15zdnd00an1n01x5 FILLER_150_152 ();
 b15zdnd11an1n04x5 FILLER_150_169 ();
 b15zdnd11an1n32x5 FILLER_150_179 ();
 b15zdnd11an1n08x5 FILLER_150_211 ();
 b15zdnd00an1n02x5 FILLER_150_219 ();
 b15zdnd11an1n32x5 FILLER_150_227 ();
 b15zdnd11an1n08x5 FILLER_150_259 ();
 b15zdnd11an1n32x5 FILLER_150_274 ();
 b15zdnd11an1n04x5 FILLER_150_306 ();
 b15zdnd00an1n02x5 FILLER_150_310 ();
 b15zdnd11an1n64x5 FILLER_150_321 ();
 b15zdnd11an1n32x5 FILLER_150_385 ();
 b15zdnd11an1n16x5 FILLER_150_417 ();
 b15zdnd11an1n32x5 FILLER_150_445 ();
 b15zdnd11an1n16x5 FILLER_150_477 ();
 b15zdnd00an1n02x5 FILLER_150_493 ();
 b15zdnd00an1n01x5 FILLER_150_495 ();
 b15zdnd11an1n04x5 FILLER_150_501 ();
 b15zdnd11an1n04x5 FILLER_150_513 ();
 b15zdnd11an1n16x5 FILLER_150_523 ();
 b15zdnd11an1n08x5 FILLER_150_539 ();
 b15zdnd11an1n04x5 FILLER_150_547 ();
 b15zdnd00an1n02x5 FILLER_150_551 ();
 b15zdnd00an1n01x5 FILLER_150_553 ();
 b15zdnd11an1n08x5 FILLER_150_566 ();
 b15zdnd11an1n04x5 FILLER_150_574 ();
 b15zdnd00an1n01x5 FILLER_150_578 ();
 b15zdnd11an1n04x5 FILLER_150_591 ();
 b15zdnd00an1n02x5 FILLER_150_595 ();
 b15zdnd11an1n64x5 FILLER_150_609 ();
 b15zdnd11an1n08x5 FILLER_150_673 ();
 b15zdnd11an1n04x5 FILLER_150_681 ();
 b15zdnd00an1n02x5 FILLER_150_685 ();
 b15zdnd00an1n01x5 FILLER_150_687 ();
 b15zdnd11an1n16x5 FILLER_150_700 ();
 b15zdnd00an1n02x5 FILLER_150_716 ();
 b15zdnd11an1n16x5 FILLER_150_726 ();
 b15zdnd00an1n02x5 FILLER_150_742 ();
 b15zdnd00an1n01x5 FILLER_150_744 ();
 b15zdnd11an1n64x5 FILLER_150_771 ();
 b15zdnd11an1n64x5 FILLER_150_841 ();
 b15zdnd11an1n16x5 FILLER_150_905 ();
 b15zdnd11an1n04x5 FILLER_150_921 ();
 b15zdnd00an1n02x5 FILLER_150_925 ();
 b15zdnd00an1n01x5 FILLER_150_927 ();
 b15zdnd11an1n08x5 FILLER_150_950 ();
 b15zdnd00an1n01x5 FILLER_150_958 ();
 b15zdnd11an1n04x5 FILLER_150_965 ();
 b15zdnd11an1n64x5 FILLER_150_974 ();
 b15zdnd11an1n16x5 FILLER_150_1038 ();
 b15zdnd11an1n08x5 FILLER_150_1054 ();
 b15zdnd11an1n04x5 FILLER_150_1072 ();
 b15zdnd11an1n04x5 FILLER_150_1085 ();
 b15zdnd00an1n01x5 FILLER_150_1089 ();
 b15zdnd11an1n04x5 FILLER_150_1101 ();
 b15zdnd11an1n04x5 FILLER_150_1125 ();
 b15zdnd00an1n01x5 FILLER_150_1129 ();
 b15zdnd11an1n32x5 FILLER_150_1161 ();
 b15zdnd11an1n16x5 FILLER_150_1193 ();
 b15zdnd11an1n08x5 FILLER_150_1209 ();
 b15zdnd11an1n04x5 FILLER_150_1217 ();
 b15zdnd00an1n02x5 FILLER_150_1221 ();
 b15zdnd00an1n01x5 FILLER_150_1223 ();
 b15zdnd11an1n04x5 FILLER_150_1236 ();
 b15zdnd11an1n64x5 FILLER_150_1250 ();
 b15zdnd11an1n32x5 FILLER_150_1314 ();
 b15zdnd11an1n16x5 FILLER_150_1346 ();
 b15zdnd11an1n04x5 FILLER_150_1362 ();
 b15zdnd00an1n02x5 FILLER_150_1366 ();
 b15zdnd00an1n01x5 FILLER_150_1368 ();
 b15zdnd11an1n08x5 FILLER_150_1373 ();
 b15zdnd00an1n02x5 FILLER_150_1381 ();
 b15zdnd00an1n01x5 FILLER_150_1383 ();
 b15zdnd11an1n64x5 FILLER_150_1400 ();
 b15zdnd11an1n32x5 FILLER_150_1464 ();
 b15zdnd11an1n16x5 FILLER_150_1496 ();
 b15zdnd11an1n04x5 FILLER_150_1512 ();
 b15zdnd00an1n02x5 FILLER_150_1516 ();
 b15zdnd11an1n16x5 FILLER_150_1528 ();
 b15zdnd11an1n04x5 FILLER_150_1544 ();
 b15zdnd00an1n02x5 FILLER_150_1548 ();
 b15zdnd00an1n01x5 FILLER_150_1550 ();
 b15zdnd11an1n32x5 FILLER_150_1557 ();
 b15zdnd11an1n16x5 FILLER_150_1589 ();
 b15zdnd11an1n08x5 FILLER_150_1605 ();
 b15zdnd11an1n04x5 FILLER_150_1613 ();
 b15zdnd00an1n01x5 FILLER_150_1617 ();
 b15zdnd11an1n04x5 FILLER_150_1644 ();
 b15zdnd11an1n32x5 FILLER_150_1668 ();
 b15zdnd00an1n02x5 FILLER_150_1700 ();
 b15zdnd11an1n16x5 FILLER_150_1707 ();
 b15zdnd00an1n02x5 FILLER_150_1723 ();
 b15zdnd00an1n01x5 FILLER_150_1725 ();
 b15zdnd11an1n04x5 FILLER_150_1737 ();
 b15zdnd11an1n32x5 FILLER_150_1761 ();
 b15zdnd11an1n08x5 FILLER_150_1793 ();
 b15zdnd11an1n04x5 FILLER_150_1801 ();
 b15zdnd11an1n16x5 FILLER_150_1836 ();
 b15zdnd11an1n08x5 FILLER_150_1852 ();
 b15zdnd00an1n02x5 FILLER_150_1860 ();
 b15zdnd00an1n01x5 FILLER_150_1862 ();
 b15zdnd11an1n64x5 FILLER_150_1902 ();
 b15zdnd11an1n08x5 FILLER_150_1966 ();
 b15zdnd11an1n64x5 FILLER_150_2005 ();
 b15zdnd11an1n64x5 FILLER_150_2069 ();
 b15zdnd11an1n04x5 FILLER_150_2133 ();
 b15zdnd00an1n02x5 FILLER_150_2137 ();
 b15zdnd00an1n01x5 FILLER_150_2139 ();
 b15zdnd11an1n08x5 FILLER_150_2145 ();
 b15zdnd00an1n01x5 FILLER_150_2153 ();
 b15zdnd11an1n32x5 FILLER_150_2162 ();
 b15zdnd11an1n08x5 FILLER_150_2194 ();
 b15zdnd00an1n01x5 FILLER_150_2202 ();
 b15zdnd11an1n16x5 FILLER_150_2223 ();
 b15zdnd00an1n02x5 FILLER_150_2239 ();
 b15zdnd00an1n01x5 FILLER_150_2241 ();
 b15zdnd11an1n04x5 FILLER_150_2253 ();
 b15zdnd00an1n02x5 FILLER_150_2257 ();
 b15zdnd00an1n01x5 FILLER_150_2259 ();
 b15zdnd11an1n04x5 FILLER_150_2265 ();
 b15zdnd00an1n02x5 FILLER_150_2273 ();
 b15zdnd00an1n01x5 FILLER_150_2275 ();
 b15zdnd11an1n64x5 FILLER_151_0 ();
 b15zdnd11an1n04x5 FILLER_151_77 ();
 b15zdnd11an1n16x5 FILLER_151_85 ();
 b15zdnd11an1n32x5 FILLER_151_107 ();
 b15zdnd11an1n16x5 FILLER_151_139 ();
 b15zdnd11an1n08x5 FILLER_151_155 ();
 b15zdnd11an1n04x5 FILLER_151_172 ();
 b15zdnd11an1n64x5 FILLER_151_181 ();
 b15zdnd11an1n32x5 FILLER_151_245 ();
 b15zdnd11an1n08x5 FILLER_151_277 ();
 b15zdnd11an1n04x5 FILLER_151_285 ();
 b15zdnd00an1n02x5 FILLER_151_289 ();
 b15zdnd00an1n01x5 FILLER_151_291 ();
 b15zdnd11an1n04x5 FILLER_151_296 ();
 b15zdnd11an1n32x5 FILLER_151_312 ();
 b15zdnd11an1n08x5 FILLER_151_344 ();
 b15zdnd00an1n02x5 FILLER_151_352 ();
 b15zdnd11an1n04x5 FILLER_151_358 ();
 b15zdnd11an1n64x5 FILLER_151_366 ();
 b15zdnd11an1n64x5 FILLER_151_430 ();
 b15zdnd11an1n16x5 FILLER_151_505 ();
 b15zdnd11an1n08x5 FILLER_151_521 ();
 b15zdnd00an1n02x5 FILLER_151_529 ();
 b15zdnd00an1n01x5 FILLER_151_531 ();
 b15zdnd11an1n16x5 FILLER_151_548 ();
 b15zdnd11an1n04x5 FILLER_151_564 ();
 b15zdnd00an1n01x5 FILLER_151_568 ();
 b15zdnd11an1n04x5 FILLER_151_579 ();
 b15zdnd11an1n16x5 FILLER_151_588 ();
 b15zdnd11an1n08x5 FILLER_151_604 ();
 b15zdnd11an1n04x5 FILLER_151_612 ();
 b15zdnd11an1n32x5 FILLER_151_626 ();
 b15zdnd11an1n04x5 FILLER_151_658 ();
 b15zdnd00an1n01x5 FILLER_151_662 ();
 b15zdnd11an1n08x5 FILLER_151_669 ();
 b15zdnd11an1n04x5 FILLER_151_677 ();
 b15zdnd00an1n02x5 FILLER_151_681 ();
 b15zdnd00an1n01x5 FILLER_151_683 ();
 b15zdnd11an1n32x5 FILLER_151_689 ();
 b15zdnd11an1n16x5 FILLER_151_721 ();
 b15zdnd11an1n08x5 FILLER_151_737 ();
 b15zdnd00an1n01x5 FILLER_151_745 ();
 b15zdnd11an1n04x5 FILLER_151_777 ();
 b15zdnd00an1n02x5 FILLER_151_781 ();
 b15zdnd11an1n64x5 FILLER_151_803 ();
 b15zdnd11an1n04x5 FILLER_151_867 ();
 b15zdnd11an1n32x5 FILLER_151_882 ();
 b15zdnd11an1n16x5 FILLER_151_914 ();
 b15zdnd11an1n04x5 FILLER_151_930 ();
 b15zdnd00an1n02x5 FILLER_151_934 ();
 b15zdnd00an1n01x5 FILLER_151_936 ();
 b15zdnd11an1n08x5 FILLER_151_968 ();
 b15zdnd11an1n04x5 FILLER_151_976 ();
 b15zdnd00an1n01x5 FILLER_151_980 ();
 b15zdnd11an1n16x5 FILLER_151_1001 ();
 b15zdnd11an1n04x5 FILLER_151_1017 ();
 b15zdnd00an1n01x5 FILLER_151_1021 ();
 b15zdnd11an1n04x5 FILLER_151_1031 ();
 b15zdnd11an1n64x5 FILLER_151_1055 ();
 b15zdnd11an1n16x5 FILLER_151_1119 ();
 b15zdnd11an1n08x5 FILLER_151_1135 ();
 b15zdnd00an1n02x5 FILLER_151_1143 ();
 b15zdnd11an1n08x5 FILLER_151_1160 ();
 b15zdnd11an1n04x5 FILLER_151_1168 ();
 b15zdnd11an1n16x5 FILLER_151_1198 ();
 b15zdnd11an1n08x5 FILLER_151_1214 ();
 b15zdnd11an1n04x5 FILLER_151_1222 ();
 b15zdnd11an1n64x5 FILLER_151_1254 ();
 b15zdnd11an1n32x5 FILLER_151_1318 ();
 b15zdnd11an1n04x5 FILLER_151_1356 ();
 b15zdnd00an1n02x5 FILLER_151_1360 ();
 b15zdnd00an1n01x5 FILLER_151_1362 ();
 b15zdnd11an1n16x5 FILLER_151_1375 ();
 b15zdnd11an1n08x5 FILLER_151_1391 ();
 b15zdnd00an1n02x5 FILLER_151_1399 ();
 b15zdnd11an1n16x5 FILLER_151_1407 ();
 b15zdnd11an1n08x5 FILLER_151_1423 ();
 b15zdnd11an1n16x5 FILLER_151_1441 ();
 b15zdnd11an1n04x5 FILLER_151_1457 ();
 b15zdnd11an1n32x5 FILLER_151_1471 ();
 b15zdnd11an1n16x5 FILLER_151_1503 ();
 b15zdnd00an1n02x5 FILLER_151_1519 ();
 b15zdnd11an1n08x5 FILLER_151_1541 ();
 b15zdnd00an1n02x5 FILLER_151_1549 ();
 b15zdnd00an1n01x5 FILLER_151_1551 ();
 b15zdnd11an1n16x5 FILLER_151_1568 ();
 b15zdnd00an1n01x5 FILLER_151_1584 ();
 b15zdnd11an1n04x5 FILLER_151_1601 ();
 b15zdnd11an1n08x5 FILLER_151_1617 ();
 b15zdnd00an1n01x5 FILLER_151_1625 ();
 b15zdnd11an1n32x5 FILLER_151_1657 ();
 b15zdnd11an1n16x5 FILLER_151_1689 ();
 b15zdnd11an1n08x5 FILLER_151_1705 ();
 b15zdnd00an1n01x5 FILLER_151_1713 ();
 b15zdnd11an1n16x5 FILLER_151_1734 ();
 b15zdnd11an1n08x5 FILLER_151_1750 ();
 b15zdnd00an1n01x5 FILLER_151_1758 ();
 b15zdnd11an1n32x5 FILLER_151_1770 ();
 b15zdnd11an1n08x5 FILLER_151_1802 ();
 b15zdnd00an1n01x5 FILLER_151_1810 ();
 b15zdnd11an1n64x5 FILLER_151_1831 ();
 b15zdnd11an1n64x5 FILLER_151_1895 ();
 b15zdnd11an1n64x5 FILLER_151_1959 ();
 b15zdnd11an1n64x5 FILLER_151_2023 ();
 b15zdnd11an1n16x5 FILLER_151_2087 ();
 b15zdnd11an1n04x5 FILLER_151_2103 ();
 b15zdnd00an1n02x5 FILLER_151_2107 ();
 b15zdnd11an1n08x5 FILLER_151_2129 ();
 b15zdnd11an1n04x5 FILLER_151_2137 ();
 b15zdnd11an1n04x5 FILLER_151_2151 ();
 b15zdnd11an1n04x5 FILLER_151_2164 ();
 b15zdnd00an1n02x5 FILLER_151_2168 ();
 b15zdnd00an1n01x5 FILLER_151_2170 ();
 b15zdnd11an1n32x5 FILLER_151_2191 ();
 b15zdnd11an1n16x5 FILLER_151_2223 ();
 b15zdnd11an1n04x5 FILLER_151_2239 ();
 b15zdnd00an1n02x5 FILLER_151_2243 ();
 b15zdnd00an1n01x5 FILLER_151_2245 ();
 b15zdnd11an1n04x5 FILLER_151_2257 ();
 b15zdnd11an1n04x5 FILLER_151_2265 ();
 b15zdnd11an1n08x5 FILLER_151_2273 ();
 b15zdnd00an1n02x5 FILLER_151_2281 ();
 b15zdnd00an1n01x5 FILLER_151_2283 ();
 b15zdnd11an1n32x5 FILLER_152_8 ();
 b15zdnd11an1n04x5 FILLER_152_40 ();
 b15zdnd00an1n01x5 FILLER_152_44 ();
 b15zdnd11an1n04x5 FILLER_152_50 ();
 b15zdnd00an1n01x5 FILLER_152_54 ();
 b15zdnd11an1n64x5 FILLER_152_59 ();
 b15zdnd11an1n32x5 FILLER_152_123 ();
 b15zdnd00an1n02x5 FILLER_152_155 ();
 b15zdnd11an1n16x5 FILLER_152_167 ();
 b15zdnd00an1n02x5 FILLER_152_183 ();
 b15zdnd11an1n08x5 FILLER_152_193 ();
 b15zdnd11an1n32x5 FILLER_152_227 ();
 b15zdnd11an1n16x5 FILLER_152_259 ();
 b15zdnd00an1n01x5 FILLER_152_275 ();
 b15zdnd11an1n04x5 FILLER_152_289 ();
 b15zdnd11an1n04x5 FILLER_152_299 ();
 b15zdnd11an1n16x5 FILLER_152_312 ();
 b15zdnd11an1n08x5 FILLER_152_328 ();
 b15zdnd11an1n04x5 FILLER_152_336 ();
 b15zdnd00an1n01x5 FILLER_152_340 ();
 b15zdnd11an1n04x5 FILLER_152_348 ();
 b15zdnd00an1n01x5 FILLER_152_352 ();
 b15zdnd11an1n32x5 FILLER_152_360 ();
 b15zdnd11an1n16x5 FILLER_152_392 ();
 b15zdnd11an1n08x5 FILLER_152_408 ();
 b15zdnd11an1n08x5 FILLER_152_422 ();
 b15zdnd11an1n04x5 FILLER_152_430 ();
 b15zdnd00an1n01x5 FILLER_152_434 ();
 b15zdnd11an1n16x5 FILLER_152_440 ();
 b15zdnd11an1n08x5 FILLER_152_456 ();
 b15zdnd11an1n04x5 FILLER_152_464 ();
 b15zdnd00an1n01x5 FILLER_152_468 ();
 b15zdnd11an1n64x5 FILLER_152_473 ();
 b15zdnd11an1n16x5 FILLER_152_537 ();
 b15zdnd00an1n02x5 FILLER_152_553 ();
 b15zdnd00an1n01x5 FILLER_152_555 ();
 b15zdnd11an1n04x5 FILLER_152_568 ();
 b15zdnd11an1n16x5 FILLER_152_592 ();
 b15zdnd11an1n08x5 FILLER_152_608 ();
 b15zdnd11an1n04x5 FILLER_152_632 ();
 b15zdnd11an1n16x5 FILLER_152_640 ();
 b15zdnd11an1n04x5 FILLER_152_656 ();
 b15zdnd00an1n02x5 FILLER_152_660 ();
 b15zdnd00an1n01x5 FILLER_152_662 ();
 b15zdnd11an1n16x5 FILLER_152_668 ();
 b15zdnd11an1n04x5 FILLER_152_684 ();
 b15zdnd00an1n02x5 FILLER_152_688 ();
 b15zdnd11an1n08x5 FILLER_152_708 ();
 b15zdnd00an1n02x5 FILLER_152_716 ();
 b15zdnd11an1n64x5 FILLER_152_726 ();
 b15zdnd11an1n64x5 FILLER_152_790 ();
 b15zdnd11an1n16x5 FILLER_152_854 ();
 b15zdnd11an1n04x5 FILLER_152_870 ();
 b15zdnd11an1n08x5 FILLER_152_894 ();
 b15zdnd11an1n16x5 FILLER_152_906 ();
 b15zdnd11an1n08x5 FILLER_152_922 ();
 b15zdnd11an1n04x5 FILLER_152_930 ();
 b15zdnd00an1n02x5 FILLER_152_934 ();
 b15zdnd00an1n01x5 FILLER_152_936 ();
 b15zdnd11an1n64x5 FILLER_152_968 ();
 b15zdnd11an1n32x5 FILLER_152_1032 ();
 b15zdnd11an1n04x5 FILLER_152_1064 ();
 b15zdnd00an1n02x5 FILLER_152_1068 ();
 b15zdnd11an1n64x5 FILLER_152_1082 ();
 b15zdnd11an1n64x5 FILLER_152_1146 ();
 b15zdnd11an1n32x5 FILLER_152_1210 ();
 b15zdnd11an1n08x5 FILLER_152_1254 ();
 b15zdnd00an1n01x5 FILLER_152_1262 ();
 b15zdnd11an1n04x5 FILLER_152_1274 ();
 b15zdnd11an1n08x5 FILLER_152_1285 ();
 b15zdnd00an1n02x5 FILLER_152_1293 ();
 b15zdnd11an1n32x5 FILLER_152_1301 ();
 b15zdnd11an1n16x5 FILLER_152_1333 ();
 b15zdnd11an1n04x5 FILLER_152_1349 ();
 b15zdnd11an1n64x5 FILLER_152_1358 ();
 b15zdnd11an1n16x5 FILLER_152_1422 ();
 b15zdnd11an1n08x5 FILLER_152_1438 ();
 b15zdnd11an1n04x5 FILLER_152_1446 ();
 b15zdnd00an1n02x5 FILLER_152_1450 ();
 b15zdnd00an1n01x5 FILLER_152_1452 ();
 b15zdnd11an1n64x5 FILLER_152_1458 ();
 b15zdnd11an1n16x5 FILLER_152_1522 ();
 b15zdnd11an1n04x5 FILLER_152_1538 ();
 b15zdnd11an1n16x5 FILLER_152_1565 ();
 b15zdnd11an1n08x5 FILLER_152_1581 ();
 b15zdnd11an1n04x5 FILLER_152_1589 ();
 b15zdnd00an1n02x5 FILLER_152_1593 ();
 b15zdnd00an1n01x5 FILLER_152_1595 ();
 b15zdnd11an1n16x5 FILLER_152_1622 ();
 b15zdnd11an1n08x5 FILLER_152_1638 ();
 b15zdnd11an1n04x5 FILLER_152_1646 ();
 b15zdnd11an1n32x5 FILLER_152_1655 ();
 b15zdnd11an1n04x5 FILLER_152_1687 ();
 b15zdnd00an1n02x5 FILLER_152_1691 ();
 b15zdnd11an1n04x5 FILLER_152_1724 ();
 b15zdnd11an1n64x5 FILLER_152_1733 ();
 b15zdnd11an1n04x5 FILLER_152_1797 ();
 b15zdnd00an1n02x5 FILLER_152_1801 ();
 b15zdnd11an1n04x5 FILLER_152_1807 ();
 b15zdnd11an1n64x5 FILLER_152_1816 ();
 b15zdnd11an1n32x5 FILLER_152_1880 ();
 b15zdnd11an1n16x5 FILLER_152_1912 ();
 b15zdnd00an1n01x5 FILLER_152_1928 ();
 b15zdnd11an1n32x5 FILLER_152_1939 ();
 b15zdnd11an1n08x5 FILLER_152_1971 ();
 b15zdnd11an1n04x5 FILLER_152_1979 ();
 b15zdnd00an1n01x5 FILLER_152_1983 ();
 b15zdnd11an1n64x5 FILLER_152_2001 ();
 b15zdnd11an1n32x5 FILLER_152_2065 ();
 b15zdnd11an1n16x5 FILLER_152_2097 ();
 b15zdnd11an1n08x5 FILLER_152_2113 ();
 b15zdnd11an1n04x5 FILLER_152_2121 ();
 b15zdnd00an1n02x5 FILLER_152_2125 ();
 b15zdnd11an1n16x5 FILLER_152_2138 ();
 b15zdnd11an1n08x5 FILLER_152_2162 ();
 b15zdnd11an1n32x5 FILLER_152_2181 ();
 b15zdnd11an1n16x5 FILLER_152_2213 ();
 b15zdnd00an1n01x5 FILLER_152_2229 ();
 b15zdnd11an1n08x5 FILLER_152_2233 ();
 b15zdnd11an1n04x5 FILLER_152_2241 ();
 b15zdnd00an1n01x5 FILLER_152_2245 ();
 b15zdnd11an1n16x5 FILLER_152_2250 ();
 b15zdnd00an1n01x5 FILLER_152_2266 ();
 b15zdnd11an1n04x5 FILLER_152_2271 ();
 b15zdnd00an1n01x5 FILLER_152_2275 ();
 b15zdnd11an1n32x5 FILLER_153_0 ();
 b15zdnd11an1n16x5 FILLER_153_32 ();
 b15zdnd00an1n02x5 FILLER_153_48 ();
 b15zdnd11an1n64x5 FILLER_153_63 ();
 b15zdnd11an1n32x5 FILLER_153_127 ();
 b15zdnd00an1n02x5 FILLER_153_159 ();
 b15zdnd11an1n16x5 FILLER_153_171 ();
 b15zdnd11an1n04x5 FILLER_153_187 ();
 b15zdnd00an1n02x5 FILLER_153_191 ();
 b15zdnd00an1n01x5 FILLER_153_193 ();
 b15zdnd11an1n16x5 FILLER_153_201 ();
 b15zdnd11an1n04x5 FILLER_153_217 ();
 b15zdnd00an1n02x5 FILLER_153_221 ();
 b15zdnd11an1n32x5 FILLER_153_228 ();
 b15zdnd11an1n04x5 FILLER_153_260 ();
 b15zdnd00an1n02x5 FILLER_153_264 ();
 b15zdnd11an1n64x5 FILLER_153_272 ();
 b15zdnd11an1n64x5 FILLER_153_336 ();
 b15zdnd11an1n08x5 FILLER_153_400 ();
 b15zdnd00an1n02x5 FILLER_153_408 ();
 b15zdnd00an1n01x5 FILLER_153_410 ();
 b15zdnd11an1n04x5 FILLER_153_427 ();
 b15zdnd11an1n08x5 FILLER_153_437 ();
 b15zdnd11an1n04x5 FILLER_153_445 ();
 b15zdnd00an1n01x5 FILLER_153_449 ();
 b15zdnd11an1n04x5 FILLER_153_456 ();
 b15zdnd00an1n01x5 FILLER_153_460 ();
 b15zdnd11an1n32x5 FILLER_153_474 ();
 b15zdnd00an1n01x5 FILLER_153_506 ();
 b15zdnd11an1n32x5 FILLER_153_529 ();
 b15zdnd11an1n16x5 FILLER_153_561 ();
 b15zdnd11an1n08x5 FILLER_153_577 ();
 b15zdnd11an1n04x5 FILLER_153_585 ();
 b15zdnd00an1n02x5 FILLER_153_589 ();
 b15zdnd11an1n16x5 FILLER_153_603 ();
 b15zdnd00an1n02x5 FILLER_153_619 ();
 b15zdnd00an1n01x5 FILLER_153_621 ();
 b15zdnd11an1n16x5 FILLER_153_643 ();
 b15zdnd11an1n04x5 FILLER_153_659 ();
 b15zdnd00an1n01x5 FILLER_153_663 ();
 b15zdnd11an1n32x5 FILLER_153_677 ();
 b15zdnd11an1n16x5 FILLER_153_709 ();
 b15zdnd11an1n04x5 FILLER_153_725 ();
 b15zdnd00an1n02x5 FILLER_153_729 ();
 b15zdnd11an1n32x5 FILLER_153_751 ();
 b15zdnd11an1n08x5 FILLER_153_783 ();
 b15zdnd11an1n04x5 FILLER_153_791 ();
 b15zdnd00an1n01x5 FILLER_153_795 ();
 b15zdnd11an1n04x5 FILLER_153_801 ();
 b15zdnd11an1n04x5 FILLER_153_825 ();
 b15zdnd11an1n64x5 FILLER_153_832 ();
 b15zdnd11an1n64x5 FILLER_153_896 ();
 b15zdnd11an1n32x5 FILLER_153_960 ();
 b15zdnd11an1n16x5 FILLER_153_992 ();
 b15zdnd11an1n08x5 FILLER_153_1008 ();
 b15zdnd11an1n04x5 FILLER_153_1016 ();
 b15zdnd00an1n01x5 FILLER_153_1020 ();
 b15zdnd11an1n64x5 FILLER_153_1047 ();
 b15zdnd11an1n64x5 FILLER_153_1111 ();
 b15zdnd11an1n08x5 FILLER_153_1175 ();
 b15zdnd11an1n04x5 FILLER_153_1183 ();
 b15zdnd00an1n01x5 FILLER_153_1187 ();
 b15zdnd11an1n32x5 FILLER_153_1197 ();
 b15zdnd11an1n08x5 FILLER_153_1229 ();
 b15zdnd11an1n04x5 FILLER_153_1237 ();
 b15zdnd11an1n16x5 FILLER_153_1251 ();
 b15zdnd00an1n02x5 FILLER_153_1267 ();
 b15zdnd11an1n04x5 FILLER_153_1276 ();
 b15zdnd11an1n04x5 FILLER_153_1296 ();
 b15zdnd11an1n32x5 FILLER_153_1307 ();
 b15zdnd11an1n08x5 FILLER_153_1339 ();
 b15zdnd11an1n04x5 FILLER_153_1347 ();
 b15zdnd00an1n01x5 FILLER_153_1351 ();
 b15zdnd11an1n64x5 FILLER_153_1366 ();
 b15zdnd11an1n08x5 FILLER_153_1430 ();
 b15zdnd00an1n02x5 FILLER_153_1438 ();
 b15zdnd00an1n01x5 FILLER_153_1440 ();
 b15zdnd11an1n04x5 FILLER_153_1463 ();
 b15zdnd11an1n08x5 FILLER_153_1471 ();
 b15zdnd11an1n64x5 FILLER_153_1491 ();
 b15zdnd11an1n08x5 FILLER_153_1555 ();
 b15zdnd11an1n04x5 FILLER_153_1563 ();
 b15zdnd00an1n02x5 FILLER_153_1567 ();
 b15zdnd11an1n04x5 FILLER_153_1579 ();
 b15zdnd11an1n08x5 FILLER_153_1599 ();
 b15zdnd00an1n01x5 FILLER_153_1607 ();
 b15zdnd11an1n64x5 FILLER_153_1634 ();
 b15zdnd11an1n32x5 FILLER_153_1698 ();
 b15zdnd11an1n16x5 FILLER_153_1730 ();
 b15zdnd00an1n02x5 FILLER_153_1746 ();
 b15zdnd00an1n01x5 FILLER_153_1748 ();
 b15zdnd11an1n16x5 FILLER_153_1780 ();
 b15zdnd11an1n08x5 FILLER_153_1796 ();
 b15zdnd00an1n02x5 FILLER_153_1804 ();
 b15zdnd00an1n01x5 FILLER_153_1806 ();
 b15zdnd11an1n64x5 FILLER_153_1822 ();
 b15zdnd11an1n32x5 FILLER_153_1886 ();
 b15zdnd11an1n08x5 FILLER_153_1918 ();
 b15zdnd11an1n04x5 FILLER_153_1926 ();
 b15zdnd11an1n16x5 FILLER_153_1953 ();
 b15zdnd11an1n08x5 FILLER_153_1969 ();
 b15zdnd00an1n02x5 FILLER_153_1977 ();
 b15zdnd11an1n16x5 FILLER_153_2010 ();
 b15zdnd11an1n04x5 FILLER_153_2026 ();
 b15zdnd00an1n02x5 FILLER_153_2030 ();
 b15zdnd00an1n01x5 FILLER_153_2032 ();
 b15zdnd11an1n04x5 FILLER_153_2045 ();
 b15zdnd00an1n01x5 FILLER_153_2049 ();
 b15zdnd11an1n08x5 FILLER_153_2076 ();
 b15zdnd00an1n01x5 FILLER_153_2084 ();
 b15zdnd11an1n64x5 FILLER_153_2107 ();
 b15zdnd11an1n32x5 FILLER_153_2171 ();
 b15zdnd00an1n02x5 FILLER_153_2203 ();
 b15zdnd11an1n08x5 FILLER_153_2225 ();
 b15zdnd11an1n08x5 FILLER_153_2237 ();
 b15zdnd00an1n01x5 FILLER_153_2245 ();
 b15zdnd11an1n04x5 FILLER_153_2249 ();
 b15zdnd11an1n04x5 FILLER_153_2257 ();
 b15zdnd11an1n04x5 FILLER_153_2265 ();
 b15zdnd11an1n08x5 FILLER_153_2273 ();
 b15zdnd00an1n02x5 FILLER_153_2281 ();
 b15zdnd00an1n01x5 FILLER_153_2283 ();
 b15zdnd11an1n64x5 FILLER_154_8 ();
 b15zdnd00an1n02x5 FILLER_154_72 ();
 b15zdnd00an1n01x5 FILLER_154_74 ();
 b15zdnd11an1n16x5 FILLER_154_88 ();
 b15zdnd00an1n02x5 FILLER_154_104 ();
 b15zdnd11an1n64x5 FILLER_154_110 ();
 b15zdnd11an1n32x5 FILLER_154_174 ();
 b15zdnd11an1n08x5 FILLER_154_206 ();
 b15zdnd11an1n04x5 FILLER_154_214 ();
 b15zdnd00an1n01x5 FILLER_154_218 ();
 b15zdnd11an1n08x5 FILLER_154_224 ();
 b15zdnd11an1n04x5 FILLER_154_232 ();
 b15zdnd11an1n08x5 FILLER_154_242 ();
 b15zdnd11an1n04x5 FILLER_154_250 ();
 b15zdnd00an1n02x5 FILLER_154_254 ();
 b15zdnd00an1n01x5 FILLER_154_256 ();
 b15zdnd11an1n32x5 FILLER_154_261 ();
 b15zdnd11an1n08x5 FILLER_154_293 ();
 b15zdnd00an1n01x5 FILLER_154_301 ();
 b15zdnd11an1n04x5 FILLER_154_314 ();
 b15zdnd00an1n02x5 FILLER_154_318 ();
 b15zdnd11an1n64x5 FILLER_154_333 ();
 b15zdnd11an1n04x5 FILLER_154_397 ();
 b15zdnd00an1n02x5 FILLER_154_401 ();
 b15zdnd00an1n01x5 FILLER_154_403 ();
 b15zdnd11an1n32x5 FILLER_154_413 ();
 b15zdnd11an1n08x5 FILLER_154_445 ();
 b15zdnd11an1n04x5 FILLER_154_453 ();
 b15zdnd00an1n02x5 FILLER_154_457 ();
 b15zdnd00an1n01x5 FILLER_154_459 ();
 b15zdnd11an1n32x5 FILLER_154_481 ();
 b15zdnd11an1n16x5 FILLER_154_513 ();
 b15zdnd11an1n08x5 FILLER_154_529 ();
 b15zdnd11an1n04x5 FILLER_154_537 ();
 b15zdnd00an1n01x5 FILLER_154_541 ();
 b15zdnd11an1n64x5 FILLER_154_553 ();
 b15zdnd11an1n64x5 FILLER_154_617 ();
 b15zdnd11an1n04x5 FILLER_154_681 ();
 b15zdnd11an1n16x5 FILLER_154_691 ();
 b15zdnd11an1n08x5 FILLER_154_707 ();
 b15zdnd00an1n02x5 FILLER_154_715 ();
 b15zdnd00an1n01x5 FILLER_154_717 ();
 b15zdnd11an1n04x5 FILLER_154_726 ();
 b15zdnd00an1n02x5 FILLER_154_730 ();
 b15zdnd11an1n64x5 FILLER_154_748 ();
 b15zdnd11an1n64x5 FILLER_154_812 ();
 b15zdnd11an1n32x5 FILLER_154_876 ();
 b15zdnd11an1n16x5 FILLER_154_908 ();
 b15zdnd11an1n08x5 FILLER_154_924 ();
 b15zdnd11an1n04x5 FILLER_154_932 ();
 b15zdnd00an1n02x5 FILLER_154_936 ();
 b15zdnd11an1n64x5 FILLER_154_964 ();
 b15zdnd11an1n64x5 FILLER_154_1028 ();
 b15zdnd11an1n64x5 FILLER_154_1092 ();
 b15zdnd11an1n16x5 FILLER_154_1156 ();
 b15zdnd11an1n04x5 FILLER_154_1172 ();
 b15zdnd00an1n02x5 FILLER_154_1176 ();
 b15zdnd00an1n01x5 FILLER_154_1178 ();
 b15zdnd11an1n64x5 FILLER_154_1188 ();
 b15zdnd11an1n32x5 FILLER_154_1252 ();
 b15zdnd11an1n08x5 FILLER_154_1284 ();
 b15zdnd11an1n04x5 FILLER_154_1292 ();
 b15zdnd00an1n02x5 FILLER_154_1296 ();
 b15zdnd00an1n01x5 FILLER_154_1298 ();
 b15zdnd11an1n04x5 FILLER_154_1305 ();
 b15zdnd11an1n16x5 FILLER_154_1315 ();
 b15zdnd11an1n08x5 FILLER_154_1331 ();
 b15zdnd00an1n02x5 FILLER_154_1339 ();
 b15zdnd00an1n01x5 FILLER_154_1341 ();
 b15zdnd11an1n64x5 FILLER_154_1363 ();
 b15zdnd11an1n64x5 FILLER_154_1427 ();
 b15zdnd11an1n16x5 FILLER_154_1491 ();
 b15zdnd11an1n08x5 FILLER_154_1507 ();
 b15zdnd11an1n04x5 FILLER_154_1515 ();
 b15zdnd00an1n01x5 FILLER_154_1519 ();
 b15zdnd11an1n04x5 FILLER_154_1526 ();
 b15zdnd11an1n32x5 FILLER_154_1536 ();
 b15zdnd11an1n08x5 FILLER_154_1568 ();
 b15zdnd00an1n01x5 FILLER_154_1576 ();
 b15zdnd11an1n32x5 FILLER_154_1593 ();
 b15zdnd11an1n04x5 FILLER_154_1625 ();
 b15zdnd11an1n04x5 FILLER_154_1655 ();
 b15zdnd11an1n64x5 FILLER_154_1679 ();
 b15zdnd11an1n08x5 FILLER_154_1743 ();
 b15zdnd11an1n64x5 FILLER_154_1769 ();
 b15zdnd11an1n32x5 FILLER_154_1833 ();
 b15zdnd11an1n16x5 FILLER_154_1865 ();
 b15zdnd11an1n04x5 FILLER_154_1881 ();
 b15zdnd00an1n02x5 FILLER_154_1885 ();
 b15zdnd11an1n64x5 FILLER_154_1905 ();
 b15zdnd11an1n64x5 FILLER_154_1969 ();
 b15zdnd00an1n02x5 FILLER_154_2033 ();
 b15zdnd00an1n01x5 FILLER_154_2035 ();
 b15zdnd11an1n16x5 FILLER_154_2061 ();
 b15zdnd11an1n08x5 FILLER_154_2077 ();
 b15zdnd00an1n01x5 FILLER_154_2085 ();
 b15zdnd11an1n08x5 FILLER_154_2117 ();
 b15zdnd11an1n04x5 FILLER_154_2125 ();
 b15zdnd00an1n02x5 FILLER_154_2129 ();
 b15zdnd00an1n02x5 FILLER_154_2152 ();
 b15zdnd11an1n32x5 FILLER_154_2162 ();
 b15zdnd11an1n16x5 FILLER_154_2194 ();
 b15zdnd11an1n08x5 FILLER_154_2210 ();
 b15zdnd11an1n04x5 FILLER_154_2218 ();
 b15zdnd00an1n02x5 FILLER_154_2222 ();
 b15zdnd11an1n08x5 FILLER_154_2228 ();
 b15zdnd11an1n04x5 FILLER_154_2236 ();
 b15zdnd11an1n16x5 FILLER_154_2250 ();
 b15zdnd11an1n04x5 FILLER_154_2266 ();
 b15zdnd00an1n02x5 FILLER_154_2274 ();
 b15zdnd11an1n64x5 FILLER_155_0 ();
 b15zdnd11an1n08x5 FILLER_155_64 ();
 b15zdnd11an1n04x5 FILLER_155_72 ();
 b15zdnd11an1n08x5 FILLER_155_89 ();
 b15zdnd00an1n02x5 FILLER_155_97 ();
 b15zdnd00an1n01x5 FILLER_155_99 ();
 b15zdnd11an1n04x5 FILLER_155_105 ();
 b15zdnd00an1n01x5 FILLER_155_109 ();
 b15zdnd11an1n16x5 FILLER_155_123 ();
 b15zdnd11an1n08x5 FILLER_155_139 ();
 b15zdnd00an1n02x5 FILLER_155_147 ();
 b15zdnd00an1n01x5 FILLER_155_149 ();
 b15zdnd11an1n32x5 FILLER_155_160 ();
 b15zdnd11an1n04x5 FILLER_155_192 ();
 b15zdnd00an1n01x5 FILLER_155_196 ();
 b15zdnd11an1n04x5 FILLER_155_209 ();
 b15zdnd00an1n01x5 FILLER_155_213 ();
 b15zdnd11an1n04x5 FILLER_155_228 ();
 b15zdnd11an1n08x5 FILLER_155_238 ();
 b15zdnd11an1n04x5 FILLER_155_246 ();
 b15zdnd00an1n02x5 FILLER_155_250 ();
 b15zdnd00an1n01x5 FILLER_155_252 ();
 b15zdnd11an1n08x5 FILLER_155_260 ();
 b15zdnd11an1n04x5 FILLER_155_268 ();
 b15zdnd11an1n32x5 FILLER_155_279 ();
 b15zdnd11an1n08x5 FILLER_155_311 ();
 b15zdnd00an1n01x5 FILLER_155_319 ();
 b15zdnd11an1n04x5 FILLER_155_328 ();
 b15zdnd11an1n64x5 FILLER_155_336 ();
 b15zdnd11an1n64x5 FILLER_155_400 ();
 b15zdnd11an1n32x5 FILLER_155_464 ();
 b15zdnd11an1n08x5 FILLER_155_496 ();
 b15zdnd11an1n04x5 FILLER_155_504 ();
 b15zdnd00an1n02x5 FILLER_155_508 ();
 b15zdnd00an1n01x5 FILLER_155_510 ();
 b15zdnd11an1n16x5 FILLER_155_520 ();
 b15zdnd11an1n08x5 FILLER_155_536 ();
 b15zdnd00an1n02x5 FILLER_155_544 ();
 b15zdnd00an1n01x5 FILLER_155_546 ();
 b15zdnd11an1n08x5 FILLER_155_555 ();
 b15zdnd11an1n04x5 FILLER_155_563 ();
 b15zdnd11an1n08x5 FILLER_155_571 ();
 b15zdnd11an1n04x5 FILLER_155_579 ();
 b15zdnd00an1n02x5 FILLER_155_583 ();
 b15zdnd00an1n01x5 FILLER_155_585 ();
 b15zdnd11an1n04x5 FILLER_155_595 ();
 b15zdnd11an1n64x5 FILLER_155_604 ();
 b15zdnd11an1n16x5 FILLER_155_668 ();
 b15zdnd11an1n08x5 FILLER_155_691 ();
 b15zdnd11an1n04x5 FILLER_155_699 ();
 b15zdnd00an1n02x5 FILLER_155_703 ();
 b15zdnd00an1n01x5 FILLER_155_705 ();
 b15zdnd11an1n16x5 FILLER_155_712 ();
 b15zdnd11an1n04x5 FILLER_155_728 ();
 b15zdnd00an1n01x5 FILLER_155_732 ();
 b15zdnd11an1n32x5 FILLER_155_751 ();
 b15zdnd11an1n04x5 FILLER_155_783 ();
 b15zdnd11an1n64x5 FILLER_155_791 ();
 b15zdnd11an1n08x5 FILLER_155_855 ();
 b15zdnd00an1n01x5 FILLER_155_863 ();
 b15zdnd11an1n32x5 FILLER_155_867 ();
 b15zdnd11an1n16x5 FILLER_155_899 ();
 b15zdnd11an1n04x5 FILLER_155_915 ();
 b15zdnd00an1n02x5 FILLER_155_919 ();
 b15zdnd11an1n16x5 FILLER_155_953 ();
 b15zdnd11an1n04x5 FILLER_155_969 ();
 b15zdnd11an1n04x5 FILLER_155_980 ();
 b15zdnd11an1n64x5 FILLER_155_1010 ();
 b15zdnd11an1n16x5 FILLER_155_1074 ();
 b15zdnd11an1n04x5 FILLER_155_1090 ();
 b15zdnd00an1n02x5 FILLER_155_1094 ();
 b15zdnd00an1n01x5 FILLER_155_1096 ();
 b15zdnd11an1n04x5 FILLER_155_1122 ();
 b15zdnd11an1n16x5 FILLER_155_1152 ();
 b15zdnd11an1n04x5 FILLER_155_1168 ();
 b15zdnd11an1n64x5 FILLER_155_1183 ();
 b15zdnd11an1n32x5 FILLER_155_1247 ();
 b15zdnd00an1n01x5 FILLER_155_1279 ();
 b15zdnd11an1n04x5 FILLER_155_1296 ();
 b15zdnd11an1n64x5 FILLER_155_1305 ();
 b15zdnd11an1n16x5 FILLER_155_1369 ();
 b15zdnd11an1n04x5 FILLER_155_1385 ();
 b15zdnd00an1n01x5 FILLER_155_1389 ();
 b15zdnd11an1n16x5 FILLER_155_1399 ();
 b15zdnd11an1n16x5 FILLER_155_1426 ();
 b15zdnd11an1n04x5 FILLER_155_1442 ();
 b15zdnd00an1n02x5 FILLER_155_1446 ();
 b15zdnd11an1n04x5 FILLER_155_1462 ();
 b15zdnd11an1n04x5 FILLER_155_1473 ();
 b15zdnd11an1n04x5 FILLER_155_1481 ();
 b15zdnd11an1n16x5 FILLER_155_1490 ();
 b15zdnd11an1n04x5 FILLER_155_1506 ();
 b15zdnd00an1n01x5 FILLER_155_1510 ();
 b15zdnd11an1n04x5 FILLER_155_1523 ();
 b15zdnd11an1n04x5 FILLER_155_1537 ();
 b15zdnd11an1n04x5 FILLER_155_1566 ();
 b15zdnd11an1n64x5 FILLER_155_1602 ();
 b15zdnd11an1n32x5 FILLER_155_1666 ();
 b15zdnd11an1n04x5 FILLER_155_1698 ();
 b15zdnd11an1n04x5 FILLER_155_1706 ();
 b15zdnd11an1n64x5 FILLER_155_1730 ();
 b15zdnd11an1n16x5 FILLER_155_1794 ();
 b15zdnd00an1n02x5 FILLER_155_1810 ();
 b15zdnd00an1n01x5 FILLER_155_1812 ();
 b15zdnd11an1n32x5 FILLER_155_1824 ();
 b15zdnd11an1n04x5 FILLER_155_1856 ();
 b15zdnd00an1n02x5 FILLER_155_1860 ();
 b15zdnd11an1n04x5 FILLER_155_1882 ();
 b15zdnd11an1n32x5 FILLER_155_1917 ();
 b15zdnd11an1n04x5 FILLER_155_1949 ();
 b15zdnd00an1n02x5 FILLER_155_1953 ();
 b15zdnd00an1n01x5 FILLER_155_1955 ();
 b15zdnd11an1n32x5 FILLER_155_1996 ();
 b15zdnd00an1n02x5 FILLER_155_2028 ();
 b15zdnd00an1n01x5 FILLER_155_2030 ();
 b15zdnd11an1n04x5 FILLER_155_2040 ();
 b15zdnd11an1n64x5 FILLER_155_2054 ();
 b15zdnd11an1n64x5 FILLER_155_2118 ();
 b15zdnd11an1n32x5 FILLER_155_2182 ();
 b15zdnd11an1n04x5 FILLER_155_2214 ();
 b15zdnd00an1n02x5 FILLER_155_2218 ();
 b15zdnd11an1n04x5 FILLER_155_2240 ();
 b15zdnd11an1n04x5 FILLER_155_2248 ();
 b15zdnd11an1n04x5 FILLER_155_2256 ();
 b15zdnd11an1n04x5 FILLER_155_2264 ();
 b15zdnd11an1n04x5 FILLER_155_2274 ();
 b15zdnd00an1n02x5 FILLER_155_2282 ();
 b15zdnd11an1n16x5 FILLER_156_8 ();
 b15zdnd11an1n08x5 FILLER_156_24 ();
 b15zdnd11an1n04x5 FILLER_156_32 ();
 b15zdnd11an1n04x5 FILLER_156_45 ();
 b15zdnd11an1n32x5 FILLER_156_61 ();
 b15zdnd11an1n04x5 FILLER_156_93 ();
 b15zdnd11an1n04x5 FILLER_156_112 ();
 b15zdnd00an1n02x5 FILLER_156_116 ();
 b15zdnd11an1n64x5 FILLER_156_124 ();
 b15zdnd11an1n64x5 FILLER_156_188 ();
 b15zdnd11an1n16x5 FILLER_156_252 ();
 b15zdnd11an1n04x5 FILLER_156_268 ();
 b15zdnd00an1n02x5 FILLER_156_272 ();
 b15zdnd11an1n32x5 FILLER_156_294 ();
 b15zdnd00an1n01x5 FILLER_156_326 ();
 b15zdnd11an1n08x5 FILLER_156_334 ();
 b15zdnd11an1n04x5 FILLER_156_342 ();
 b15zdnd11an1n04x5 FILLER_156_351 ();
 b15zdnd11an1n32x5 FILLER_156_360 ();
 b15zdnd11an1n08x5 FILLER_156_392 ();
 b15zdnd00an1n01x5 FILLER_156_400 ();
 b15zdnd11an1n32x5 FILLER_156_410 ();
 b15zdnd11an1n08x5 FILLER_156_442 ();
 b15zdnd11an1n04x5 FILLER_156_450 ();
 b15zdnd11an1n16x5 FILLER_156_460 ();
 b15zdnd11an1n04x5 FILLER_156_476 ();
 b15zdnd11an1n16x5 FILLER_156_496 ();
 b15zdnd00an1n02x5 FILLER_156_512 ();
 b15zdnd11an1n32x5 FILLER_156_520 ();
 b15zdnd11an1n04x5 FILLER_156_552 ();
 b15zdnd00an1n01x5 FILLER_156_556 ();
 b15zdnd11an1n16x5 FILLER_156_569 ();
 b15zdnd00an1n02x5 FILLER_156_585 ();
 b15zdnd11an1n32x5 FILLER_156_600 ();
 b15zdnd11an1n16x5 FILLER_156_632 ();
 b15zdnd11an1n08x5 FILLER_156_648 ();
 b15zdnd11an1n04x5 FILLER_156_656 ();
 b15zdnd11an1n16x5 FILLER_156_670 ();
 b15zdnd11an1n04x5 FILLER_156_686 ();
 b15zdnd11an1n04x5 FILLER_156_697 ();
 b15zdnd11an1n04x5 FILLER_156_706 ();
 b15zdnd00an1n02x5 FILLER_156_716 ();
 b15zdnd11an1n16x5 FILLER_156_726 ();
 b15zdnd11an1n08x5 FILLER_156_742 ();
 b15zdnd00an1n02x5 FILLER_156_750 ();
 b15zdnd11an1n64x5 FILLER_156_770 ();
 b15zdnd11an1n32x5 FILLER_156_834 ();
 b15zdnd11an1n08x5 FILLER_156_866 ();
 b15zdnd11an1n32x5 FILLER_156_884 ();
 b15zdnd11an1n16x5 FILLER_156_916 ();
 b15zdnd11an1n08x5 FILLER_156_932 ();
 b15zdnd11an1n04x5 FILLER_156_940 ();
 b15zdnd00an1n02x5 FILLER_156_944 ();
 b15zdnd00an1n01x5 FILLER_156_946 ();
 b15zdnd11an1n64x5 FILLER_156_973 ();
 b15zdnd11an1n04x5 FILLER_156_1037 ();
 b15zdnd00an1n02x5 FILLER_156_1041 ();
 b15zdnd00an1n01x5 FILLER_156_1043 ();
 b15zdnd11an1n08x5 FILLER_156_1048 ();
 b15zdnd11an1n04x5 FILLER_156_1056 ();
 b15zdnd00an1n02x5 FILLER_156_1060 ();
 b15zdnd00an1n01x5 FILLER_156_1062 ();
 b15zdnd11an1n04x5 FILLER_156_1069 ();
 b15zdnd11an1n16x5 FILLER_156_1084 ();
 b15zdnd11an1n08x5 FILLER_156_1100 ();
 b15zdnd11an1n04x5 FILLER_156_1108 ();
 b15zdnd11an1n16x5 FILLER_156_1121 ();
 b15zdnd11an1n04x5 FILLER_156_1137 ();
 b15zdnd00an1n02x5 FILLER_156_1141 ();
 b15zdnd00an1n01x5 FILLER_156_1143 ();
 b15zdnd11an1n64x5 FILLER_156_1150 ();
 b15zdnd11an1n04x5 FILLER_156_1214 ();
 b15zdnd00an1n02x5 FILLER_156_1218 ();
 b15zdnd00an1n01x5 FILLER_156_1220 ();
 b15zdnd11an1n64x5 FILLER_156_1231 ();
 b15zdnd11an1n04x5 FILLER_156_1295 ();
 b15zdnd00an1n02x5 FILLER_156_1299 ();
 b15zdnd00an1n01x5 FILLER_156_1301 ();
 b15zdnd11an1n16x5 FILLER_156_1314 ();
 b15zdnd11an1n08x5 FILLER_156_1330 ();
 b15zdnd00an1n01x5 FILLER_156_1338 ();
 b15zdnd11an1n04x5 FILLER_156_1348 ();
 b15zdnd00an1n01x5 FILLER_156_1352 ();
 b15zdnd11an1n04x5 FILLER_156_1357 ();
 b15zdnd00an1n02x5 FILLER_156_1361 ();
 b15zdnd11an1n04x5 FILLER_156_1376 ();
 b15zdnd11an1n04x5 FILLER_156_1385 ();
 b15zdnd11an1n08x5 FILLER_156_1398 ();
 b15zdnd11an1n04x5 FILLER_156_1406 ();
 b15zdnd00an1n02x5 FILLER_156_1410 ();
 b15zdnd11an1n32x5 FILLER_156_1422 ();
 b15zdnd11an1n08x5 FILLER_156_1454 ();
 b15zdnd11an1n04x5 FILLER_156_1462 ();
 b15zdnd11an1n64x5 FILLER_156_1476 ();
 b15zdnd00an1n01x5 FILLER_156_1540 ();
 b15zdnd11an1n64x5 FILLER_156_1559 ();
 b15zdnd11an1n64x5 FILLER_156_1623 ();
 b15zdnd11an1n64x5 FILLER_156_1687 ();
 b15zdnd11an1n04x5 FILLER_156_1751 ();
 b15zdnd00an1n02x5 FILLER_156_1755 ();
 b15zdnd11an1n04x5 FILLER_156_1777 ();
 b15zdnd11an1n16x5 FILLER_156_1786 ();
 b15zdnd11an1n08x5 FILLER_156_1802 ();
 b15zdnd11an1n04x5 FILLER_156_1810 ();
 b15zdnd00an1n01x5 FILLER_156_1814 ();
 b15zdnd11an1n64x5 FILLER_156_1835 ();
 b15zdnd11an1n08x5 FILLER_156_1899 ();
 b15zdnd11an1n04x5 FILLER_156_1907 ();
 b15zdnd00an1n02x5 FILLER_156_1911 ();
 b15zdnd11an1n64x5 FILLER_156_1944 ();
 b15zdnd11an1n64x5 FILLER_156_2008 ();
 b15zdnd11an1n08x5 FILLER_156_2072 ();
 b15zdnd11an1n04x5 FILLER_156_2080 ();
 b15zdnd11an1n08x5 FILLER_156_2099 ();
 b15zdnd11an1n04x5 FILLER_156_2107 ();
 b15zdnd00an1n01x5 FILLER_156_2111 ();
 b15zdnd11an1n16x5 FILLER_156_2130 ();
 b15zdnd11an1n08x5 FILLER_156_2146 ();
 b15zdnd11an1n64x5 FILLER_156_2162 ();
 b15zdnd11an1n16x5 FILLER_156_2226 ();
 b15zdnd00an1n02x5 FILLER_156_2242 ();
 b15zdnd11an1n08x5 FILLER_156_2248 ();
 b15zdnd11an1n04x5 FILLER_156_2256 ();
 b15zdnd11an1n08x5 FILLER_156_2264 ();
 b15zdnd11an1n04x5 FILLER_156_2272 ();
 b15zdnd11an1n32x5 FILLER_157_0 ();
 b15zdnd00an1n01x5 FILLER_157_32 ();
 b15zdnd11an1n16x5 FILLER_157_39 ();
 b15zdnd00an1n01x5 FILLER_157_55 ();
 b15zdnd11an1n04x5 FILLER_157_61 ();
 b15zdnd11an1n04x5 FILLER_157_83 ();
 b15zdnd11an1n08x5 FILLER_157_92 ();
 b15zdnd00an1n02x5 FILLER_157_100 ();
 b15zdnd00an1n01x5 FILLER_157_102 ();
 b15zdnd11an1n08x5 FILLER_157_108 ();
 b15zdnd11an1n04x5 FILLER_157_116 ();
 b15zdnd00an1n02x5 FILLER_157_120 ();
 b15zdnd00an1n01x5 FILLER_157_122 ();
 b15zdnd11an1n32x5 FILLER_157_128 ();
 b15zdnd11an1n08x5 FILLER_157_160 ();
 b15zdnd11an1n04x5 FILLER_157_168 ();
 b15zdnd00an1n02x5 FILLER_157_172 ();
 b15zdnd11an1n32x5 FILLER_157_179 ();
 b15zdnd11an1n16x5 FILLER_157_211 ();
 b15zdnd11an1n04x5 FILLER_157_227 ();
 b15zdnd11an1n32x5 FILLER_157_238 ();
 b15zdnd00an1n02x5 FILLER_157_270 ();
 b15zdnd00an1n01x5 FILLER_157_272 ();
 b15zdnd11an1n04x5 FILLER_157_288 ();
 b15zdnd11an1n32x5 FILLER_157_298 ();
 b15zdnd11an1n16x5 FILLER_157_330 ();
 b15zdnd00an1n01x5 FILLER_157_346 ();
 b15zdnd11an1n32x5 FILLER_157_352 ();
 b15zdnd11an1n16x5 FILLER_157_384 ();
 b15zdnd11an1n08x5 FILLER_157_400 ();
 b15zdnd00an1n02x5 FILLER_157_408 ();
 b15zdnd00an1n01x5 FILLER_157_410 ();
 b15zdnd11an1n16x5 FILLER_157_419 ();
 b15zdnd11an1n08x5 FILLER_157_435 ();
 b15zdnd00an1n01x5 FILLER_157_443 ();
 b15zdnd11an1n08x5 FILLER_157_449 ();
 b15zdnd00an1n02x5 FILLER_157_457 ();
 b15zdnd11an1n32x5 FILLER_157_468 ();
 b15zdnd11an1n08x5 FILLER_157_500 ();
 b15zdnd11an1n04x5 FILLER_157_508 ();
 b15zdnd00an1n02x5 FILLER_157_512 ();
 b15zdnd00an1n01x5 FILLER_157_514 ();
 b15zdnd11an1n16x5 FILLER_157_520 ();
 b15zdnd11an1n04x5 FILLER_157_536 ();
 b15zdnd00an1n02x5 FILLER_157_540 ();
 b15zdnd11an1n08x5 FILLER_157_548 ();
 b15zdnd00an1n01x5 FILLER_157_556 ();
 b15zdnd11an1n16x5 FILLER_157_574 ();
 b15zdnd11an1n08x5 FILLER_157_590 ();
 b15zdnd11an1n04x5 FILLER_157_598 ();
 b15zdnd11an1n16x5 FILLER_157_616 ();
 b15zdnd11an1n16x5 FILLER_157_644 ();
 b15zdnd11an1n04x5 FILLER_157_660 ();
 b15zdnd11an1n32x5 FILLER_157_669 ();
 b15zdnd11an1n16x5 FILLER_157_701 ();
 b15zdnd00an1n01x5 FILLER_157_717 ();
 b15zdnd11an1n04x5 FILLER_157_734 ();
 b15zdnd00an1n01x5 FILLER_157_738 ();
 b15zdnd11an1n08x5 FILLER_157_762 ();
 b15zdnd00an1n02x5 FILLER_157_770 ();
 b15zdnd11an1n08x5 FILLER_157_790 ();
 b15zdnd11an1n04x5 FILLER_157_798 ();
 b15zdnd00an1n02x5 FILLER_157_802 ();
 b15zdnd11an1n32x5 FILLER_157_824 ();
 b15zdnd11an1n08x5 FILLER_157_856 ();
 b15zdnd11an1n04x5 FILLER_157_864 ();
 b15zdnd11an1n08x5 FILLER_157_888 ();
 b15zdnd11an1n04x5 FILLER_157_896 ();
 b15zdnd00an1n01x5 FILLER_157_900 ();
 b15zdnd11an1n04x5 FILLER_157_915 ();
 b15zdnd00an1n02x5 FILLER_157_919 ();
 b15zdnd11an1n04x5 FILLER_157_944 ();
 b15zdnd00an1n02x5 FILLER_157_948 ();
 b15zdnd11an1n04x5 FILLER_157_976 ();
 b15zdnd00an1n01x5 FILLER_157_980 ();
 b15zdnd11an1n04x5 FILLER_157_990 ();
 b15zdnd11an1n16x5 FILLER_157_1006 ();
 b15zdnd11an1n08x5 FILLER_157_1022 ();
 b15zdnd11an1n04x5 FILLER_157_1030 ();
 b15zdnd00an1n02x5 FILLER_157_1034 ();
 b15zdnd00an1n01x5 FILLER_157_1036 ();
 b15zdnd11an1n16x5 FILLER_157_1047 ();
 b15zdnd11an1n08x5 FILLER_157_1063 ();
 b15zdnd11an1n04x5 FILLER_157_1071 ();
 b15zdnd00an1n01x5 FILLER_157_1075 ();
 b15zdnd11an1n16x5 FILLER_157_1082 ();
 b15zdnd11an1n08x5 FILLER_157_1098 ();
 b15zdnd11an1n04x5 FILLER_157_1106 ();
 b15zdnd00an1n02x5 FILLER_157_1110 ();
 b15zdnd00an1n01x5 FILLER_157_1112 ();
 b15zdnd11an1n16x5 FILLER_157_1127 ();
 b15zdnd11an1n16x5 FILLER_157_1149 ();
 b15zdnd11an1n08x5 FILLER_157_1165 ();
 b15zdnd00an1n02x5 FILLER_157_1173 ();
 b15zdnd00an1n01x5 FILLER_157_1175 ();
 b15zdnd11an1n64x5 FILLER_157_1188 ();
 b15zdnd11an1n04x5 FILLER_157_1252 ();
 b15zdnd11an1n16x5 FILLER_157_1266 ();
 b15zdnd11an1n04x5 FILLER_157_1282 ();
 b15zdnd00an1n01x5 FILLER_157_1286 ();
 b15zdnd11an1n32x5 FILLER_157_1305 ();
 b15zdnd11an1n16x5 FILLER_157_1337 ();
 b15zdnd00an1n02x5 FILLER_157_1353 ();
 b15zdnd00an1n01x5 FILLER_157_1355 ();
 b15zdnd11an1n16x5 FILLER_157_1365 ();
 b15zdnd11an1n04x5 FILLER_157_1381 ();
 b15zdnd11an1n16x5 FILLER_157_1393 ();
 b15zdnd11an1n08x5 FILLER_157_1409 ();
 b15zdnd00an1n02x5 FILLER_157_1417 ();
 b15zdnd11an1n16x5 FILLER_157_1429 ();
 b15zdnd11an1n08x5 FILLER_157_1445 ();
 b15zdnd00an1n02x5 FILLER_157_1453 ();
 b15zdnd00an1n01x5 FILLER_157_1455 ();
 b15zdnd11an1n04x5 FILLER_157_1460 ();
 b15zdnd11an1n08x5 FILLER_157_1496 ();
 b15zdnd00an1n02x5 FILLER_157_1504 ();
 b15zdnd11an1n04x5 FILLER_157_1522 ();
 b15zdnd11an1n64x5 FILLER_157_1557 ();
 b15zdnd11an1n08x5 FILLER_157_1621 ();
 b15zdnd11an1n04x5 FILLER_157_1629 ();
 b15zdnd00an1n01x5 FILLER_157_1633 ();
 b15zdnd11an1n04x5 FILLER_157_1654 ();
 b15zdnd11an1n64x5 FILLER_157_1663 ();
 b15zdnd11an1n32x5 FILLER_157_1727 ();
 b15zdnd11an1n04x5 FILLER_157_1759 ();
 b15zdnd11an1n64x5 FILLER_157_1789 ();
 b15zdnd11an1n64x5 FILLER_157_1853 ();
 b15zdnd11an1n16x5 FILLER_157_1917 ();
 b15zdnd11an1n08x5 FILLER_157_1933 ();
 b15zdnd00an1n02x5 FILLER_157_1941 ();
 b15zdnd00an1n01x5 FILLER_157_1943 ();
 b15zdnd11an1n16x5 FILLER_157_2001 ();
 b15zdnd00an1n02x5 FILLER_157_2017 ();
 b15zdnd11an1n32x5 FILLER_157_2050 ();
 b15zdnd11an1n08x5 FILLER_157_2082 ();
 b15zdnd11an1n04x5 FILLER_157_2090 ();
 b15zdnd00an1n02x5 FILLER_157_2094 ();
 b15zdnd00an1n01x5 FILLER_157_2096 ();
 b15zdnd11an1n16x5 FILLER_157_2119 ();
 b15zdnd11an1n08x5 FILLER_157_2135 ();
 b15zdnd11an1n16x5 FILLER_157_2149 ();
 b15zdnd11an1n08x5 FILLER_157_2165 ();
 b15zdnd11an1n04x5 FILLER_157_2173 ();
 b15zdnd11an1n64x5 FILLER_157_2182 ();
 b15zdnd11an1n32x5 FILLER_157_2246 ();
 b15zdnd11an1n04x5 FILLER_157_2278 ();
 b15zdnd00an1n02x5 FILLER_157_2282 ();
 b15zdnd11an1n64x5 FILLER_158_8 ();
 b15zdnd11an1n64x5 FILLER_158_72 ();
 b15zdnd11an1n08x5 FILLER_158_136 ();
 b15zdnd11an1n04x5 FILLER_158_144 ();
 b15zdnd11an1n16x5 FILLER_158_155 ();
 b15zdnd11an1n04x5 FILLER_158_171 ();
 b15zdnd11an1n08x5 FILLER_158_180 ();
 b15zdnd11an1n04x5 FILLER_158_188 ();
 b15zdnd11an1n32x5 FILLER_158_196 ();
 b15zdnd11an1n04x5 FILLER_158_228 ();
 b15zdnd00an1n02x5 FILLER_158_232 ();
 b15zdnd00an1n01x5 FILLER_158_234 ();
 b15zdnd11an1n16x5 FILLER_158_240 ();
 b15zdnd11an1n08x5 FILLER_158_256 ();
 b15zdnd11an1n04x5 FILLER_158_264 ();
 b15zdnd00an1n01x5 FILLER_158_268 ();
 b15zdnd11an1n16x5 FILLER_158_276 ();
 b15zdnd11an1n08x5 FILLER_158_292 ();
 b15zdnd11an1n04x5 FILLER_158_300 ();
 b15zdnd00an1n02x5 FILLER_158_304 ();
 b15zdnd00an1n01x5 FILLER_158_306 ();
 b15zdnd11an1n64x5 FILLER_158_326 ();
 b15zdnd11an1n08x5 FILLER_158_390 ();
 b15zdnd11an1n04x5 FILLER_158_398 ();
 b15zdnd00an1n02x5 FILLER_158_402 ();
 b15zdnd11an1n04x5 FILLER_158_410 ();
 b15zdnd11an1n16x5 FILLER_158_422 ();
 b15zdnd11an1n08x5 FILLER_158_438 ();
 b15zdnd00an1n01x5 FILLER_158_446 ();
 b15zdnd11an1n04x5 FILLER_158_453 ();
 b15zdnd11an1n08x5 FILLER_158_465 ();
 b15zdnd00an1n02x5 FILLER_158_473 ();
 b15zdnd11an1n08x5 FILLER_158_483 ();
 b15zdnd00an1n02x5 FILLER_158_491 ();
 b15zdnd11an1n64x5 FILLER_158_500 ();
 b15zdnd11an1n16x5 FILLER_158_564 ();
 b15zdnd11an1n04x5 FILLER_158_580 ();
 b15zdnd00an1n02x5 FILLER_158_584 ();
 b15zdnd11an1n16x5 FILLER_158_592 ();
 b15zdnd00an1n02x5 FILLER_158_608 ();
 b15zdnd00an1n01x5 FILLER_158_610 ();
 b15zdnd11an1n32x5 FILLER_158_615 ();
 b15zdnd11an1n04x5 FILLER_158_659 ();
 b15zdnd11an1n04x5 FILLER_158_672 ();
 b15zdnd00an1n02x5 FILLER_158_676 ();
 b15zdnd00an1n01x5 FILLER_158_678 ();
 b15zdnd11an1n08x5 FILLER_158_695 ();
 b15zdnd11an1n04x5 FILLER_158_703 ();
 b15zdnd11an1n04x5 FILLER_158_714 ();
 b15zdnd11an1n64x5 FILLER_158_726 ();
 b15zdnd11an1n64x5 FILLER_158_790 ();
 b15zdnd11an1n04x5 FILLER_158_854 ();
 b15zdnd00an1n01x5 FILLER_158_858 ();
 b15zdnd11an1n04x5 FILLER_158_882 ();
 b15zdnd11an1n04x5 FILLER_158_904 ();
 b15zdnd11an1n16x5 FILLER_158_925 ();
 b15zdnd00an1n02x5 FILLER_158_941 ();
 b15zdnd11an1n08x5 FILLER_158_974 ();
 b15zdnd11an1n04x5 FILLER_158_982 ();
 b15zdnd00an1n02x5 FILLER_158_986 ();
 b15zdnd00an1n01x5 FILLER_158_988 ();
 b15zdnd11an1n08x5 FILLER_158_995 ();
 b15zdnd11an1n04x5 FILLER_158_1003 ();
 b15zdnd00an1n01x5 FILLER_158_1007 ();
 b15zdnd11an1n04x5 FILLER_158_1015 ();
 b15zdnd11an1n08x5 FILLER_158_1025 ();
 b15zdnd11an1n04x5 FILLER_158_1033 ();
 b15zdnd00an1n02x5 FILLER_158_1037 ();
 b15zdnd11an1n04x5 FILLER_158_1045 ();
 b15zdnd11an1n64x5 FILLER_158_1059 ();
 b15zdnd11an1n08x5 FILLER_158_1123 ();
 b15zdnd11an1n04x5 FILLER_158_1131 ();
 b15zdnd00an1n02x5 FILLER_158_1135 ();
 b15zdnd00an1n01x5 FILLER_158_1137 ();
 b15zdnd11an1n04x5 FILLER_158_1143 ();
 b15zdnd00an1n02x5 FILLER_158_1147 ();
 b15zdnd00an1n01x5 FILLER_158_1149 ();
 b15zdnd11an1n04x5 FILLER_158_1156 ();
 b15zdnd11an1n16x5 FILLER_158_1176 ();
 b15zdnd00an1n02x5 FILLER_158_1192 ();
 b15zdnd00an1n01x5 FILLER_158_1194 ();
 b15zdnd11an1n16x5 FILLER_158_1212 ();
 b15zdnd11an1n04x5 FILLER_158_1228 ();
 b15zdnd00an1n02x5 FILLER_158_1232 ();
 b15zdnd11an1n64x5 FILLER_158_1256 ();
 b15zdnd11an1n64x5 FILLER_158_1320 ();
 b15zdnd11an1n08x5 FILLER_158_1384 ();
 b15zdnd00an1n01x5 FILLER_158_1392 ();
 b15zdnd11an1n04x5 FILLER_158_1409 ();
 b15zdnd00an1n02x5 FILLER_158_1413 ();
 b15zdnd00an1n01x5 FILLER_158_1415 ();
 b15zdnd11an1n16x5 FILLER_158_1436 ();
 b15zdnd11an1n08x5 FILLER_158_1452 ();
 b15zdnd11an1n04x5 FILLER_158_1466 ();
 b15zdnd11an1n64x5 FILLER_158_1475 ();
 b15zdnd11an1n64x5 FILLER_158_1539 ();
 b15zdnd11an1n64x5 FILLER_158_1603 ();
 b15zdnd11an1n64x5 FILLER_158_1667 ();
 b15zdnd11an1n64x5 FILLER_158_1731 ();
 b15zdnd11an1n08x5 FILLER_158_1795 ();
 b15zdnd00an1n01x5 FILLER_158_1803 ();
 b15zdnd11an1n32x5 FILLER_158_1808 ();
 b15zdnd11an1n16x5 FILLER_158_1840 ();
 b15zdnd11an1n08x5 FILLER_158_1856 ();
 b15zdnd11an1n04x5 FILLER_158_1864 ();
 b15zdnd00an1n02x5 FILLER_158_1868 ();
 b15zdnd00an1n01x5 FILLER_158_1870 ();
 b15zdnd11an1n04x5 FILLER_158_1876 ();
 b15zdnd11an1n64x5 FILLER_158_1900 ();
 b15zdnd11an1n64x5 FILLER_158_1964 ();
 b15zdnd11an1n32x5 FILLER_158_2028 ();
 b15zdnd11an1n04x5 FILLER_158_2060 ();
 b15zdnd00an1n01x5 FILLER_158_2064 ();
 b15zdnd11an1n16x5 FILLER_158_2083 ();
 b15zdnd11an1n04x5 FILLER_158_2099 ();
 b15zdnd00an1n01x5 FILLER_158_2103 ();
 b15zdnd11an1n16x5 FILLER_158_2135 ();
 b15zdnd00an1n02x5 FILLER_158_2151 ();
 b15zdnd00an1n01x5 FILLER_158_2153 ();
 b15zdnd11an1n08x5 FILLER_158_2162 ();
 b15zdnd00an1n02x5 FILLER_158_2170 ();
 b15zdnd11an1n32x5 FILLER_158_2192 ();
 b15zdnd11an1n16x5 FILLER_158_2224 ();
 b15zdnd11an1n04x5 FILLER_158_2240 ();
 b15zdnd00an1n02x5 FILLER_158_2244 ();
 b15zdnd11an1n16x5 FILLER_158_2250 ();
 b15zdnd11an1n04x5 FILLER_158_2266 ();
 b15zdnd00an1n02x5 FILLER_158_2274 ();
 b15zdnd11an1n32x5 FILLER_159_0 ();
 b15zdnd11an1n16x5 FILLER_159_32 ();
 b15zdnd11an1n04x5 FILLER_159_48 ();
 b15zdnd00an1n01x5 FILLER_159_52 ();
 b15zdnd11an1n64x5 FILLER_159_59 ();
 b15zdnd11an1n32x5 FILLER_159_123 ();
 b15zdnd11an1n04x5 FILLER_159_155 ();
 b15zdnd11an1n08x5 FILLER_159_168 ();
 b15zdnd11an1n04x5 FILLER_159_176 ();
 b15zdnd00an1n01x5 FILLER_159_180 ();
 b15zdnd11an1n08x5 FILLER_159_187 ();
 b15zdnd00an1n01x5 FILLER_159_195 ();
 b15zdnd11an1n32x5 FILLER_159_206 ();
 b15zdnd11an1n16x5 FILLER_159_238 ();
 b15zdnd11an1n08x5 FILLER_159_254 ();
 b15zdnd11an1n04x5 FILLER_159_262 ();
 b15zdnd11an1n64x5 FILLER_159_273 ();
 b15zdnd11an1n64x5 FILLER_159_337 ();
 b15zdnd11an1n64x5 FILLER_159_401 ();
 b15zdnd11an1n08x5 FILLER_159_474 ();
 b15zdnd11an1n04x5 FILLER_159_482 ();
 b15zdnd00an1n01x5 FILLER_159_486 ();
 b15zdnd11an1n04x5 FILLER_159_496 ();
 b15zdnd11an1n32x5 FILLER_159_514 ();
 b15zdnd11an1n16x5 FILLER_159_546 ();
 b15zdnd11an1n64x5 FILLER_159_567 ();
 b15zdnd11an1n32x5 FILLER_159_631 ();
 b15zdnd11an1n04x5 FILLER_159_663 ();
 b15zdnd00an1n02x5 FILLER_159_667 ();
 b15zdnd00an1n01x5 FILLER_159_669 ();
 b15zdnd11an1n64x5 FILLER_159_682 ();
 b15zdnd11an1n64x5 FILLER_159_746 ();
 b15zdnd11an1n64x5 FILLER_159_810 ();
 b15zdnd11an1n64x5 FILLER_159_874 ();
 b15zdnd00an1n02x5 FILLER_159_938 ();
 b15zdnd11an1n04x5 FILLER_159_952 ();
 b15zdnd00an1n02x5 FILLER_159_956 ();
 b15zdnd11an1n08x5 FILLER_159_976 ();
 b15zdnd00an1n02x5 FILLER_159_984 ();
 b15zdnd11an1n08x5 FILLER_159_991 ();
 b15zdnd11an1n04x5 FILLER_159_999 ();
 b15zdnd00an1n02x5 FILLER_159_1003 ();
 b15zdnd00an1n01x5 FILLER_159_1005 ();
 b15zdnd11an1n64x5 FILLER_159_1012 ();
 b15zdnd11an1n64x5 FILLER_159_1076 ();
 b15zdnd11an1n16x5 FILLER_159_1140 ();
 b15zdnd11an1n04x5 FILLER_159_1156 ();
 b15zdnd00an1n02x5 FILLER_159_1160 ();
 b15zdnd11an1n04x5 FILLER_159_1170 ();
 b15zdnd11an1n64x5 FILLER_159_1194 ();
 b15zdnd11an1n16x5 FILLER_159_1258 ();
 b15zdnd11an1n08x5 FILLER_159_1274 ();
 b15zdnd00an1n02x5 FILLER_159_1282 ();
 b15zdnd00an1n01x5 FILLER_159_1284 ();
 b15zdnd11an1n64x5 FILLER_159_1305 ();
 b15zdnd11an1n64x5 FILLER_159_1369 ();
 b15zdnd11an1n64x5 FILLER_159_1433 ();
 b15zdnd11an1n64x5 FILLER_159_1497 ();
 b15zdnd11an1n32x5 FILLER_159_1561 ();
 b15zdnd11an1n16x5 FILLER_159_1593 ();
 b15zdnd11an1n64x5 FILLER_159_1629 ();
 b15zdnd11an1n16x5 FILLER_159_1693 ();
 b15zdnd11an1n08x5 FILLER_159_1709 ();
 b15zdnd11an1n04x5 FILLER_159_1717 ();
 b15zdnd00an1n01x5 FILLER_159_1721 ();
 b15zdnd11an1n32x5 FILLER_159_1742 ();
 b15zdnd11an1n08x5 FILLER_159_1774 ();
 b15zdnd11an1n04x5 FILLER_159_1782 ();
 b15zdnd11an1n16x5 FILLER_159_1817 ();
 b15zdnd00an1n01x5 FILLER_159_1833 ();
 b15zdnd11an1n08x5 FILLER_159_1865 ();
 b15zdnd11an1n04x5 FILLER_159_1873 ();
 b15zdnd11an1n64x5 FILLER_159_1895 ();
 b15zdnd11an1n64x5 FILLER_159_1959 ();
 b15zdnd11an1n32x5 FILLER_159_2023 ();
 b15zdnd11an1n08x5 FILLER_159_2055 ();
 b15zdnd11an1n04x5 FILLER_159_2063 ();
 b15zdnd00an1n01x5 FILLER_159_2067 ();
 b15zdnd11an1n32x5 FILLER_159_2086 ();
 b15zdnd11an1n04x5 FILLER_159_2118 ();
 b15zdnd00an1n01x5 FILLER_159_2122 ();
 b15zdnd11an1n08x5 FILLER_159_2133 ();
 b15zdnd11an1n04x5 FILLER_159_2141 ();
 b15zdnd11an1n08x5 FILLER_159_2164 ();
 b15zdnd11an1n04x5 FILLER_159_2172 ();
 b15zdnd00an1n02x5 FILLER_159_2176 ();
 b15zdnd11an1n16x5 FILLER_159_2181 ();
 b15zdnd11an1n08x5 FILLER_159_2197 ();
 b15zdnd11an1n04x5 FILLER_159_2205 ();
 b15zdnd00an1n02x5 FILLER_159_2209 ();
 b15zdnd00an1n01x5 FILLER_159_2211 ();
 b15zdnd11an1n04x5 FILLER_159_2232 ();
 b15zdnd11an1n04x5 FILLER_159_2256 ();
 b15zdnd11an1n04x5 FILLER_159_2264 ();
 b15zdnd00an1n01x5 FILLER_159_2268 ();
 b15zdnd11an1n04x5 FILLER_159_2273 ();
 b15zdnd00an1n01x5 FILLER_159_2277 ();
 b15zdnd00an1n02x5 FILLER_159_2282 ();
 b15zdnd11an1n64x5 FILLER_160_8 ();
 b15zdnd11an1n16x5 FILLER_160_72 ();
 b15zdnd11an1n08x5 FILLER_160_88 ();
 b15zdnd11an1n32x5 FILLER_160_102 ();
 b15zdnd11an1n16x5 FILLER_160_134 ();
 b15zdnd00an1n02x5 FILLER_160_150 ();
 b15zdnd11an1n16x5 FILLER_160_156 ();
 b15zdnd00an1n01x5 FILLER_160_172 ();
 b15zdnd11an1n16x5 FILLER_160_177 ();
 b15zdnd11an1n08x5 FILLER_160_193 ();
 b15zdnd00an1n01x5 FILLER_160_201 ();
 b15zdnd11an1n16x5 FILLER_160_209 ();
 b15zdnd11an1n08x5 FILLER_160_225 ();
 b15zdnd00an1n01x5 FILLER_160_233 ();
 b15zdnd11an1n16x5 FILLER_160_241 ();
 b15zdnd11an1n04x5 FILLER_160_257 ();
 b15zdnd00an1n01x5 FILLER_160_261 ();
 b15zdnd11an1n04x5 FILLER_160_269 ();
 b15zdnd11an1n64x5 FILLER_160_284 ();
 b15zdnd11an1n64x5 FILLER_160_348 ();
 b15zdnd11an1n64x5 FILLER_160_412 ();
 b15zdnd00an1n01x5 FILLER_160_476 ();
 b15zdnd11an1n04x5 FILLER_160_495 ();
 b15zdnd11an1n04x5 FILLER_160_513 ();
 b15zdnd00an1n02x5 FILLER_160_517 ();
 b15zdnd11an1n64x5 FILLER_160_529 ();
 b15zdnd11an1n04x5 FILLER_160_593 ();
 b15zdnd00an1n02x5 FILLER_160_597 ();
 b15zdnd00an1n01x5 FILLER_160_599 ();
 b15zdnd11an1n08x5 FILLER_160_604 ();
 b15zdnd11an1n04x5 FILLER_160_612 ();
 b15zdnd00an1n02x5 FILLER_160_616 ();
 b15zdnd11an1n16x5 FILLER_160_622 ();
 b15zdnd00an1n02x5 FILLER_160_638 ();
 b15zdnd11an1n64x5 FILLER_160_650 ();
 b15zdnd11an1n04x5 FILLER_160_714 ();
 b15zdnd11an1n32x5 FILLER_160_726 ();
 b15zdnd00an1n02x5 FILLER_160_758 ();
 b15zdnd00an1n01x5 FILLER_160_760 ();
 b15zdnd11an1n64x5 FILLER_160_769 ();
 b15zdnd11an1n04x5 FILLER_160_833 ();
 b15zdnd00an1n01x5 FILLER_160_837 ();
 b15zdnd11an1n16x5 FILLER_160_858 ();
 b15zdnd11an1n08x5 FILLER_160_874 ();
 b15zdnd11an1n08x5 FILLER_160_900 ();
 b15zdnd11an1n32x5 FILLER_160_913 ();
 b15zdnd11an1n08x5 FILLER_160_945 ();
 b15zdnd00an1n02x5 FILLER_160_953 ();
 b15zdnd00an1n01x5 FILLER_160_955 ();
 b15zdnd11an1n08x5 FILLER_160_965 ();
 b15zdnd11an1n04x5 FILLER_160_973 ();
 b15zdnd00an1n01x5 FILLER_160_977 ();
 b15zdnd11an1n04x5 FILLER_160_987 ();
 b15zdnd11an1n16x5 FILLER_160_997 ();
 b15zdnd11an1n04x5 FILLER_160_1013 ();
 b15zdnd00an1n02x5 FILLER_160_1017 ();
 b15zdnd11an1n32x5 FILLER_160_1025 ();
 b15zdnd11an1n16x5 FILLER_160_1057 ();
 b15zdnd11an1n08x5 FILLER_160_1073 ();
 b15zdnd00an1n01x5 FILLER_160_1081 ();
 b15zdnd11an1n32x5 FILLER_160_1088 ();
 b15zdnd11an1n08x5 FILLER_160_1120 ();
 b15zdnd00an1n02x5 FILLER_160_1128 ();
 b15zdnd11an1n64x5 FILLER_160_1135 ();
 b15zdnd11an1n16x5 FILLER_160_1199 ();
 b15zdnd11an1n64x5 FILLER_160_1229 ();
 b15zdnd11an1n64x5 FILLER_160_1293 ();
 b15zdnd11an1n64x5 FILLER_160_1357 ();
 b15zdnd11an1n64x5 FILLER_160_1421 ();
 b15zdnd11an1n64x5 FILLER_160_1485 ();
 b15zdnd11an1n04x5 FILLER_160_1549 ();
 b15zdnd00an1n01x5 FILLER_160_1553 ();
 b15zdnd11an1n04x5 FILLER_160_1573 ();
 b15zdnd11an1n04x5 FILLER_160_1608 ();
 b15zdnd11an1n32x5 FILLER_160_1621 ();
 b15zdnd11an1n16x5 FILLER_160_1653 ();
 b15zdnd00an1n02x5 FILLER_160_1669 ();
 b15zdnd11an1n16x5 FILLER_160_1691 ();
 b15zdnd00an1n02x5 FILLER_160_1707 ();
 b15zdnd11an1n16x5 FILLER_160_1729 ();
 b15zdnd00an1n02x5 FILLER_160_1745 ();
 b15zdnd00an1n01x5 FILLER_160_1747 ();
 b15zdnd11an1n16x5 FILLER_160_1757 ();
 b15zdnd11an1n64x5 FILLER_160_1788 ();
 b15zdnd11an1n32x5 FILLER_160_1852 ();
 b15zdnd11an1n04x5 FILLER_160_1884 ();
 b15zdnd00an1n02x5 FILLER_160_1888 ();
 b15zdnd00an1n01x5 FILLER_160_1890 ();
 b15zdnd11an1n04x5 FILLER_160_1922 ();
 b15zdnd00an1n01x5 FILLER_160_1926 ();
 b15zdnd11an1n16x5 FILLER_160_1947 ();
 b15zdnd11an1n08x5 FILLER_160_1963 ();
 b15zdnd11an1n04x5 FILLER_160_1971 ();
 b15zdnd00an1n02x5 FILLER_160_1975 ();
 b15zdnd00an1n01x5 FILLER_160_1977 ();
 b15zdnd11an1n16x5 FILLER_160_1989 ();
 b15zdnd11an1n04x5 FILLER_160_2005 ();
 b15zdnd11an1n16x5 FILLER_160_2021 ();
 b15zdnd00an1n02x5 FILLER_160_2037 ();
 b15zdnd11an1n64x5 FILLER_160_2070 ();
 b15zdnd11an1n16x5 FILLER_160_2134 ();
 b15zdnd11an1n04x5 FILLER_160_2150 ();
 b15zdnd11an1n64x5 FILLER_160_2162 ();
 b15zdnd11an1n16x5 FILLER_160_2226 ();
 b15zdnd11an1n08x5 FILLER_160_2242 ();
 b15zdnd00an1n02x5 FILLER_160_2250 ();
 b15zdnd00an1n01x5 FILLER_160_2252 ();
 b15zdnd11an1n04x5 FILLER_160_2257 ();
 b15zdnd11an1n04x5 FILLER_160_2265 ();
 b15zdnd00an1n02x5 FILLER_160_2273 ();
 b15zdnd00an1n01x5 FILLER_160_2275 ();
 b15zdnd11an1n64x5 FILLER_161_0 ();
 b15zdnd11an1n32x5 FILLER_161_64 ();
 b15zdnd11an1n08x5 FILLER_161_105 ();
 b15zdnd11an1n04x5 FILLER_161_113 ();
 b15zdnd00an1n02x5 FILLER_161_117 ();
 b15zdnd11an1n04x5 FILLER_161_128 ();
 b15zdnd00an1n02x5 FILLER_161_132 ();
 b15zdnd11an1n32x5 FILLER_161_139 ();
 b15zdnd00an1n01x5 FILLER_161_171 ();
 b15zdnd11an1n16x5 FILLER_161_179 ();
 b15zdnd11an1n04x5 FILLER_161_195 ();
 b15zdnd11an1n08x5 FILLER_161_206 ();
 b15zdnd00an1n01x5 FILLER_161_214 ();
 b15zdnd11an1n32x5 FILLER_161_235 ();
 b15zdnd11an1n16x5 FILLER_161_267 ();
 b15zdnd00an1n02x5 FILLER_161_283 ();
 b15zdnd00an1n01x5 FILLER_161_285 ();
 b15zdnd11an1n04x5 FILLER_161_292 ();
 b15zdnd11an1n04x5 FILLER_161_302 ();
 b15zdnd00an1n02x5 FILLER_161_306 ();
 b15zdnd00an1n01x5 FILLER_161_308 ();
 b15zdnd11an1n16x5 FILLER_161_314 ();
 b15zdnd00an1n01x5 FILLER_161_330 ();
 b15zdnd11an1n32x5 FILLER_161_351 ();
 b15zdnd11an1n16x5 FILLER_161_383 ();
 b15zdnd11an1n08x5 FILLER_161_399 ();
 b15zdnd00an1n02x5 FILLER_161_407 ();
 b15zdnd11an1n64x5 FILLER_161_432 ();
 b15zdnd00an1n01x5 FILLER_161_496 ();
 b15zdnd11an1n04x5 FILLER_161_512 ();
 b15zdnd11an1n32x5 FILLER_161_523 ();
 b15zdnd11an1n08x5 FILLER_161_555 ();
 b15zdnd11an1n04x5 FILLER_161_563 ();
 b15zdnd00an1n02x5 FILLER_161_567 ();
 b15zdnd11an1n16x5 FILLER_161_573 ();
 b15zdnd11an1n04x5 FILLER_161_589 ();
 b15zdnd00an1n01x5 FILLER_161_593 ();
 b15zdnd11an1n08x5 FILLER_161_599 ();
 b15zdnd11an1n64x5 FILLER_161_613 ();
 b15zdnd11an1n04x5 FILLER_161_677 ();
 b15zdnd00an1n02x5 FILLER_161_681 ();
 b15zdnd00an1n01x5 FILLER_161_683 ();
 b15zdnd11an1n32x5 FILLER_161_691 ();
 b15zdnd11an1n08x5 FILLER_161_723 ();
 b15zdnd11an1n04x5 FILLER_161_731 ();
 b15zdnd11an1n04x5 FILLER_161_742 ();
 b15zdnd11an1n04x5 FILLER_161_752 ();
 b15zdnd11an1n64x5 FILLER_161_764 ();
 b15zdnd11an1n64x5 FILLER_161_828 ();
 b15zdnd11an1n08x5 FILLER_161_892 ();
 b15zdnd11an1n04x5 FILLER_161_900 ();
 b15zdnd11an1n16x5 FILLER_161_916 ();
 b15zdnd11an1n08x5 FILLER_161_932 ();
 b15zdnd11an1n04x5 FILLER_161_940 ();
 b15zdnd00an1n02x5 FILLER_161_944 ();
 b15zdnd11an1n64x5 FILLER_161_953 ();
 b15zdnd11an1n16x5 FILLER_161_1017 ();
 b15zdnd11an1n04x5 FILLER_161_1033 ();
 b15zdnd00an1n02x5 FILLER_161_1037 ();
 b15zdnd11an1n16x5 FILLER_161_1050 ();
 b15zdnd11an1n04x5 FILLER_161_1066 ();
 b15zdnd11an1n16x5 FILLER_161_1083 ();
 b15zdnd00an1n02x5 FILLER_161_1099 ();
 b15zdnd11an1n08x5 FILLER_161_1107 ();
 b15zdnd11an1n04x5 FILLER_161_1115 ();
 b15zdnd00an1n02x5 FILLER_161_1119 ();
 b15zdnd11an1n04x5 FILLER_161_1130 ();
 b15zdnd11an1n32x5 FILLER_161_1141 ();
 b15zdnd11an1n16x5 FILLER_161_1173 ();
 b15zdnd11an1n04x5 FILLER_161_1189 ();
 b15zdnd11an1n64x5 FILLER_161_1207 ();
 b15zdnd11an1n16x5 FILLER_161_1271 ();
 b15zdnd00an1n02x5 FILLER_161_1287 ();
 b15zdnd00an1n01x5 FILLER_161_1289 ();
 b15zdnd11an1n16x5 FILLER_161_1310 ();
 b15zdnd11an1n08x5 FILLER_161_1326 ();
 b15zdnd11an1n04x5 FILLER_161_1334 ();
 b15zdnd11an1n64x5 FILLER_161_1369 ();
 b15zdnd11an1n64x5 FILLER_161_1433 ();
 b15zdnd11an1n64x5 FILLER_161_1497 ();
 b15zdnd11an1n32x5 FILLER_161_1561 ();
 b15zdnd11an1n16x5 FILLER_161_1593 ();
 b15zdnd00an1n01x5 FILLER_161_1609 ();
 b15zdnd11an1n08x5 FILLER_161_1619 ();
 b15zdnd11an1n04x5 FILLER_161_1627 ();
 b15zdnd00an1n02x5 FILLER_161_1631 ();
 b15zdnd00an1n01x5 FILLER_161_1633 ();
 b15zdnd11an1n04x5 FILLER_161_1665 ();
 b15zdnd11an1n04x5 FILLER_161_1674 ();
 b15zdnd11an1n64x5 FILLER_161_1709 ();
 b15zdnd11an1n04x5 FILLER_161_1773 ();
 b15zdnd00an1n02x5 FILLER_161_1777 ();
 b15zdnd00an1n01x5 FILLER_161_1779 ();
 b15zdnd11an1n64x5 FILLER_161_1800 ();
 b15zdnd11an1n32x5 FILLER_161_1864 ();
 b15zdnd11an1n04x5 FILLER_161_1896 ();
 b15zdnd00an1n02x5 FILLER_161_1900 ();
 b15zdnd11an1n16x5 FILLER_161_1906 ();
 b15zdnd11an1n04x5 FILLER_161_1922 ();
 b15zdnd11an1n64x5 FILLER_161_1931 ();
 b15zdnd11an1n16x5 FILLER_161_1995 ();
 b15zdnd11an1n04x5 FILLER_161_2011 ();
 b15zdnd00an1n02x5 FILLER_161_2015 ();
 b15zdnd11an1n04x5 FILLER_161_2021 ();
 b15zdnd11an1n64x5 FILLER_161_2046 ();
 b15zdnd11an1n16x5 FILLER_161_2110 ();
 b15zdnd11an1n04x5 FILLER_161_2126 ();
 b15zdnd11an1n64x5 FILLER_161_2135 ();
 b15zdnd11an1n16x5 FILLER_161_2199 ();
 b15zdnd11an1n08x5 FILLER_161_2215 ();
 b15zdnd11an1n04x5 FILLER_161_2223 ();
 b15zdnd00an1n02x5 FILLER_161_2227 ();
 b15zdnd11an1n16x5 FILLER_161_2233 ();
 b15zdnd11an1n04x5 FILLER_161_2249 ();
 b15zdnd00an1n01x5 FILLER_161_2253 ();
 b15zdnd11an1n04x5 FILLER_161_2258 ();
 b15zdnd11an1n08x5 FILLER_161_2266 ();
 b15zdnd11an1n04x5 FILLER_161_2278 ();
 b15zdnd00an1n02x5 FILLER_161_2282 ();
 b15zdnd11an1n32x5 FILLER_162_8 ();
 b15zdnd11an1n16x5 FILLER_162_40 ();
 b15zdnd11an1n32x5 FILLER_162_72 ();
 b15zdnd11an1n16x5 FILLER_162_104 ();
 b15zdnd00an1n01x5 FILLER_162_120 ();
 b15zdnd11an1n64x5 FILLER_162_126 ();
 b15zdnd00an1n02x5 FILLER_162_190 ();
 b15zdnd00an1n01x5 FILLER_162_192 ();
 b15zdnd11an1n64x5 FILLER_162_198 ();
 b15zdnd11an1n32x5 FILLER_162_262 ();
 b15zdnd11an1n16x5 FILLER_162_294 ();
 b15zdnd11an1n16x5 FILLER_162_324 ();
 b15zdnd00an1n02x5 FILLER_162_340 ();
 b15zdnd00an1n01x5 FILLER_162_342 ();
 b15zdnd11an1n04x5 FILLER_162_347 ();
 b15zdnd11an1n64x5 FILLER_162_361 ();
 b15zdnd11an1n16x5 FILLER_162_425 ();
 b15zdnd11an1n04x5 FILLER_162_441 ();
 b15zdnd00an1n02x5 FILLER_162_445 ();
 b15zdnd11an1n64x5 FILLER_162_459 ();
 b15zdnd11an1n08x5 FILLER_162_523 ();
 b15zdnd11an1n04x5 FILLER_162_531 ();
 b15zdnd00an1n01x5 FILLER_162_535 ();
 b15zdnd11an1n04x5 FILLER_162_560 ();
 b15zdnd11an1n08x5 FILLER_162_579 ();
 b15zdnd11an1n04x5 FILLER_162_587 ();
 b15zdnd00an1n02x5 FILLER_162_591 ();
 b15zdnd00an1n01x5 FILLER_162_593 ();
 b15zdnd11an1n04x5 FILLER_162_614 ();
 b15zdnd11an1n08x5 FILLER_162_644 ();
 b15zdnd11an1n04x5 FILLER_162_652 ();
 b15zdnd00an1n02x5 FILLER_162_656 ();
 b15zdnd11an1n16x5 FILLER_162_663 ();
 b15zdnd11an1n04x5 FILLER_162_679 ();
 b15zdnd00an1n01x5 FILLER_162_683 ();
 b15zdnd11an1n08x5 FILLER_162_694 ();
 b15zdnd00an1n02x5 FILLER_162_716 ();
 b15zdnd11an1n08x5 FILLER_162_726 ();
 b15zdnd00an1n02x5 FILLER_162_734 ();
 b15zdnd00an1n01x5 FILLER_162_736 ();
 b15zdnd11an1n32x5 FILLER_162_745 ();
 b15zdnd00an1n02x5 FILLER_162_777 ();
 b15zdnd00an1n01x5 FILLER_162_779 ();
 b15zdnd11an1n04x5 FILLER_162_800 ();
 b15zdnd11an1n16x5 FILLER_162_828 ();
 b15zdnd11an1n08x5 FILLER_162_844 ();
 b15zdnd11an1n04x5 FILLER_162_852 ();
 b15zdnd00an1n02x5 FILLER_162_856 ();
 b15zdnd00an1n01x5 FILLER_162_858 ();
 b15zdnd11an1n08x5 FILLER_162_877 ();
 b15zdnd11an1n04x5 FILLER_162_885 ();
 b15zdnd00an1n02x5 FILLER_162_889 ();
 b15zdnd11an1n16x5 FILLER_162_914 ();
 b15zdnd11an1n04x5 FILLER_162_930 ();
 b15zdnd00an1n02x5 FILLER_162_934 ();
 b15zdnd11an1n64x5 FILLER_162_960 ();
 b15zdnd11an1n64x5 FILLER_162_1024 ();
 b15zdnd11an1n16x5 FILLER_162_1088 ();
 b15zdnd11an1n08x5 FILLER_162_1104 ();
 b15zdnd11an1n04x5 FILLER_162_1112 ();
 b15zdnd00an1n01x5 FILLER_162_1116 ();
 b15zdnd11an1n16x5 FILLER_162_1129 ();
 b15zdnd11an1n08x5 FILLER_162_1145 ();
 b15zdnd11an1n04x5 FILLER_162_1153 ();
 b15zdnd00an1n01x5 FILLER_162_1157 ();
 b15zdnd11an1n16x5 FILLER_162_1163 ();
 b15zdnd11an1n08x5 FILLER_162_1179 ();
 b15zdnd11an1n04x5 FILLER_162_1187 ();
 b15zdnd00an1n02x5 FILLER_162_1191 ();
 b15zdnd00an1n01x5 FILLER_162_1193 ();
 b15zdnd11an1n64x5 FILLER_162_1210 ();
 b15zdnd11an1n16x5 FILLER_162_1274 ();
 b15zdnd00an1n01x5 FILLER_162_1290 ();
 b15zdnd11an1n32x5 FILLER_162_1295 ();
 b15zdnd11an1n16x5 FILLER_162_1327 ();
 b15zdnd11an1n04x5 FILLER_162_1343 ();
 b15zdnd00an1n02x5 FILLER_162_1347 ();
 b15zdnd11an1n64x5 FILLER_162_1375 ();
 b15zdnd11an1n64x5 FILLER_162_1439 ();
 b15zdnd11an1n04x5 FILLER_162_1503 ();
 b15zdnd11an1n08x5 FILLER_162_1514 ();
 b15zdnd11an1n16x5 FILLER_162_1526 ();
 b15zdnd11an1n04x5 FILLER_162_1542 ();
 b15zdnd00an1n02x5 FILLER_162_1546 ();
 b15zdnd00an1n01x5 FILLER_162_1548 ();
 b15zdnd11an1n64x5 FILLER_162_1553 ();
 b15zdnd11an1n64x5 FILLER_162_1617 ();
 b15zdnd11an1n64x5 FILLER_162_1681 ();
 b15zdnd11an1n64x5 FILLER_162_1745 ();
 b15zdnd11an1n32x5 FILLER_162_1809 ();
 b15zdnd11an1n08x5 FILLER_162_1841 ();
 b15zdnd00an1n02x5 FILLER_162_1849 ();
 b15zdnd11an1n64x5 FILLER_162_1871 ();
 b15zdnd11an1n08x5 FILLER_162_1935 ();
 b15zdnd11an1n64x5 FILLER_162_1969 ();
 b15zdnd11an1n08x5 FILLER_162_2033 ();
 b15zdnd11an1n04x5 FILLER_162_2041 ();
 b15zdnd00an1n02x5 FILLER_162_2045 ();
 b15zdnd00an1n01x5 FILLER_162_2047 ();
 b15zdnd11an1n32x5 FILLER_162_2080 ();
 b15zdnd11an1n08x5 FILLER_162_2112 ();
 b15zdnd00an1n01x5 FILLER_162_2120 ();
 b15zdnd11an1n16x5 FILLER_162_2131 ();
 b15zdnd11an1n04x5 FILLER_162_2147 ();
 b15zdnd00an1n02x5 FILLER_162_2151 ();
 b15zdnd00an1n01x5 FILLER_162_2153 ();
 b15zdnd11an1n16x5 FILLER_162_2162 ();
 b15zdnd11an1n08x5 FILLER_162_2178 ();
 b15zdnd11an1n04x5 FILLER_162_2186 ();
 b15zdnd11an1n04x5 FILLER_162_2194 ();
 b15zdnd11an1n64x5 FILLER_162_2203 ();
 b15zdnd00an1n02x5 FILLER_162_2267 ();
 b15zdnd00an1n01x5 FILLER_162_2269 ();
 b15zdnd00an1n02x5 FILLER_162_2274 ();
 b15zdnd11an1n32x5 FILLER_163_0 ();
 b15zdnd11an1n04x5 FILLER_163_32 ();
 b15zdnd11an1n04x5 FILLER_163_43 ();
 b15zdnd11an1n04x5 FILLER_163_53 ();
 b15zdnd11an1n16x5 FILLER_163_67 ();
 b15zdnd11an1n08x5 FILLER_163_83 ();
 b15zdnd00an1n01x5 FILLER_163_91 ();
 b15zdnd11an1n32x5 FILLER_163_99 ();
 b15zdnd11an1n16x5 FILLER_163_131 ();
 b15zdnd00an1n02x5 FILLER_163_147 ();
 b15zdnd00an1n01x5 FILLER_163_149 ();
 b15zdnd11an1n64x5 FILLER_163_169 ();
 b15zdnd11an1n08x5 FILLER_163_233 ();
 b15zdnd11an1n04x5 FILLER_163_241 ();
 b15zdnd11an1n32x5 FILLER_163_253 ();
 b15zdnd00an1n02x5 FILLER_163_285 ();
 b15zdnd00an1n01x5 FILLER_163_287 ();
 b15zdnd11an1n04x5 FILLER_163_293 ();
 b15zdnd11an1n08x5 FILLER_163_303 ();
 b15zdnd11an1n04x5 FILLER_163_311 ();
 b15zdnd00an1n01x5 FILLER_163_315 ();
 b15zdnd11an1n04x5 FILLER_163_327 ();
 b15zdnd11an1n08x5 FILLER_163_337 ();
 b15zdnd00an1n02x5 FILLER_163_345 ();
 b15zdnd00an1n01x5 FILLER_163_347 ();
 b15zdnd11an1n32x5 FILLER_163_360 ();
 b15zdnd11an1n16x5 FILLER_163_392 ();
 b15zdnd00an1n02x5 FILLER_163_408 ();
 b15zdnd11an1n64x5 FILLER_163_417 ();
 b15zdnd11an1n64x5 FILLER_163_481 ();
 b15zdnd11an1n32x5 FILLER_163_545 ();
 b15zdnd11an1n16x5 FILLER_163_577 ();
 b15zdnd00an1n02x5 FILLER_163_593 ();
 b15zdnd11an1n04x5 FILLER_163_605 ();
 b15zdnd11an1n32x5 FILLER_163_613 ();
 b15zdnd11an1n08x5 FILLER_163_645 ();
 b15zdnd11an1n04x5 FILLER_163_653 ();
 b15zdnd00an1n01x5 FILLER_163_657 ();
 b15zdnd11an1n32x5 FILLER_163_664 ();
 b15zdnd11an1n16x5 FILLER_163_696 ();
 b15zdnd11an1n08x5 FILLER_163_712 ();
 b15zdnd11an1n04x5 FILLER_163_720 ();
 b15zdnd00an1n02x5 FILLER_163_724 ();
 b15zdnd11an1n32x5 FILLER_163_730 ();
 b15zdnd11an1n04x5 FILLER_163_762 ();
 b15zdnd00an1n01x5 FILLER_163_766 ();
 b15zdnd11an1n32x5 FILLER_163_785 ();
 b15zdnd00an1n02x5 FILLER_163_817 ();
 b15zdnd00an1n01x5 FILLER_163_819 ();
 b15zdnd11an1n32x5 FILLER_163_825 ();
 b15zdnd11an1n08x5 FILLER_163_857 ();
 b15zdnd00an1n01x5 FILLER_163_865 ();
 b15zdnd11an1n08x5 FILLER_163_871 ();
 b15zdnd11an1n04x5 FILLER_163_879 ();
 b15zdnd00an1n02x5 FILLER_163_883 ();
 b15zdnd11an1n08x5 FILLER_163_890 ();
 b15zdnd11an1n04x5 FILLER_163_898 ();
 b15zdnd00an1n01x5 FILLER_163_902 ();
 b15zdnd11an1n16x5 FILLER_163_917 ();
 b15zdnd11an1n04x5 FILLER_163_933 ();
 b15zdnd00an1n01x5 FILLER_163_937 ();
 b15zdnd11an1n16x5 FILLER_163_950 ();
 b15zdnd11an1n08x5 FILLER_163_966 ();
 b15zdnd00an1n02x5 FILLER_163_974 ();
 b15zdnd11an1n08x5 FILLER_163_997 ();
 b15zdnd00an1n02x5 FILLER_163_1005 ();
 b15zdnd00an1n01x5 FILLER_163_1007 ();
 b15zdnd11an1n04x5 FILLER_163_1022 ();
 b15zdnd11an1n08x5 FILLER_163_1038 ();
 b15zdnd11an1n04x5 FILLER_163_1052 ();
 b15zdnd00an1n02x5 FILLER_163_1056 ();
 b15zdnd00an1n01x5 FILLER_163_1058 ();
 b15zdnd11an1n32x5 FILLER_163_1064 ();
 b15zdnd11an1n04x5 FILLER_163_1096 ();
 b15zdnd00an1n02x5 FILLER_163_1100 ();
 b15zdnd00an1n01x5 FILLER_163_1102 ();
 b15zdnd11an1n16x5 FILLER_163_1113 ();
 b15zdnd11an1n08x5 FILLER_163_1129 ();
 b15zdnd11an1n08x5 FILLER_163_1143 ();
 b15zdnd11an1n04x5 FILLER_163_1151 ();
 b15zdnd00an1n02x5 FILLER_163_1155 ();
 b15zdnd11an1n32x5 FILLER_163_1164 ();
 b15zdnd11an1n04x5 FILLER_163_1206 ();
 b15zdnd11an1n32x5 FILLER_163_1228 ();
 b15zdnd00an1n02x5 FILLER_163_1260 ();
 b15zdnd00an1n01x5 FILLER_163_1262 ();
 b15zdnd11an1n04x5 FILLER_163_1283 ();
 b15zdnd11an1n08x5 FILLER_163_1292 ();
 b15zdnd00an1n02x5 FILLER_163_1300 ();
 b15zdnd11an1n04x5 FILLER_163_1322 ();
 b15zdnd11an1n08x5 FILLER_163_1344 ();
 b15zdnd11an1n32x5 FILLER_163_1364 ();
 b15zdnd11an1n16x5 FILLER_163_1396 ();
 b15zdnd11an1n04x5 FILLER_163_1412 ();
 b15zdnd11an1n08x5 FILLER_163_1447 ();
 b15zdnd11an1n04x5 FILLER_163_1455 ();
 b15zdnd00an1n02x5 FILLER_163_1459 ();
 b15zdnd11an1n04x5 FILLER_163_1482 ();
 b15zdnd11an1n04x5 FILLER_163_1511 ();
 b15zdnd11an1n16x5 FILLER_163_1520 ();
 b15zdnd11an1n08x5 FILLER_163_1536 ();
 b15zdnd00an1n01x5 FILLER_163_1544 ();
 b15zdnd11an1n04x5 FILLER_163_1550 ();
 b15zdnd11an1n32x5 FILLER_163_1559 ();
 b15zdnd11an1n08x5 FILLER_163_1591 ();
 b15zdnd11an1n04x5 FILLER_163_1599 ();
 b15zdnd00an1n02x5 FILLER_163_1603 ();
 b15zdnd00an1n01x5 FILLER_163_1605 ();
 b15zdnd11an1n64x5 FILLER_163_1617 ();
 b15zdnd11an1n32x5 FILLER_163_1681 ();
 b15zdnd00an1n01x5 FILLER_163_1713 ();
 b15zdnd11an1n64x5 FILLER_163_1739 ();
 b15zdnd11an1n64x5 FILLER_163_1803 ();
 b15zdnd11an1n16x5 FILLER_163_1867 ();
 b15zdnd11an1n08x5 FILLER_163_1883 ();
 b15zdnd11an1n04x5 FILLER_163_1891 ();
 b15zdnd00an1n01x5 FILLER_163_1895 ();
 b15zdnd11an1n04x5 FILLER_163_1916 ();
 b15zdnd00an1n02x5 FILLER_163_1920 ();
 b15zdnd11an1n64x5 FILLER_163_1953 ();
 b15zdnd11an1n64x5 FILLER_163_2017 ();
 b15zdnd11an1n16x5 FILLER_163_2081 ();
 b15zdnd11an1n04x5 FILLER_163_2097 ();
 b15zdnd00an1n01x5 FILLER_163_2101 ();
 b15zdnd11an1n32x5 FILLER_163_2133 ();
 b15zdnd11an1n16x5 FILLER_163_2165 ();
 b15zdnd11an1n08x5 FILLER_163_2181 ();
 b15zdnd00an1n01x5 FILLER_163_2189 ();
 b15zdnd11an1n04x5 FILLER_163_2194 ();
 b15zdnd11an1n08x5 FILLER_163_2218 ();
 b15zdnd00an1n02x5 FILLER_163_2226 ();
 b15zdnd00an1n01x5 FILLER_163_2228 ();
 b15zdnd11an1n04x5 FILLER_163_2239 ();
 b15zdnd11an1n32x5 FILLER_163_2247 ();
 b15zdnd11an1n04x5 FILLER_163_2279 ();
 b15zdnd00an1n01x5 FILLER_163_2283 ();
 b15zdnd11an1n16x5 FILLER_164_8 ();
 b15zdnd11an1n08x5 FILLER_164_24 ();
 b15zdnd00an1n01x5 FILLER_164_32 ();
 b15zdnd11an1n04x5 FILLER_164_38 ();
 b15zdnd11an1n32x5 FILLER_164_47 ();
 b15zdnd00an1n02x5 FILLER_164_79 ();
 b15zdnd11an1n04x5 FILLER_164_86 ();
 b15zdnd11an1n16x5 FILLER_164_98 ();
 b15zdnd00an1n01x5 FILLER_164_114 ();
 b15zdnd11an1n04x5 FILLER_164_120 ();
 b15zdnd11an1n16x5 FILLER_164_132 ();
 b15zdnd11an1n08x5 FILLER_164_148 ();
 b15zdnd11an1n04x5 FILLER_164_156 ();
 b15zdnd00an1n01x5 FILLER_164_160 ();
 b15zdnd11an1n64x5 FILLER_164_167 ();
 b15zdnd11an1n32x5 FILLER_164_231 ();
 b15zdnd11an1n16x5 FILLER_164_270 ();
 b15zdnd11an1n08x5 FILLER_164_286 ();
 b15zdnd11an1n04x5 FILLER_164_294 ();
 b15zdnd00an1n01x5 FILLER_164_298 ();
 b15zdnd11an1n04x5 FILLER_164_325 ();
 b15zdnd00an1n01x5 FILLER_164_329 ();
 b15zdnd11an1n64x5 FILLER_164_340 ();
 b15zdnd11an1n04x5 FILLER_164_404 ();
 b15zdnd00an1n01x5 FILLER_164_408 ();
 b15zdnd11an1n32x5 FILLER_164_413 ();
 b15zdnd00an1n01x5 FILLER_164_445 ();
 b15zdnd11an1n08x5 FILLER_164_456 ();
 b15zdnd00an1n01x5 FILLER_164_464 ();
 b15zdnd11an1n08x5 FILLER_164_481 ();
 b15zdnd11an1n04x5 FILLER_164_489 ();
 b15zdnd11an1n32x5 FILLER_164_503 ();
 b15zdnd11an1n04x5 FILLER_164_535 ();
 b15zdnd00an1n02x5 FILLER_164_539 ();
 b15zdnd00an1n01x5 FILLER_164_541 ();
 b15zdnd11an1n08x5 FILLER_164_551 ();
 b15zdnd00an1n01x5 FILLER_164_559 ();
 b15zdnd11an1n04x5 FILLER_164_571 ();
 b15zdnd11an1n08x5 FILLER_164_580 ();
 b15zdnd11an1n04x5 FILLER_164_588 ();
 b15zdnd00an1n02x5 FILLER_164_592 ();
 b15zdnd00an1n01x5 FILLER_164_594 ();
 b15zdnd11an1n08x5 FILLER_164_615 ();
 b15zdnd00an1n02x5 FILLER_164_623 ();
 b15zdnd00an1n01x5 FILLER_164_625 ();
 b15zdnd11an1n04x5 FILLER_164_640 ();
 b15zdnd11an1n16x5 FILLER_164_665 ();
 b15zdnd11an1n32x5 FILLER_164_686 ();
 b15zdnd11an1n04x5 FILLER_164_726 ();
 b15zdnd00an1n01x5 FILLER_164_730 ();
 b15zdnd11an1n64x5 FILLER_164_736 ();
 b15zdnd11an1n16x5 FILLER_164_800 ();
 b15zdnd11an1n04x5 FILLER_164_816 ();
 b15zdnd00an1n01x5 FILLER_164_820 ();
 b15zdnd11an1n16x5 FILLER_164_825 ();
 b15zdnd11an1n08x5 FILLER_164_841 ();
 b15zdnd11an1n04x5 FILLER_164_849 ();
 b15zdnd00an1n02x5 FILLER_164_853 ();
 b15zdnd00an1n01x5 FILLER_164_855 ();
 b15zdnd11an1n04x5 FILLER_164_861 ();
 b15zdnd11an1n04x5 FILLER_164_871 ();
 b15zdnd11an1n32x5 FILLER_164_906 ();
 b15zdnd11an1n08x5 FILLER_164_951 ();
 b15zdnd11an1n04x5 FILLER_164_959 ();
 b15zdnd00an1n02x5 FILLER_164_963 ();
 b15zdnd11an1n08x5 FILLER_164_973 ();
 b15zdnd11an1n04x5 FILLER_164_981 ();
 b15zdnd00an1n01x5 FILLER_164_985 ();
 b15zdnd11an1n04x5 FILLER_164_998 ();
 b15zdnd00an1n02x5 FILLER_164_1002 ();
 b15zdnd11an1n04x5 FILLER_164_1016 ();
 b15zdnd11an1n32x5 FILLER_164_1025 ();
 b15zdnd00an1n02x5 FILLER_164_1057 ();
 b15zdnd11an1n04x5 FILLER_164_1071 ();
 b15zdnd00an1n02x5 FILLER_164_1075 ();
 b15zdnd11an1n16x5 FILLER_164_1093 ();
 b15zdnd11an1n32x5 FILLER_164_1133 ();
 b15zdnd00an1n02x5 FILLER_164_1165 ();
 b15zdnd11an1n16x5 FILLER_164_1174 ();
 b15zdnd00an1n01x5 FILLER_164_1190 ();
 b15zdnd11an1n04x5 FILLER_164_1199 ();
 b15zdnd11an1n64x5 FILLER_164_1217 ();
 b15zdnd11an1n64x5 FILLER_164_1281 ();
 b15zdnd11an1n04x5 FILLER_164_1345 ();
 b15zdnd00an1n01x5 FILLER_164_1349 ();
 b15zdnd11an1n08x5 FILLER_164_1376 ();
 b15zdnd00an1n02x5 FILLER_164_1384 ();
 b15zdnd00an1n01x5 FILLER_164_1386 ();
 b15zdnd11an1n64x5 FILLER_164_1418 ();
 b15zdnd11an1n64x5 FILLER_164_1482 ();
 b15zdnd11an1n08x5 FILLER_164_1546 ();
 b15zdnd11an1n04x5 FILLER_164_1554 ();
 b15zdnd00an1n02x5 FILLER_164_1558 ();
 b15zdnd11an1n64x5 FILLER_164_1566 ();
 b15zdnd11an1n64x5 FILLER_164_1630 ();
 b15zdnd11an1n16x5 FILLER_164_1694 ();
 b15zdnd11an1n04x5 FILLER_164_1710 ();
 b15zdnd11an1n08x5 FILLER_164_1745 ();
 b15zdnd11an1n04x5 FILLER_164_1758 ();
 b15zdnd11an1n32x5 FILLER_164_1782 ();
 b15zdnd11an1n08x5 FILLER_164_1814 ();
 b15zdnd11an1n64x5 FILLER_164_1842 ();
 b15zdnd11an1n64x5 FILLER_164_1906 ();
 b15zdnd11an1n08x5 FILLER_164_1970 ();
 b15zdnd00an1n02x5 FILLER_164_1978 ();
 b15zdnd00an1n01x5 FILLER_164_1980 ();
 b15zdnd11an1n32x5 FILLER_164_1991 ();
 b15zdnd11an1n04x5 FILLER_164_2023 ();
 b15zdnd00an1n02x5 FILLER_164_2027 ();
 b15zdnd00an1n01x5 FILLER_164_2029 ();
 b15zdnd11an1n32x5 FILLER_164_2040 ();
 b15zdnd11an1n08x5 FILLER_164_2072 ();
 b15zdnd11an1n04x5 FILLER_164_2106 ();
 b15zdnd11an1n04x5 FILLER_164_2127 ();
 b15zdnd00an1n02x5 FILLER_164_2151 ();
 b15zdnd00an1n01x5 FILLER_164_2153 ();
 b15zdnd11an1n32x5 FILLER_164_2162 ();
 b15zdnd00an1n02x5 FILLER_164_2194 ();
 b15zdnd11an1n16x5 FILLER_164_2216 ();
 b15zdnd11an1n08x5 FILLER_164_2232 ();
 b15zdnd00an1n02x5 FILLER_164_2240 ();
 b15zdnd11an1n04x5 FILLER_164_2252 ();
 b15zdnd11an1n04x5 FILLER_164_2260 ();
 b15zdnd11an1n08x5 FILLER_164_2268 ();
 b15zdnd11an1n64x5 FILLER_165_0 ();
 b15zdnd11an1n64x5 FILLER_165_64 ();
 b15zdnd11an1n64x5 FILLER_165_128 ();
 b15zdnd11an1n08x5 FILLER_165_192 ();
 b15zdnd11an1n64x5 FILLER_165_206 ();
 b15zdnd11an1n64x5 FILLER_165_270 ();
 b15zdnd11an1n64x5 FILLER_165_334 ();
 b15zdnd11an1n08x5 FILLER_165_398 ();
 b15zdnd00an1n01x5 FILLER_165_406 ();
 b15zdnd11an1n16x5 FILLER_165_412 ();
 b15zdnd11an1n04x5 FILLER_165_428 ();
 b15zdnd11an1n04x5 FILLER_165_448 ();
 b15zdnd11an1n04x5 FILLER_165_458 ();
 b15zdnd11an1n08x5 FILLER_165_468 ();
 b15zdnd00an1n02x5 FILLER_165_476 ();
 b15zdnd11an1n04x5 FILLER_165_492 ();
 b15zdnd00an1n01x5 FILLER_165_496 ();
 b15zdnd11an1n32x5 FILLER_165_507 ();
 b15zdnd11an1n08x5 FILLER_165_539 ();
 b15zdnd11an1n32x5 FILLER_165_553 ();
 b15zdnd11an1n08x5 FILLER_165_585 ();
 b15zdnd11an1n04x5 FILLER_165_593 ();
 b15zdnd11an1n16x5 FILLER_165_601 ();
 b15zdnd11an1n04x5 FILLER_165_617 ();
 b15zdnd00an1n02x5 FILLER_165_621 ();
 b15zdnd11an1n32x5 FILLER_165_649 ();
 b15zdnd11an1n08x5 FILLER_165_686 ();
 b15zdnd00an1n02x5 FILLER_165_694 ();
 b15zdnd00an1n01x5 FILLER_165_696 ();
 b15zdnd11an1n64x5 FILLER_165_711 ();
 b15zdnd11an1n64x5 FILLER_165_775 ();
 b15zdnd11an1n64x5 FILLER_165_839 ();
 b15zdnd11an1n16x5 FILLER_165_903 ();
 b15zdnd00an1n02x5 FILLER_165_919 ();
 b15zdnd00an1n01x5 FILLER_165_921 ();
 b15zdnd11an1n16x5 FILLER_165_938 ();
 b15zdnd11an1n08x5 FILLER_165_954 ();
 b15zdnd00an1n02x5 FILLER_165_962 ();
 b15zdnd00an1n01x5 FILLER_165_964 ();
 b15zdnd11an1n64x5 FILLER_165_972 ();
 b15zdnd11an1n04x5 FILLER_165_1036 ();
 b15zdnd00an1n02x5 FILLER_165_1040 ();
 b15zdnd11an1n04x5 FILLER_165_1047 ();
 b15zdnd11an1n64x5 FILLER_165_1063 ();
 b15zdnd11an1n64x5 FILLER_165_1127 ();
 b15zdnd11an1n04x5 FILLER_165_1191 ();
 b15zdnd00an1n02x5 FILLER_165_1195 ();
 b15zdnd11an1n32x5 FILLER_165_1209 ();
 b15zdnd11an1n16x5 FILLER_165_1241 ();
 b15zdnd11an1n08x5 FILLER_165_1257 ();
 b15zdnd11an1n04x5 FILLER_165_1265 ();
 b15zdnd11an1n04x5 FILLER_165_1300 ();
 b15zdnd11an1n04x5 FILLER_165_1326 ();
 b15zdnd00an1n02x5 FILLER_165_1330 ();
 b15zdnd00an1n01x5 FILLER_165_1332 ();
 b15zdnd11an1n04x5 FILLER_165_1344 ();
 b15zdnd11an1n04x5 FILLER_165_1374 ();
 b15zdnd11an1n16x5 FILLER_165_1404 ();
 b15zdnd11an1n04x5 FILLER_165_1420 ();
 b15zdnd00an1n02x5 FILLER_165_1424 ();
 b15zdnd00an1n01x5 FILLER_165_1426 ();
 b15zdnd11an1n04x5 FILLER_165_1433 ();
 b15zdnd11an1n08x5 FILLER_165_1441 ();
 b15zdnd11an1n04x5 FILLER_165_1449 ();
 b15zdnd00an1n01x5 FILLER_165_1453 ();
 b15zdnd11an1n16x5 FILLER_165_1461 ();
 b15zdnd11an1n04x5 FILLER_165_1477 ();
 b15zdnd00an1n02x5 FILLER_165_1481 ();
 b15zdnd11an1n32x5 FILLER_165_1514 ();
 b15zdnd11an1n08x5 FILLER_165_1546 ();
 b15zdnd11an1n04x5 FILLER_165_1554 ();
 b15zdnd00an1n02x5 FILLER_165_1558 ();
 b15zdnd00an1n01x5 FILLER_165_1560 ();
 b15zdnd11an1n64x5 FILLER_165_1581 ();
 b15zdnd11an1n64x5 FILLER_165_1645 ();
 b15zdnd11an1n16x5 FILLER_165_1709 ();
 b15zdnd11an1n04x5 FILLER_165_1725 ();
 b15zdnd00an1n02x5 FILLER_165_1729 ();
 b15zdnd00an1n01x5 FILLER_165_1731 ();
 b15zdnd11an1n04x5 FILLER_165_1763 ();
 b15zdnd11an1n04x5 FILLER_165_1798 ();
 b15zdnd00an1n02x5 FILLER_165_1802 ();
 b15zdnd11an1n08x5 FILLER_165_1808 ();
 b15zdnd11an1n16x5 FILLER_165_1821 ();
 b15zdnd00an1n02x5 FILLER_165_1837 ();
 b15zdnd11an1n08x5 FILLER_165_1864 ();
 b15zdnd11an1n04x5 FILLER_165_1872 ();
 b15zdnd11an1n64x5 FILLER_165_1881 ();
 b15zdnd11an1n32x5 FILLER_165_1945 ();
 b15zdnd11an1n08x5 FILLER_165_1977 ();
 b15zdnd00an1n02x5 FILLER_165_1985 ();
 b15zdnd00an1n01x5 FILLER_165_1987 ();
 b15zdnd11an1n16x5 FILLER_165_1997 ();
 b15zdnd11an1n04x5 FILLER_165_2013 ();
 b15zdnd11an1n64x5 FILLER_165_2049 ();
 b15zdnd11an1n64x5 FILLER_165_2113 ();
 b15zdnd11an1n64x5 FILLER_165_2177 ();
 b15zdnd11an1n32x5 FILLER_165_2241 ();
 b15zdnd11an1n08x5 FILLER_165_2273 ();
 b15zdnd00an1n02x5 FILLER_165_2281 ();
 b15zdnd00an1n01x5 FILLER_165_2283 ();
 b15zdnd11an1n64x5 FILLER_166_8 ();
 b15zdnd11an1n04x5 FILLER_166_72 ();
 b15zdnd00an1n02x5 FILLER_166_76 ();
 b15zdnd00an1n01x5 FILLER_166_78 ();
 b15zdnd11an1n16x5 FILLER_166_89 ();
 b15zdnd11an1n08x5 FILLER_166_105 ();
 b15zdnd00an1n02x5 FILLER_166_113 ();
 b15zdnd00an1n01x5 FILLER_166_115 ();
 b15zdnd11an1n04x5 FILLER_166_124 ();
 b15zdnd11an1n16x5 FILLER_166_140 ();
 b15zdnd11an1n08x5 FILLER_166_156 ();
 b15zdnd11an1n08x5 FILLER_166_172 ();
 b15zdnd11an1n04x5 FILLER_166_180 ();
 b15zdnd00an1n02x5 FILLER_166_184 ();
 b15zdnd00an1n01x5 FILLER_166_186 ();
 b15zdnd11an1n04x5 FILLER_166_195 ();
 b15zdnd11an1n08x5 FILLER_166_211 ();
 b15zdnd11an1n04x5 FILLER_166_219 ();
 b15zdnd00an1n02x5 FILLER_166_223 ();
 b15zdnd00an1n01x5 FILLER_166_225 ();
 b15zdnd11an1n08x5 FILLER_166_231 ();
 b15zdnd00an1n02x5 FILLER_166_239 ();
 b15zdnd00an1n01x5 FILLER_166_241 ();
 b15zdnd11an1n04x5 FILLER_166_249 ();
 b15zdnd11an1n04x5 FILLER_166_260 ();
 b15zdnd00an1n01x5 FILLER_166_264 ();
 b15zdnd11an1n08x5 FILLER_166_272 ();
 b15zdnd00an1n02x5 FILLER_166_280 ();
 b15zdnd11an1n64x5 FILLER_166_289 ();
 b15zdnd11an1n32x5 FILLER_166_353 ();
 b15zdnd11an1n16x5 FILLER_166_385 ();
 b15zdnd11an1n04x5 FILLER_166_401 ();
 b15zdnd00an1n02x5 FILLER_166_405 ();
 b15zdnd11an1n32x5 FILLER_166_419 ();
 b15zdnd11an1n04x5 FILLER_166_451 ();
 b15zdnd00an1n02x5 FILLER_166_455 ();
 b15zdnd00an1n01x5 FILLER_166_457 ();
 b15zdnd11an1n32x5 FILLER_166_465 ();
 b15zdnd11an1n16x5 FILLER_166_497 ();
 b15zdnd00an1n02x5 FILLER_166_513 ();
 b15zdnd00an1n01x5 FILLER_166_515 ();
 b15zdnd11an1n08x5 FILLER_166_538 ();
 b15zdnd00an1n01x5 FILLER_166_546 ();
 b15zdnd11an1n32x5 FILLER_166_553 ();
 b15zdnd11an1n08x5 FILLER_166_585 ();
 b15zdnd00an1n02x5 FILLER_166_593 ();
 b15zdnd00an1n01x5 FILLER_166_595 ();
 b15zdnd11an1n08x5 FILLER_166_610 ();
 b15zdnd11an1n16x5 FILLER_166_630 ();
 b15zdnd11an1n08x5 FILLER_166_646 ();
 b15zdnd11an1n04x5 FILLER_166_654 ();
 b15zdnd11an1n04x5 FILLER_166_665 ();
 b15zdnd00an1n01x5 FILLER_166_669 ();
 b15zdnd11an1n08x5 FILLER_166_676 ();
 b15zdnd11an1n04x5 FILLER_166_692 ();
 b15zdnd11an1n08x5 FILLER_166_704 ();
 b15zdnd11an1n04x5 FILLER_166_712 ();
 b15zdnd00an1n02x5 FILLER_166_716 ();
 b15zdnd11an1n16x5 FILLER_166_726 ();
 b15zdnd11an1n04x5 FILLER_166_742 ();
 b15zdnd11an1n04x5 FILLER_166_778 ();
 b15zdnd11an1n64x5 FILLER_166_802 ();
 b15zdnd00an1n01x5 FILLER_166_866 ();
 b15zdnd11an1n16x5 FILLER_166_871 ();
 b15zdnd11an1n08x5 FILLER_166_887 ();
 b15zdnd11an1n04x5 FILLER_166_902 ();
 b15zdnd11an1n64x5 FILLER_166_932 ();
 b15zdnd11an1n64x5 FILLER_166_996 ();
 b15zdnd11an1n32x5 FILLER_166_1060 ();
 b15zdnd11an1n16x5 FILLER_166_1092 ();
 b15zdnd11an1n08x5 FILLER_166_1108 ();
 b15zdnd00an1n02x5 FILLER_166_1116 ();
 b15zdnd00an1n01x5 FILLER_166_1118 ();
 b15zdnd11an1n32x5 FILLER_166_1123 ();
 b15zdnd11an1n08x5 FILLER_166_1155 ();
 b15zdnd00an1n02x5 FILLER_166_1163 ();
 b15zdnd00an1n01x5 FILLER_166_1165 ();
 b15zdnd11an1n64x5 FILLER_166_1172 ();
 b15zdnd11an1n64x5 FILLER_166_1236 ();
 b15zdnd11an1n16x5 FILLER_166_1300 ();
 b15zdnd00an1n02x5 FILLER_166_1316 ();
 b15zdnd11an1n08x5 FILLER_166_1340 ();
 b15zdnd00an1n02x5 FILLER_166_1348 ();
 b15zdnd11an1n32x5 FILLER_166_1363 ();
 b15zdnd00an1n02x5 FILLER_166_1395 ();
 b15zdnd11an1n08x5 FILLER_166_1409 ();
 b15zdnd11an1n04x5 FILLER_166_1417 ();
 b15zdnd00an1n02x5 FILLER_166_1421 ();
 b15zdnd11an1n04x5 FILLER_166_1433 ();
 b15zdnd11an1n64x5 FILLER_166_1442 ();
 b15zdnd00an1n02x5 FILLER_166_1506 ();
 b15zdnd11an1n16x5 FILLER_166_1513 ();
 b15zdnd11an1n04x5 FILLER_166_1529 ();
 b15zdnd00an1n02x5 FILLER_166_1533 ();
 b15zdnd00an1n01x5 FILLER_166_1535 ();
 b15zdnd11an1n04x5 FILLER_166_1545 ();
 b15zdnd11an1n08x5 FILLER_166_1553 ();
 b15zdnd11an1n64x5 FILLER_166_1567 ();
 b15zdnd00an1n02x5 FILLER_166_1631 ();
 b15zdnd11an1n04x5 FILLER_166_1665 ();
 b15zdnd11an1n64x5 FILLER_166_1687 ();
 b15zdnd11an1n08x5 FILLER_166_1751 ();
 b15zdnd11an1n04x5 FILLER_166_1759 ();
 b15zdnd11an1n64x5 FILLER_166_1794 ();
 b15zdnd11an1n08x5 FILLER_166_1858 ();
 b15zdnd11an1n04x5 FILLER_166_1866 ();
 b15zdnd00an1n02x5 FILLER_166_1870 ();
 b15zdnd11an1n64x5 FILLER_166_1878 ();
 b15zdnd11an1n08x5 FILLER_166_1942 ();
 b15zdnd00an1n02x5 FILLER_166_1950 ();
 b15zdnd11an1n16x5 FILLER_166_1964 ();
 b15zdnd11an1n04x5 FILLER_166_1980 ();
 b15zdnd00an1n01x5 FILLER_166_1984 ();
 b15zdnd11an1n32x5 FILLER_166_1997 ();
 b15zdnd11an1n16x5 FILLER_166_2029 ();
 b15zdnd11an1n08x5 FILLER_166_2045 ();
 b15zdnd00an1n01x5 FILLER_166_2053 ();
 b15zdnd11an1n64x5 FILLER_166_2086 ();
 b15zdnd11an1n04x5 FILLER_166_2150 ();
 b15zdnd11an1n64x5 FILLER_166_2162 ();
 b15zdnd11an1n08x5 FILLER_166_2226 ();
 b15zdnd00an1n02x5 FILLER_166_2234 ();
 b15zdnd00an1n01x5 FILLER_166_2236 ();
 b15zdnd11an1n04x5 FILLER_166_2247 ();
 b15zdnd11an1n04x5 FILLER_166_2255 ();
 b15zdnd11an1n04x5 FILLER_166_2263 ();
 b15zdnd00an1n02x5 FILLER_166_2267 ();
 b15zdnd00an1n01x5 FILLER_166_2269 ();
 b15zdnd00an1n02x5 FILLER_166_2274 ();
 b15zdnd11an1n64x5 FILLER_167_0 ();
 b15zdnd11an1n08x5 FILLER_167_64 ();
 b15zdnd11an1n32x5 FILLER_167_78 ();
 b15zdnd11an1n04x5 FILLER_167_124 ();
 b15zdnd00an1n02x5 FILLER_167_128 ();
 b15zdnd00an1n01x5 FILLER_167_130 ();
 b15zdnd11an1n16x5 FILLER_167_144 ();
 b15zdnd11an1n04x5 FILLER_167_160 ();
 b15zdnd00an1n02x5 FILLER_167_164 ();
 b15zdnd00an1n01x5 FILLER_167_166 ();
 b15zdnd11an1n16x5 FILLER_167_179 ();
 b15zdnd11an1n08x5 FILLER_167_199 ();
 b15zdnd11an1n04x5 FILLER_167_207 ();
 b15zdnd11an1n04x5 FILLER_167_217 ();
 b15zdnd11an1n16x5 FILLER_167_226 ();
 b15zdnd11an1n08x5 FILLER_167_242 ();
 b15zdnd11an1n04x5 FILLER_167_250 ();
 b15zdnd00an1n02x5 FILLER_167_254 ();
 b15zdnd11an1n04x5 FILLER_167_261 ();
 b15zdnd00an1n02x5 FILLER_167_265 ();
 b15zdnd11an1n16x5 FILLER_167_293 ();
 b15zdnd11an1n04x5 FILLER_167_321 ();
 b15zdnd00an1n02x5 FILLER_167_325 ();
 b15zdnd11an1n64x5 FILLER_167_337 ();
 b15zdnd11an1n32x5 FILLER_167_401 ();
 b15zdnd11an1n16x5 FILLER_167_433 ();
 b15zdnd00an1n02x5 FILLER_167_449 ();
 b15zdnd11an1n32x5 FILLER_167_467 ();
 b15zdnd11an1n04x5 FILLER_167_499 ();
 b15zdnd00an1n01x5 FILLER_167_503 ();
 b15zdnd11an1n32x5 FILLER_167_508 ();
 b15zdnd11an1n16x5 FILLER_167_540 ();
 b15zdnd11an1n08x5 FILLER_167_556 ();
 b15zdnd11an1n04x5 FILLER_167_564 ();
 b15zdnd00an1n01x5 FILLER_167_568 ();
 b15zdnd11an1n08x5 FILLER_167_576 ();
 b15zdnd00an1n01x5 FILLER_167_584 ();
 b15zdnd11an1n64x5 FILLER_167_594 ();
 b15zdnd11an1n16x5 FILLER_167_658 ();
 b15zdnd11an1n08x5 FILLER_167_674 ();
 b15zdnd11an1n64x5 FILLER_167_689 ();
 b15zdnd11an1n16x5 FILLER_167_753 ();
 b15zdnd11an1n08x5 FILLER_167_769 ();
 b15zdnd00an1n01x5 FILLER_167_777 ();
 b15zdnd11an1n08x5 FILLER_167_783 ();
 b15zdnd11an1n04x5 FILLER_167_791 ();
 b15zdnd00an1n02x5 FILLER_167_795 ();
 b15zdnd00an1n01x5 FILLER_167_797 ();
 b15zdnd11an1n32x5 FILLER_167_801 ();
 b15zdnd11an1n16x5 FILLER_167_833 ();
 b15zdnd11an1n04x5 FILLER_167_849 ();
 b15zdnd00an1n01x5 FILLER_167_853 ();
 b15zdnd11an1n32x5 FILLER_167_861 ();
 b15zdnd11an1n08x5 FILLER_167_893 ();
 b15zdnd00an1n01x5 FILLER_167_901 ();
 b15zdnd11an1n32x5 FILLER_167_914 ();
 b15zdnd11an1n16x5 FILLER_167_946 ();
 b15zdnd11an1n08x5 FILLER_167_962 ();
 b15zdnd11an1n04x5 FILLER_167_970 ();
 b15zdnd00an1n01x5 FILLER_167_974 ();
 b15zdnd11an1n64x5 FILLER_167_980 ();
 b15zdnd11an1n16x5 FILLER_167_1044 ();
 b15zdnd11an1n08x5 FILLER_167_1060 ();
 b15zdnd11an1n04x5 FILLER_167_1068 ();
 b15zdnd00an1n01x5 FILLER_167_1072 ();
 b15zdnd11an1n08x5 FILLER_167_1078 ();
 b15zdnd11an1n08x5 FILLER_167_1090 ();
 b15zdnd11an1n04x5 FILLER_167_1098 ();
 b15zdnd00an1n02x5 FILLER_167_1102 ();
 b15zdnd00an1n01x5 FILLER_167_1104 ();
 b15zdnd11an1n04x5 FILLER_167_1121 ();
 b15zdnd11an1n16x5 FILLER_167_1131 ();
 b15zdnd11an1n64x5 FILLER_167_1160 ();
 b15zdnd11an1n64x5 FILLER_167_1224 ();
 b15zdnd11an1n32x5 FILLER_167_1288 ();
 b15zdnd11an1n04x5 FILLER_167_1351 ();
 b15zdnd11an1n32x5 FILLER_167_1361 ();
 b15zdnd11an1n16x5 FILLER_167_1393 ();
 b15zdnd11an1n08x5 FILLER_167_1409 ();
 b15zdnd11an1n04x5 FILLER_167_1417 ();
 b15zdnd00an1n02x5 FILLER_167_1421 ();
 b15zdnd00an1n01x5 FILLER_167_1423 ();
 b15zdnd11an1n16x5 FILLER_167_1428 ();
 b15zdnd11an1n08x5 FILLER_167_1444 ();
 b15zdnd11an1n04x5 FILLER_167_1452 ();
 b15zdnd00an1n01x5 FILLER_167_1456 ();
 b15zdnd11an1n32x5 FILLER_167_1467 ();
 b15zdnd11an1n04x5 FILLER_167_1499 ();
 b15zdnd11an1n08x5 FILLER_167_1518 ();
 b15zdnd00an1n02x5 FILLER_167_1526 ();
 b15zdnd00an1n01x5 FILLER_167_1528 ();
 b15zdnd11an1n16x5 FILLER_167_1543 ();
 b15zdnd00an1n01x5 FILLER_167_1559 ();
 b15zdnd11an1n08x5 FILLER_167_1566 ();
 b15zdnd11an1n04x5 FILLER_167_1574 ();
 b15zdnd00an1n01x5 FILLER_167_1578 ();
 b15zdnd11an1n16x5 FILLER_167_1582 ();
 b15zdnd11an1n08x5 FILLER_167_1598 ();
 b15zdnd11an1n04x5 FILLER_167_1606 ();
 b15zdnd00an1n02x5 FILLER_167_1610 ();
 b15zdnd00an1n01x5 FILLER_167_1612 ();
 b15zdnd11an1n08x5 FILLER_167_1618 ();
 b15zdnd11an1n04x5 FILLER_167_1634 ();
 b15zdnd11an1n32x5 FILLER_167_1643 ();
 b15zdnd11an1n08x5 FILLER_167_1675 ();
 b15zdnd00an1n01x5 FILLER_167_1683 ();
 b15zdnd11an1n16x5 FILLER_167_1709 ();
 b15zdnd11an1n08x5 FILLER_167_1725 ();
 b15zdnd11an1n04x5 FILLER_167_1733 ();
 b15zdnd00an1n02x5 FILLER_167_1737 ();
 b15zdnd11an1n64x5 FILLER_167_1750 ();
 b15zdnd11an1n16x5 FILLER_167_1814 ();
 b15zdnd11an1n08x5 FILLER_167_1830 ();
 b15zdnd11an1n04x5 FILLER_167_1838 ();
 b15zdnd00an1n02x5 FILLER_167_1842 ();
 b15zdnd11an1n04x5 FILLER_167_1864 ();
 b15zdnd11an1n08x5 FILLER_167_1875 ();
 b15zdnd00an1n02x5 FILLER_167_1883 ();
 b15zdnd11an1n04x5 FILLER_167_1892 ();
 b15zdnd11an1n64x5 FILLER_167_1901 ();
 b15zdnd11an1n64x5 FILLER_167_1965 ();
 b15zdnd11an1n64x5 FILLER_167_2029 ();
 b15zdnd11an1n64x5 FILLER_167_2093 ();
 b15zdnd11an1n64x5 FILLER_167_2157 ();
 b15zdnd00an1n01x5 FILLER_167_2221 ();
 b15zdnd11an1n16x5 FILLER_167_2227 ();
 b15zdnd11an1n04x5 FILLER_167_2243 ();
 b15zdnd00an1n01x5 FILLER_167_2247 ();
 b15zdnd11an1n08x5 FILLER_167_2252 ();
 b15zdnd11an1n16x5 FILLER_167_2266 ();
 b15zdnd00an1n02x5 FILLER_167_2282 ();
 b15zdnd11an1n16x5 FILLER_168_8 ();
 b15zdnd11an1n08x5 FILLER_168_24 ();
 b15zdnd00an1n02x5 FILLER_168_32 ();
 b15zdnd00an1n01x5 FILLER_168_34 ();
 b15zdnd11an1n08x5 FILLER_168_40 ();
 b15zdnd11an1n64x5 FILLER_168_62 ();
 b15zdnd11an1n04x5 FILLER_168_126 ();
 b15zdnd00an1n02x5 FILLER_168_130 ();
 b15zdnd00an1n01x5 FILLER_168_132 ();
 b15zdnd11an1n16x5 FILLER_168_141 ();
 b15zdnd11an1n08x5 FILLER_168_157 ();
 b15zdnd00an1n02x5 FILLER_168_165 ();
 b15zdnd00an1n01x5 FILLER_168_167 ();
 b15zdnd11an1n32x5 FILLER_168_174 ();
 b15zdnd11an1n16x5 FILLER_168_206 ();
 b15zdnd00an1n01x5 FILLER_168_222 ();
 b15zdnd11an1n64x5 FILLER_168_229 ();
 b15zdnd11an1n04x5 FILLER_168_305 ();
 b15zdnd00an1n01x5 FILLER_168_309 ();
 b15zdnd11an1n04x5 FILLER_168_324 ();
 b15zdnd00an1n01x5 FILLER_168_328 ();
 b15zdnd11an1n64x5 FILLER_168_341 ();
 b15zdnd11an1n08x5 FILLER_168_405 ();
 b15zdnd11an1n04x5 FILLER_168_413 ();
 b15zdnd00an1n02x5 FILLER_168_417 ();
 b15zdnd00an1n01x5 FILLER_168_419 ();
 b15zdnd11an1n04x5 FILLER_168_426 ();
 b15zdnd11an1n32x5 FILLER_168_437 ();
 b15zdnd11an1n16x5 FILLER_168_469 ();
 b15zdnd11an1n08x5 FILLER_168_485 ();
 b15zdnd11an1n04x5 FILLER_168_493 ();
 b15zdnd00an1n02x5 FILLER_168_497 ();
 b15zdnd00an1n01x5 FILLER_168_499 ();
 b15zdnd11an1n04x5 FILLER_168_512 ();
 b15zdnd11an1n16x5 FILLER_168_521 ();
 b15zdnd11an1n04x5 FILLER_168_537 ();
 b15zdnd00an1n02x5 FILLER_168_541 ();
 b15zdnd00an1n01x5 FILLER_168_543 ();
 b15zdnd11an1n08x5 FILLER_168_550 ();
 b15zdnd11an1n04x5 FILLER_168_558 ();
 b15zdnd00an1n02x5 FILLER_168_562 ();
 b15zdnd00an1n01x5 FILLER_168_564 ();
 b15zdnd11an1n08x5 FILLER_168_577 ();
 b15zdnd00an1n01x5 FILLER_168_585 ();
 b15zdnd11an1n64x5 FILLER_168_591 ();
 b15zdnd11an1n32x5 FILLER_168_655 ();
 b15zdnd11an1n16x5 FILLER_168_687 ();
 b15zdnd11an1n08x5 FILLER_168_703 ();
 b15zdnd11an1n04x5 FILLER_168_711 ();
 b15zdnd00an1n02x5 FILLER_168_715 ();
 b15zdnd00an1n01x5 FILLER_168_717 ();
 b15zdnd11an1n08x5 FILLER_168_726 ();
 b15zdnd11an1n04x5 FILLER_168_734 ();
 b15zdnd11an1n64x5 FILLER_168_744 ();
 b15zdnd11an1n32x5 FILLER_168_808 ();
 b15zdnd11an1n08x5 FILLER_168_840 ();
 b15zdnd11an1n04x5 FILLER_168_848 ();
 b15zdnd11an1n16x5 FILLER_168_857 ();
 b15zdnd11an1n08x5 FILLER_168_873 ();
 b15zdnd11an1n04x5 FILLER_168_889 ();
 b15zdnd11an1n32x5 FILLER_168_919 ();
 b15zdnd11an1n16x5 FILLER_168_951 ();
 b15zdnd00an1n02x5 FILLER_168_967 ();
 b15zdnd00an1n01x5 FILLER_168_969 ();
 b15zdnd11an1n32x5 FILLER_168_980 ();
 b15zdnd11an1n04x5 FILLER_168_1012 ();
 b15zdnd00an1n01x5 FILLER_168_1016 ();
 b15zdnd11an1n32x5 FILLER_168_1026 ();
 b15zdnd11an1n04x5 FILLER_168_1058 ();
 b15zdnd00an1n02x5 FILLER_168_1062 ();
 b15zdnd00an1n01x5 FILLER_168_1064 ();
 b15zdnd11an1n32x5 FILLER_168_1097 ();
 b15zdnd11an1n08x5 FILLER_168_1129 ();
 b15zdnd11an1n04x5 FILLER_168_1137 ();
 b15zdnd11an1n04x5 FILLER_168_1161 ();
 b15zdnd00an1n02x5 FILLER_168_1165 ();
 b15zdnd00an1n01x5 FILLER_168_1167 ();
 b15zdnd11an1n16x5 FILLER_168_1178 ();
 b15zdnd11an1n04x5 FILLER_168_1194 ();
 b15zdnd11an1n32x5 FILLER_168_1202 ();
 b15zdnd11an1n16x5 FILLER_168_1234 ();
 b15zdnd00an1n02x5 FILLER_168_1250 ();
 b15zdnd11an1n32x5 FILLER_168_1272 ();
 b15zdnd00an1n02x5 FILLER_168_1304 ();
 b15zdnd11an1n16x5 FILLER_168_1324 ();
 b15zdnd11an1n04x5 FILLER_168_1340 ();
 b15zdnd00an1n02x5 FILLER_168_1344 ();
 b15zdnd11an1n16x5 FILLER_168_1361 ();
 b15zdnd00an1n01x5 FILLER_168_1377 ();
 b15zdnd11an1n04x5 FILLER_168_1388 ();
 b15zdnd00an1n02x5 FILLER_168_1392 ();
 b15zdnd11an1n16x5 FILLER_168_1402 ();
 b15zdnd00an1n01x5 FILLER_168_1418 ();
 b15zdnd11an1n16x5 FILLER_168_1427 ();
 b15zdnd11an1n08x5 FILLER_168_1443 ();
 b15zdnd00an1n01x5 FILLER_168_1451 ();
 b15zdnd11an1n16x5 FILLER_168_1458 ();
 b15zdnd00an1n01x5 FILLER_168_1474 ();
 b15zdnd11an1n04x5 FILLER_168_1487 ();
 b15zdnd11an1n16x5 FILLER_168_1497 ();
 b15zdnd11an1n64x5 FILLER_168_1522 ();
 b15zdnd11an1n64x5 FILLER_168_1586 ();
 b15zdnd11an1n32x5 FILLER_168_1650 ();
 b15zdnd00an1n02x5 FILLER_168_1682 ();
 b15zdnd00an1n01x5 FILLER_168_1684 ();
 b15zdnd11an1n64x5 FILLER_168_1700 ();
 b15zdnd11an1n32x5 FILLER_168_1764 ();
 b15zdnd11an1n16x5 FILLER_168_1796 ();
 b15zdnd11an1n08x5 FILLER_168_1812 ();
 b15zdnd11an1n04x5 FILLER_168_1820 ();
 b15zdnd00an1n02x5 FILLER_168_1824 ();
 b15zdnd11an1n16x5 FILLER_168_1848 ();
 b15zdnd11an1n04x5 FILLER_168_1864 ();
 b15zdnd00an1n01x5 FILLER_168_1868 ();
 b15zdnd11an1n04x5 FILLER_168_1878 ();
 b15zdnd00an1n02x5 FILLER_168_1882 ();
 b15zdnd11an1n04x5 FILLER_168_1889 ();
 b15zdnd00an1n02x5 FILLER_168_1893 ();
 b15zdnd00an1n01x5 FILLER_168_1895 ();
 b15zdnd11an1n16x5 FILLER_168_1899 ();
 b15zdnd11an1n04x5 FILLER_168_1915 ();
 b15zdnd00an1n02x5 FILLER_168_1919 ();
 b15zdnd11an1n64x5 FILLER_168_1941 ();
 b15zdnd11an1n16x5 FILLER_168_2005 ();
 b15zdnd11an1n04x5 FILLER_168_2021 ();
 b15zdnd00an1n02x5 FILLER_168_2025 ();
 b15zdnd00an1n01x5 FILLER_168_2027 ();
 b15zdnd11an1n64x5 FILLER_168_2039 ();
 b15zdnd11an1n32x5 FILLER_168_2103 ();
 b15zdnd11an1n16x5 FILLER_168_2135 ();
 b15zdnd00an1n02x5 FILLER_168_2151 ();
 b15zdnd00an1n01x5 FILLER_168_2153 ();
 b15zdnd11an1n08x5 FILLER_168_2162 ();
 b15zdnd11an1n16x5 FILLER_168_2190 ();
 b15zdnd00an1n02x5 FILLER_168_2206 ();
 b15zdnd11an1n04x5 FILLER_168_2212 ();
 b15zdnd11an1n04x5 FILLER_168_2220 ();
 b15zdnd11an1n08x5 FILLER_168_2244 ();
 b15zdnd11an1n08x5 FILLER_168_2256 ();
 b15zdnd11an1n04x5 FILLER_168_2264 ();
 b15zdnd00an1n02x5 FILLER_168_2268 ();
 b15zdnd00an1n02x5 FILLER_168_2274 ();
 b15zdnd11an1n16x5 FILLER_169_0 ();
 b15zdnd11an1n04x5 FILLER_169_20 ();
 b15zdnd00an1n01x5 FILLER_169_24 ();
 b15zdnd11an1n08x5 FILLER_169_31 ();
 b15zdnd11an1n04x5 FILLER_169_43 ();
 b15zdnd00an1n02x5 FILLER_169_47 ();
 b15zdnd11an1n08x5 FILLER_169_55 ();
 b15zdnd11an1n04x5 FILLER_169_63 ();
 b15zdnd11an1n04x5 FILLER_169_79 ();
 b15zdnd00an1n02x5 FILLER_169_83 ();
 b15zdnd11an1n16x5 FILLER_169_91 ();
 b15zdnd00an1n02x5 FILLER_169_107 ();
 b15zdnd11an1n16x5 FILLER_169_119 ();
 b15zdnd11an1n04x5 FILLER_169_140 ();
 b15zdnd11an1n64x5 FILLER_169_153 ();
 b15zdnd11an1n64x5 FILLER_169_217 ();
 b15zdnd11an1n16x5 FILLER_169_281 ();
 b15zdnd11an1n08x5 FILLER_169_297 ();
 b15zdnd00an1n02x5 FILLER_169_305 ();
 b15zdnd11an1n04x5 FILLER_169_322 ();
 b15zdnd11an1n32x5 FILLER_169_335 ();
 b15zdnd11an1n16x5 FILLER_169_367 ();
 b15zdnd11an1n08x5 FILLER_169_383 ();
 b15zdnd11an1n04x5 FILLER_169_391 ();
 b15zdnd00an1n02x5 FILLER_169_395 ();
 b15zdnd11an1n08x5 FILLER_169_404 ();
 b15zdnd00an1n01x5 FILLER_169_412 ();
 b15zdnd11an1n32x5 FILLER_169_421 ();
 b15zdnd00an1n01x5 FILLER_169_453 ();
 b15zdnd11an1n32x5 FILLER_169_463 ();
 b15zdnd11an1n04x5 FILLER_169_495 ();
 b15zdnd11an1n32x5 FILLER_169_513 ();
 b15zdnd00an1n02x5 FILLER_169_545 ();
 b15zdnd00an1n01x5 FILLER_169_547 ();
 b15zdnd11an1n32x5 FILLER_169_562 ();
 b15zdnd11an1n16x5 FILLER_169_594 ();
 b15zdnd11an1n04x5 FILLER_169_610 ();
 b15zdnd00an1n02x5 FILLER_169_614 ();
 b15zdnd00an1n01x5 FILLER_169_616 ();
 b15zdnd11an1n16x5 FILLER_169_624 ();
 b15zdnd11an1n08x5 FILLER_169_640 ();
 b15zdnd11an1n04x5 FILLER_169_648 ();
 b15zdnd00an1n02x5 FILLER_169_652 ();
 b15zdnd11an1n16x5 FILLER_169_661 ();
 b15zdnd11an1n04x5 FILLER_169_677 ();
 b15zdnd00an1n01x5 FILLER_169_681 ();
 b15zdnd11an1n16x5 FILLER_169_686 ();
 b15zdnd11an1n32x5 FILLER_169_713 ();
 b15zdnd11an1n16x5 FILLER_169_745 ();
 b15zdnd00an1n02x5 FILLER_169_761 ();
 b15zdnd00an1n01x5 FILLER_169_763 ();
 b15zdnd11an1n64x5 FILLER_169_768 ();
 b15zdnd11an1n16x5 FILLER_169_832 ();
 b15zdnd11an1n04x5 FILLER_169_848 ();
 b15zdnd00an1n02x5 FILLER_169_852 ();
 b15zdnd00an1n01x5 FILLER_169_854 ();
 b15zdnd11an1n32x5 FILLER_169_864 ();
 b15zdnd00an1n02x5 FILLER_169_896 ();
 b15zdnd00an1n01x5 FILLER_169_898 ();
 b15zdnd11an1n04x5 FILLER_169_904 ();
 b15zdnd11an1n08x5 FILLER_169_916 ();
 b15zdnd11an1n04x5 FILLER_169_924 ();
 b15zdnd00an1n02x5 FILLER_169_928 ();
 b15zdnd11an1n08x5 FILLER_169_936 ();
 b15zdnd11an1n04x5 FILLER_169_975 ();
 b15zdnd00an1n02x5 FILLER_169_979 ();
 b15zdnd00an1n01x5 FILLER_169_981 ();
 b15zdnd11an1n04x5 FILLER_169_988 ();
 b15zdnd11an1n16x5 FILLER_169_999 ();
 b15zdnd11an1n04x5 FILLER_169_1015 ();
 b15zdnd00an1n01x5 FILLER_169_1019 ();
 b15zdnd11an1n16x5 FILLER_169_1035 ();
 b15zdnd11an1n08x5 FILLER_169_1051 ();
 b15zdnd11an1n08x5 FILLER_169_1063 ();
 b15zdnd11an1n04x5 FILLER_169_1071 ();
 b15zdnd00an1n02x5 FILLER_169_1075 ();
 b15zdnd11an1n32x5 FILLER_169_1082 ();
 b15zdnd11an1n08x5 FILLER_169_1114 ();
 b15zdnd11an1n04x5 FILLER_169_1122 ();
 b15zdnd11an1n64x5 FILLER_169_1133 ();
 b15zdnd11an1n64x5 FILLER_169_1197 ();
 b15zdnd11an1n16x5 FILLER_169_1261 ();
 b15zdnd11an1n04x5 FILLER_169_1277 ();
 b15zdnd00an1n02x5 FILLER_169_1281 ();
 b15zdnd11an1n04x5 FILLER_169_1301 ();
 b15zdnd11an1n16x5 FILLER_169_1328 ();
 b15zdnd11an1n08x5 FILLER_169_1344 ();
 b15zdnd11an1n64x5 FILLER_169_1362 ();
 b15zdnd11an1n16x5 FILLER_169_1432 ();
 b15zdnd11an1n04x5 FILLER_169_1448 ();
 b15zdnd00an1n01x5 FILLER_169_1452 ();
 b15zdnd11an1n16x5 FILLER_169_1459 ();
 b15zdnd00an1n02x5 FILLER_169_1475 ();
 b15zdnd11an1n32x5 FILLER_169_1481 ();
 b15zdnd11an1n08x5 FILLER_169_1513 ();
 b15zdnd11an1n04x5 FILLER_169_1521 ();
 b15zdnd00an1n02x5 FILLER_169_1525 ();
 b15zdnd11an1n04x5 FILLER_169_1545 ();
 b15zdnd11an1n08x5 FILLER_169_1567 ();
 b15zdnd11an1n04x5 FILLER_169_1575 ();
 b15zdnd00an1n02x5 FILLER_169_1579 ();
 b15zdnd11an1n16x5 FILLER_169_1593 ();
 b15zdnd00an1n01x5 FILLER_169_1609 ();
 b15zdnd11an1n16x5 FILLER_169_1627 ();
 b15zdnd11an1n04x5 FILLER_169_1643 ();
 b15zdnd00an1n02x5 FILLER_169_1647 ();
 b15zdnd11an1n64x5 FILLER_169_1673 ();
 b15zdnd00an1n01x5 FILLER_169_1737 ();
 b15zdnd11an1n64x5 FILLER_169_1758 ();
 b15zdnd11an1n64x5 FILLER_169_1822 ();
 b15zdnd11an1n08x5 FILLER_169_1886 ();
 b15zdnd11an1n04x5 FILLER_169_1894 ();
 b15zdnd00an1n02x5 FILLER_169_1898 ();
 b15zdnd00an1n01x5 FILLER_169_1900 ();
 b15zdnd11an1n32x5 FILLER_169_1910 ();
 b15zdnd11an1n08x5 FILLER_169_1942 ();
 b15zdnd11an1n04x5 FILLER_169_1950 ();
 b15zdnd00an1n02x5 FILLER_169_1954 ();
 b15zdnd00an1n01x5 FILLER_169_1956 ();
 b15zdnd11an1n64x5 FILLER_169_1975 ();
 b15zdnd11an1n08x5 FILLER_169_2039 ();
 b15zdnd00an1n01x5 FILLER_169_2047 ();
 b15zdnd11an1n16x5 FILLER_169_2073 ();
 b15zdnd00an1n02x5 FILLER_169_2089 ();
 b15zdnd11an1n32x5 FILLER_169_2119 ();
 b15zdnd11an1n04x5 FILLER_169_2156 ();
 b15zdnd11an1n08x5 FILLER_169_2180 ();
 b15zdnd00an1n02x5 FILLER_169_2188 ();
 b15zdnd00an1n01x5 FILLER_169_2190 ();
 b15zdnd11an1n64x5 FILLER_169_2196 ();
 b15zdnd11an1n16x5 FILLER_169_2260 ();
 b15zdnd11an1n08x5 FILLER_169_2276 ();
 b15zdnd11an1n16x5 FILLER_170_8 ();
 b15zdnd00an1n02x5 FILLER_170_24 ();
 b15zdnd11an1n16x5 FILLER_170_33 ();
 b15zdnd11an1n04x5 FILLER_170_49 ();
 b15zdnd11an1n04x5 FILLER_170_59 ();
 b15zdnd00an1n01x5 FILLER_170_63 ();
 b15zdnd11an1n04x5 FILLER_170_73 ();
 b15zdnd00an1n02x5 FILLER_170_77 ();
 b15zdnd11an1n08x5 FILLER_170_83 ();
 b15zdnd11an1n16x5 FILLER_170_105 ();
 b15zdnd11an1n64x5 FILLER_170_130 ();
 b15zdnd11an1n16x5 FILLER_170_194 ();
 b15zdnd11an1n64x5 FILLER_170_215 ();
 b15zdnd11an1n32x5 FILLER_170_279 ();
 b15zdnd11an1n16x5 FILLER_170_311 ();
 b15zdnd00an1n02x5 FILLER_170_327 ();
 b15zdnd00an1n01x5 FILLER_170_329 ();
 b15zdnd11an1n32x5 FILLER_170_343 ();
 b15zdnd11an1n16x5 FILLER_170_375 ();
 b15zdnd11an1n08x5 FILLER_170_391 ();
 b15zdnd00an1n02x5 FILLER_170_399 ();
 b15zdnd00an1n01x5 FILLER_170_401 ();
 b15zdnd11an1n32x5 FILLER_170_408 ();
 b15zdnd11an1n16x5 FILLER_170_440 ();
 b15zdnd00an1n02x5 FILLER_170_456 ();
 b15zdnd11an1n16x5 FILLER_170_478 ();
 b15zdnd11an1n04x5 FILLER_170_494 ();
 b15zdnd11an1n04x5 FILLER_170_510 ();
 b15zdnd11an1n64x5 FILLER_170_520 ();
 b15zdnd11an1n16x5 FILLER_170_584 ();
 b15zdnd11an1n08x5 FILLER_170_600 ();
 b15zdnd00an1n02x5 FILLER_170_608 ();
 b15zdnd11an1n16x5 FILLER_170_623 ();
 b15zdnd00an1n02x5 FILLER_170_639 ();
 b15zdnd11an1n04x5 FILLER_170_646 ();
 b15zdnd11an1n16x5 FILLER_170_657 ();
 b15zdnd00an1n02x5 FILLER_170_673 ();
 b15zdnd11an1n08x5 FILLER_170_690 ();
 b15zdnd11an1n04x5 FILLER_170_698 ();
 b15zdnd11an1n08x5 FILLER_170_709 ();
 b15zdnd00an1n01x5 FILLER_170_717 ();
 b15zdnd11an1n16x5 FILLER_170_726 ();
 b15zdnd11an1n08x5 FILLER_170_742 ();
 b15zdnd11an1n04x5 FILLER_170_750 ();
 b15zdnd11an1n64x5 FILLER_170_758 ();
 b15zdnd11an1n32x5 FILLER_170_822 ();
 b15zdnd11an1n16x5 FILLER_170_854 ();
 b15zdnd11an1n08x5 FILLER_170_870 ();
 b15zdnd00an1n01x5 FILLER_170_878 ();
 b15zdnd11an1n32x5 FILLER_170_891 ();
 b15zdnd11an1n04x5 FILLER_170_923 ();
 b15zdnd00an1n02x5 FILLER_170_927 ();
 b15zdnd11an1n16x5 FILLER_170_933 ();
 b15zdnd11an1n08x5 FILLER_170_949 ();
 b15zdnd11an1n32x5 FILLER_170_973 ();
 b15zdnd11an1n04x5 FILLER_170_1005 ();
 b15zdnd00an1n02x5 FILLER_170_1009 ();
 b15zdnd00an1n01x5 FILLER_170_1011 ();
 b15zdnd11an1n32x5 FILLER_170_1024 ();
 b15zdnd00an1n02x5 FILLER_170_1056 ();
 b15zdnd11an1n04x5 FILLER_170_1070 ();
 b15zdnd11an1n64x5 FILLER_170_1090 ();
 b15zdnd00an1n02x5 FILLER_170_1154 ();
 b15zdnd11an1n04x5 FILLER_170_1160 ();
 b15zdnd11an1n04x5 FILLER_170_1170 ();
 b15zdnd11an1n16x5 FILLER_170_1180 ();
 b15zdnd00an1n02x5 FILLER_170_1196 ();
 b15zdnd11an1n64x5 FILLER_170_1204 ();
 b15zdnd11an1n64x5 FILLER_170_1268 ();
 b15zdnd11an1n16x5 FILLER_170_1332 ();
 b15zdnd11an1n32x5 FILLER_170_1362 ();
 b15zdnd00an1n02x5 FILLER_170_1394 ();
 b15zdnd00an1n01x5 FILLER_170_1396 ();
 b15zdnd11an1n32x5 FILLER_170_1406 ();
 b15zdnd11an1n04x5 FILLER_170_1438 ();
 b15zdnd00an1n01x5 FILLER_170_1442 ();
 b15zdnd11an1n08x5 FILLER_170_1450 ();
 b15zdnd11an1n64x5 FILLER_170_1478 ();
 b15zdnd11an1n64x5 FILLER_170_1542 ();
 b15zdnd11an1n64x5 FILLER_170_1606 ();
 b15zdnd11an1n64x5 FILLER_170_1670 ();
 b15zdnd11an1n32x5 FILLER_170_1734 ();
 b15zdnd11an1n16x5 FILLER_170_1766 ();
 b15zdnd00an1n02x5 FILLER_170_1782 ();
 b15zdnd11an1n08x5 FILLER_170_1803 ();
 b15zdnd00an1n02x5 FILLER_170_1811 ();
 b15zdnd00an1n01x5 FILLER_170_1813 ();
 b15zdnd11an1n64x5 FILLER_170_1834 ();
 b15zdnd11an1n64x5 FILLER_170_1898 ();
 b15zdnd11an1n64x5 FILLER_170_1962 ();
 b15zdnd11an1n32x5 FILLER_170_2026 ();
 b15zdnd11an1n16x5 FILLER_170_2058 ();
 b15zdnd11an1n04x5 FILLER_170_2074 ();
 b15zdnd00an1n02x5 FILLER_170_2078 ();
 b15zdnd11an1n04x5 FILLER_170_2090 ();
 b15zdnd11an1n04x5 FILLER_170_2112 ();
 b15zdnd11an1n16x5 FILLER_170_2134 ();
 b15zdnd11an1n04x5 FILLER_170_2150 ();
 b15zdnd11an1n16x5 FILLER_170_2162 ();
 b15zdnd11an1n08x5 FILLER_170_2178 ();
 b15zdnd11an1n04x5 FILLER_170_2186 ();
 b15zdnd11an1n64x5 FILLER_170_2210 ();
 b15zdnd00an1n02x5 FILLER_170_2274 ();
 b15zdnd11an1n64x5 FILLER_171_0 ();
 b15zdnd11an1n64x5 FILLER_171_64 ();
 b15zdnd11an1n32x5 FILLER_171_128 ();
 b15zdnd11an1n16x5 FILLER_171_160 ();
 b15zdnd11an1n04x5 FILLER_171_176 ();
 b15zdnd00an1n01x5 FILLER_171_180 ();
 b15zdnd11an1n16x5 FILLER_171_186 ();
 b15zdnd11an1n04x5 FILLER_171_202 ();
 b15zdnd00an1n02x5 FILLER_171_206 ();
 b15zdnd00an1n01x5 FILLER_171_208 ();
 b15zdnd11an1n16x5 FILLER_171_214 ();
 b15zdnd11an1n08x5 FILLER_171_230 ();
 b15zdnd00an1n02x5 FILLER_171_238 ();
 b15zdnd00an1n01x5 FILLER_171_240 ();
 b15zdnd11an1n04x5 FILLER_171_253 ();
 b15zdnd00an1n02x5 FILLER_171_257 ();
 b15zdnd11an1n08x5 FILLER_171_279 ();
 b15zdnd11an1n04x5 FILLER_171_293 ();
 b15zdnd11an1n64x5 FILLER_171_303 ();
 b15zdnd11an1n32x5 FILLER_171_367 ();
 b15zdnd11an1n16x5 FILLER_171_399 ();
 b15zdnd11an1n08x5 FILLER_171_415 ();
 b15zdnd11an1n04x5 FILLER_171_423 ();
 b15zdnd00an1n02x5 FILLER_171_427 ();
 b15zdnd00an1n01x5 FILLER_171_429 ();
 b15zdnd11an1n04x5 FILLER_171_436 ();
 b15zdnd11an1n04x5 FILLER_171_447 ();
 b15zdnd11an1n32x5 FILLER_171_457 ();
 b15zdnd11an1n16x5 FILLER_171_489 ();
 b15zdnd11an1n08x5 FILLER_171_505 ();
 b15zdnd00an1n02x5 FILLER_171_513 ();
 b15zdnd00an1n01x5 FILLER_171_515 ();
 b15zdnd11an1n64x5 FILLER_171_523 ();
 b15zdnd11an1n32x5 FILLER_171_587 ();
 b15zdnd11an1n16x5 FILLER_171_619 ();
 b15zdnd00an1n01x5 FILLER_171_635 ();
 b15zdnd11an1n04x5 FILLER_171_642 ();
 b15zdnd11an1n04x5 FILLER_171_674 ();
 b15zdnd00an1n02x5 FILLER_171_678 ();
 b15zdnd00an1n01x5 FILLER_171_680 ();
 b15zdnd11an1n16x5 FILLER_171_686 ();
 b15zdnd00an1n02x5 FILLER_171_702 ();
 b15zdnd11an1n04x5 FILLER_171_716 ();
 b15zdnd11an1n64x5 FILLER_171_729 ();
 b15zdnd11an1n32x5 FILLER_171_793 ();
 b15zdnd11an1n08x5 FILLER_171_825 ();
 b15zdnd11an1n04x5 FILLER_171_833 ();
 b15zdnd00an1n02x5 FILLER_171_837 ();
 b15zdnd11an1n32x5 FILLER_171_845 ();
 b15zdnd11an1n16x5 FILLER_171_890 ();
 b15zdnd00an1n02x5 FILLER_171_906 ();
 b15zdnd00an1n01x5 FILLER_171_908 ();
 b15zdnd11an1n04x5 FILLER_171_913 ();
 b15zdnd11an1n64x5 FILLER_171_930 ();
 b15zdnd11an1n64x5 FILLER_171_994 ();
 b15zdnd00an1n01x5 FILLER_171_1058 ();
 b15zdnd11an1n64x5 FILLER_171_1066 ();
 b15zdnd11an1n32x5 FILLER_171_1130 ();
 b15zdnd11an1n16x5 FILLER_171_1162 ();
 b15zdnd11an1n08x5 FILLER_171_1178 ();
 b15zdnd11an1n04x5 FILLER_171_1186 ();
 b15zdnd11an1n32x5 FILLER_171_1222 ();
 b15zdnd11an1n16x5 FILLER_171_1254 ();
 b15zdnd11an1n08x5 FILLER_171_1270 ();
 b15zdnd11an1n04x5 FILLER_171_1278 ();
 b15zdnd00an1n02x5 FILLER_171_1282 ();
 b15zdnd11an1n04x5 FILLER_171_1302 ();
 b15zdnd11an1n64x5 FILLER_171_1332 ();
 b15zdnd11an1n64x5 FILLER_171_1396 ();
 b15zdnd11an1n32x5 FILLER_171_1460 ();
 b15zdnd11an1n08x5 FILLER_171_1492 ();
 b15zdnd00an1n02x5 FILLER_171_1500 ();
 b15zdnd11an1n32x5 FILLER_171_1506 ();
 b15zdnd11an1n08x5 FILLER_171_1538 ();
 b15zdnd11an1n04x5 FILLER_171_1546 ();
 b15zdnd00an1n02x5 FILLER_171_1550 ();
 b15zdnd00an1n01x5 FILLER_171_1552 ();
 b15zdnd11an1n08x5 FILLER_171_1557 ();
 b15zdnd00an1n01x5 FILLER_171_1565 ();
 b15zdnd11an1n32x5 FILLER_171_1572 ();
 b15zdnd11an1n08x5 FILLER_171_1604 ();
 b15zdnd11an1n04x5 FILLER_171_1612 ();
 b15zdnd00an1n02x5 FILLER_171_1616 ();
 b15zdnd11an1n04x5 FILLER_171_1631 ();
 b15zdnd11an1n64x5 FILLER_171_1661 ();
 b15zdnd11an1n32x5 FILLER_171_1725 ();
 b15zdnd11an1n08x5 FILLER_171_1757 ();
 b15zdnd11an1n04x5 FILLER_171_1765 ();
 b15zdnd00an1n02x5 FILLER_171_1769 ();
 b15zdnd11an1n16x5 FILLER_171_1797 ();
 b15zdnd11an1n04x5 FILLER_171_1813 ();
 b15zdnd00an1n01x5 FILLER_171_1817 ();
 b15zdnd11an1n64x5 FILLER_171_1823 ();
 b15zdnd11an1n64x5 FILLER_171_1887 ();
 b15zdnd11an1n32x5 FILLER_171_1951 ();
 b15zdnd11an1n08x5 FILLER_171_2009 ();
 b15zdnd11an1n04x5 FILLER_171_2017 ();
 b15zdnd00an1n02x5 FILLER_171_2021 ();
 b15zdnd11an1n04x5 FILLER_171_2054 ();
 b15zdnd11an1n16x5 FILLER_171_2067 ();
 b15zdnd11an1n04x5 FILLER_171_2083 ();
 b15zdnd00an1n01x5 FILLER_171_2087 ();
 b15zdnd11an1n16x5 FILLER_171_2112 ();
 b15zdnd11an1n04x5 FILLER_171_2128 ();
 b15zdnd00an1n01x5 FILLER_171_2132 ();
 b15zdnd11an1n32x5 FILLER_171_2148 ();
 b15zdnd11an1n08x5 FILLER_171_2180 ();
 b15zdnd11an1n04x5 FILLER_171_2188 ();
 b15zdnd00an1n01x5 FILLER_171_2192 ();
 b15zdnd11an1n32x5 FILLER_171_2197 ();
 b15zdnd11an1n16x5 FILLER_171_2229 ();
 b15zdnd11an1n16x5 FILLER_171_2249 ();
 b15zdnd11an1n04x5 FILLER_171_2265 ();
 b15zdnd00an1n01x5 FILLER_171_2269 ();
 b15zdnd11an1n04x5 FILLER_171_2274 ();
 b15zdnd00an1n02x5 FILLER_171_2282 ();
 b15zdnd11an1n64x5 FILLER_172_8 ();
 b15zdnd11an1n32x5 FILLER_172_72 ();
 b15zdnd11an1n08x5 FILLER_172_104 ();
 b15zdnd00an1n02x5 FILLER_172_112 ();
 b15zdnd11an1n16x5 FILLER_172_123 ();
 b15zdnd11an1n04x5 FILLER_172_139 ();
 b15zdnd00an1n02x5 FILLER_172_143 ();
 b15zdnd11an1n16x5 FILLER_172_158 ();
 b15zdnd00an1n02x5 FILLER_172_174 ();
 b15zdnd11an1n16x5 FILLER_172_182 ();
 b15zdnd11an1n04x5 FILLER_172_198 ();
 b15zdnd11an1n16x5 FILLER_172_207 ();
 b15zdnd11an1n08x5 FILLER_172_223 ();
 b15zdnd11an1n04x5 FILLER_172_231 ();
 b15zdnd11an1n04x5 FILLER_172_246 ();
 b15zdnd00an1n02x5 FILLER_172_250 ();
 b15zdnd11an1n08x5 FILLER_172_272 ();
 b15zdnd11an1n04x5 FILLER_172_280 ();
 b15zdnd00an1n02x5 FILLER_172_284 ();
 b15zdnd11an1n64x5 FILLER_172_302 ();
 b15zdnd11an1n32x5 FILLER_172_366 ();
 b15zdnd11an1n64x5 FILLER_172_405 ();
 b15zdnd11an1n16x5 FILLER_172_469 ();
 b15zdnd11an1n08x5 FILLER_172_485 ();
 b15zdnd00an1n02x5 FILLER_172_493 ();
 b15zdnd11an1n32x5 FILLER_172_516 ();
 b15zdnd11an1n08x5 FILLER_172_548 ();
 b15zdnd11an1n04x5 FILLER_172_556 ();
 b15zdnd11an1n08x5 FILLER_172_565 ();
 b15zdnd11an1n04x5 FILLER_172_573 ();
 b15zdnd11an1n64x5 FILLER_172_591 ();
 b15zdnd11an1n16x5 FILLER_172_655 ();
 b15zdnd11an1n04x5 FILLER_172_671 ();
 b15zdnd00an1n02x5 FILLER_172_675 ();
 b15zdnd00an1n01x5 FILLER_172_677 ();
 b15zdnd11an1n16x5 FILLER_172_687 ();
 b15zdnd11an1n08x5 FILLER_172_703 ();
 b15zdnd11an1n04x5 FILLER_172_711 ();
 b15zdnd00an1n02x5 FILLER_172_715 ();
 b15zdnd00an1n01x5 FILLER_172_717 ();
 b15zdnd11an1n04x5 FILLER_172_726 ();
 b15zdnd00an1n02x5 FILLER_172_730 ();
 b15zdnd11an1n08x5 FILLER_172_752 ();
 b15zdnd11an1n04x5 FILLER_172_780 ();
 b15zdnd11an1n32x5 FILLER_172_789 ();
 b15zdnd11an1n16x5 FILLER_172_821 ();
 b15zdnd00an1n01x5 FILLER_172_837 ();
 b15zdnd11an1n16x5 FILLER_172_842 ();
 b15zdnd11an1n04x5 FILLER_172_858 ();
 b15zdnd00an1n02x5 FILLER_172_862 ();
 b15zdnd11an1n32x5 FILLER_172_876 ();
 b15zdnd11an1n16x5 FILLER_172_908 ();
 b15zdnd11an1n04x5 FILLER_172_924 ();
 b15zdnd00an1n02x5 FILLER_172_928 ();
 b15zdnd11an1n04x5 FILLER_172_935 ();
 b15zdnd00an1n02x5 FILLER_172_939 ();
 b15zdnd00an1n01x5 FILLER_172_941 ();
 b15zdnd11an1n32x5 FILLER_172_954 ();
 b15zdnd00an1n01x5 FILLER_172_986 ();
 b15zdnd11an1n04x5 FILLER_172_992 ();
 b15zdnd11an1n08x5 FILLER_172_1000 ();
 b15zdnd00an1n02x5 FILLER_172_1008 ();
 b15zdnd11an1n04x5 FILLER_172_1016 ();
 b15zdnd11an1n64x5 FILLER_172_1024 ();
 b15zdnd11an1n32x5 FILLER_172_1088 ();
 b15zdnd11an1n08x5 FILLER_172_1120 ();
 b15zdnd11an1n04x5 FILLER_172_1128 ();
 b15zdnd00an1n02x5 FILLER_172_1132 ();
 b15zdnd11an1n64x5 FILLER_172_1138 ();
 b15zdnd00an1n01x5 FILLER_172_1202 ();
 b15zdnd11an1n32x5 FILLER_172_1217 ();
 b15zdnd11an1n16x5 FILLER_172_1249 ();
 b15zdnd11an1n08x5 FILLER_172_1285 ();
 b15zdnd11an1n16x5 FILLER_172_1317 ();
 b15zdnd11an1n08x5 FILLER_172_1333 ();
 b15zdnd11an1n04x5 FILLER_172_1341 ();
 b15zdnd11an1n16x5 FILLER_172_1360 ();
 b15zdnd00an1n01x5 FILLER_172_1376 ();
 b15zdnd11an1n04x5 FILLER_172_1389 ();
 b15zdnd11an1n04x5 FILLER_172_1418 ();
 b15zdnd11an1n32x5 FILLER_172_1426 ();
 b15zdnd11an1n32x5 FILLER_172_1463 ();
 b15zdnd00an1n01x5 FILLER_172_1495 ();
 b15zdnd11an1n04x5 FILLER_172_1500 ();
 b15zdnd11an1n04x5 FILLER_172_1513 ();
 b15zdnd11an1n16x5 FILLER_172_1533 ();
 b15zdnd00an1n02x5 FILLER_172_1549 ();
 b15zdnd00an1n01x5 FILLER_172_1551 ();
 b15zdnd11an1n04x5 FILLER_172_1562 ();
 b15zdnd00an1n02x5 FILLER_172_1566 ();
 b15zdnd11an1n04x5 FILLER_172_1573 ();
 b15zdnd11an1n16x5 FILLER_172_1586 ();
 b15zdnd00an1n02x5 FILLER_172_1602 ();
 b15zdnd00an1n01x5 FILLER_172_1604 ();
 b15zdnd11an1n16x5 FILLER_172_1611 ();
 b15zdnd11an1n08x5 FILLER_172_1627 ();
 b15zdnd11an1n64x5 FILLER_172_1661 ();
 b15zdnd11an1n32x5 FILLER_172_1725 ();
 b15zdnd11an1n04x5 FILLER_172_1757 ();
 b15zdnd11an1n32x5 FILLER_172_1772 ();
 b15zdnd11an1n08x5 FILLER_172_1804 ();
 b15zdnd00an1n01x5 FILLER_172_1812 ();
 b15zdnd11an1n16x5 FILLER_172_1819 ();
 b15zdnd11an1n08x5 FILLER_172_1835 ();
 b15zdnd11an1n04x5 FILLER_172_1843 ();
 b15zdnd00an1n01x5 FILLER_172_1847 ();
 b15zdnd11an1n16x5 FILLER_172_1853 ();
 b15zdnd11an1n08x5 FILLER_172_1869 ();
 b15zdnd11an1n04x5 FILLER_172_1877 ();
 b15zdnd00an1n01x5 FILLER_172_1881 ();
 b15zdnd11an1n32x5 FILLER_172_1886 ();
 b15zdnd00an1n01x5 FILLER_172_1918 ();
 b15zdnd11an1n04x5 FILLER_172_1923 ();
 b15zdnd11an1n16x5 FILLER_172_1947 ();
 b15zdnd11an1n08x5 FILLER_172_1963 ();
 b15zdnd00an1n02x5 FILLER_172_1971 ();
 b15zdnd00an1n01x5 FILLER_172_1973 ();
 b15zdnd11an1n32x5 FILLER_172_1985 ();
 b15zdnd11an1n08x5 FILLER_172_2017 ();
 b15zdnd00an1n02x5 FILLER_172_2025 ();
 b15zdnd11an1n64x5 FILLER_172_2045 ();
 b15zdnd00an1n02x5 FILLER_172_2109 ();
 b15zdnd00an1n01x5 FILLER_172_2111 ();
 b15zdnd11an1n04x5 FILLER_172_2132 ();
 b15zdnd11an1n04x5 FILLER_172_2147 ();
 b15zdnd00an1n02x5 FILLER_172_2151 ();
 b15zdnd00an1n01x5 FILLER_172_2153 ();
 b15zdnd11an1n64x5 FILLER_172_2162 ();
 b15zdnd00an1n02x5 FILLER_172_2226 ();
 b15zdnd00an1n01x5 FILLER_172_2228 ();
 b15zdnd11an1n04x5 FILLER_172_2232 ();
 b15zdnd11an1n08x5 FILLER_172_2239 ();
 b15zdnd00an1n02x5 FILLER_172_2247 ();
 b15zdnd00an1n01x5 FILLER_172_2249 ();
 b15zdnd11an1n04x5 FILLER_172_2261 ();
 b15zdnd11an1n04x5 FILLER_172_2269 ();
 b15zdnd00an1n02x5 FILLER_172_2273 ();
 b15zdnd00an1n01x5 FILLER_172_2275 ();
 b15zdnd11an1n16x5 FILLER_173_0 ();
 b15zdnd11an1n04x5 FILLER_173_16 ();
 b15zdnd00an1n01x5 FILLER_173_20 ();
 b15zdnd11an1n32x5 FILLER_173_25 ();
 b15zdnd11an1n08x5 FILLER_173_57 ();
 b15zdnd00an1n02x5 FILLER_173_65 ();
 b15zdnd00an1n01x5 FILLER_173_67 ();
 b15zdnd11an1n16x5 FILLER_173_73 ();
 b15zdnd11an1n08x5 FILLER_173_89 ();
 b15zdnd11an1n04x5 FILLER_173_97 ();
 b15zdnd00an1n01x5 FILLER_173_101 ();
 b15zdnd11an1n08x5 FILLER_173_132 ();
 b15zdnd11an1n04x5 FILLER_173_140 ();
 b15zdnd00an1n02x5 FILLER_173_144 ();
 b15zdnd00an1n01x5 FILLER_173_146 ();
 b15zdnd11an1n08x5 FILLER_173_167 ();
 b15zdnd00an1n02x5 FILLER_173_175 ();
 b15zdnd11an1n04x5 FILLER_173_198 ();
 b15zdnd11an1n32x5 FILLER_173_208 ();
 b15zdnd11an1n16x5 FILLER_173_240 ();
 b15zdnd00an1n02x5 FILLER_173_256 ();
 b15zdnd00an1n01x5 FILLER_173_258 ();
 b15zdnd11an1n64x5 FILLER_173_281 ();
 b15zdnd11an1n32x5 FILLER_173_345 ();
 b15zdnd11an1n16x5 FILLER_173_377 ();
 b15zdnd11an1n04x5 FILLER_173_393 ();
 b15zdnd11an1n04x5 FILLER_173_409 ();
 b15zdnd00an1n01x5 FILLER_173_413 ();
 b15zdnd11an1n04x5 FILLER_173_430 ();
 b15zdnd11an1n64x5 FILLER_173_440 ();
 b15zdnd11an1n32x5 FILLER_173_504 ();
 b15zdnd11an1n04x5 FILLER_173_536 ();
 b15zdnd00an1n01x5 FILLER_173_540 ();
 b15zdnd11an1n08x5 FILLER_173_547 ();
 b15zdnd11an1n04x5 FILLER_173_555 ();
 b15zdnd11an1n16x5 FILLER_173_566 ();
 b15zdnd11an1n16x5 FILLER_173_587 ();
 b15zdnd00an1n02x5 FILLER_173_603 ();
 b15zdnd00an1n01x5 FILLER_173_605 ();
 b15zdnd11an1n04x5 FILLER_173_612 ();
 b15zdnd11an1n64x5 FILLER_173_620 ();
 b15zdnd11an1n32x5 FILLER_173_684 ();
 b15zdnd11an1n16x5 FILLER_173_716 ();
 b15zdnd11an1n08x5 FILLER_173_732 ();
 b15zdnd00an1n01x5 FILLER_173_740 ();
 b15zdnd11an1n04x5 FILLER_173_756 ();
 b15zdnd11an1n04x5 FILLER_173_772 ();
 b15zdnd11an1n64x5 FILLER_173_782 ();
 b15zdnd11an1n32x5 FILLER_173_846 ();
 b15zdnd11an1n08x5 FILLER_173_878 ();
 b15zdnd00an1n02x5 FILLER_173_886 ();
 b15zdnd00an1n01x5 FILLER_173_888 ();
 b15zdnd11an1n04x5 FILLER_173_912 ();
 b15zdnd11an1n16x5 FILLER_173_927 ();
 b15zdnd00an1n02x5 FILLER_173_943 ();
 b15zdnd00an1n01x5 FILLER_173_945 ();
 b15zdnd11an1n16x5 FILLER_173_958 ();
 b15zdnd11an1n08x5 FILLER_173_974 ();
 b15zdnd00an1n02x5 FILLER_173_982 ();
 b15zdnd00an1n01x5 FILLER_173_984 ();
 b15zdnd11an1n32x5 FILLER_173_999 ();
 b15zdnd11an1n16x5 FILLER_173_1031 ();
 b15zdnd11an1n08x5 FILLER_173_1047 ();
 b15zdnd11an1n04x5 FILLER_173_1055 ();
 b15zdnd00an1n01x5 FILLER_173_1059 ();
 b15zdnd11an1n08x5 FILLER_173_1068 ();
 b15zdnd00an1n01x5 FILLER_173_1076 ();
 b15zdnd11an1n04x5 FILLER_173_1083 ();
 b15zdnd11an1n16x5 FILLER_173_1093 ();
 b15zdnd00an1n02x5 FILLER_173_1109 ();
 b15zdnd11an1n16x5 FILLER_173_1122 ();
 b15zdnd11an1n04x5 FILLER_173_1143 ();
 b15zdnd11an1n16x5 FILLER_173_1153 ();
 b15zdnd11an1n04x5 FILLER_173_1169 ();
 b15zdnd11an1n64x5 FILLER_173_1179 ();
 b15zdnd11an1n32x5 FILLER_173_1243 ();
 b15zdnd00an1n02x5 FILLER_173_1275 ();
 b15zdnd11an1n04x5 FILLER_173_1281 ();
 b15zdnd11an1n16x5 FILLER_173_1291 ();
 b15zdnd11an1n04x5 FILLER_173_1307 ();
 b15zdnd00an1n01x5 FILLER_173_1311 ();
 b15zdnd11an1n04x5 FILLER_173_1332 ();
 b15zdnd00an1n02x5 FILLER_173_1336 ();
 b15zdnd00an1n01x5 FILLER_173_1338 ();
 b15zdnd11an1n16x5 FILLER_173_1358 ();
 b15zdnd11an1n08x5 FILLER_173_1374 ();
 b15zdnd00an1n02x5 FILLER_173_1382 ();
 b15zdnd00an1n01x5 FILLER_173_1384 ();
 b15zdnd11an1n16x5 FILLER_173_1392 ();
 b15zdnd11an1n08x5 FILLER_173_1414 ();
 b15zdnd11an1n08x5 FILLER_173_1434 ();
 b15zdnd11an1n08x5 FILLER_173_1446 ();
 b15zdnd11an1n04x5 FILLER_173_1454 ();
 b15zdnd00an1n02x5 FILLER_173_1458 ();
 b15zdnd00an1n01x5 FILLER_173_1460 ();
 b15zdnd11an1n16x5 FILLER_173_1468 ();
 b15zdnd00an1n02x5 FILLER_173_1484 ();
 b15zdnd11an1n04x5 FILLER_173_1490 ();
 b15zdnd00an1n02x5 FILLER_173_1494 ();
 b15zdnd00an1n01x5 FILLER_173_1496 ();
 b15zdnd11an1n32x5 FILLER_173_1505 ();
 b15zdnd11an1n16x5 FILLER_173_1537 ();
 b15zdnd00an1n01x5 FILLER_173_1553 ();
 b15zdnd11an1n16x5 FILLER_173_1561 ();
 b15zdnd11an1n08x5 FILLER_173_1577 ();
 b15zdnd11an1n04x5 FILLER_173_1585 ();
 b15zdnd11an1n08x5 FILLER_173_1605 ();
 b15zdnd00an1n02x5 FILLER_173_1613 ();
 b15zdnd00an1n01x5 FILLER_173_1615 ();
 b15zdnd11an1n16x5 FILLER_173_1626 ();
 b15zdnd11an1n04x5 FILLER_173_1642 ();
 b15zdnd00an1n02x5 FILLER_173_1646 ();
 b15zdnd00an1n01x5 FILLER_173_1648 ();
 b15zdnd11an1n16x5 FILLER_173_1657 ();
 b15zdnd11an1n04x5 FILLER_173_1673 ();
 b15zdnd00an1n01x5 FILLER_173_1677 ();
 b15zdnd11an1n64x5 FILLER_173_1694 ();
 b15zdnd11an1n16x5 FILLER_173_1758 ();
 b15zdnd00an1n02x5 FILLER_173_1774 ();
 b15zdnd11an1n32x5 FILLER_173_1796 ();
 b15zdnd11an1n16x5 FILLER_173_1828 ();
 b15zdnd00an1n02x5 FILLER_173_1844 ();
 b15zdnd11an1n08x5 FILLER_173_1866 ();
 b15zdnd11an1n04x5 FILLER_173_1874 ();
 b15zdnd11an1n16x5 FILLER_173_1889 ();
 b15zdnd11an1n08x5 FILLER_173_1905 ();
 b15zdnd11an1n04x5 FILLER_173_1913 ();
 b15zdnd11an1n04x5 FILLER_173_1924 ();
 b15zdnd11an1n32x5 FILLER_173_1937 ();
 b15zdnd11an1n16x5 FILLER_173_1989 ();
 b15zdnd11an1n08x5 FILLER_173_2005 ();
 b15zdnd11an1n04x5 FILLER_173_2013 ();
 b15zdnd00an1n02x5 FILLER_173_2017 ();
 b15zdnd11an1n08x5 FILLER_173_2031 ();
 b15zdnd00an1n02x5 FILLER_173_2039 ();
 b15zdnd11an1n64x5 FILLER_173_2051 ();
 b15zdnd11an1n16x5 FILLER_173_2115 ();
 b15zdnd11an1n08x5 FILLER_173_2131 ();
 b15zdnd11an1n04x5 FILLER_173_2139 ();
 b15zdnd00an1n02x5 FILLER_173_2143 ();
 b15zdnd00an1n01x5 FILLER_173_2145 ();
 b15zdnd11an1n32x5 FILLER_173_2164 ();
 b15zdnd11an1n16x5 FILLER_173_2196 ();
 b15zdnd11an1n08x5 FILLER_173_2212 ();
 b15zdnd00an1n02x5 FILLER_173_2220 ();
 b15zdnd11an1n04x5 FILLER_173_2242 ();
 b15zdnd00an1n01x5 FILLER_173_2246 ();
 b15zdnd11an1n32x5 FILLER_173_2251 ();
 b15zdnd00an1n01x5 FILLER_173_2283 ();
 b15zdnd11an1n16x5 FILLER_174_8 ();
 b15zdnd11an1n08x5 FILLER_174_24 ();
 b15zdnd11an1n04x5 FILLER_174_32 ();
 b15zdnd11an1n16x5 FILLER_174_46 ();
 b15zdnd11an1n04x5 FILLER_174_62 ();
 b15zdnd00an1n01x5 FILLER_174_66 ();
 b15zdnd11an1n16x5 FILLER_174_75 ();
 b15zdnd11an1n08x5 FILLER_174_91 ();
 b15zdnd00an1n01x5 FILLER_174_99 ();
 b15zdnd11an1n16x5 FILLER_174_123 ();
 b15zdnd11an1n08x5 FILLER_174_139 ();
 b15zdnd11an1n04x5 FILLER_174_157 ();
 b15zdnd11an1n16x5 FILLER_174_167 ();
 b15zdnd11an1n08x5 FILLER_174_183 ();
 b15zdnd00an1n01x5 FILLER_174_191 ();
 b15zdnd11an1n64x5 FILLER_174_199 ();
 b15zdnd11an1n32x5 FILLER_174_263 ();
 b15zdnd11an1n04x5 FILLER_174_295 ();
 b15zdnd00an1n01x5 FILLER_174_299 ();
 b15zdnd11an1n04x5 FILLER_174_321 ();
 b15zdnd11an1n64x5 FILLER_174_331 ();
 b15zdnd11an1n04x5 FILLER_174_395 ();
 b15zdnd00an1n02x5 FILLER_174_399 ();
 b15zdnd11an1n64x5 FILLER_174_406 ();
 b15zdnd11an1n04x5 FILLER_174_470 ();
 b15zdnd00an1n01x5 FILLER_174_474 ();
 b15zdnd11an1n04x5 FILLER_174_482 ();
 b15zdnd11an1n16x5 FILLER_174_492 ();
 b15zdnd11an1n08x5 FILLER_174_508 ();
 b15zdnd00an1n02x5 FILLER_174_516 ();
 b15zdnd00an1n01x5 FILLER_174_518 ();
 b15zdnd11an1n16x5 FILLER_174_524 ();
 b15zdnd00an1n02x5 FILLER_174_540 ();
 b15zdnd11an1n04x5 FILLER_174_547 ();
 b15zdnd11an1n64x5 FILLER_174_567 ();
 b15zdnd11an1n08x5 FILLER_174_631 ();
 b15zdnd11an1n04x5 FILLER_174_639 ();
 b15zdnd00an1n01x5 FILLER_174_643 ();
 b15zdnd11an1n64x5 FILLER_174_648 ();
 b15zdnd11an1n04x5 FILLER_174_712 ();
 b15zdnd00an1n02x5 FILLER_174_716 ();
 b15zdnd11an1n08x5 FILLER_174_726 ();
 b15zdnd00an1n02x5 FILLER_174_734 ();
 b15zdnd00an1n01x5 FILLER_174_736 ();
 b15zdnd11an1n64x5 FILLER_174_747 ();
 b15zdnd11an1n32x5 FILLER_174_811 ();
 b15zdnd11an1n16x5 FILLER_174_843 ();
 b15zdnd11an1n08x5 FILLER_174_859 ();
 b15zdnd11an1n04x5 FILLER_174_867 ();
 b15zdnd00an1n01x5 FILLER_174_871 ();
 b15zdnd11an1n64x5 FILLER_174_878 ();
 b15zdnd00an1n02x5 FILLER_174_942 ();
 b15zdnd00an1n01x5 FILLER_174_944 ();
 b15zdnd11an1n32x5 FILLER_174_949 ();
 b15zdnd11an1n16x5 FILLER_174_981 ();
 b15zdnd11an1n08x5 FILLER_174_997 ();
 b15zdnd11an1n04x5 FILLER_174_1005 ();
 b15zdnd00an1n02x5 FILLER_174_1009 ();
 b15zdnd00an1n01x5 FILLER_174_1011 ();
 b15zdnd11an1n04x5 FILLER_174_1018 ();
 b15zdnd11an1n16x5 FILLER_174_1030 ();
 b15zdnd11an1n08x5 FILLER_174_1046 ();
 b15zdnd11an1n04x5 FILLER_174_1054 ();
 b15zdnd00an1n02x5 FILLER_174_1058 ();
 b15zdnd11an1n08x5 FILLER_174_1065 ();
 b15zdnd11an1n04x5 FILLER_174_1073 ();
 b15zdnd11an1n64x5 FILLER_174_1081 ();
 b15zdnd00an1n02x5 FILLER_174_1145 ();
 b15zdnd00an1n01x5 FILLER_174_1147 ();
 b15zdnd11an1n16x5 FILLER_174_1155 ();
 b15zdnd11an1n04x5 FILLER_174_1171 ();
 b15zdnd00an1n02x5 FILLER_174_1175 ();
 b15zdnd11an1n04x5 FILLER_174_1184 ();
 b15zdnd11an1n04x5 FILLER_174_1192 ();
 b15zdnd00an1n02x5 FILLER_174_1196 ();
 b15zdnd11an1n64x5 FILLER_174_1204 ();
 b15zdnd11an1n16x5 FILLER_174_1268 ();
 b15zdnd00an1n02x5 FILLER_174_1284 ();
 b15zdnd11an1n04x5 FILLER_174_1312 ();
 b15zdnd11an1n04x5 FILLER_174_1322 ();
 b15zdnd11an1n32x5 FILLER_174_1344 ();
 b15zdnd11an1n04x5 FILLER_174_1376 ();
 b15zdnd00an1n02x5 FILLER_174_1380 ();
 b15zdnd00an1n01x5 FILLER_174_1382 ();
 b15zdnd11an1n32x5 FILLER_174_1393 ();
 b15zdnd11an1n08x5 FILLER_174_1425 ();
 b15zdnd11an1n04x5 FILLER_174_1433 ();
 b15zdnd00an1n02x5 FILLER_174_1437 ();
 b15zdnd11an1n08x5 FILLER_174_1446 ();
 b15zdnd11an1n04x5 FILLER_174_1454 ();
 b15zdnd11an1n16x5 FILLER_174_1474 ();
 b15zdnd00an1n01x5 FILLER_174_1490 ();
 b15zdnd11an1n16x5 FILLER_174_1503 ();
 b15zdnd11an1n04x5 FILLER_174_1519 ();
 b15zdnd00an1n02x5 FILLER_174_1523 ();
 b15zdnd11an1n32x5 FILLER_174_1530 ();
 b15zdnd11an1n16x5 FILLER_174_1562 ();
 b15zdnd11an1n08x5 FILLER_174_1578 ();
 b15zdnd11an1n04x5 FILLER_174_1586 ();
 b15zdnd00an1n02x5 FILLER_174_1590 ();
 b15zdnd00an1n01x5 FILLER_174_1592 ();
 b15zdnd11an1n16x5 FILLER_174_1597 ();
 b15zdnd11an1n04x5 FILLER_174_1613 ();
 b15zdnd11an1n04x5 FILLER_174_1627 ();
 b15zdnd11an1n04x5 FILLER_174_1640 ();
 b15zdnd00an1n02x5 FILLER_174_1644 ();
 b15zdnd00an1n01x5 FILLER_174_1646 ();
 b15zdnd11an1n04x5 FILLER_174_1652 ();
 b15zdnd11an1n16x5 FILLER_174_1669 ();
 b15zdnd11an1n04x5 FILLER_174_1685 ();
 b15zdnd11an1n64x5 FILLER_174_1713 ();
 b15zdnd11an1n64x5 FILLER_174_1777 ();
 b15zdnd11an1n32x5 FILLER_174_1841 ();
 b15zdnd11an1n08x5 FILLER_174_1873 ();
 b15zdnd00an1n02x5 FILLER_174_1881 ();
 b15zdnd11an1n16x5 FILLER_174_1903 ();
 b15zdnd11an1n08x5 FILLER_174_1919 ();
 b15zdnd00an1n02x5 FILLER_174_1927 ();
 b15zdnd11an1n04x5 FILLER_174_1933 ();
 b15zdnd11an1n64x5 FILLER_174_1957 ();
 b15zdnd11an1n32x5 FILLER_174_2021 ();
 b15zdnd11an1n16x5 FILLER_174_2053 ();
 b15zdnd11an1n04x5 FILLER_174_2069 ();
 b15zdnd00an1n01x5 FILLER_174_2073 ();
 b15zdnd11an1n16x5 FILLER_174_2105 ();
 b15zdnd11an1n08x5 FILLER_174_2121 ();
 b15zdnd11an1n04x5 FILLER_174_2129 ();
 b15zdnd00an1n02x5 FILLER_174_2133 ();
 b15zdnd11an1n04x5 FILLER_174_2149 ();
 b15zdnd00an1n01x5 FILLER_174_2153 ();
 b15zdnd11an1n04x5 FILLER_174_2162 ();
 b15zdnd00an1n02x5 FILLER_174_2166 ();
 b15zdnd00an1n01x5 FILLER_174_2168 ();
 b15zdnd11an1n16x5 FILLER_174_2189 ();
 b15zdnd11an1n04x5 FILLER_174_2205 ();
 b15zdnd11an1n16x5 FILLER_174_2217 ();
 b15zdnd11an1n04x5 FILLER_174_2233 ();
 b15zdnd00an1n02x5 FILLER_174_2237 ();
 b15zdnd00an1n01x5 FILLER_174_2239 ();
 b15zdnd11an1n08x5 FILLER_174_2244 ();
 b15zdnd11an1n04x5 FILLER_174_2252 ();
 b15zdnd00an1n02x5 FILLER_174_2256 ();
 b15zdnd11an1n08x5 FILLER_174_2263 ();
 b15zdnd11an1n04x5 FILLER_174_2271 ();
 b15zdnd00an1n01x5 FILLER_174_2275 ();
 b15zdnd11an1n32x5 FILLER_175_0 ();
 b15zdnd11an1n08x5 FILLER_175_32 ();
 b15zdnd11an1n04x5 FILLER_175_40 ();
 b15zdnd00an1n01x5 FILLER_175_44 ();
 b15zdnd11an1n04x5 FILLER_175_61 ();
 b15zdnd11an1n04x5 FILLER_175_79 ();
 b15zdnd11an1n16x5 FILLER_175_91 ();
 b15zdnd11an1n64x5 FILLER_175_117 ();
 b15zdnd11an1n08x5 FILLER_175_181 ();
 b15zdnd00an1n01x5 FILLER_175_189 ();
 b15zdnd11an1n16x5 FILLER_175_196 ();
 b15zdnd11an1n04x5 FILLER_175_212 ();
 b15zdnd00an1n02x5 FILLER_175_216 ();
 b15zdnd11an1n04x5 FILLER_175_224 ();
 b15zdnd11an1n08x5 FILLER_175_238 ();
 b15zdnd11an1n04x5 FILLER_175_246 ();
 b15zdnd11an1n32x5 FILLER_175_263 ();
 b15zdnd11an1n04x5 FILLER_175_295 ();
 b15zdnd00an1n02x5 FILLER_175_299 ();
 b15zdnd00an1n01x5 FILLER_175_301 ();
 b15zdnd11an1n16x5 FILLER_175_310 ();
 b15zdnd11an1n64x5 FILLER_175_332 ();
 b15zdnd11an1n64x5 FILLER_175_396 ();
 b15zdnd11an1n16x5 FILLER_175_460 ();
 b15zdnd11an1n04x5 FILLER_175_476 ();
 b15zdnd00an1n01x5 FILLER_175_480 ();
 b15zdnd11an1n16x5 FILLER_175_492 ();
 b15zdnd11an1n04x5 FILLER_175_508 ();
 b15zdnd00an1n02x5 FILLER_175_512 ();
 b15zdnd00an1n01x5 FILLER_175_514 ();
 b15zdnd11an1n64x5 FILLER_175_530 ();
 b15zdnd11an1n08x5 FILLER_175_594 ();
 b15zdnd11an1n04x5 FILLER_175_602 ();
 b15zdnd11an1n16x5 FILLER_175_611 ();
 b15zdnd11an1n08x5 FILLER_175_627 ();
 b15zdnd00an1n02x5 FILLER_175_635 ();
 b15zdnd00an1n01x5 FILLER_175_637 ();
 b15zdnd11an1n04x5 FILLER_175_647 ();
 b15zdnd11an1n64x5 FILLER_175_658 ();
 b15zdnd11an1n32x5 FILLER_175_722 ();
 b15zdnd11an1n04x5 FILLER_175_754 ();
 b15zdnd00an1n02x5 FILLER_175_758 ();
 b15zdnd11an1n64x5 FILLER_175_791 ();
 b15zdnd11an1n32x5 FILLER_175_855 ();
 b15zdnd00an1n02x5 FILLER_175_887 ();
 b15zdnd11an1n64x5 FILLER_175_905 ();
 b15zdnd00an1n01x5 FILLER_175_969 ();
 b15zdnd11an1n32x5 FILLER_175_983 ();
 b15zdnd11an1n04x5 FILLER_175_1015 ();
 b15zdnd00an1n02x5 FILLER_175_1019 ();
 b15zdnd11an1n32x5 FILLER_175_1029 ();
 b15zdnd00an1n02x5 FILLER_175_1061 ();
 b15zdnd00an1n01x5 FILLER_175_1063 ();
 b15zdnd11an1n16x5 FILLER_175_1071 ();
 b15zdnd11an1n08x5 FILLER_175_1087 ();
 b15zdnd11an1n04x5 FILLER_175_1095 ();
 b15zdnd00an1n02x5 FILLER_175_1099 ();
 b15zdnd00an1n01x5 FILLER_175_1101 ();
 b15zdnd11an1n64x5 FILLER_175_1107 ();
 b15zdnd11an1n16x5 FILLER_175_1171 ();
 b15zdnd11an1n08x5 FILLER_175_1187 ();
 b15zdnd11an1n08x5 FILLER_175_1202 ();
 b15zdnd00an1n01x5 FILLER_175_1210 ();
 b15zdnd11an1n16x5 FILLER_175_1221 ();
 b15zdnd00an1n02x5 FILLER_175_1237 ();
 b15zdnd11an1n32x5 FILLER_175_1252 ();
 b15zdnd11an1n04x5 FILLER_175_1302 ();
 b15zdnd11an1n08x5 FILLER_175_1315 ();
 b15zdnd11an1n04x5 FILLER_175_1323 ();
 b15zdnd11an1n04x5 FILLER_175_1350 ();
 b15zdnd11an1n08x5 FILLER_175_1361 ();
 b15zdnd00an1n02x5 FILLER_175_1369 ();
 b15zdnd00an1n01x5 FILLER_175_1371 ();
 b15zdnd11an1n32x5 FILLER_175_1379 ();
 b15zdnd11an1n08x5 FILLER_175_1411 ();
 b15zdnd00an1n02x5 FILLER_175_1419 ();
 b15zdnd00an1n01x5 FILLER_175_1421 ();
 b15zdnd11an1n32x5 FILLER_175_1436 ();
 b15zdnd11an1n16x5 FILLER_175_1468 ();
 b15zdnd11an1n08x5 FILLER_175_1484 ();
 b15zdnd11an1n04x5 FILLER_175_1492 ();
 b15zdnd00an1n01x5 FILLER_175_1496 ();
 b15zdnd11an1n16x5 FILLER_175_1501 ();
 b15zdnd11an1n08x5 FILLER_175_1517 ();
 b15zdnd00an1n02x5 FILLER_175_1525 ();
 b15zdnd00an1n01x5 FILLER_175_1527 ();
 b15zdnd11an1n32x5 FILLER_175_1535 ();
 b15zdnd00an1n02x5 FILLER_175_1567 ();
 b15zdnd11an1n64x5 FILLER_175_1575 ();
 b15zdnd11an1n64x5 FILLER_175_1639 ();
 b15zdnd11an1n08x5 FILLER_175_1703 ();
 b15zdnd11an1n04x5 FILLER_175_1711 ();
 b15zdnd00an1n02x5 FILLER_175_1715 ();
 b15zdnd00an1n01x5 FILLER_175_1717 ();
 b15zdnd11an1n04x5 FILLER_175_1733 ();
 b15zdnd00an1n02x5 FILLER_175_1737 ();
 b15zdnd00an1n01x5 FILLER_175_1739 ();
 b15zdnd11an1n16x5 FILLER_175_1750 ();
 b15zdnd11an1n04x5 FILLER_175_1766 ();
 b15zdnd00an1n02x5 FILLER_175_1770 ();
 b15zdnd11an1n32x5 FILLER_175_1792 ();
 b15zdnd11an1n16x5 FILLER_175_1824 ();
 b15zdnd11an1n04x5 FILLER_175_1840 ();
 b15zdnd00an1n01x5 FILLER_175_1844 ();
 b15zdnd11an1n64x5 FILLER_175_1854 ();
 b15zdnd11an1n32x5 FILLER_175_1918 ();
 b15zdnd11an1n16x5 FILLER_175_1950 ();
 b15zdnd11an1n08x5 FILLER_175_1966 ();
 b15zdnd00an1n02x5 FILLER_175_1974 ();
 b15zdnd00an1n01x5 FILLER_175_1976 ();
 b15zdnd11an1n32x5 FILLER_175_1986 ();
 b15zdnd11an1n16x5 FILLER_175_2018 ();
 b15zdnd00an1n02x5 FILLER_175_2034 ();
 b15zdnd11an1n08x5 FILLER_175_2054 ();
 b15zdnd00an1n02x5 FILLER_175_2062 ();
 b15zdnd11an1n04x5 FILLER_175_2074 ();
 b15zdnd11an1n64x5 FILLER_175_2088 ();
 b15zdnd11an1n16x5 FILLER_175_2152 ();
 b15zdnd00an1n01x5 FILLER_175_2168 ();
 b15zdnd11an1n08x5 FILLER_175_2174 ();
 b15zdnd00an1n01x5 FILLER_175_2182 ();
 b15zdnd11an1n32x5 FILLER_175_2187 ();
 b15zdnd11an1n08x5 FILLER_175_2219 ();
 b15zdnd00an1n02x5 FILLER_175_2227 ();
 b15zdnd11an1n04x5 FILLER_175_2233 ();
 b15zdnd11an1n04x5 FILLER_175_2241 ();
 b15zdnd11an1n04x5 FILLER_175_2249 ();
 b15zdnd00an1n01x5 FILLER_175_2253 ();
 b15zdnd11an1n16x5 FILLER_175_2258 ();
 b15zdnd11an1n08x5 FILLER_175_2274 ();
 b15zdnd00an1n02x5 FILLER_175_2282 ();
 b15zdnd00an1n02x5 FILLER_176_8 ();
 b15zdnd00an1n01x5 FILLER_176_10 ();
 b15zdnd11an1n32x5 FILLER_176_19 ();
 b15zdnd11an1n08x5 FILLER_176_51 ();
 b15zdnd11an1n04x5 FILLER_176_59 ();
 b15zdnd00an1n02x5 FILLER_176_63 ();
 b15zdnd11an1n04x5 FILLER_176_72 ();
 b15zdnd00an1n02x5 FILLER_176_76 ();
 b15zdnd11an1n08x5 FILLER_176_84 ();
 b15zdnd00an1n02x5 FILLER_176_92 ();
 b15zdnd11an1n32x5 FILLER_176_104 ();
 b15zdnd11an1n08x5 FILLER_176_136 ();
 b15zdnd11an1n64x5 FILLER_176_153 ();
 b15zdnd11an1n16x5 FILLER_176_217 ();
 b15zdnd11an1n08x5 FILLER_176_233 ();
 b15zdnd11an1n04x5 FILLER_176_241 ();
 b15zdnd00an1n02x5 FILLER_176_245 ();
 b15zdnd11an1n08x5 FILLER_176_253 ();
 b15zdnd00an1n02x5 FILLER_176_261 ();
 b15zdnd00an1n01x5 FILLER_176_263 ();
 b15zdnd11an1n16x5 FILLER_176_278 ();
 b15zdnd11an1n08x5 FILLER_176_294 ();
 b15zdnd11an1n08x5 FILLER_176_314 ();
 b15zdnd11an1n04x5 FILLER_176_322 ();
 b15zdnd11an1n64x5 FILLER_176_338 ();
 b15zdnd11an1n04x5 FILLER_176_402 ();
 b15zdnd11an1n16x5 FILLER_176_411 ();
 b15zdnd11an1n04x5 FILLER_176_427 ();
 b15zdnd00an1n02x5 FILLER_176_431 ();
 b15zdnd11an1n16x5 FILLER_176_442 ();
 b15zdnd11an1n08x5 FILLER_176_458 ();
 b15zdnd11an1n04x5 FILLER_176_466 ();
 b15zdnd11an1n08x5 FILLER_176_475 ();
 b15zdnd11an1n04x5 FILLER_176_483 ();
 b15zdnd00an1n02x5 FILLER_176_487 ();
 b15zdnd00an1n01x5 FILLER_176_489 ();
 b15zdnd11an1n16x5 FILLER_176_494 ();
 b15zdnd11an1n32x5 FILLER_176_525 ();
 b15zdnd11an1n16x5 FILLER_176_557 ();
 b15zdnd11an1n08x5 FILLER_176_573 ();
 b15zdnd11an1n04x5 FILLER_176_581 ();
 b15zdnd11an1n16x5 FILLER_176_600 ();
 b15zdnd11an1n04x5 FILLER_176_616 ();
 b15zdnd00an1n02x5 FILLER_176_620 ();
 b15zdnd11an1n04x5 FILLER_176_633 ();
 b15zdnd11an1n32x5 FILLER_176_649 ();
 b15zdnd11an1n08x5 FILLER_176_681 ();
 b15zdnd11an1n04x5 FILLER_176_689 ();
 b15zdnd00an1n02x5 FILLER_176_693 ();
 b15zdnd00an1n01x5 FILLER_176_695 ();
 b15zdnd11an1n04x5 FILLER_176_714 ();
 b15zdnd11an1n08x5 FILLER_176_726 ();
 b15zdnd11an1n04x5 FILLER_176_734 ();
 b15zdnd00an1n02x5 FILLER_176_738 ();
 b15zdnd00an1n01x5 FILLER_176_740 ();
 b15zdnd11an1n04x5 FILLER_176_747 ();
 b15zdnd11an1n32x5 FILLER_176_783 ();
 b15zdnd11an1n16x5 FILLER_176_815 ();
 b15zdnd11an1n08x5 FILLER_176_831 ();
 b15zdnd11an1n16x5 FILLER_176_848 ();
 b15zdnd00an1n01x5 FILLER_176_864 ();
 b15zdnd11an1n04x5 FILLER_176_869 ();
 b15zdnd00an1n01x5 FILLER_176_873 ();
 b15zdnd11an1n08x5 FILLER_176_880 ();
 b15zdnd11an1n04x5 FILLER_176_888 ();
 b15zdnd00an1n01x5 FILLER_176_892 ();
 b15zdnd11an1n04x5 FILLER_176_900 ();
 b15zdnd11an1n32x5 FILLER_176_909 ();
 b15zdnd11an1n04x5 FILLER_176_941 ();
 b15zdnd00an1n01x5 FILLER_176_945 ();
 b15zdnd11an1n04x5 FILLER_176_962 ();
 b15zdnd11an1n16x5 FILLER_176_997 ();
 b15zdnd00an1n01x5 FILLER_176_1013 ();
 b15zdnd11an1n64x5 FILLER_176_1023 ();
 b15zdnd11an1n16x5 FILLER_176_1087 ();
 b15zdnd00an1n01x5 FILLER_176_1103 ();
 b15zdnd11an1n04x5 FILLER_176_1109 ();
 b15zdnd11an1n16x5 FILLER_176_1125 ();
 b15zdnd11an1n32x5 FILLER_176_1150 ();
 b15zdnd11an1n04x5 FILLER_176_1182 ();
 b15zdnd00an1n01x5 FILLER_176_1186 ();
 b15zdnd11an1n64x5 FILLER_176_1219 ();
 b15zdnd11an1n64x5 FILLER_176_1283 ();
 b15zdnd11an1n16x5 FILLER_176_1353 ();
 b15zdnd00an1n02x5 FILLER_176_1369 ();
 b15zdnd11an1n04x5 FILLER_176_1377 ();
 b15zdnd11an1n64x5 FILLER_176_1405 ();
 b15zdnd11an1n32x5 FILLER_176_1469 ();
 b15zdnd11an1n16x5 FILLER_176_1501 ();
 b15zdnd11an1n08x5 FILLER_176_1517 ();
 b15zdnd00an1n02x5 FILLER_176_1525 ();
 b15zdnd11an1n08x5 FILLER_176_1539 ();
 b15zdnd11an1n04x5 FILLER_176_1547 ();
 b15zdnd00an1n02x5 FILLER_176_1551 ();
 b15zdnd00an1n01x5 FILLER_176_1553 ();
 b15zdnd11an1n16x5 FILLER_176_1580 ();
 b15zdnd11an1n04x5 FILLER_176_1596 ();
 b15zdnd00an1n02x5 FILLER_176_1600 ();
 b15zdnd11an1n16x5 FILLER_176_1606 ();
 b15zdnd00an1n01x5 FILLER_176_1622 ();
 b15zdnd11an1n64x5 FILLER_176_1637 ();
 b15zdnd00an1n02x5 FILLER_176_1701 ();
 b15zdnd00an1n01x5 FILLER_176_1703 ();
 b15zdnd11an1n64x5 FILLER_176_1715 ();
 b15zdnd11an1n32x5 FILLER_176_1779 ();
 b15zdnd11an1n16x5 FILLER_176_1811 ();
 b15zdnd11an1n08x5 FILLER_176_1827 ();
 b15zdnd11an1n64x5 FILLER_176_1846 ();
 b15zdnd11an1n32x5 FILLER_176_1910 ();
 b15zdnd11an1n08x5 FILLER_176_1942 ();
 b15zdnd11an1n04x5 FILLER_176_1950 ();
 b15zdnd00an1n02x5 FILLER_176_1954 ();
 b15zdnd00an1n01x5 FILLER_176_1956 ();
 b15zdnd11an1n16x5 FILLER_176_1968 ();
 b15zdnd11an1n08x5 FILLER_176_1984 ();
 b15zdnd00an1n01x5 FILLER_176_1992 ();
 b15zdnd11an1n16x5 FILLER_176_1998 ();
 b15zdnd11an1n04x5 FILLER_176_2014 ();
 b15zdnd00an1n02x5 FILLER_176_2018 ();
 b15zdnd11an1n64x5 FILLER_176_2044 ();
 b15zdnd11an1n32x5 FILLER_176_2108 ();
 b15zdnd11an1n08x5 FILLER_176_2140 ();
 b15zdnd11an1n04x5 FILLER_176_2148 ();
 b15zdnd00an1n02x5 FILLER_176_2152 ();
 b15zdnd11an1n32x5 FILLER_176_2162 ();
 b15zdnd11an1n08x5 FILLER_176_2194 ();
 b15zdnd11an1n32x5 FILLER_176_2207 ();
 b15zdnd11an1n04x5 FILLER_176_2239 ();
 b15zdnd00an1n02x5 FILLER_176_2243 ();
 b15zdnd00an1n01x5 FILLER_176_2245 ();
 b15zdnd11an1n08x5 FILLER_176_2250 ();
 b15zdnd11an1n04x5 FILLER_176_2258 ();
 b15zdnd11an1n08x5 FILLER_176_2266 ();
 b15zdnd00an1n02x5 FILLER_176_2274 ();
 b15zdnd11an1n16x5 FILLER_177_0 ();
 b15zdnd11an1n64x5 FILLER_177_23 ();
 b15zdnd00an1n02x5 FILLER_177_87 ();
 b15zdnd11an1n64x5 FILLER_177_95 ();
 b15zdnd11an1n04x5 FILLER_177_159 ();
 b15zdnd00an1n01x5 FILLER_177_163 ();
 b15zdnd11an1n04x5 FILLER_177_172 ();
 b15zdnd00an1n02x5 FILLER_177_176 ();
 b15zdnd11an1n32x5 FILLER_177_190 ();
 b15zdnd11an1n16x5 FILLER_177_222 ();
 b15zdnd11an1n04x5 FILLER_177_238 ();
 b15zdnd00an1n02x5 FILLER_177_242 ();
 b15zdnd11an1n32x5 FILLER_177_253 ();
 b15zdnd11an1n16x5 FILLER_177_285 ();
 b15zdnd00an1n02x5 FILLER_177_301 ();
 b15zdnd11an1n16x5 FILLER_177_307 ();
 b15zdnd00an1n02x5 FILLER_177_323 ();
 b15zdnd00an1n01x5 FILLER_177_325 ();
 b15zdnd11an1n04x5 FILLER_177_332 ();
 b15zdnd11an1n64x5 FILLER_177_340 ();
 b15zdnd11an1n08x5 FILLER_177_404 ();
 b15zdnd00an1n01x5 FILLER_177_412 ();
 b15zdnd11an1n16x5 FILLER_177_433 ();
 b15zdnd11an1n08x5 FILLER_177_449 ();
 b15zdnd11an1n04x5 FILLER_177_463 ();
 b15zdnd00an1n02x5 FILLER_177_467 ();
 b15zdnd11an1n32x5 FILLER_177_475 ();
 b15zdnd11an1n08x5 FILLER_177_507 ();
 b15zdnd11an1n04x5 FILLER_177_515 ();
 b15zdnd11an1n16x5 FILLER_177_524 ();
 b15zdnd11an1n04x5 FILLER_177_540 ();
 b15zdnd00an1n01x5 FILLER_177_544 ();
 b15zdnd11an1n08x5 FILLER_177_552 ();
 b15zdnd00an1n01x5 FILLER_177_560 ();
 b15zdnd11an1n64x5 FILLER_177_567 ();
 b15zdnd11an1n16x5 FILLER_177_631 ();
 b15zdnd11an1n04x5 FILLER_177_647 ();
 b15zdnd00an1n02x5 FILLER_177_651 ();
 b15zdnd11an1n04x5 FILLER_177_663 ();
 b15zdnd11an1n16x5 FILLER_177_673 ();
 b15zdnd00an1n01x5 FILLER_177_689 ();
 b15zdnd11an1n04x5 FILLER_177_694 ();
 b15zdnd00an1n01x5 FILLER_177_698 ();
 b15zdnd11an1n64x5 FILLER_177_705 ();
 b15zdnd11an1n32x5 FILLER_177_769 ();
 b15zdnd11an1n16x5 FILLER_177_801 ();
 b15zdnd11an1n08x5 FILLER_177_817 ();
 b15zdnd11an1n04x5 FILLER_177_825 ();
 b15zdnd00an1n02x5 FILLER_177_829 ();
 b15zdnd00an1n01x5 FILLER_177_831 ();
 b15zdnd11an1n16x5 FILLER_177_845 ();
 b15zdnd00an1n01x5 FILLER_177_861 ();
 b15zdnd11an1n04x5 FILLER_177_869 ();
 b15zdnd11an1n16x5 FILLER_177_882 ();
 b15zdnd11an1n08x5 FILLER_177_898 ();
 b15zdnd11an1n32x5 FILLER_177_915 ();
 b15zdnd11an1n08x5 FILLER_177_947 ();
 b15zdnd00an1n01x5 FILLER_177_955 ();
 b15zdnd11an1n64x5 FILLER_177_962 ();
 b15zdnd11an1n08x5 FILLER_177_1026 ();
 b15zdnd00an1n02x5 FILLER_177_1034 ();
 b15zdnd00an1n01x5 FILLER_177_1036 ();
 b15zdnd11an1n08x5 FILLER_177_1042 ();
 b15zdnd11an1n04x5 FILLER_177_1050 ();
 b15zdnd11an1n08x5 FILLER_177_1059 ();
 b15zdnd11an1n04x5 FILLER_177_1067 ();
 b15zdnd00an1n01x5 FILLER_177_1071 ();
 b15zdnd11an1n32x5 FILLER_177_1077 ();
 b15zdnd11an1n08x5 FILLER_177_1109 ();
 b15zdnd00an1n02x5 FILLER_177_1117 ();
 b15zdnd00an1n01x5 FILLER_177_1119 ();
 b15zdnd11an1n16x5 FILLER_177_1128 ();
 b15zdnd11an1n04x5 FILLER_177_1144 ();
 b15zdnd00an1n02x5 FILLER_177_1148 ();
 b15zdnd00an1n01x5 FILLER_177_1150 ();
 b15zdnd11an1n04x5 FILLER_177_1167 ();
 b15zdnd11an1n64x5 FILLER_177_1176 ();
 b15zdnd11an1n64x5 FILLER_177_1240 ();
 b15zdnd11an1n64x5 FILLER_177_1304 ();
 b15zdnd11an1n64x5 FILLER_177_1368 ();
 b15zdnd11an1n16x5 FILLER_177_1432 ();
 b15zdnd11an1n04x5 FILLER_177_1448 ();
 b15zdnd00an1n02x5 FILLER_177_1452 ();
 b15zdnd00an1n01x5 FILLER_177_1454 ();
 b15zdnd11an1n16x5 FILLER_177_1467 ();
 b15zdnd11an1n08x5 FILLER_177_1483 ();
 b15zdnd11an1n04x5 FILLER_177_1491 ();
 b15zdnd11an1n16x5 FILLER_177_1503 ();
 b15zdnd11an1n04x5 FILLER_177_1519 ();
 b15zdnd00an1n01x5 FILLER_177_1523 ();
 b15zdnd11an1n32x5 FILLER_177_1529 ();
 b15zdnd11an1n04x5 FILLER_177_1566 ();
 b15zdnd11an1n04x5 FILLER_177_1576 ();
 b15zdnd00an1n02x5 FILLER_177_1580 ();
 b15zdnd11an1n04x5 FILLER_177_1594 ();
 b15zdnd11an1n08x5 FILLER_177_1605 ();
 b15zdnd00an1n02x5 FILLER_177_1613 ();
 b15zdnd11an1n16x5 FILLER_177_1621 ();
 b15zdnd11an1n08x5 FILLER_177_1637 ();
 b15zdnd00an1n02x5 FILLER_177_1645 ();
 b15zdnd11an1n04x5 FILLER_177_1656 ();
 b15zdnd11an1n64x5 FILLER_177_1667 ();
 b15zdnd11an1n16x5 FILLER_177_1731 ();
 b15zdnd11an1n04x5 FILLER_177_1747 ();
 b15zdnd00an1n01x5 FILLER_177_1751 ();
 b15zdnd11an1n08x5 FILLER_177_1762 ();
 b15zdnd11an1n04x5 FILLER_177_1770 ();
 b15zdnd11an1n08x5 FILLER_177_1779 ();
 b15zdnd11an1n04x5 FILLER_177_1787 ();
 b15zdnd11an1n04x5 FILLER_177_1806 ();
 b15zdnd11an1n08x5 FILLER_177_1830 ();
 b15zdnd11an1n64x5 FILLER_177_1843 ();
 b15zdnd11an1n64x5 FILLER_177_1907 ();
 b15zdnd11an1n16x5 FILLER_177_1971 ();
 b15zdnd11an1n04x5 FILLER_177_1987 ();
 b15zdnd11an1n32x5 FILLER_177_2011 ();
 b15zdnd11an1n16x5 FILLER_177_2043 ();
 b15zdnd11an1n08x5 FILLER_177_2059 ();
 b15zdnd00an1n02x5 FILLER_177_2067 ();
 b15zdnd11an1n16x5 FILLER_177_2094 ();
 b15zdnd11an1n04x5 FILLER_177_2110 ();
 b15zdnd11an1n64x5 FILLER_177_2120 ();
 b15zdnd11an1n16x5 FILLER_177_2184 ();
 b15zdnd11an1n16x5 FILLER_177_2220 ();
 b15zdnd11an1n04x5 FILLER_177_2236 ();
 b15zdnd00an1n02x5 FILLER_177_2240 ();
 b15zdnd00an1n01x5 FILLER_177_2242 ();
 b15zdnd11an1n04x5 FILLER_177_2251 ();
 b15zdnd11an1n04x5 FILLER_177_2259 ();
 b15zdnd00an1n02x5 FILLER_177_2263 ();
 b15zdnd00an1n01x5 FILLER_177_2265 ();
 b15zdnd11an1n08x5 FILLER_177_2270 ();
 b15zdnd00an1n02x5 FILLER_177_2282 ();
 b15zdnd11an1n32x5 FILLER_178_8 ();
 b15zdnd00an1n02x5 FILLER_178_40 ();
 b15zdnd00an1n01x5 FILLER_178_42 ();
 b15zdnd11an1n08x5 FILLER_178_47 ();
 b15zdnd00an1n02x5 FILLER_178_55 ();
 b15zdnd11an1n32x5 FILLER_178_64 ();
 b15zdnd11an1n16x5 FILLER_178_96 ();
 b15zdnd11an1n04x5 FILLER_178_112 ();
 b15zdnd00an1n01x5 FILLER_178_116 ();
 b15zdnd11an1n32x5 FILLER_178_125 ();
 b15zdnd11an1n08x5 FILLER_178_157 ();
 b15zdnd11an1n04x5 FILLER_178_165 ();
 b15zdnd00an1n02x5 FILLER_178_169 ();
 b15zdnd11an1n16x5 FILLER_178_181 ();
 b15zdnd11an1n04x5 FILLER_178_197 ();
 b15zdnd11an1n04x5 FILLER_178_211 ();
 b15zdnd11an1n32x5 FILLER_178_235 ();
 b15zdnd11an1n16x5 FILLER_178_267 ();
 b15zdnd11an1n08x5 FILLER_178_283 ();
 b15zdnd00an1n02x5 FILLER_178_291 ();
 b15zdnd00an1n01x5 FILLER_178_293 ();
 b15zdnd11an1n64x5 FILLER_178_310 ();
 b15zdnd11an1n16x5 FILLER_178_374 ();
 b15zdnd11an1n08x5 FILLER_178_390 ();
 b15zdnd00an1n01x5 FILLER_178_398 ();
 b15zdnd11an1n16x5 FILLER_178_407 ();
 b15zdnd11an1n08x5 FILLER_178_423 ();
 b15zdnd00an1n02x5 FILLER_178_431 ();
 b15zdnd00an1n01x5 FILLER_178_433 ();
 b15zdnd11an1n32x5 FILLER_178_440 ();
 b15zdnd11an1n16x5 FILLER_178_472 ();
 b15zdnd11an1n04x5 FILLER_178_488 ();
 b15zdnd00an1n01x5 FILLER_178_492 ();
 b15zdnd11an1n32x5 FILLER_178_499 ();
 b15zdnd11an1n16x5 FILLER_178_531 ();
 b15zdnd00an1n01x5 FILLER_178_547 ();
 b15zdnd11an1n32x5 FILLER_178_554 ();
 b15zdnd11an1n16x5 FILLER_178_591 ();
 b15zdnd11an1n04x5 FILLER_178_607 ();
 b15zdnd00an1n01x5 FILLER_178_611 ();
 b15zdnd11an1n16x5 FILLER_178_627 ();
 b15zdnd00an1n01x5 FILLER_178_643 ();
 b15zdnd11an1n04x5 FILLER_178_659 ();
 b15zdnd00an1n01x5 FILLER_178_663 ();
 b15zdnd11an1n04x5 FILLER_178_688 ();
 b15zdnd11an1n16x5 FILLER_178_700 ();
 b15zdnd00an1n02x5 FILLER_178_716 ();
 b15zdnd11an1n64x5 FILLER_178_726 ();
 b15zdnd11an1n32x5 FILLER_178_790 ();
 b15zdnd11an1n08x5 FILLER_178_822 ();
 b15zdnd11an1n04x5 FILLER_178_830 ();
 b15zdnd00an1n02x5 FILLER_178_834 ();
 b15zdnd00an1n01x5 FILLER_178_836 ();
 b15zdnd11an1n16x5 FILLER_178_843 ();
 b15zdnd00an1n02x5 FILLER_178_859 ();
 b15zdnd00an1n01x5 FILLER_178_861 ();
 b15zdnd11an1n08x5 FILLER_178_867 ();
 b15zdnd11an1n04x5 FILLER_178_875 ();
 b15zdnd00an1n01x5 FILLER_178_879 ();
 b15zdnd11an1n16x5 FILLER_178_893 ();
 b15zdnd11an1n32x5 FILLER_178_916 ();
 b15zdnd00an1n01x5 FILLER_178_948 ();
 b15zdnd11an1n32x5 FILLER_178_959 ();
 b15zdnd11an1n16x5 FILLER_178_991 ();
 b15zdnd11an1n08x5 FILLER_178_1007 ();
 b15zdnd11an1n04x5 FILLER_178_1015 ();
 b15zdnd11an1n04x5 FILLER_178_1026 ();
 b15zdnd11an1n08x5 FILLER_178_1042 ();
 b15zdnd11an1n04x5 FILLER_178_1050 ();
 b15zdnd11an1n32x5 FILLER_178_1066 ();
 b15zdnd11an1n16x5 FILLER_178_1098 ();
 b15zdnd00an1n02x5 FILLER_178_1114 ();
 b15zdnd00an1n01x5 FILLER_178_1116 ();
 b15zdnd11an1n16x5 FILLER_178_1129 ();
 b15zdnd11an1n08x5 FILLER_178_1145 ();
 b15zdnd00an1n02x5 FILLER_178_1153 ();
 b15zdnd11an1n08x5 FILLER_178_1159 ();
 b15zdnd11an1n64x5 FILLER_178_1176 ();
 b15zdnd11an1n32x5 FILLER_178_1240 ();
 b15zdnd11an1n16x5 FILLER_178_1272 ();
 b15zdnd11an1n08x5 FILLER_178_1288 ();
 b15zdnd11an1n04x5 FILLER_178_1296 ();
 b15zdnd00an1n01x5 FILLER_178_1300 ();
 b15zdnd11an1n04x5 FILLER_178_1308 ();
 b15zdnd00an1n01x5 FILLER_178_1312 ();
 b15zdnd11an1n16x5 FILLER_178_1317 ();
 b15zdnd11an1n04x5 FILLER_178_1337 ();
 b15zdnd11an1n04x5 FILLER_178_1346 ();
 b15zdnd11an1n64x5 FILLER_178_1358 ();
 b15zdnd11an1n32x5 FILLER_178_1422 ();
 b15zdnd11an1n04x5 FILLER_178_1454 ();
 b15zdnd11an1n32x5 FILLER_178_1464 ();
 b15zdnd11an1n32x5 FILLER_178_1511 ();
 b15zdnd11an1n04x5 FILLER_178_1543 ();
 b15zdnd00an1n01x5 FILLER_178_1547 ();
 b15zdnd11an1n32x5 FILLER_178_1553 ();
 b15zdnd11an1n16x5 FILLER_178_1585 ();
 b15zdnd11an1n08x5 FILLER_178_1601 ();
 b15zdnd11an1n04x5 FILLER_178_1609 ();
 b15zdnd00an1n02x5 FILLER_178_1613 ();
 b15zdnd11an1n64x5 FILLER_178_1631 ();
 b15zdnd11an1n08x5 FILLER_178_1695 ();
 b15zdnd11an1n04x5 FILLER_178_1703 ();
 b15zdnd00an1n01x5 FILLER_178_1707 ();
 b15zdnd11an1n08x5 FILLER_178_1713 ();
 b15zdnd00an1n01x5 FILLER_178_1721 ();
 b15zdnd11an1n32x5 FILLER_178_1726 ();
 b15zdnd11an1n04x5 FILLER_178_1758 ();
 b15zdnd00an1n02x5 FILLER_178_1762 ();
 b15zdnd11an1n32x5 FILLER_178_1790 ();
 b15zdnd11an1n16x5 FILLER_178_1822 ();
 b15zdnd11an1n04x5 FILLER_178_1838 ();
 b15zdnd11an1n16x5 FILLER_178_1863 ();
 b15zdnd00an1n02x5 FILLER_178_1879 ();
 b15zdnd11an1n16x5 FILLER_178_1885 ();
 b15zdnd11an1n08x5 FILLER_178_1901 ();
 b15zdnd11an1n04x5 FILLER_178_1909 ();
 b15zdnd00an1n02x5 FILLER_178_1913 ();
 b15zdnd11an1n32x5 FILLER_178_1919 ();
 b15zdnd11an1n16x5 FILLER_178_1951 ();
 b15zdnd00an1n02x5 FILLER_178_1967 ();
 b15zdnd00an1n01x5 FILLER_178_1969 ();
 b15zdnd11an1n04x5 FILLER_178_1981 ();
 b15zdnd11an1n32x5 FILLER_178_1997 ();
 b15zdnd11an1n16x5 FILLER_178_2029 ();
 b15zdnd11an1n08x5 FILLER_178_2045 ();
 b15zdnd11an1n08x5 FILLER_178_2079 ();
 b15zdnd00an1n02x5 FILLER_178_2087 ();
 b15zdnd00an1n01x5 FILLER_178_2089 ();
 b15zdnd11an1n04x5 FILLER_178_2110 ();
 b15zdnd11an1n32x5 FILLER_178_2119 ();
 b15zdnd00an1n02x5 FILLER_178_2151 ();
 b15zdnd00an1n01x5 FILLER_178_2153 ();
 b15zdnd11an1n64x5 FILLER_178_2162 ();
 b15zdnd11an1n08x5 FILLER_178_2226 ();
 b15zdnd11an1n04x5 FILLER_178_2234 ();
 b15zdnd11an1n04x5 FILLER_178_2242 ();
 b15zdnd11an1n04x5 FILLER_178_2254 ();
 b15zdnd00an1n02x5 FILLER_178_2258 ();
 b15zdnd00an1n01x5 FILLER_178_2260 ();
 b15zdnd11an1n08x5 FILLER_178_2265 ();
 b15zdnd00an1n02x5 FILLER_178_2273 ();
 b15zdnd00an1n01x5 FILLER_178_2275 ();
 b15zdnd11an1n08x5 FILLER_179_0 ();
 b15zdnd11an1n04x5 FILLER_179_8 ();
 b15zdnd00an1n02x5 FILLER_179_12 ();
 b15zdnd11an1n64x5 FILLER_179_18 ();
 b15zdnd11an1n64x5 FILLER_179_82 ();
 b15zdnd11an1n16x5 FILLER_179_151 ();
 b15zdnd00an1n01x5 FILLER_179_167 ();
 b15zdnd11an1n16x5 FILLER_179_180 ();
 b15zdnd11an1n08x5 FILLER_179_196 ();
 b15zdnd11an1n04x5 FILLER_179_210 ();
 b15zdnd11an1n16x5 FILLER_179_228 ();
 b15zdnd11an1n08x5 FILLER_179_244 ();
 b15zdnd00an1n02x5 FILLER_179_252 ();
 b15zdnd00an1n01x5 FILLER_179_254 ();
 b15zdnd11an1n04x5 FILLER_179_265 ();
 b15zdnd00an1n02x5 FILLER_179_269 ();
 b15zdnd00an1n01x5 FILLER_179_271 ();
 b15zdnd11an1n16x5 FILLER_179_278 ();
 b15zdnd11an1n08x5 FILLER_179_294 ();
 b15zdnd11an1n04x5 FILLER_179_302 ();
 b15zdnd00an1n01x5 FILLER_179_306 ();
 b15zdnd11an1n64x5 FILLER_179_313 ();
 b15zdnd11an1n16x5 FILLER_179_377 ();
 b15zdnd11an1n04x5 FILLER_179_393 ();
 b15zdnd00an1n01x5 FILLER_179_397 ();
 b15zdnd11an1n16x5 FILLER_179_405 ();
 b15zdnd11an1n08x5 FILLER_179_421 ();
 b15zdnd11an1n64x5 FILLER_179_439 ();
 b15zdnd11an1n08x5 FILLER_179_503 ();
 b15zdnd00an1n02x5 FILLER_179_511 ();
 b15zdnd11an1n16x5 FILLER_179_518 ();
 b15zdnd11an1n04x5 FILLER_179_534 ();
 b15zdnd00an1n02x5 FILLER_179_538 ();
 b15zdnd11an1n64x5 FILLER_179_544 ();
 b15zdnd11an1n04x5 FILLER_179_608 ();
 b15zdnd00an1n01x5 FILLER_179_612 ();
 b15zdnd11an1n08x5 FILLER_179_619 ();
 b15zdnd11an1n04x5 FILLER_179_627 ();
 b15zdnd11an1n04x5 FILLER_179_641 ();
 b15zdnd11an1n16x5 FILLER_179_661 ();
 b15zdnd11an1n08x5 FILLER_179_677 ();
 b15zdnd11an1n04x5 FILLER_179_685 ();
 b15zdnd11an1n16x5 FILLER_179_707 ();
 b15zdnd11an1n04x5 FILLER_179_723 ();
 b15zdnd00an1n01x5 FILLER_179_727 ();
 b15zdnd11an1n16x5 FILLER_179_744 ();
 b15zdnd11an1n64x5 FILLER_179_766 ();
 b15zdnd11an1n32x5 FILLER_179_830 ();
 b15zdnd11an1n16x5 FILLER_179_862 ();
 b15zdnd11an1n08x5 FILLER_179_878 ();
 b15zdnd11an1n04x5 FILLER_179_886 ();
 b15zdnd00an1n02x5 FILLER_179_890 ();
 b15zdnd00an1n01x5 FILLER_179_892 ();
 b15zdnd11an1n32x5 FILLER_179_909 ();
 b15zdnd11an1n04x5 FILLER_179_941 ();
 b15zdnd00an1n02x5 FILLER_179_945 ();
 b15zdnd00an1n01x5 FILLER_179_947 ();
 b15zdnd11an1n08x5 FILLER_179_964 ();
 b15zdnd11an1n32x5 FILLER_179_992 ();
 b15zdnd11an1n08x5 FILLER_179_1024 ();
 b15zdnd11an1n04x5 FILLER_179_1032 ();
 b15zdnd00an1n01x5 FILLER_179_1036 ();
 b15zdnd11an1n08x5 FILLER_179_1042 ();
 b15zdnd11an1n16x5 FILLER_179_1054 ();
 b15zdnd11an1n04x5 FILLER_179_1070 ();
 b15zdnd00an1n02x5 FILLER_179_1074 ();
 b15zdnd11an1n16x5 FILLER_179_1082 ();
 b15zdnd11an1n08x5 FILLER_179_1098 ();
 b15zdnd11an1n04x5 FILLER_179_1106 ();
 b15zdnd00an1n02x5 FILLER_179_1110 ();
 b15zdnd11an1n04x5 FILLER_179_1133 ();
 b15zdnd00an1n02x5 FILLER_179_1137 ();
 b15zdnd11an1n04x5 FILLER_179_1145 ();
 b15zdnd11an1n04x5 FILLER_179_1156 ();
 b15zdnd00an1n02x5 FILLER_179_1160 ();
 b15zdnd11an1n64x5 FILLER_179_1166 ();
 b15zdnd11an1n64x5 FILLER_179_1230 ();
 b15zdnd11an1n04x5 FILLER_179_1294 ();
 b15zdnd11an1n08x5 FILLER_179_1305 ();
 b15zdnd00an1n02x5 FILLER_179_1313 ();
 b15zdnd11an1n16x5 FILLER_179_1331 ();
 b15zdnd00an1n01x5 FILLER_179_1347 ();
 b15zdnd11an1n32x5 FILLER_179_1356 ();
 b15zdnd00an1n02x5 FILLER_179_1388 ();
 b15zdnd11an1n04x5 FILLER_179_1397 ();
 b15zdnd11an1n32x5 FILLER_179_1406 ();
 b15zdnd11an1n04x5 FILLER_179_1438 ();
 b15zdnd00an1n02x5 FILLER_179_1442 ();
 b15zdnd11an1n08x5 FILLER_179_1450 ();
 b15zdnd11an1n16x5 FILLER_179_1472 ();
 b15zdnd11an1n08x5 FILLER_179_1488 ();
 b15zdnd00an1n01x5 FILLER_179_1496 ();
 b15zdnd11an1n64x5 FILLER_179_1503 ();
 b15zdnd00an1n01x5 FILLER_179_1567 ();
 b15zdnd11an1n04x5 FILLER_179_1574 ();
 b15zdnd11an1n32x5 FILLER_179_1588 ();
 b15zdnd11an1n16x5 FILLER_179_1620 ();
 b15zdnd11an1n08x5 FILLER_179_1636 ();
 b15zdnd11an1n32x5 FILLER_179_1650 ();
 b15zdnd11an1n16x5 FILLER_179_1682 ();
 b15zdnd11an1n08x5 FILLER_179_1698 ();
 b15zdnd00an1n02x5 FILLER_179_1706 ();
 b15zdnd00an1n01x5 FILLER_179_1708 ();
 b15zdnd11an1n64x5 FILLER_179_1718 ();
 b15zdnd11an1n64x5 FILLER_179_1782 ();
 b15zdnd11an1n08x5 FILLER_179_1846 ();
 b15zdnd00an1n02x5 FILLER_179_1854 ();
 b15zdnd00an1n01x5 FILLER_179_1856 ();
 b15zdnd11an1n16x5 FILLER_179_1862 ();
 b15zdnd00an1n02x5 FILLER_179_1878 ();
 b15zdnd00an1n01x5 FILLER_179_1880 ();
 b15zdnd11an1n08x5 FILLER_179_1901 ();
 b15zdnd00an1n02x5 FILLER_179_1909 ();
 b15zdnd00an1n01x5 FILLER_179_1911 ();
 b15zdnd11an1n04x5 FILLER_179_1917 ();
 b15zdnd11an1n64x5 FILLER_179_1932 ();
 b15zdnd11an1n64x5 FILLER_179_1996 ();
 b15zdnd11an1n64x5 FILLER_179_2060 ();
 b15zdnd00an1n02x5 FILLER_179_2124 ();
 b15zdnd00an1n01x5 FILLER_179_2126 ();
 b15zdnd11an1n04x5 FILLER_179_2147 ();
 b15zdnd11an1n32x5 FILLER_179_2156 ();
 b15zdnd11an1n08x5 FILLER_179_2206 ();
 b15zdnd11an1n04x5 FILLER_179_2214 ();
 b15zdnd00an1n02x5 FILLER_179_2218 ();
 b15zdnd11an1n04x5 FILLER_179_2240 ();
 b15zdnd11an1n08x5 FILLER_179_2248 ();
 b15zdnd11an1n08x5 FILLER_179_2264 ();
 b15zdnd11an1n08x5 FILLER_179_2276 ();
 b15zdnd11an1n32x5 FILLER_180_8 ();
 b15zdnd11an1n08x5 FILLER_180_40 ();
 b15zdnd00an1n01x5 FILLER_180_48 ();
 b15zdnd11an1n08x5 FILLER_180_58 ();
 b15zdnd11an1n16x5 FILLER_180_75 ();
 b15zdnd00an1n02x5 FILLER_180_91 ();
 b15zdnd11an1n64x5 FILLER_180_102 ();
 b15zdnd11an1n16x5 FILLER_180_166 ();
 b15zdnd11an1n08x5 FILLER_180_182 ();
 b15zdnd11an1n04x5 FILLER_180_190 ();
 b15zdnd00an1n01x5 FILLER_180_194 ();
 b15zdnd11an1n32x5 FILLER_180_200 ();
 b15zdnd11an1n08x5 FILLER_180_232 ();
 b15zdnd11an1n04x5 FILLER_180_240 ();
 b15zdnd00an1n02x5 FILLER_180_244 ();
 b15zdnd00an1n01x5 FILLER_180_246 ();
 b15zdnd11an1n16x5 FILLER_180_252 ();
 b15zdnd11an1n04x5 FILLER_180_268 ();
 b15zdnd00an1n01x5 FILLER_180_272 ();
 b15zdnd11an1n04x5 FILLER_180_283 ();
 b15zdnd11an1n16x5 FILLER_180_292 ();
 b15zdnd11an1n04x5 FILLER_180_308 ();
 b15zdnd00an1n01x5 FILLER_180_312 ();
 b15zdnd11an1n64x5 FILLER_180_321 ();
 b15zdnd11an1n64x5 FILLER_180_385 ();
 b15zdnd00an1n01x5 FILLER_180_449 ();
 b15zdnd11an1n32x5 FILLER_180_454 ();
 b15zdnd11an1n08x5 FILLER_180_486 ();
 b15zdnd11an1n04x5 FILLER_180_494 ();
 b15zdnd00an1n02x5 FILLER_180_498 ();
 b15zdnd00an1n01x5 FILLER_180_500 ();
 b15zdnd11an1n32x5 FILLER_180_514 ();
 b15zdnd11an1n04x5 FILLER_180_546 ();
 b15zdnd00an1n01x5 FILLER_180_550 ();
 b15zdnd11an1n32x5 FILLER_180_559 ();
 b15zdnd00an1n01x5 FILLER_180_591 ();
 b15zdnd11an1n16x5 FILLER_180_604 ();
 b15zdnd11an1n08x5 FILLER_180_620 ();
 b15zdnd00an1n02x5 FILLER_180_628 ();
 b15zdnd11an1n08x5 FILLER_180_636 ();
 b15zdnd11an1n32x5 FILLER_180_658 ();
 b15zdnd11an1n16x5 FILLER_180_690 ();
 b15zdnd11an1n08x5 FILLER_180_706 ();
 b15zdnd11an1n04x5 FILLER_180_714 ();
 b15zdnd11an1n32x5 FILLER_180_726 ();
 b15zdnd11an1n04x5 FILLER_180_758 ();
 b15zdnd00an1n02x5 FILLER_180_762 ();
 b15zdnd00an1n01x5 FILLER_180_764 ();
 b15zdnd11an1n64x5 FILLER_180_770 ();
 b15zdnd11an1n64x5 FILLER_180_834 ();
 b15zdnd11an1n64x5 FILLER_180_898 ();
 b15zdnd11an1n16x5 FILLER_180_962 ();
 b15zdnd11an1n04x5 FILLER_180_978 ();
 b15zdnd00an1n01x5 FILLER_180_982 ();
 b15zdnd11an1n04x5 FILLER_180_988 ();
 b15zdnd11an1n32x5 FILLER_180_1001 ();
 b15zdnd11an1n08x5 FILLER_180_1033 ();
 b15zdnd11an1n04x5 FILLER_180_1041 ();
 b15zdnd00an1n02x5 FILLER_180_1045 ();
 b15zdnd00an1n01x5 FILLER_180_1047 ();
 b15zdnd11an1n32x5 FILLER_180_1053 ();
 b15zdnd11an1n16x5 FILLER_180_1085 ();
 b15zdnd11an1n08x5 FILLER_180_1101 ();
 b15zdnd00an1n02x5 FILLER_180_1109 ();
 b15zdnd00an1n01x5 FILLER_180_1111 ();
 b15zdnd11an1n32x5 FILLER_180_1118 ();
 b15zdnd11an1n04x5 FILLER_180_1150 ();
 b15zdnd00an1n02x5 FILLER_180_1154 ();
 b15zdnd00an1n01x5 FILLER_180_1156 ();
 b15zdnd11an1n04x5 FILLER_180_1177 ();
 b15zdnd11an1n64x5 FILLER_180_1186 ();
 b15zdnd11an1n16x5 FILLER_180_1250 ();
 b15zdnd11an1n08x5 FILLER_180_1266 ();
 b15zdnd11an1n04x5 FILLER_180_1274 ();
 b15zdnd00an1n02x5 FILLER_180_1278 ();
 b15zdnd00an1n01x5 FILLER_180_1280 ();
 b15zdnd11an1n32x5 FILLER_180_1295 ();
 b15zdnd11an1n16x5 FILLER_180_1327 ();
 b15zdnd11an1n04x5 FILLER_180_1343 ();
 b15zdnd00an1n01x5 FILLER_180_1347 ();
 b15zdnd11an1n32x5 FILLER_180_1354 ();
 b15zdnd11an1n04x5 FILLER_180_1386 ();
 b15zdnd00an1n01x5 FILLER_180_1390 ();
 b15zdnd11an1n04x5 FILLER_180_1398 ();
 b15zdnd11an1n08x5 FILLER_180_1407 ();
 b15zdnd11an1n04x5 FILLER_180_1415 ();
 b15zdnd00an1n02x5 FILLER_180_1419 ();
 b15zdnd11an1n32x5 FILLER_180_1437 ();
 b15zdnd11an1n16x5 FILLER_180_1469 ();
 b15zdnd11an1n08x5 FILLER_180_1485 ();
 b15zdnd11an1n64x5 FILLER_180_1501 ();
 b15zdnd11an1n32x5 FILLER_180_1565 ();
 b15zdnd11an1n16x5 FILLER_180_1597 ();
 b15zdnd11an1n04x5 FILLER_180_1613 ();
 b15zdnd11an1n32x5 FILLER_180_1624 ();
 b15zdnd11an1n08x5 FILLER_180_1656 ();
 b15zdnd11an1n64x5 FILLER_180_1680 ();
 b15zdnd11an1n32x5 FILLER_180_1744 ();
 b15zdnd00an1n02x5 FILLER_180_1776 ();
 b15zdnd00an1n01x5 FILLER_180_1778 ();
 b15zdnd11an1n64x5 FILLER_180_1788 ();
 b15zdnd11an1n32x5 FILLER_180_1852 ();
 b15zdnd11an1n16x5 FILLER_180_1884 ();
 b15zdnd11an1n08x5 FILLER_180_1900 ();
 b15zdnd11an1n04x5 FILLER_180_1908 ();
 b15zdnd00an1n02x5 FILLER_180_1912 ();
 b15zdnd00an1n01x5 FILLER_180_1914 ();
 b15zdnd11an1n08x5 FILLER_180_1921 ();
 b15zdnd11an1n08x5 FILLER_180_1935 ();
 b15zdnd11an1n04x5 FILLER_180_1943 ();
 b15zdnd00an1n01x5 FILLER_180_1947 ();
 b15zdnd11an1n64x5 FILLER_180_1968 ();
 b15zdnd11an1n16x5 FILLER_180_2032 ();
 b15zdnd11an1n08x5 FILLER_180_2048 ();
 b15zdnd00an1n02x5 FILLER_180_2056 ();
 b15zdnd11an1n64x5 FILLER_180_2079 ();
 b15zdnd11an1n08x5 FILLER_180_2143 ();
 b15zdnd00an1n02x5 FILLER_180_2151 ();
 b15zdnd00an1n01x5 FILLER_180_2153 ();
 b15zdnd11an1n16x5 FILLER_180_2162 ();
 b15zdnd11an1n04x5 FILLER_180_2178 ();
 b15zdnd11an1n32x5 FILLER_180_2193 ();
 b15zdnd11an1n04x5 FILLER_180_2225 ();
 b15zdnd00an1n02x5 FILLER_180_2229 ();
 b15zdnd11an1n08x5 FILLER_180_2234 ();
 b15zdnd11an1n04x5 FILLER_180_2242 ();
 b15zdnd11an1n04x5 FILLER_180_2250 ();
 b15zdnd11an1n16x5 FILLER_180_2258 ();
 b15zdnd00an1n02x5 FILLER_180_2274 ();
 b15zdnd11an1n32x5 FILLER_181_0 ();
 b15zdnd11an1n04x5 FILLER_181_32 ();
 b15zdnd00an1n02x5 FILLER_181_36 ();
 b15zdnd11an1n04x5 FILLER_181_43 ();
 b15zdnd11an1n32x5 FILLER_181_52 ();
 b15zdnd11an1n04x5 FILLER_181_84 ();
 b15zdnd00an1n02x5 FILLER_181_88 ();
 b15zdnd11an1n16x5 FILLER_181_97 ();
 b15zdnd00an1n02x5 FILLER_181_113 ();
 b15zdnd11an1n16x5 FILLER_181_119 ();
 b15zdnd11an1n08x5 FILLER_181_135 ();
 b15zdnd11an1n04x5 FILLER_181_143 ();
 b15zdnd11an1n16x5 FILLER_181_154 ();
 b15zdnd00an1n01x5 FILLER_181_170 ();
 b15zdnd11an1n16x5 FILLER_181_183 ();
 b15zdnd11an1n32x5 FILLER_181_204 ();
 b15zdnd11an1n04x5 FILLER_181_236 ();
 b15zdnd00an1n02x5 FILLER_181_240 ();
 b15zdnd11an1n16x5 FILLER_181_247 ();
 b15zdnd11an1n04x5 FILLER_181_263 ();
 b15zdnd00an1n01x5 FILLER_181_267 ();
 b15zdnd11an1n64x5 FILLER_181_274 ();
 b15zdnd11an1n32x5 FILLER_181_338 ();
 b15zdnd11an1n16x5 FILLER_181_370 ();
 b15zdnd11an1n04x5 FILLER_181_386 ();
 b15zdnd00an1n02x5 FILLER_181_390 ();
 b15zdnd11an1n16x5 FILLER_181_420 ();
 b15zdnd11an1n08x5 FILLER_181_436 ();
 b15zdnd00an1n02x5 FILLER_181_444 ();
 b15zdnd00an1n01x5 FILLER_181_446 ();
 b15zdnd11an1n04x5 FILLER_181_463 ();
 b15zdnd11an1n04x5 FILLER_181_483 ();
 b15zdnd11an1n04x5 FILLER_181_493 ();
 b15zdnd11an1n04x5 FILLER_181_513 ();
 b15zdnd11an1n16x5 FILLER_181_526 ();
 b15zdnd11an1n08x5 FILLER_181_542 ();
 b15zdnd11an1n04x5 FILLER_181_550 ();
 b15zdnd00an1n02x5 FILLER_181_554 ();
 b15zdnd00an1n01x5 FILLER_181_556 ();
 b15zdnd11an1n16x5 FILLER_181_565 ();
 b15zdnd11an1n32x5 FILLER_181_602 ();
 b15zdnd11an1n04x5 FILLER_181_634 ();
 b15zdnd00an1n01x5 FILLER_181_638 ();
 b15zdnd11an1n64x5 FILLER_181_645 ();
 b15zdnd11an1n08x5 FILLER_181_719 ();
 b15zdnd00an1n02x5 FILLER_181_727 ();
 b15zdnd11an1n04x5 FILLER_181_736 ();
 b15zdnd11an1n64x5 FILLER_181_744 ();
 b15zdnd11an1n64x5 FILLER_181_808 ();
 b15zdnd11an1n32x5 FILLER_181_872 ();
 b15zdnd11an1n08x5 FILLER_181_904 ();
 b15zdnd00an1n01x5 FILLER_181_912 ();
 b15zdnd11an1n32x5 FILLER_181_929 ();
 b15zdnd11an1n08x5 FILLER_181_961 ();
 b15zdnd11an1n04x5 FILLER_181_969 ();
 b15zdnd00an1n01x5 FILLER_181_973 ();
 b15zdnd11an1n16x5 FILLER_181_992 ();
 b15zdnd11an1n08x5 FILLER_181_1008 ();
 b15zdnd11an1n04x5 FILLER_181_1016 ();
 b15zdnd00an1n02x5 FILLER_181_1020 ();
 b15zdnd00an1n01x5 FILLER_181_1022 ();
 b15zdnd11an1n64x5 FILLER_181_1028 ();
 b15zdnd11an1n16x5 FILLER_181_1092 ();
 b15zdnd11an1n04x5 FILLER_181_1108 ();
 b15zdnd00an1n02x5 FILLER_181_1112 ();
 b15zdnd00an1n01x5 FILLER_181_1114 ();
 b15zdnd11an1n32x5 FILLER_181_1122 ();
 b15zdnd11an1n16x5 FILLER_181_1154 ();
 b15zdnd11an1n08x5 FILLER_181_1170 ();
 b15zdnd11an1n04x5 FILLER_181_1178 ();
 b15zdnd11an1n04x5 FILLER_181_1192 ();
 b15zdnd11an1n08x5 FILLER_181_1210 ();
 b15zdnd11an1n04x5 FILLER_181_1218 ();
 b15zdnd00an1n01x5 FILLER_181_1222 ();
 b15zdnd11an1n04x5 FILLER_181_1239 ();
 b15zdnd11an1n32x5 FILLER_181_1268 ();
 b15zdnd11an1n04x5 FILLER_181_1300 ();
 b15zdnd00an1n02x5 FILLER_181_1304 ();
 b15zdnd00an1n01x5 FILLER_181_1306 ();
 b15zdnd11an1n04x5 FILLER_181_1315 ();
 b15zdnd11an1n04x5 FILLER_181_1333 ();
 b15zdnd00an1n01x5 FILLER_181_1337 ();
 b15zdnd11an1n64x5 FILLER_181_1352 ();
 b15zdnd11an1n32x5 FILLER_181_1416 ();
 b15zdnd11an1n04x5 FILLER_181_1453 ();
 b15zdnd11an1n32x5 FILLER_181_1463 ();
 b15zdnd11an1n16x5 FILLER_181_1495 ();
 b15zdnd11an1n08x5 FILLER_181_1511 ();
 b15zdnd00an1n02x5 FILLER_181_1519 ();
 b15zdnd11an1n08x5 FILLER_181_1528 ();
 b15zdnd11an1n04x5 FILLER_181_1536 ();
 b15zdnd00an1n02x5 FILLER_181_1540 ();
 b15zdnd00an1n01x5 FILLER_181_1542 ();
 b15zdnd11an1n32x5 FILLER_181_1550 ();
 b15zdnd11an1n16x5 FILLER_181_1582 ();
 b15zdnd11an1n04x5 FILLER_181_1598 ();
 b15zdnd00an1n02x5 FILLER_181_1602 ();
 b15zdnd11an1n04x5 FILLER_181_1608 ();
 b15zdnd11an1n04x5 FILLER_181_1617 ();
 b15zdnd11an1n08x5 FILLER_181_1639 ();
 b15zdnd11an1n04x5 FILLER_181_1647 ();
 b15zdnd00an1n01x5 FILLER_181_1651 ();
 b15zdnd11an1n32x5 FILLER_181_1683 ();
 b15zdnd11an1n08x5 FILLER_181_1715 ();
 b15zdnd00an1n01x5 FILLER_181_1723 ();
 b15zdnd11an1n04x5 FILLER_181_1735 ();
 b15zdnd00an1n02x5 FILLER_181_1739 ();
 b15zdnd11an1n08x5 FILLER_181_1761 ();
 b15zdnd11an1n04x5 FILLER_181_1769 ();
 b15zdnd11an1n32x5 FILLER_181_1793 ();
 b15zdnd11an1n16x5 FILLER_181_1825 ();
 b15zdnd11an1n08x5 FILLER_181_1841 ();
 b15zdnd00an1n01x5 FILLER_181_1849 ();
 b15zdnd11an1n64x5 FILLER_181_1870 ();
 b15zdnd11an1n64x5 FILLER_181_1934 ();
 b15zdnd11an1n32x5 FILLER_181_1998 ();
 b15zdnd11an1n08x5 FILLER_181_2030 ();
 b15zdnd00an1n01x5 FILLER_181_2038 ();
 b15zdnd11an1n04x5 FILLER_181_2071 ();
 b15zdnd00an1n01x5 FILLER_181_2075 ();
 b15zdnd11an1n16x5 FILLER_181_2085 ();
 b15zdnd11an1n08x5 FILLER_181_2101 ();
 b15zdnd11an1n04x5 FILLER_181_2109 ();
 b15zdnd11an1n08x5 FILLER_181_2138 ();
 b15zdnd11an1n04x5 FILLER_181_2146 ();
 b15zdnd00an1n02x5 FILLER_181_2150 ();
 b15zdnd00an1n01x5 FILLER_181_2152 ();
 b15zdnd11an1n04x5 FILLER_181_2184 ();
 b15zdnd11an1n32x5 FILLER_181_2208 ();
 b15zdnd11an1n04x5 FILLER_181_2240 ();
 b15zdnd00an1n02x5 FILLER_181_2244 ();
 b15zdnd11an1n04x5 FILLER_181_2254 ();
 b15zdnd00an1n02x5 FILLER_181_2258 ();
 b15zdnd11an1n08x5 FILLER_181_2264 ();
 b15zdnd11an1n04x5 FILLER_181_2272 ();
 b15zdnd11an1n04x5 FILLER_181_2280 ();
 b15zdnd11an1n64x5 FILLER_182_8 ();
 b15zdnd11an1n04x5 FILLER_182_72 ();
 b15zdnd00an1n01x5 FILLER_182_76 ();
 b15zdnd11an1n16x5 FILLER_182_93 ();
 b15zdnd11an1n04x5 FILLER_182_109 ();
 b15zdnd00an1n01x5 FILLER_182_113 ();
 b15zdnd11an1n64x5 FILLER_182_121 ();
 b15zdnd11an1n64x5 FILLER_182_185 ();
 b15zdnd11an1n08x5 FILLER_182_249 ();
 b15zdnd11an1n04x5 FILLER_182_257 ();
 b15zdnd11an1n64x5 FILLER_182_266 ();
 b15zdnd11an1n04x5 FILLER_182_330 ();
 b15zdnd00an1n02x5 FILLER_182_334 ();
 b15zdnd11an1n16x5 FILLER_182_368 ();
 b15zdnd11an1n08x5 FILLER_182_384 ();
 b15zdnd11an1n04x5 FILLER_182_406 ();
 b15zdnd00an1n01x5 FILLER_182_410 ();
 b15zdnd11an1n08x5 FILLER_182_442 ();
 b15zdnd00an1n02x5 FILLER_182_450 ();
 b15zdnd11an1n16x5 FILLER_182_462 ();
 b15zdnd11an1n04x5 FILLER_182_478 ();
 b15zdnd00an1n02x5 FILLER_182_482 ();
 b15zdnd11an1n64x5 FILLER_182_489 ();
 b15zdnd11an1n64x5 FILLER_182_553 ();
 b15zdnd11an1n16x5 FILLER_182_617 ();
 b15zdnd11an1n08x5 FILLER_182_633 ();
 b15zdnd00an1n02x5 FILLER_182_641 ();
 b15zdnd11an1n04x5 FILLER_182_649 ();
 b15zdnd00an1n02x5 FILLER_182_653 ();
 b15zdnd00an1n01x5 FILLER_182_655 ();
 b15zdnd11an1n04x5 FILLER_182_676 ();
 b15zdnd11an1n08x5 FILLER_182_696 ();
 b15zdnd11an1n04x5 FILLER_182_714 ();
 b15zdnd11an1n08x5 FILLER_182_726 ();
 b15zdnd11an1n04x5 FILLER_182_734 ();
 b15zdnd00an1n01x5 FILLER_182_738 ();
 b15zdnd11an1n04x5 FILLER_182_765 ();
 b15zdnd11an1n32x5 FILLER_182_773 ();
 b15zdnd11an1n16x5 FILLER_182_805 ();
 b15zdnd11an1n08x5 FILLER_182_821 ();
 b15zdnd00an1n02x5 FILLER_182_829 ();
 b15zdnd00an1n01x5 FILLER_182_831 ();
 b15zdnd11an1n04x5 FILLER_182_837 ();
 b15zdnd11an1n32x5 FILLER_182_850 ();
 b15zdnd11an1n04x5 FILLER_182_882 ();
 b15zdnd11an1n16x5 FILLER_182_892 ();
 b15zdnd11an1n08x5 FILLER_182_908 ();
 b15zdnd11an1n04x5 FILLER_182_916 ();
 b15zdnd00an1n02x5 FILLER_182_920 ();
 b15zdnd11an1n08x5 FILLER_182_942 ();
 b15zdnd00an1n02x5 FILLER_182_950 ();
 b15zdnd00an1n01x5 FILLER_182_952 ();
 b15zdnd11an1n04x5 FILLER_182_960 ();
 b15zdnd11an1n08x5 FILLER_182_973 ();
 b15zdnd00an1n01x5 FILLER_182_981 ();
 b15zdnd11an1n32x5 FILLER_182_987 ();
 b15zdnd00an1n02x5 FILLER_182_1019 ();
 b15zdnd00an1n01x5 FILLER_182_1021 ();
 b15zdnd11an1n08x5 FILLER_182_1029 ();
 b15zdnd11an1n04x5 FILLER_182_1037 ();
 b15zdnd00an1n02x5 FILLER_182_1041 ();
 b15zdnd11an1n16x5 FILLER_182_1053 ();
 b15zdnd11an1n04x5 FILLER_182_1069 ();
 b15zdnd11an1n16x5 FILLER_182_1078 ();
 b15zdnd00an1n01x5 FILLER_182_1094 ();
 b15zdnd11an1n64x5 FILLER_182_1106 ();
 b15zdnd11an1n08x5 FILLER_182_1170 ();
 b15zdnd11an1n04x5 FILLER_182_1178 ();
 b15zdnd11an1n04x5 FILLER_182_1187 ();
 b15zdnd11an1n64x5 FILLER_182_1211 ();
 b15zdnd11an1n32x5 FILLER_182_1275 ();
 b15zdnd11an1n16x5 FILLER_182_1307 ();
 b15zdnd11an1n04x5 FILLER_182_1323 ();
 b15zdnd00an1n02x5 FILLER_182_1327 ();
 b15zdnd00an1n01x5 FILLER_182_1329 ();
 b15zdnd11an1n04x5 FILLER_182_1340 ();
 b15zdnd00an1n02x5 FILLER_182_1344 ();
 b15zdnd11an1n16x5 FILLER_182_1352 ();
 b15zdnd11an1n08x5 FILLER_182_1368 ();
 b15zdnd11an1n64x5 FILLER_182_1394 ();
 b15zdnd11an1n32x5 FILLER_182_1462 ();
 b15zdnd11an1n16x5 FILLER_182_1494 ();
 b15zdnd11an1n08x5 FILLER_182_1510 ();
 b15zdnd11an1n04x5 FILLER_182_1518 ();
 b15zdnd00an1n02x5 FILLER_182_1522 ();
 b15zdnd11an1n08x5 FILLER_182_1530 ();
 b15zdnd11an1n04x5 FILLER_182_1538 ();
 b15zdnd00an1n02x5 FILLER_182_1542 ();
 b15zdnd11an1n16x5 FILLER_182_1556 ();
 b15zdnd11an1n08x5 FILLER_182_1572 ();
 b15zdnd11an1n08x5 FILLER_182_1592 ();
 b15zdnd11an1n04x5 FILLER_182_1600 ();
 b15zdnd11an1n64x5 FILLER_182_1610 ();
 b15zdnd11an1n64x5 FILLER_182_1674 ();
 b15zdnd11an1n16x5 FILLER_182_1738 ();
 b15zdnd11an1n08x5 FILLER_182_1754 ();
 b15zdnd00an1n02x5 FILLER_182_1762 ();
 b15zdnd00an1n01x5 FILLER_182_1764 ();
 b15zdnd11an1n04x5 FILLER_182_1774 ();
 b15zdnd11an1n16x5 FILLER_182_1783 ();
 b15zdnd11an1n08x5 FILLER_182_1799 ();
 b15zdnd00an1n02x5 FILLER_182_1807 ();
 b15zdnd11an1n04x5 FILLER_182_1829 ();
 b15zdnd11an1n64x5 FILLER_182_1838 ();
 b15zdnd11an1n32x5 FILLER_182_1902 ();
 b15zdnd11an1n16x5 FILLER_182_1934 ();
 b15zdnd11an1n04x5 FILLER_182_1950 ();
 b15zdnd00an1n02x5 FILLER_182_1954 ();
 b15zdnd11an1n64x5 FILLER_182_1974 ();
 b15zdnd11an1n64x5 FILLER_182_2038 ();
 b15zdnd11an1n32x5 FILLER_182_2102 ();
 b15zdnd11an1n16x5 FILLER_182_2134 ();
 b15zdnd11an1n04x5 FILLER_182_2150 ();
 b15zdnd11an1n64x5 FILLER_182_2162 ();
 b15zdnd11an1n16x5 FILLER_182_2226 ();
 b15zdnd00an1n01x5 FILLER_182_2242 ();
 b15zdnd11an1n08x5 FILLER_182_2251 ();
 b15zdnd00an1n02x5 FILLER_182_2259 ();
 b15zdnd11an1n08x5 FILLER_182_2265 ();
 b15zdnd00an1n02x5 FILLER_182_2273 ();
 b15zdnd00an1n01x5 FILLER_182_2275 ();
 b15zdnd11an1n32x5 FILLER_183_0 ();
 b15zdnd11an1n04x5 FILLER_183_32 ();
 b15zdnd00an1n02x5 FILLER_183_36 ();
 b15zdnd11an1n16x5 FILLER_183_56 ();
 b15zdnd11an1n04x5 FILLER_183_72 ();
 b15zdnd00an1n02x5 FILLER_183_76 ();
 b15zdnd00an1n01x5 FILLER_183_78 ();
 b15zdnd11an1n04x5 FILLER_183_83 ();
 b15zdnd11an1n16x5 FILLER_183_93 ();
 b15zdnd11an1n08x5 FILLER_183_109 ();
 b15zdnd11an1n04x5 FILLER_183_117 ();
 b15zdnd00an1n01x5 FILLER_183_121 ();
 b15zdnd11an1n08x5 FILLER_183_130 ();
 b15zdnd11an1n04x5 FILLER_183_138 ();
 b15zdnd00an1n02x5 FILLER_183_142 ();
 b15zdnd11an1n32x5 FILLER_183_150 ();
 b15zdnd00an1n02x5 FILLER_183_182 ();
 b15zdnd00an1n01x5 FILLER_183_184 ();
 b15zdnd11an1n64x5 FILLER_183_205 ();
 b15zdnd11an1n64x5 FILLER_183_269 ();
 b15zdnd11an1n32x5 FILLER_183_333 ();
 b15zdnd11an1n16x5 FILLER_183_365 ();
 b15zdnd11an1n08x5 FILLER_183_381 ();
 b15zdnd11an1n04x5 FILLER_183_389 ();
 b15zdnd00an1n02x5 FILLER_183_393 ();
 b15zdnd11an1n32x5 FILLER_183_405 ();
 b15zdnd11an1n16x5 FILLER_183_437 ();
 b15zdnd00an1n02x5 FILLER_183_453 ();
 b15zdnd11an1n04x5 FILLER_183_468 ();
 b15zdnd11an1n32x5 FILLER_183_497 ();
 b15zdnd11an1n04x5 FILLER_183_529 ();
 b15zdnd11an1n04x5 FILLER_183_543 ();
 b15zdnd00an1n01x5 FILLER_183_547 ();
 b15zdnd11an1n04x5 FILLER_183_552 ();
 b15zdnd11an1n08x5 FILLER_183_564 ();
 b15zdnd00an1n02x5 FILLER_183_572 ();
 b15zdnd11an1n64x5 FILLER_183_580 ();
 b15zdnd11an1n04x5 FILLER_183_644 ();
 b15zdnd00an1n02x5 FILLER_183_648 ();
 b15zdnd11an1n08x5 FILLER_183_655 ();
 b15zdnd11an1n04x5 FILLER_183_663 ();
 b15zdnd00an1n01x5 FILLER_183_667 ();
 b15zdnd11an1n04x5 FILLER_183_679 ();
 b15zdnd11an1n08x5 FILLER_183_693 ();
 b15zdnd11an1n04x5 FILLER_183_701 ();
 b15zdnd00an1n02x5 FILLER_183_705 ();
 b15zdnd11an1n16x5 FILLER_183_714 ();
 b15zdnd11an1n08x5 FILLER_183_730 ();
 b15zdnd00an1n01x5 FILLER_183_738 ();
 b15zdnd11an1n08x5 FILLER_183_765 ();
 b15zdnd11an1n32x5 FILLER_183_782 ();
 b15zdnd11an1n08x5 FILLER_183_814 ();
 b15zdnd11an1n04x5 FILLER_183_822 ();
 b15zdnd00an1n01x5 FILLER_183_826 ();
 b15zdnd11an1n08x5 FILLER_183_839 ();
 b15zdnd11an1n08x5 FILLER_183_856 ();
 b15zdnd11an1n04x5 FILLER_183_864 ();
 b15zdnd11an1n04x5 FILLER_183_876 ();
 b15zdnd11an1n08x5 FILLER_183_887 ();
 b15zdnd11an1n04x5 FILLER_183_895 ();
 b15zdnd11an1n04x5 FILLER_183_907 ();
 b15zdnd11an1n64x5 FILLER_183_920 ();
 b15zdnd11an1n64x5 FILLER_183_984 ();
 b15zdnd11an1n16x5 FILLER_183_1048 ();
 b15zdnd11an1n04x5 FILLER_183_1064 ();
 b15zdnd00an1n01x5 FILLER_183_1068 ();
 b15zdnd11an1n64x5 FILLER_183_1084 ();
 b15zdnd11an1n64x5 FILLER_183_1148 ();
 b15zdnd11an1n32x5 FILLER_183_1212 ();
 b15zdnd11an1n16x5 FILLER_183_1244 ();
 b15zdnd11an1n04x5 FILLER_183_1260 ();
 b15zdnd00an1n02x5 FILLER_183_1264 ();
 b15zdnd11an1n08x5 FILLER_183_1298 ();
 b15zdnd11an1n04x5 FILLER_183_1306 ();
 b15zdnd00an1n02x5 FILLER_183_1310 ();
 b15zdnd11an1n16x5 FILLER_183_1320 ();
 b15zdnd11an1n04x5 FILLER_183_1340 ();
 b15zdnd00an1n01x5 FILLER_183_1344 ();
 b15zdnd11an1n16x5 FILLER_183_1354 ();
 b15zdnd11an1n08x5 FILLER_183_1370 ();
 b15zdnd11an1n16x5 FILLER_183_1392 ();
 b15zdnd11an1n04x5 FILLER_183_1408 ();
 b15zdnd11an1n08x5 FILLER_183_1433 ();
 b15zdnd00an1n01x5 FILLER_183_1441 ();
 b15zdnd11an1n64x5 FILLER_183_1452 ();
 b15zdnd11an1n32x5 FILLER_183_1516 ();
 b15zdnd11an1n16x5 FILLER_183_1548 ();
 b15zdnd11an1n08x5 FILLER_183_1564 ();
 b15zdnd00an1n02x5 FILLER_183_1572 ();
 b15zdnd00an1n01x5 FILLER_183_1574 ();
 b15zdnd11an1n16x5 FILLER_183_1601 ();
 b15zdnd00an1n01x5 FILLER_183_1617 ();
 b15zdnd11an1n16x5 FILLER_183_1625 ();
 b15zdnd11an1n08x5 FILLER_183_1641 ();
 b15zdnd00an1n02x5 FILLER_183_1649 ();
 b15zdnd11an1n32x5 FILLER_183_1666 ();
 b15zdnd11an1n08x5 FILLER_183_1698 ();
 b15zdnd00an1n02x5 FILLER_183_1706 ();
 b15zdnd00an1n01x5 FILLER_183_1708 ();
 b15zdnd11an1n32x5 FILLER_183_1729 ();
 b15zdnd11an1n08x5 FILLER_183_1761 ();
 b15zdnd11an1n04x5 FILLER_183_1769 ();
 b15zdnd00an1n02x5 FILLER_183_1773 ();
 b15zdnd00an1n01x5 FILLER_183_1775 ();
 b15zdnd11an1n64x5 FILLER_183_1802 ();
 b15zdnd11an1n64x5 FILLER_183_1866 ();
 b15zdnd11an1n64x5 FILLER_183_1930 ();
 b15zdnd11an1n64x5 FILLER_183_1994 ();
 b15zdnd11an1n64x5 FILLER_183_2058 ();
 b15zdnd11an1n16x5 FILLER_183_2122 ();
 b15zdnd11an1n08x5 FILLER_183_2138 ();
 b15zdnd11an1n64x5 FILLER_183_2166 ();
 b15zdnd11an1n08x5 FILLER_183_2230 ();
 b15zdnd11an1n04x5 FILLER_183_2238 ();
 b15zdnd11an1n16x5 FILLER_183_2246 ();
 b15zdnd11an1n04x5 FILLER_183_2262 ();
 b15zdnd11an1n08x5 FILLER_183_2271 ();
 b15zdnd11an1n04x5 FILLER_183_2279 ();
 b15zdnd00an1n01x5 FILLER_183_2283 ();
 b15zdnd11an1n32x5 FILLER_184_8 ();
 b15zdnd11an1n04x5 FILLER_184_40 ();
 b15zdnd00an1n02x5 FILLER_184_44 ();
 b15zdnd00an1n01x5 FILLER_184_46 ();
 b15zdnd11an1n16x5 FILLER_184_59 ();
 b15zdnd11an1n08x5 FILLER_184_75 ();
 b15zdnd11an1n04x5 FILLER_184_83 ();
 b15zdnd00an1n01x5 FILLER_184_87 ();
 b15zdnd11an1n16x5 FILLER_184_94 ();
 b15zdnd11an1n08x5 FILLER_184_110 ();
 b15zdnd00an1n02x5 FILLER_184_118 ();
 b15zdnd11an1n16x5 FILLER_184_124 ();
 b15zdnd11an1n04x5 FILLER_184_140 ();
 b15zdnd00an1n02x5 FILLER_184_144 ();
 b15zdnd00an1n01x5 FILLER_184_146 ();
 b15zdnd11an1n64x5 FILLER_184_155 ();
 b15zdnd11an1n04x5 FILLER_184_219 ();
 b15zdnd11an1n16x5 FILLER_184_231 ();
 b15zdnd11an1n04x5 FILLER_184_247 ();
 b15zdnd00an1n01x5 FILLER_184_251 ();
 b15zdnd11an1n04x5 FILLER_184_278 ();
 b15zdnd11an1n08x5 FILLER_184_298 ();
 b15zdnd00an1n02x5 FILLER_184_306 ();
 b15zdnd11an1n32x5 FILLER_184_334 ();
 b15zdnd11an1n08x5 FILLER_184_366 ();
 b15zdnd11an1n04x5 FILLER_184_374 ();
 b15zdnd00an1n02x5 FILLER_184_378 ();
 b15zdnd00an1n01x5 FILLER_184_380 ();
 b15zdnd11an1n32x5 FILLER_184_387 ();
 b15zdnd11an1n16x5 FILLER_184_419 ();
 b15zdnd11an1n04x5 FILLER_184_435 ();
 b15zdnd11an1n16x5 FILLER_184_459 ();
 b15zdnd00an1n01x5 FILLER_184_475 ();
 b15zdnd11an1n16x5 FILLER_184_488 ();
 b15zdnd00an1n02x5 FILLER_184_504 ();
 b15zdnd11an1n08x5 FILLER_184_521 ();
 b15zdnd00an1n01x5 FILLER_184_529 ();
 b15zdnd11an1n16x5 FILLER_184_546 ();
 b15zdnd11an1n08x5 FILLER_184_562 ();
 b15zdnd00an1n02x5 FILLER_184_570 ();
 b15zdnd11an1n08x5 FILLER_184_585 ();
 b15zdnd00an1n02x5 FILLER_184_593 ();
 b15zdnd00an1n01x5 FILLER_184_595 ();
 b15zdnd11an1n16x5 FILLER_184_606 ();
 b15zdnd11an1n32x5 FILLER_184_627 ();
 b15zdnd11an1n16x5 FILLER_184_659 ();
 b15zdnd00an1n01x5 FILLER_184_675 ();
 b15zdnd11an1n08x5 FILLER_184_686 ();
 b15zdnd11an1n04x5 FILLER_184_694 ();
 b15zdnd00an1n02x5 FILLER_184_698 ();
 b15zdnd11an1n08x5 FILLER_184_704 ();
 b15zdnd11an1n04x5 FILLER_184_712 ();
 b15zdnd00an1n02x5 FILLER_184_716 ();
 b15zdnd11an1n64x5 FILLER_184_726 ();
 b15zdnd11an1n32x5 FILLER_184_790 ();
 b15zdnd11an1n16x5 FILLER_184_822 ();
 b15zdnd00an1n02x5 FILLER_184_838 ();
 b15zdnd11an1n32x5 FILLER_184_848 ();
 b15zdnd11an1n04x5 FILLER_184_880 ();
 b15zdnd00an1n01x5 FILLER_184_884 ();
 b15zdnd11an1n64x5 FILLER_184_892 ();
 b15zdnd11an1n32x5 FILLER_184_956 ();
 b15zdnd11an1n16x5 FILLER_184_988 ();
 b15zdnd11an1n04x5 FILLER_184_1004 ();
 b15zdnd00an1n02x5 FILLER_184_1008 ();
 b15zdnd00an1n01x5 FILLER_184_1010 ();
 b15zdnd11an1n16x5 FILLER_184_1016 ();
 b15zdnd00an1n02x5 FILLER_184_1032 ();
 b15zdnd11an1n32x5 FILLER_184_1054 ();
 b15zdnd11an1n08x5 FILLER_184_1086 ();
 b15zdnd11an1n04x5 FILLER_184_1094 ();
 b15zdnd00an1n02x5 FILLER_184_1098 ();
 b15zdnd11an1n32x5 FILLER_184_1112 ();
 b15zdnd11an1n04x5 FILLER_184_1160 ();
 b15zdnd00an1n01x5 FILLER_184_1164 ();
 b15zdnd11an1n32x5 FILLER_184_1179 ();
 b15zdnd11an1n08x5 FILLER_184_1211 ();
 b15zdnd00an1n02x5 FILLER_184_1219 ();
 b15zdnd11an1n64x5 FILLER_184_1247 ();
 b15zdnd11an1n16x5 FILLER_184_1311 ();
 b15zdnd11an1n04x5 FILLER_184_1327 ();
 b15zdnd00an1n02x5 FILLER_184_1331 ();
 b15zdnd00an1n01x5 FILLER_184_1333 ();
 b15zdnd11an1n64x5 FILLER_184_1345 ();
 b15zdnd11an1n64x5 FILLER_184_1409 ();
 b15zdnd11an1n32x5 FILLER_184_1473 ();
 b15zdnd11an1n16x5 FILLER_184_1505 ();
 b15zdnd11an1n04x5 FILLER_184_1521 ();
 b15zdnd00an1n01x5 FILLER_184_1525 ();
 b15zdnd11an1n16x5 FILLER_184_1531 ();
 b15zdnd11an1n08x5 FILLER_184_1547 ();
 b15zdnd11an1n04x5 FILLER_184_1555 ();
 b15zdnd11an1n32x5 FILLER_184_1565 ();
 b15zdnd00an1n02x5 FILLER_184_1597 ();
 b15zdnd00an1n01x5 FILLER_184_1599 ();
 b15zdnd11an1n64x5 FILLER_184_1607 ();
 b15zdnd11an1n64x5 FILLER_184_1671 ();
 b15zdnd11an1n64x5 FILLER_184_1735 ();
 b15zdnd11an1n08x5 FILLER_184_1799 ();
 b15zdnd00an1n02x5 FILLER_184_1807 ();
 b15zdnd11an1n32x5 FILLER_184_1840 ();
 b15zdnd11an1n04x5 FILLER_184_1872 ();
 b15zdnd00an1n02x5 FILLER_184_1876 ();
 b15zdnd11an1n08x5 FILLER_184_1883 ();
 b15zdnd11an1n04x5 FILLER_184_1891 ();
 b15zdnd00an1n02x5 FILLER_184_1895 ();
 b15zdnd00an1n01x5 FILLER_184_1897 ();
 b15zdnd11an1n04x5 FILLER_184_1909 ();
 b15zdnd11an1n04x5 FILLER_184_1917 ();
 b15zdnd11an1n32x5 FILLER_184_1927 ();
 b15zdnd11an1n04x5 FILLER_184_1984 ();
 b15zdnd00an1n02x5 FILLER_184_1988 ();
 b15zdnd00an1n01x5 FILLER_184_1990 ();
 b15zdnd11an1n08x5 FILLER_184_2003 ();
 b15zdnd11an1n04x5 FILLER_184_2011 ();
 b15zdnd00an1n01x5 FILLER_184_2015 ();
 b15zdnd11an1n32x5 FILLER_184_2036 ();
 b15zdnd00an1n02x5 FILLER_184_2068 ();
 b15zdnd11an1n64x5 FILLER_184_2082 ();
 b15zdnd11an1n08x5 FILLER_184_2146 ();
 b15zdnd11an1n32x5 FILLER_184_2162 ();
 b15zdnd11an1n16x5 FILLER_184_2194 ();
 b15zdnd11an1n08x5 FILLER_184_2210 ();
 b15zdnd11an1n04x5 FILLER_184_2218 ();
 b15zdnd00an1n02x5 FILLER_184_2222 ();
 b15zdnd00an1n01x5 FILLER_184_2224 ();
 b15zdnd11an1n16x5 FILLER_184_2231 ();
 b15zdnd11an1n04x5 FILLER_184_2250 ();
 b15zdnd11an1n08x5 FILLER_184_2262 ();
 b15zdnd11an1n04x5 FILLER_184_2270 ();
 b15zdnd00an1n02x5 FILLER_184_2274 ();
 b15zdnd11an1n08x5 FILLER_185_0 ();
 b15zdnd11an1n04x5 FILLER_185_8 ();
 b15zdnd00an1n02x5 FILLER_185_12 ();
 b15zdnd00an1n01x5 FILLER_185_14 ();
 b15zdnd11an1n32x5 FILLER_185_23 ();
 b15zdnd11an1n04x5 FILLER_185_61 ();
 b15zdnd11an1n08x5 FILLER_185_71 ();
 b15zdnd11an1n04x5 FILLER_185_79 ();
 b15zdnd00an1n01x5 FILLER_185_83 ();
 b15zdnd11an1n32x5 FILLER_185_89 ();
 b15zdnd11an1n16x5 FILLER_185_121 ();
 b15zdnd11an1n08x5 FILLER_185_137 ();
 b15zdnd00an1n02x5 FILLER_185_145 ();
 b15zdnd00an1n01x5 FILLER_185_147 ();
 b15zdnd11an1n04x5 FILLER_185_156 ();
 b15zdnd00an1n01x5 FILLER_185_160 ();
 b15zdnd11an1n32x5 FILLER_185_187 ();
 b15zdnd00an1n01x5 FILLER_185_219 ();
 b15zdnd11an1n16x5 FILLER_185_236 ();
 b15zdnd00an1n01x5 FILLER_185_252 ();
 b15zdnd11an1n04x5 FILLER_185_260 ();
 b15zdnd11an1n16x5 FILLER_185_280 ();
 b15zdnd11an1n04x5 FILLER_185_296 ();
 b15zdnd11an1n32x5 FILLER_185_312 ();
 b15zdnd11an1n16x5 FILLER_185_344 ();
 b15zdnd11an1n08x5 FILLER_185_360 ();
 b15zdnd11an1n04x5 FILLER_185_374 ();
 b15zdnd11an1n32x5 FILLER_185_392 ();
 b15zdnd11an1n08x5 FILLER_185_424 ();
 b15zdnd00an1n01x5 FILLER_185_432 ();
 b15zdnd11an1n32x5 FILLER_185_447 ();
 b15zdnd11an1n04x5 FILLER_185_479 ();
 b15zdnd11an1n16x5 FILLER_185_487 ();
 b15zdnd11an1n08x5 FILLER_185_503 ();
 b15zdnd11an1n04x5 FILLER_185_511 ();
 b15zdnd00an1n02x5 FILLER_185_515 ();
 b15zdnd11an1n32x5 FILLER_185_523 ();
 b15zdnd11an1n16x5 FILLER_185_555 ();
 b15zdnd11an1n08x5 FILLER_185_571 ();
 b15zdnd11an1n04x5 FILLER_185_579 ();
 b15zdnd00an1n01x5 FILLER_185_583 ();
 b15zdnd11an1n04x5 FILLER_185_605 ();
 b15zdnd11an1n04x5 FILLER_185_615 ();
 b15zdnd00an1n02x5 FILLER_185_619 ();
 b15zdnd11an1n32x5 FILLER_185_630 ();
 b15zdnd11an1n16x5 FILLER_185_662 ();
 b15zdnd11an1n04x5 FILLER_185_678 ();
 b15zdnd00an1n02x5 FILLER_185_682 ();
 b15zdnd00an1n01x5 FILLER_185_684 ();
 b15zdnd11an1n32x5 FILLER_185_691 ();
 b15zdnd11an1n16x5 FILLER_185_723 ();
 b15zdnd11an1n04x5 FILLER_185_739 ();
 b15zdnd00an1n02x5 FILLER_185_743 ();
 b15zdnd11an1n64x5 FILLER_185_749 ();
 b15zdnd11an1n32x5 FILLER_185_813 ();
 b15zdnd11an1n16x5 FILLER_185_845 ();
 b15zdnd00an1n01x5 FILLER_185_861 ();
 b15zdnd11an1n64x5 FILLER_185_866 ();
 b15zdnd11an1n32x5 FILLER_185_930 ();
 b15zdnd11an1n04x5 FILLER_185_962 ();
 b15zdnd00an1n02x5 FILLER_185_966 ();
 b15zdnd00an1n01x5 FILLER_185_968 ();
 b15zdnd11an1n32x5 FILLER_185_977 ();
 b15zdnd00an1n02x5 FILLER_185_1009 ();
 b15zdnd00an1n01x5 FILLER_185_1011 ();
 b15zdnd11an1n16x5 FILLER_185_1021 ();
 b15zdnd11an1n04x5 FILLER_185_1037 ();
 b15zdnd00an1n01x5 FILLER_185_1041 ();
 b15zdnd11an1n08x5 FILLER_185_1055 ();
 b15zdnd11an1n16x5 FILLER_185_1073 ();
 b15zdnd11an1n08x5 FILLER_185_1089 ();
 b15zdnd00an1n01x5 FILLER_185_1097 ();
 b15zdnd11an1n32x5 FILLER_185_1105 ();
 b15zdnd11an1n04x5 FILLER_185_1137 ();
 b15zdnd00an1n02x5 FILLER_185_1141 ();
 b15zdnd11an1n04x5 FILLER_185_1164 ();
 b15zdnd11an1n08x5 FILLER_185_1175 ();
 b15zdnd11an1n08x5 FILLER_185_1190 ();
 b15zdnd00an1n02x5 FILLER_185_1198 ();
 b15zdnd11an1n64x5 FILLER_185_1207 ();
 b15zdnd11an1n16x5 FILLER_185_1271 ();
 b15zdnd11an1n08x5 FILLER_185_1287 ();
 b15zdnd11an1n04x5 FILLER_185_1295 ();
 b15zdnd00an1n01x5 FILLER_185_1299 ();
 b15zdnd11an1n64x5 FILLER_185_1320 ();
 b15zdnd11an1n16x5 FILLER_185_1384 ();
 b15zdnd11an1n08x5 FILLER_185_1400 ();
 b15zdnd11an1n04x5 FILLER_185_1408 ();
 b15zdnd00an1n02x5 FILLER_185_1412 ();
 b15zdnd11an1n16x5 FILLER_185_1418 ();
 b15zdnd00an1n01x5 FILLER_185_1434 ();
 b15zdnd11an1n16x5 FILLER_185_1440 ();
 b15zdnd00an1n02x5 FILLER_185_1456 ();
 b15zdnd00an1n01x5 FILLER_185_1458 ();
 b15zdnd11an1n04x5 FILLER_185_1468 ();
 b15zdnd00an1n02x5 FILLER_185_1472 ();
 b15zdnd11an1n16x5 FILLER_185_1478 ();
 b15zdnd11an1n08x5 FILLER_185_1494 ();
 b15zdnd11an1n08x5 FILLER_185_1508 ();
 b15zdnd11an1n04x5 FILLER_185_1516 ();
 b15zdnd11an1n32x5 FILLER_185_1525 ();
 b15zdnd11an1n04x5 FILLER_185_1557 ();
 b15zdnd00an1n02x5 FILLER_185_1561 ();
 b15zdnd11an1n04x5 FILLER_185_1573 ();
 b15zdnd00an1n01x5 FILLER_185_1577 ();
 b15zdnd11an1n16x5 FILLER_185_1584 ();
 b15zdnd11an1n08x5 FILLER_185_1600 ();
 b15zdnd11an1n04x5 FILLER_185_1608 ();
 b15zdnd00an1n02x5 FILLER_185_1612 ();
 b15zdnd11an1n32x5 FILLER_185_1623 ();
 b15zdnd11an1n08x5 FILLER_185_1655 ();
 b15zdnd11an1n04x5 FILLER_185_1663 ();
 b15zdnd00an1n02x5 FILLER_185_1667 ();
 b15zdnd00an1n01x5 FILLER_185_1669 ();
 b15zdnd11an1n16x5 FILLER_185_1696 ();
 b15zdnd00an1n01x5 FILLER_185_1712 ();
 b15zdnd11an1n64x5 FILLER_185_1733 ();
 b15zdnd11an1n64x5 FILLER_185_1797 ();
 b15zdnd11an1n16x5 FILLER_185_1861 ();
 b15zdnd00an1n02x5 FILLER_185_1877 ();
 b15zdnd11an1n08x5 FILLER_185_1899 ();
 b15zdnd00an1n02x5 FILLER_185_1907 ();
 b15zdnd11an1n04x5 FILLER_185_1914 ();
 b15zdnd11an1n04x5 FILLER_185_1924 ();
 b15zdnd11an1n64x5 FILLER_185_1948 ();
 b15zdnd11an1n08x5 FILLER_185_2012 ();
 b15zdnd11an1n04x5 FILLER_185_2020 ();
 b15zdnd00an1n01x5 FILLER_185_2024 ();
 b15zdnd11an1n64x5 FILLER_185_2042 ();
 b15zdnd11an1n08x5 FILLER_185_2106 ();
 b15zdnd11an1n04x5 FILLER_185_2117 ();
 b15zdnd11an1n04x5 FILLER_185_2141 ();
 b15zdnd11an1n64x5 FILLER_185_2150 ();
 b15zdnd00an1n02x5 FILLER_185_2214 ();
 b15zdnd00an1n01x5 FILLER_185_2216 ();
 b15zdnd11an1n16x5 FILLER_185_2237 ();
 b15zdnd00an1n01x5 FILLER_185_2253 ();
 b15zdnd11an1n04x5 FILLER_185_2258 ();
 b15zdnd11an1n16x5 FILLER_185_2266 ();
 b15zdnd00an1n02x5 FILLER_185_2282 ();
 b15zdnd11an1n16x5 FILLER_186_8 ();
 b15zdnd11an1n08x5 FILLER_186_24 ();
 b15zdnd11an1n04x5 FILLER_186_32 ();
 b15zdnd00an1n02x5 FILLER_186_36 ();
 b15zdnd00an1n01x5 FILLER_186_38 ();
 b15zdnd11an1n04x5 FILLER_186_51 ();
 b15zdnd11an1n16x5 FILLER_186_67 ();
 b15zdnd11an1n08x5 FILLER_186_83 ();
 b15zdnd11an1n04x5 FILLER_186_91 ();
 b15zdnd00an1n01x5 FILLER_186_95 ();
 b15zdnd11an1n32x5 FILLER_186_106 ();
 b15zdnd11an1n08x5 FILLER_186_138 ();
 b15zdnd11an1n04x5 FILLER_186_146 ();
 b15zdnd00an1n01x5 FILLER_186_150 ();
 b15zdnd11an1n04x5 FILLER_186_156 ();
 b15zdnd11an1n04x5 FILLER_186_165 ();
 b15zdnd00an1n02x5 FILLER_186_169 ();
 b15zdnd11an1n04x5 FILLER_186_196 ();
 b15zdnd11an1n16x5 FILLER_186_210 ();
 b15zdnd11an1n04x5 FILLER_186_226 ();
 b15zdnd00an1n01x5 FILLER_186_230 ();
 b15zdnd11an1n08x5 FILLER_186_243 ();
 b15zdnd00an1n02x5 FILLER_186_251 ();
 b15zdnd11an1n04x5 FILLER_186_259 ();
 b15zdnd11an1n16x5 FILLER_186_273 ();
 b15zdnd11an1n04x5 FILLER_186_289 ();
 b15zdnd00an1n02x5 FILLER_186_293 ();
 b15zdnd11an1n16x5 FILLER_186_302 ();
 b15zdnd11an1n08x5 FILLER_186_318 ();
 b15zdnd11an1n04x5 FILLER_186_326 ();
 b15zdnd00an1n01x5 FILLER_186_330 ();
 b15zdnd11an1n64x5 FILLER_186_363 ();
 b15zdnd00an1n01x5 FILLER_186_427 ();
 b15zdnd11an1n64x5 FILLER_186_432 ();
 b15zdnd00an1n02x5 FILLER_186_496 ();
 b15zdnd11an1n04x5 FILLER_186_502 ();
 b15zdnd11an1n64x5 FILLER_186_516 ();
 b15zdnd11an1n32x5 FILLER_186_580 ();
 b15zdnd11an1n04x5 FILLER_186_612 ();
 b15zdnd00an1n01x5 FILLER_186_616 ();
 b15zdnd11an1n16x5 FILLER_186_629 ();
 b15zdnd11an1n04x5 FILLER_186_645 ();
 b15zdnd00an1n01x5 FILLER_186_649 ();
 b15zdnd11an1n32x5 FILLER_186_662 ();
 b15zdnd11an1n16x5 FILLER_186_694 ();
 b15zdnd11an1n08x5 FILLER_186_710 ();
 b15zdnd00an1n02x5 FILLER_186_726 ();
 b15zdnd00an1n01x5 FILLER_186_728 ();
 b15zdnd11an1n04x5 FILLER_186_757 ();
 b15zdnd11an1n08x5 FILLER_186_768 ();
 b15zdnd00an1n02x5 FILLER_186_776 ();
 b15zdnd00an1n01x5 FILLER_186_778 ();
 b15zdnd11an1n64x5 FILLER_186_794 ();
 b15zdnd11an1n64x5 FILLER_186_858 ();
 b15zdnd00an1n02x5 FILLER_186_922 ();
 b15zdnd00an1n01x5 FILLER_186_924 ();
 b15zdnd11an1n32x5 FILLER_186_937 ();
 b15zdnd11an1n16x5 FILLER_186_969 ();
 b15zdnd00an1n02x5 FILLER_186_985 ();
 b15zdnd11an1n32x5 FILLER_186_991 ();
 b15zdnd11an1n16x5 FILLER_186_1023 ();
 b15zdnd11an1n08x5 FILLER_186_1039 ();
 b15zdnd00an1n02x5 FILLER_186_1047 ();
 b15zdnd11an1n08x5 FILLER_186_1053 ();
 b15zdnd00an1n02x5 FILLER_186_1061 ();
 b15zdnd11an1n04x5 FILLER_186_1078 ();
 b15zdnd00an1n01x5 FILLER_186_1082 ();
 b15zdnd11an1n04x5 FILLER_186_1115 ();
 b15zdnd11an1n04x5 FILLER_186_1139 ();
 b15zdnd11an1n16x5 FILLER_186_1152 ();
 b15zdnd11an1n04x5 FILLER_186_1173 ();
 b15zdnd11an1n64x5 FILLER_186_1187 ();
 b15zdnd11an1n32x5 FILLER_186_1251 ();
 b15zdnd00an1n01x5 FILLER_186_1283 ();
 b15zdnd11an1n04x5 FILLER_186_1305 ();
 b15zdnd11an1n32x5 FILLER_186_1325 ();
 b15zdnd11an1n16x5 FILLER_186_1357 ();
 b15zdnd11an1n08x5 FILLER_186_1377 ();
 b15zdnd00an1n02x5 FILLER_186_1385 ();
 b15zdnd11an1n04x5 FILLER_186_1393 ();
 b15zdnd11an1n08x5 FILLER_186_1403 ();
 b15zdnd00an1n02x5 FILLER_186_1411 ();
 b15zdnd11an1n16x5 FILLER_186_1418 ();
 b15zdnd11an1n04x5 FILLER_186_1434 ();
 b15zdnd00an1n02x5 FILLER_186_1438 ();
 b15zdnd11an1n16x5 FILLER_186_1447 ();
 b15zdnd11an1n04x5 FILLER_186_1463 ();
 b15zdnd11an1n04x5 FILLER_186_1481 ();
 b15zdnd11an1n04x5 FILLER_186_1495 ();
 b15zdnd11an1n04x5 FILLER_186_1509 ();
 b15zdnd00an1n01x5 FILLER_186_1513 ();
 b15zdnd11an1n32x5 FILLER_186_1535 ();
 b15zdnd11an1n08x5 FILLER_186_1567 ();
 b15zdnd11an1n32x5 FILLER_186_1585 ();
 b15zdnd11an1n04x5 FILLER_186_1617 ();
 b15zdnd00an1n01x5 FILLER_186_1621 ();
 b15zdnd11an1n16x5 FILLER_186_1631 ();
 b15zdnd11an1n08x5 FILLER_186_1647 ();
 b15zdnd11an1n04x5 FILLER_186_1655 ();
 b15zdnd11an1n32x5 FILLER_186_1671 ();
 b15zdnd11an1n16x5 FILLER_186_1703 ();
 b15zdnd11an1n04x5 FILLER_186_1719 ();
 b15zdnd00an1n02x5 FILLER_186_1723 ();
 b15zdnd11an1n16x5 FILLER_186_1737 ();
 b15zdnd11an1n08x5 FILLER_186_1753 ();
 b15zdnd00an1n02x5 FILLER_186_1761 ();
 b15zdnd00an1n01x5 FILLER_186_1763 ();
 b15zdnd11an1n32x5 FILLER_186_1779 ();
 b15zdnd11an1n16x5 FILLER_186_1811 ();
 b15zdnd11an1n04x5 FILLER_186_1827 ();
 b15zdnd00an1n01x5 FILLER_186_1831 ();
 b15zdnd11an1n64x5 FILLER_186_1850 ();
 b15zdnd11an1n64x5 FILLER_186_1914 ();
 b15zdnd11an1n64x5 FILLER_186_1978 ();
 b15zdnd11an1n04x5 FILLER_186_2042 ();
 b15zdnd00an1n01x5 FILLER_186_2046 ();
 b15zdnd11an1n04x5 FILLER_186_2052 ();
 b15zdnd11an1n16x5 FILLER_186_2076 ();
 b15zdnd00an1n02x5 FILLER_186_2092 ();
 b15zdnd00an1n01x5 FILLER_186_2094 ();
 b15zdnd11an1n16x5 FILLER_186_2104 ();
 b15zdnd11an1n08x5 FILLER_186_2140 ();
 b15zdnd11an1n04x5 FILLER_186_2148 ();
 b15zdnd00an1n02x5 FILLER_186_2152 ();
 b15zdnd11an1n32x5 FILLER_186_2162 ();
 b15zdnd11an1n08x5 FILLER_186_2194 ();
 b15zdnd11an1n04x5 FILLER_186_2222 ();
 b15zdnd11an1n16x5 FILLER_186_2231 ();
 b15zdnd00an1n02x5 FILLER_186_2247 ();
 b15zdnd11an1n04x5 FILLER_186_2254 ();
 b15zdnd11an1n08x5 FILLER_186_2262 ();
 b15zdnd00an1n02x5 FILLER_186_2274 ();
 b15zdnd11an1n64x5 FILLER_187_0 ();
 b15zdnd11an1n16x5 FILLER_187_64 ();
 b15zdnd00an1n02x5 FILLER_187_80 ();
 b15zdnd11an1n04x5 FILLER_187_86 ();
 b15zdnd11an1n04x5 FILLER_187_95 ();
 b15zdnd11an1n32x5 FILLER_187_108 ();
 b15zdnd00an1n02x5 FILLER_187_140 ();
 b15zdnd11an1n08x5 FILLER_187_155 ();
 b15zdnd11an1n04x5 FILLER_187_163 ();
 b15zdnd00an1n01x5 FILLER_187_167 ();
 b15zdnd11an1n16x5 FILLER_187_174 ();
 b15zdnd00an1n01x5 FILLER_187_190 ();
 b15zdnd11an1n16x5 FILLER_187_202 ();
 b15zdnd11an1n08x5 FILLER_187_218 ();
 b15zdnd11an1n04x5 FILLER_187_226 ();
 b15zdnd00an1n02x5 FILLER_187_230 ();
 b15zdnd11an1n04x5 FILLER_187_243 ();
 b15zdnd11an1n16x5 FILLER_187_259 ();
 b15zdnd11an1n08x5 FILLER_187_275 ();
 b15zdnd00an1n02x5 FILLER_187_283 ();
 b15zdnd11an1n64x5 FILLER_187_296 ();
 b15zdnd11an1n32x5 FILLER_187_360 ();
 b15zdnd11an1n16x5 FILLER_187_392 ();
 b15zdnd11an1n64x5 FILLER_187_418 ();
 b15zdnd11an1n32x5 FILLER_187_482 ();
 b15zdnd00an1n02x5 FILLER_187_514 ();
 b15zdnd00an1n01x5 FILLER_187_516 ();
 b15zdnd11an1n16x5 FILLER_187_521 ();
 b15zdnd11an1n08x5 FILLER_187_537 ();
 b15zdnd11an1n04x5 FILLER_187_545 ();
 b15zdnd00an1n02x5 FILLER_187_549 ();
 b15zdnd11an1n64x5 FILLER_187_556 ();
 b15zdnd11an1n16x5 FILLER_187_620 ();
 b15zdnd11an1n08x5 FILLER_187_636 ();
 b15zdnd00an1n02x5 FILLER_187_644 ();
 b15zdnd11an1n04x5 FILLER_187_652 ();
 b15zdnd11an1n32x5 FILLER_187_664 ();
 b15zdnd11an1n16x5 FILLER_187_696 ();
 b15zdnd11an1n08x5 FILLER_187_712 ();
 b15zdnd00an1n02x5 FILLER_187_720 ();
 b15zdnd11an1n04x5 FILLER_187_753 ();
 b15zdnd00an1n01x5 FILLER_187_757 ();
 b15zdnd11an1n64x5 FILLER_187_764 ();
 b15zdnd11an1n32x5 FILLER_187_828 ();
 b15zdnd11an1n08x5 FILLER_187_860 ();
 b15zdnd11an1n08x5 FILLER_187_883 ();
 b15zdnd11an1n04x5 FILLER_187_901 ();
 b15zdnd00an1n02x5 FILLER_187_905 ();
 b15zdnd00an1n01x5 FILLER_187_907 ();
 b15zdnd11an1n08x5 FILLER_187_918 ();
 b15zdnd00an1n02x5 FILLER_187_926 ();
 b15zdnd00an1n01x5 FILLER_187_928 ();
 b15zdnd11an1n16x5 FILLER_187_934 ();
 b15zdnd11an1n04x5 FILLER_187_950 ();
 b15zdnd00an1n02x5 FILLER_187_954 ();
 b15zdnd00an1n01x5 FILLER_187_956 ();
 b15zdnd11an1n04x5 FILLER_187_969 ();
 b15zdnd11an1n08x5 FILLER_187_979 ();
 b15zdnd11an1n08x5 FILLER_187_993 ();
 b15zdnd11an1n04x5 FILLER_187_1001 ();
 b15zdnd00an1n02x5 FILLER_187_1005 ();
 b15zdnd00an1n01x5 FILLER_187_1007 ();
 b15zdnd11an1n64x5 FILLER_187_1018 ();
 b15zdnd11an1n32x5 FILLER_187_1082 ();
 b15zdnd11an1n16x5 FILLER_187_1114 ();
 b15zdnd11an1n08x5 FILLER_187_1130 ();
 b15zdnd11an1n04x5 FILLER_187_1138 ();
 b15zdnd11an1n32x5 FILLER_187_1162 ();
 b15zdnd11an1n04x5 FILLER_187_1194 ();
 b15zdnd00an1n02x5 FILLER_187_1198 ();
 b15zdnd11an1n64x5 FILLER_187_1210 ();
 b15zdnd11an1n32x5 FILLER_187_1274 ();
 b15zdnd11an1n16x5 FILLER_187_1306 ();
 b15zdnd11an1n04x5 FILLER_187_1322 ();
 b15zdnd11an1n04x5 FILLER_187_1331 ();
 b15zdnd11an1n16x5 FILLER_187_1344 ();
 b15zdnd11an1n08x5 FILLER_187_1360 ();
 b15zdnd11an1n04x5 FILLER_187_1368 ();
 b15zdnd11an1n04x5 FILLER_187_1381 ();
 b15zdnd11an1n16x5 FILLER_187_1395 ();
 b15zdnd11an1n04x5 FILLER_187_1411 ();
 b15zdnd11an1n16x5 FILLER_187_1420 ();
 b15zdnd11an1n08x5 FILLER_187_1436 ();
 b15zdnd11an1n08x5 FILLER_187_1450 ();
 b15zdnd11an1n04x5 FILLER_187_1458 ();
 b15zdnd00an1n02x5 FILLER_187_1462 ();
 b15zdnd11an1n32x5 FILLER_187_1475 ();
 b15zdnd11an1n08x5 FILLER_187_1507 ();
 b15zdnd11an1n04x5 FILLER_187_1515 ();
 b15zdnd00an1n01x5 FILLER_187_1519 ();
 b15zdnd11an1n08x5 FILLER_187_1525 ();
 b15zdnd11an1n04x5 FILLER_187_1533 ();
 b15zdnd11an1n04x5 FILLER_187_1543 ();
 b15zdnd00an1n01x5 FILLER_187_1547 ();
 b15zdnd11an1n32x5 FILLER_187_1555 ();
 b15zdnd11an1n16x5 FILLER_187_1601 ();
 b15zdnd11an1n08x5 FILLER_187_1617 ();
 b15zdnd00an1n02x5 FILLER_187_1625 ();
 b15zdnd00an1n01x5 FILLER_187_1627 ();
 b15zdnd11an1n16x5 FILLER_187_1632 ();
 b15zdnd11an1n08x5 FILLER_187_1648 ();
 b15zdnd00an1n01x5 FILLER_187_1656 ();
 b15zdnd11an1n04x5 FILLER_187_1673 ();
 b15zdnd11an1n64x5 FILLER_187_1686 ();
 b15zdnd11an1n04x5 FILLER_187_1750 ();
 b15zdnd00an1n02x5 FILLER_187_1754 ();
 b15zdnd00an1n01x5 FILLER_187_1756 ();
 b15zdnd11an1n64x5 FILLER_187_1782 ();
 b15zdnd00an1n01x5 FILLER_187_1846 ();
 b15zdnd11an1n64x5 FILLER_187_1872 ();
 b15zdnd11an1n32x5 FILLER_187_1936 ();
 b15zdnd11an1n08x5 FILLER_187_1968 ();
 b15zdnd00an1n02x5 FILLER_187_1976 ();
 b15zdnd00an1n01x5 FILLER_187_1978 ();
 b15zdnd11an1n16x5 FILLER_187_1990 ();
 b15zdnd11an1n04x5 FILLER_187_2006 ();
 b15zdnd00an1n02x5 FILLER_187_2010 ();
 b15zdnd00an1n01x5 FILLER_187_2012 ();
 b15zdnd11an1n08x5 FILLER_187_2016 ();
 b15zdnd11an1n04x5 FILLER_187_2035 ();
 b15zdnd00an1n02x5 FILLER_187_2039 ();
 b15zdnd00an1n01x5 FILLER_187_2041 ();
 b15zdnd11an1n64x5 FILLER_187_2046 ();
 b15zdnd11an1n64x5 FILLER_187_2110 ();
 b15zdnd11an1n64x5 FILLER_187_2174 ();
 b15zdnd11an1n16x5 FILLER_187_2238 ();
 b15zdnd00an1n02x5 FILLER_187_2254 ();
 b15zdnd11an1n04x5 FILLER_187_2261 ();
 b15zdnd11an1n04x5 FILLER_187_2269 ();
 b15zdnd00an1n02x5 FILLER_187_2273 ();
 b15zdnd00an1n01x5 FILLER_187_2275 ();
 b15zdnd11an1n04x5 FILLER_187_2280 ();
 b15zdnd00an1n02x5 FILLER_188_8 ();
 b15zdnd11an1n08x5 FILLER_188_14 ();
 b15zdnd00an1n02x5 FILLER_188_22 ();
 b15zdnd11an1n32x5 FILLER_188_32 ();
 b15zdnd11an1n04x5 FILLER_188_64 ();
 b15zdnd00an1n02x5 FILLER_188_68 ();
 b15zdnd11an1n16x5 FILLER_188_82 ();
 b15zdnd11an1n04x5 FILLER_188_104 ();
 b15zdnd11an1n08x5 FILLER_188_115 ();
 b15zdnd00an1n02x5 FILLER_188_123 ();
 b15zdnd00an1n01x5 FILLER_188_125 ();
 b15zdnd11an1n08x5 FILLER_188_130 ();
 b15zdnd11an1n16x5 FILLER_188_146 ();
 b15zdnd11an1n04x5 FILLER_188_162 ();
 b15zdnd00an1n01x5 FILLER_188_166 ();
 b15zdnd11an1n16x5 FILLER_188_171 ();
 b15zdnd00an1n02x5 FILLER_188_187 ();
 b15zdnd00an1n01x5 FILLER_188_189 ();
 b15zdnd11an1n64x5 FILLER_188_199 ();
 b15zdnd11an1n64x5 FILLER_188_263 ();
 b15zdnd11an1n32x5 FILLER_188_327 ();
 b15zdnd11an1n16x5 FILLER_188_359 ();
 b15zdnd11an1n04x5 FILLER_188_375 ();
 b15zdnd00an1n02x5 FILLER_188_379 ();
 b15zdnd00an1n01x5 FILLER_188_381 ();
 b15zdnd11an1n08x5 FILLER_188_395 ();
 b15zdnd00an1n01x5 FILLER_188_403 ();
 b15zdnd11an1n04x5 FILLER_188_409 ();
 b15zdnd00an1n02x5 FILLER_188_413 ();
 b15zdnd11an1n16x5 FILLER_188_431 ();
 b15zdnd11an1n04x5 FILLER_188_447 ();
 b15zdnd00an1n02x5 FILLER_188_451 ();
 b15zdnd00an1n01x5 FILLER_188_453 ();
 b15zdnd11an1n04x5 FILLER_188_467 ();
 b15zdnd11an1n64x5 FILLER_188_487 ();
 b15zdnd11an1n16x5 FILLER_188_551 ();
 b15zdnd11an1n08x5 FILLER_188_567 ();
 b15zdnd00an1n01x5 FILLER_188_575 ();
 b15zdnd11an1n32x5 FILLER_188_580 ();
 b15zdnd11an1n16x5 FILLER_188_612 ();
 b15zdnd11an1n08x5 FILLER_188_628 ();
 b15zdnd00an1n02x5 FILLER_188_636 ();
 b15zdnd11an1n04x5 FILLER_188_642 ();
 b15zdnd11an1n64x5 FILLER_188_652 ();
 b15zdnd00an1n02x5 FILLER_188_716 ();
 b15zdnd11an1n32x5 FILLER_188_726 ();
 b15zdnd11an1n04x5 FILLER_188_758 ();
 b15zdnd00an1n02x5 FILLER_188_762 ();
 b15zdnd00an1n01x5 FILLER_188_764 ();
 b15zdnd11an1n08x5 FILLER_188_769 ();
 b15zdnd11an1n04x5 FILLER_188_777 ();
 b15zdnd11an1n16x5 FILLER_188_807 ();
 b15zdnd11an1n08x5 FILLER_188_823 ();
 b15zdnd11an1n04x5 FILLER_188_831 ();
 b15zdnd00an1n02x5 FILLER_188_835 ();
 b15zdnd11an1n08x5 FILLER_188_845 ();
 b15zdnd00an1n02x5 FILLER_188_853 ();
 b15zdnd00an1n01x5 FILLER_188_855 ();
 b15zdnd11an1n04x5 FILLER_188_870 ();
 b15zdnd11an1n08x5 FILLER_188_879 ();
 b15zdnd11an1n04x5 FILLER_188_887 ();
 b15zdnd00an1n01x5 FILLER_188_891 ();
 b15zdnd11an1n08x5 FILLER_188_898 ();
 b15zdnd00an1n02x5 FILLER_188_906 ();
 b15zdnd11an1n04x5 FILLER_188_913 ();
 b15zdnd00an1n02x5 FILLER_188_917 ();
 b15zdnd00an1n01x5 FILLER_188_919 ();
 b15zdnd11an1n08x5 FILLER_188_925 ();
 b15zdnd00an1n02x5 FILLER_188_933 ();
 b15zdnd11an1n04x5 FILLER_188_939 ();
 b15zdnd00an1n01x5 FILLER_188_943 ();
 b15zdnd11an1n08x5 FILLER_188_949 ();
 b15zdnd11an1n04x5 FILLER_188_957 ();
 b15zdnd00an1n02x5 FILLER_188_961 ();
 b15zdnd00an1n01x5 FILLER_188_963 ();
 b15zdnd11an1n04x5 FILLER_188_971 ();
 b15zdnd11an1n32x5 FILLER_188_982 ();
 b15zdnd11an1n16x5 FILLER_188_1014 ();
 b15zdnd11an1n04x5 FILLER_188_1030 ();
 b15zdnd00an1n02x5 FILLER_188_1034 ();
 b15zdnd00an1n01x5 FILLER_188_1036 ();
 b15zdnd11an1n16x5 FILLER_188_1042 ();
 b15zdnd11an1n08x5 FILLER_188_1058 ();
 b15zdnd00an1n02x5 FILLER_188_1066 ();
 b15zdnd11an1n64x5 FILLER_188_1094 ();
 b15zdnd11an1n32x5 FILLER_188_1158 ();
 b15zdnd11an1n08x5 FILLER_188_1190 ();
 b15zdnd00an1n02x5 FILLER_188_1198 ();
 b15zdnd11an1n64x5 FILLER_188_1210 ();
 b15zdnd11an1n04x5 FILLER_188_1274 ();
 b15zdnd00an1n02x5 FILLER_188_1278 ();
 b15zdnd11an1n08x5 FILLER_188_1291 ();
 b15zdnd11an1n04x5 FILLER_188_1299 ();
 b15zdnd11an1n08x5 FILLER_188_1321 ();
 b15zdnd11an1n04x5 FILLER_188_1329 ();
 b15zdnd00an1n02x5 FILLER_188_1333 ();
 b15zdnd00an1n01x5 FILLER_188_1335 ();
 b15zdnd11an1n32x5 FILLER_188_1340 ();
 b15zdnd11an1n04x5 FILLER_188_1372 ();
 b15zdnd00an1n01x5 FILLER_188_1376 ();
 b15zdnd11an1n64x5 FILLER_188_1387 ();
 b15zdnd11an1n64x5 FILLER_188_1451 ();
 b15zdnd11an1n32x5 FILLER_188_1515 ();
 b15zdnd00an1n02x5 FILLER_188_1547 ();
 b15zdnd11an1n32x5 FILLER_188_1555 ();
 b15zdnd11an1n16x5 FILLER_188_1587 ();
 b15zdnd11an1n08x5 FILLER_188_1603 ();
 b15zdnd00an1n02x5 FILLER_188_1611 ();
 b15zdnd11an1n08x5 FILLER_188_1619 ();
 b15zdnd11an1n04x5 FILLER_188_1627 ();
 b15zdnd11an1n16x5 FILLER_188_1637 ();
 b15zdnd11an1n04x5 FILLER_188_1653 ();
 b15zdnd00an1n02x5 FILLER_188_1657 ();
 b15zdnd00an1n01x5 FILLER_188_1659 ();
 b15zdnd11an1n04x5 FILLER_188_1686 ();
 b15zdnd11an1n32x5 FILLER_188_1705 ();
 b15zdnd11an1n08x5 FILLER_188_1737 ();
 b15zdnd11an1n04x5 FILLER_188_1745 ();
 b15zdnd00an1n02x5 FILLER_188_1749 ();
 b15zdnd11an1n16x5 FILLER_188_1771 ();
 b15zdnd11an1n04x5 FILLER_188_1787 ();
 b15zdnd00an1n02x5 FILLER_188_1791 ();
 b15zdnd00an1n01x5 FILLER_188_1793 ();
 b15zdnd11an1n16x5 FILLER_188_1814 ();
 b15zdnd11an1n08x5 FILLER_188_1830 ();
 b15zdnd11an1n04x5 FILLER_188_1838 ();
 b15zdnd11an1n64x5 FILLER_188_1853 ();
 b15zdnd11an1n32x5 FILLER_188_1917 ();
 b15zdnd11an1n16x5 FILLER_188_1949 ();
 b15zdnd11an1n08x5 FILLER_188_1965 ();
 b15zdnd11an1n04x5 FILLER_188_1973 ();
 b15zdnd00an1n02x5 FILLER_188_1977 ();
 b15zdnd00an1n01x5 FILLER_188_1979 ();
 b15zdnd11an1n16x5 FILLER_188_2000 ();
 b15zdnd11an1n08x5 FILLER_188_2016 ();
 b15zdnd00an1n02x5 FILLER_188_2024 ();
 b15zdnd11an1n64x5 FILLER_188_2041 ();
 b15zdnd11an1n32x5 FILLER_188_2105 ();
 b15zdnd11an1n16x5 FILLER_188_2137 ();
 b15zdnd00an1n01x5 FILLER_188_2153 ();
 b15zdnd11an1n64x5 FILLER_188_2162 ();
 b15zdnd11an1n04x5 FILLER_188_2226 ();
 b15zdnd11an1n04x5 FILLER_188_2250 ();
 b15zdnd11an1n16x5 FILLER_188_2258 ();
 b15zdnd00an1n02x5 FILLER_188_2274 ();
 b15zdnd11an1n32x5 FILLER_189_0 ();
 b15zdnd11an1n08x5 FILLER_189_32 ();
 b15zdnd11an1n08x5 FILLER_189_47 ();
 b15zdnd11an1n04x5 FILLER_189_55 ();
 b15zdnd00an1n02x5 FILLER_189_59 ();
 b15zdnd11an1n32x5 FILLER_189_74 ();
 b15zdnd11an1n16x5 FILLER_189_106 ();
 b15zdnd11an1n08x5 FILLER_189_122 ();
 b15zdnd11an1n04x5 FILLER_189_130 ();
 b15zdnd00an1n01x5 FILLER_189_134 ();
 b15zdnd11an1n16x5 FILLER_189_144 ();
 b15zdnd11an1n04x5 FILLER_189_164 ();
 b15zdnd11an1n32x5 FILLER_189_174 ();
 b15zdnd11an1n16x5 FILLER_189_206 ();
 b15zdnd11an1n08x5 FILLER_189_222 ();
 b15zdnd00an1n02x5 FILLER_189_230 ();
 b15zdnd11an1n64x5 FILLER_189_237 ();
 b15zdnd11an1n64x5 FILLER_189_301 ();
 b15zdnd11an1n16x5 FILLER_189_365 ();
 b15zdnd00an1n01x5 FILLER_189_381 ();
 b15zdnd11an1n16x5 FILLER_189_399 ();
 b15zdnd00an1n01x5 FILLER_189_415 ();
 b15zdnd11an1n08x5 FILLER_189_428 ();
 b15zdnd11an1n04x5 FILLER_189_436 ();
 b15zdnd11an1n04x5 FILLER_189_447 ();
 b15zdnd00an1n01x5 FILLER_189_451 ();
 b15zdnd11an1n08x5 FILLER_189_462 ();
 b15zdnd00an1n01x5 FILLER_189_470 ();
 b15zdnd11an1n16x5 FILLER_189_480 ();
 b15zdnd11an1n08x5 FILLER_189_496 ();
 b15zdnd11an1n04x5 FILLER_189_504 ();
 b15zdnd00an1n02x5 FILLER_189_508 ();
 b15zdnd11an1n16x5 FILLER_189_528 ();
 b15zdnd11an1n04x5 FILLER_189_544 ();
 b15zdnd11an1n08x5 FILLER_189_561 ();
 b15zdnd11an1n04x5 FILLER_189_569 ();
 b15zdnd11an1n32x5 FILLER_189_579 ();
 b15zdnd11an1n08x5 FILLER_189_611 ();
 b15zdnd11an1n16x5 FILLER_189_625 ();
 b15zdnd11an1n08x5 FILLER_189_641 ();
 b15zdnd00an1n02x5 FILLER_189_649 ();
 b15zdnd11an1n04x5 FILLER_189_682 ();
 b15zdnd11an1n04x5 FILLER_189_692 ();
 b15zdnd11an1n32x5 FILLER_189_701 ();
 b15zdnd11an1n08x5 FILLER_189_733 ();
 b15zdnd11an1n04x5 FILLER_189_741 ();
 b15zdnd00an1n02x5 FILLER_189_745 ();
 b15zdnd11an1n64x5 FILLER_189_757 ();
 b15zdnd11an1n08x5 FILLER_189_821 ();
 b15zdnd11an1n04x5 FILLER_189_829 ();
 b15zdnd00an1n02x5 FILLER_189_833 ();
 b15zdnd11an1n08x5 FILLER_189_841 ();
 b15zdnd11an1n04x5 FILLER_189_849 ();
 b15zdnd11an1n16x5 FILLER_189_857 ();
 b15zdnd00an1n02x5 FILLER_189_873 ();
 b15zdnd00an1n01x5 FILLER_189_875 ();
 b15zdnd11an1n16x5 FILLER_189_882 ();
 b15zdnd11an1n64x5 FILLER_189_904 ();
 b15zdnd11an1n64x5 FILLER_189_968 ();
 b15zdnd11an1n04x5 FILLER_189_1032 ();
 b15zdnd00an1n02x5 FILLER_189_1036 ();
 b15zdnd00an1n01x5 FILLER_189_1038 ();
 b15zdnd11an1n04x5 FILLER_189_1045 ();
 b15zdnd11an1n16x5 FILLER_189_1054 ();
 b15zdnd00an1n01x5 FILLER_189_1070 ();
 b15zdnd11an1n04x5 FILLER_189_1085 ();
 b15zdnd11an1n32x5 FILLER_189_1095 ();
 b15zdnd11an1n04x5 FILLER_189_1127 ();
 b15zdnd00an1n02x5 FILLER_189_1131 ();
 b15zdnd11an1n32x5 FILLER_189_1139 ();
 b15zdnd11an1n08x5 FILLER_189_1171 ();
 b15zdnd11an1n04x5 FILLER_189_1179 ();
 b15zdnd00an1n02x5 FILLER_189_1183 ();
 b15zdnd00an1n01x5 FILLER_189_1185 ();
 b15zdnd11an1n64x5 FILLER_189_1192 ();
 b15zdnd11an1n08x5 FILLER_189_1256 ();
 b15zdnd11an1n04x5 FILLER_189_1264 ();
 b15zdnd11an1n16x5 FILLER_189_1282 ();
 b15zdnd11an1n04x5 FILLER_189_1298 ();
 b15zdnd00an1n02x5 FILLER_189_1302 ();
 b15zdnd11an1n08x5 FILLER_189_1313 ();
 b15zdnd11an1n04x5 FILLER_189_1321 ();
 b15zdnd00an1n01x5 FILLER_189_1325 ();
 b15zdnd11an1n16x5 FILLER_189_1342 ();
 b15zdnd11an1n08x5 FILLER_189_1358 ();
 b15zdnd11an1n04x5 FILLER_189_1366 ();
 b15zdnd00an1n02x5 FILLER_189_1370 ();
 b15zdnd00an1n01x5 FILLER_189_1372 ();
 b15zdnd11an1n64x5 FILLER_189_1380 ();
 b15zdnd11an1n64x5 FILLER_189_1444 ();
 b15zdnd11an1n64x5 FILLER_189_1508 ();
 b15zdnd11an1n16x5 FILLER_189_1572 ();
 b15zdnd11an1n08x5 FILLER_189_1588 ();
 b15zdnd11an1n04x5 FILLER_189_1606 ();
 b15zdnd00an1n02x5 FILLER_189_1610 ();
 b15zdnd11an1n04x5 FILLER_189_1624 ();
 b15zdnd00an1n02x5 FILLER_189_1628 ();
 b15zdnd00an1n01x5 FILLER_189_1630 ();
 b15zdnd11an1n32x5 FILLER_189_1637 ();
 b15zdnd00an1n02x5 FILLER_189_1669 ();
 b15zdnd11an1n08x5 FILLER_189_1676 ();
 b15zdnd00an1n02x5 FILLER_189_1684 ();
 b15zdnd00an1n01x5 FILLER_189_1686 ();
 b15zdnd11an1n04x5 FILLER_189_1694 ();
 b15zdnd11an1n16x5 FILLER_189_1705 ();
 b15zdnd11an1n04x5 FILLER_189_1721 ();
 b15zdnd00an1n02x5 FILLER_189_1725 ();
 b15zdnd11an1n16x5 FILLER_189_1742 ();
 b15zdnd11an1n08x5 FILLER_189_1758 ();
 b15zdnd11an1n16x5 FILLER_189_1775 ();
 b15zdnd11an1n04x5 FILLER_189_1791 ();
 b15zdnd00an1n02x5 FILLER_189_1795 ();
 b15zdnd11an1n04x5 FILLER_189_1802 ();
 b15zdnd11an1n64x5 FILLER_189_1809 ();
 b15zdnd11an1n04x5 FILLER_189_1873 ();
 b15zdnd11an1n64x5 FILLER_189_1881 ();
 b15zdnd11an1n64x5 FILLER_189_1945 ();
 b15zdnd11an1n64x5 FILLER_189_2009 ();
 b15zdnd11an1n64x5 FILLER_189_2073 ();
 b15zdnd11an1n64x5 FILLER_189_2137 ();
 b15zdnd11an1n16x5 FILLER_189_2201 ();
 b15zdnd11an1n08x5 FILLER_189_2217 ();
 b15zdnd11an1n04x5 FILLER_189_2225 ();
 b15zdnd00an1n01x5 FILLER_189_2229 ();
 b15zdnd11an1n16x5 FILLER_189_2234 ();
 b15zdnd11an1n04x5 FILLER_189_2250 ();
 b15zdnd11an1n08x5 FILLER_189_2262 ();
 b15zdnd11an1n04x5 FILLER_189_2270 ();
 b15zdnd00an1n02x5 FILLER_189_2274 ();
 b15zdnd11an1n04x5 FILLER_189_2280 ();
 b15zdnd00an1n02x5 FILLER_190_8 ();
 b15zdnd00an1n01x5 FILLER_190_10 ();
 b15zdnd11an1n08x5 FILLER_190_15 ();
 b15zdnd11an1n04x5 FILLER_190_23 ();
 b15zdnd00an1n02x5 FILLER_190_27 ();
 b15zdnd00an1n01x5 FILLER_190_29 ();
 b15zdnd11an1n64x5 FILLER_190_38 ();
 b15zdnd11an1n64x5 FILLER_190_102 ();
 b15zdnd11an1n16x5 FILLER_190_166 ();
 b15zdnd11an1n08x5 FILLER_190_182 ();
 b15zdnd00an1n01x5 FILLER_190_190 ();
 b15zdnd11an1n04x5 FILLER_190_210 ();
 b15zdnd11an1n04x5 FILLER_190_221 ();
 b15zdnd11an1n64x5 FILLER_190_233 ();
 b15zdnd11an1n04x5 FILLER_190_297 ();
 b15zdnd00an1n02x5 FILLER_190_301 ();
 b15zdnd00an1n01x5 FILLER_190_303 ();
 b15zdnd11an1n04x5 FILLER_190_308 ();
 b15zdnd00an1n01x5 FILLER_190_312 ();
 b15zdnd11an1n08x5 FILLER_190_319 ();
 b15zdnd00an1n02x5 FILLER_190_327 ();
 b15zdnd00an1n01x5 FILLER_190_329 ();
 b15zdnd11an1n32x5 FILLER_190_339 ();
 b15zdnd11an1n08x5 FILLER_190_371 ();
 b15zdnd00an1n02x5 FILLER_190_379 ();
 b15zdnd11an1n32x5 FILLER_190_387 ();
 b15zdnd11an1n16x5 FILLER_190_419 ();
 b15zdnd11an1n08x5 FILLER_190_435 ();
 b15zdnd11an1n08x5 FILLER_190_448 ();
 b15zdnd11an1n32x5 FILLER_190_476 ();
 b15zdnd11an1n08x5 FILLER_190_508 ();
 b15zdnd00an1n01x5 FILLER_190_516 ();
 b15zdnd11an1n64x5 FILLER_190_524 ();
 b15zdnd11an1n16x5 FILLER_190_594 ();
 b15zdnd11an1n32x5 FILLER_190_628 ();
 b15zdnd11an1n16x5 FILLER_190_660 ();
 b15zdnd11an1n08x5 FILLER_190_676 ();
 b15zdnd11an1n04x5 FILLER_190_684 ();
 b15zdnd11an1n16x5 FILLER_190_702 ();
 b15zdnd11an1n08x5 FILLER_190_726 ();
 b15zdnd11an1n64x5 FILLER_190_744 ();
 b15zdnd11an1n32x5 FILLER_190_808 ();
 b15zdnd11an1n16x5 FILLER_190_840 ();
 b15zdnd11an1n08x5 FILLER_190_856 ();
 b15zdnd11an1n04x5 FILLER_190_864 ();
 b15zdnd00an1n02x5 FILLER_190_868 ();
 b15zdnd00an1n01x5 FILLER_190_870 ();
 b15zdnd11an1n64x5 FILLER_190_886 ();
 b15zdnd11an1n32x5 FILLER_190_950 ();
 b15zdnd00an1n02x5 FILLER_190_982 ();
 b15zdnd11an1n64x5 FILLER_190_1005 ();
 b15zdnd11an1n64x5 FILLER_190_1069 ();
 b15zdnd11an1n04x5 FILLER_190_1133 ();
 b15zdnd11an1n16x5 FILLER_190_1146 ();
 b15zdnd11an1n04x5 FILLER_190_1162 ();
 b15zdnd00an1n02x5 FILLER_190_1166 ();
 b15zdnd00an1n01x5 FILLER_190_1168 ();
 b15zdnd11an1n04x5 FILLER_190_1179 ();
 b15zdnd11an1n08x5 FILLER_190_1188 ();
 b15zdnd00an1n02x5 FILLER_190_1196 ();
 b15zdnd00an1n01x5 FILLER_190_1198 ();
 b15zdnd11an1n04x5 FILLER_190_1207 ();
 b15zdnd11an1n32x5 FILLER_190_1218 ();
 b15zdnd11an1n16x5 FILLER_190_1250 ();
 b15zdnd11an1n08x5 FILLER_190_1266 ();
 b15zdnd11an1n04x5 FILLER_190_1274 ();
 b15zdnd00an1n01x5 FILLER_190_1278 ();
 b15zdnd11an1n16x5 FILLER_190_1283 ();
 b15zdnd11an1n04x5 FILLER_190_1299 ();
 b15zdnd00an1n01x5 FILLER_190_1303 ();
 b15zdnd11an1n64x5 FILLER_190_1308 ();
 b15zdnd11an1n08x5 FILLER_190_1372 ();
 b15zdnd11an1n04x5 FILLER_190_1380 ();
 b15zdnd00an1n01x5 FILLER_190_1384 ();
 b15zdnd11an1n32x5 FILLER_190_1393 ();
 b15zdnd00an1n01x5 FILLER_190_1425 ();
 b15zdnd11an1n16x5 FILLER_190_1432 ();
 b15zdnd11an1n08x5 FILLER_190_1448 ();
 b15zdnd00an1n02x5 FILLER_190_1456 ();
 b15zdnd11an1n04x5 FILLER_190_1465 ();
 b15zdnd11an1n64x5 FILLER_190_1474 ();
 b15zdnd11an1n64x5 FILLER_190_1538 ();
 b15zdnd11an1n32x5 FILLER_190_1602 ();
 b15zdnd00an1n01x5 FILLER_190_1634 ();
 b15zdnd11an1n16x5 FILLER_190_1644 ();
 b15zdnd11an1n08x5 FILLER_190_1660 ();
 b15zdnd00an1n02x5 FILLER_190_1668 ();
 b15zdnd11an1n08x5 FILLER_190_1676 ();
 b15zdnd11an1n04x5 FILLER_190_1684 ();
 b15zdnd00an1n01x5 FILLER_190_1688 ();
 b15zdnd11an1n08x5 FILLER_190_1715 ();
 b15zdnd11an1n04x5 FILLER_190_1723 ();
 b15zdnd00an1n02x5 FILLER_190_1727 ();
 b15zdnd00an1n01x5 FILLER_190_1729 ();
 b15zdnd11an1n16x5 FILLER_190_1748 ();
 b15zdnd00an1n01x5 FILLER_190_1764 ();
 b15zdnd11an1n64x5 FILLER_190_1776 ();
 b15zdnd11an1n16x5 FILLER_190_1840 ();
 b15zdnd11an1n08x5 FILLER_190_1856 ();
 b15zdnd00an1n02x5 FILLER_190_1864 ();
 b15zdnd11an1n64x5 FILLER_190_1871 ();
 b15zdnd11an1n32x5 FILLER_190_1935 ();
 b15zdnd11an1n08x5 FILLER_190_1967 ();
 b15zdnd11an1n04x5 FILLER_190_1975 ();
 b15zdnd00an1n02x5 FILLER_190_1979 ();
 b15zdnd11an1n32x5 FILLER_190_1993 ();
 b15zdnd11an1n16x5 FILLER_190_2025 ();
 b15zdnd11an1n08x5 FILLER_190_2041 ();
 b15zdnd00an1n01x5 FILLER_190_2049 ();
 b15zdnd11an1n64x5 FILLER_190_2055 ();
 b15zdnd11an1n32x5 FILLER_190_2119 ();
 b15zdnd00an1n02x5 FILLER_190_2151 ();
 b15zdnd00an1n01x5 FILLER_190_2153 ();
 b15zdnd00an1n02x5 FILLER_190_2162 ();
 b15zdnd11an1n16x5 FILLER_190_2170 ();
 b15zdnd11an1n08x5 FILLER_190_2186 ();
 b15zdnd11an1n04x5 FILLER_190_2194 ();
 b15zdnd00an1n01x5 FILLER_190_2198 ();
 b15zdnd11an1n32x5 FILLER_190_2219 ();
 b15zdnd00an1n01x5 FILLER_190_2251 ();
 b15zdnd11an1n04x5 FILLER_190_2256 ();
 b15zdnd11an1n04x5 FILLER_190_2264 ();
 b15zdnd11an1n04x5 FILLER_190_2272 ();
 b15zdnd11an1n16x5 FILLER_191_0 ();
 b15zdnd11an1n08x5 FILLER_191_16 ();
 b15zdnd11an1n04x5 FILLER_191_24 ();
 b15zdnd11an1n16x5 FILLER_191_44 ();
 b15zdnd11an1n08x5 FILLER_191_60 ();
 b15zdnd00an1n01x5 FILLER_191_68 ();
 b15zdnd11an1n04x5 FILLER_191_85 ();
 b15zdnd00an1n02x5 FILLER_191_89 ();
 b15zdnd11an1n16x5 FILLER_191_101 ();
 b15zdnd11an1n64x5 FILLER_191_123 ();
 b15zdnd11an1n16x5 FILLER_191_187 ();
 b15zdnd11an1n08x5 FILLER_191_203 ();
 b15zdnd11an1n04x5 FILLER_191_211 ();
 b15zdnd11an1n32x5 FILLER_191_226 ();
 b15zdnd11an1n16x5 FILLER_191_258 ();
 b15zdnd11an1n08x5 FILLER_191_274 ();
 b15zdnd11an1n04x5 FILLER_191_313 ();
 b15zdnd00an1n02x5 FILLER_191_317 ();
 b15zdnd11an1n04x5 FILLER_191_328 ();
 b15zdnd11an1n04x5 FILLER_191_348 ();
 b15zdnd11an1n64x5 FILLER_191_356 ();
 b15zdnd11an1n32x5 FILLER_191_420 ();
 b15zdnd11an1n04x5 FILLER_191_452 ();
 b15zdnd00an1n02x5 FILLER_191_456 ();
 b15zdnd11an1n04x5 FILLER_191_465 ();
 b15zdnd11an1n16x5 FILLER_191_475 ();
 b15zdnd11an1n08x5 FILLER_191_491 ();
 b15zdnd11an1n04x5 FILLER_191_499 ();
 b15zdnd00an1n02x5 FILLER_191_503 ();
 b15zdnd11an1n16x5 FILLER_191_518 ();
 b15zdnd11an1n08x5 FILLER_191_534 ();
 b15zdnd00an1n01x5 FILLER_191_542 ();
 b15zdnd11an1n32x5 FILLER_191_555 ();
 b15zdnd11an1n16x5 FILLER_191_587 ();
 b15zdnd11an1n08x5 FILLER_191_603 ();
 b15zdnd00an1n02x5 FILLER_191_611 ();
 b15zdnd00an1n01x5 FILLER_191_613 ();
 b15zdnd11an1n04x5 FILLER_191_618 ();
 b15zdnd11an1n08x5 FILLER_191_628 ();
 b15zdnd11an1n04x5 FILLER_191_636 ();
 b15zdnd00an1n01x5 FILLER_191_640 ();
 b15zdnd11an1n04x5 FILLER_191_647 ();
 b15zdnd11an1n32x5 FILLER_191_657 ();
 b15zdnd11an1n08x5 FILLER_191_689 ();
 b15zdnd00an1n02x5 FILLER_191_697 ();
 b15zdnd11an1n16x5 FILLER_191_713 ();
 b15zdnd11an1n08x5 FILLER_191_729 ();
 b15zdnd00an1n01x5 FILLER_191_737 ();
 b15zdnd11an1n64x5 FILLER_191_750 ();
 b15zdnd11an1n16x5 FILLER_191_814 ();
 b15zdnd11an1n08x5 FILLER_191_830 ();
 b15zdnd11an1n64x5 FILLER_191_843 ();
 b15zdnd11an1n32x5 FILLER_191_907 ();
 b15zdnd11an1n08x5 FILLER_191_939 ();
 b15zdnd00an1n02x5 FILLER_191_947 ();
 b15zdnd11an1n04x5 FILLER_191_959 ();
 b15zdnd11an1n16x5 FILLER_191_980 ();
 b15zdnd11an1n04x5 FILLER_191_996 ();
 b15zdnd00an1n02x5 FILLER_191_1000 ();
 b15zdnd11an1n04x5 FILLER_191_1014 ();
 b15zdnd11an1n64x5 FILLER_191_1022 ();
 b15zdnd11an1n16x5 FILLER_191_1086 ();
 b15zdnd11an1n08x5 FILLER_191_1102 ();
 b15zdnd11an1n04x5 FILLER_191_1110 ();
 b15zdnd00an1n02x5 FILLER_191_1114 ();
 b15zdnd11an1n04x5 FILLER_191_1134 ();
 b15zdnd11an1n64x5 FILLER_191_1143 ();
 b15zdnd11an1n64x5 FILLER_191_1207 ();
 b15zdnd11an1n08x5 FILLER_191_1271 ();
 b15zdnd11an1n04x5 FILLER_191_1279 ();
 b15zdnd00an1n02x5 FILLER_191_1283 ();
 b15zdnd11an1n04x5 FILLER_191_1289 ();
 b15zdnd00an1n02x5 FILLER_191_1293 ();
 b15zdnd00an1n01x5 FILLER_191_1295 ();
 b15zdnd11an1n16x5 FILLER_191_1304 ();
 b15zdnd11an1n04x5 FILLER_191_1320 ();
 b15zdnd00an1n02x5 FILLER_191_1324 ();
 b15zdnd11an1n32x5 FILLER_191_1340 ();
 b15zdnd11an1n04x5 FILLER_191_1372 ();
 b15zdnd00an1n01x5 FILLER_191_1376 ();
 b15zdnd11an1n04x5 FILLER_191_1381 ();
 b15zdnd11an1n16x5 FILLER_191_1391 ();
 b15zdnd11an1n08x5 FILLER_191_1407 ();
 b15zdnd11an1n04x5 FILLER_191_1415 ();
 b15zdnd00an1n01x5 FILLER_191_1419 ();
 b15zdnd11an1n04x5 FILLER_191_1433 ();
 b15zdnd11an1n08x5 FILLER_191_1444 ();
 b15zdnd11an1n04x5 FILLER_191_1452 ();
 b15zdnd00an1n01x5 FILLER_191_1456 ();
 b15zdnd11an1n04x5 FILLER_191_1461 ();
 b15zdnd11an1n16x5 FILLER_191_1475 ();
 b15zdnd11an1n04x5 FILLER_191_1491 ();
 b15zdnd00an1n01x5 FILLER_191_1495 ();
 b15zdnd11an1n04x5 FILLER_191_1508 ();
 b15zdnd11an1n08x5 FILLER_191_1528 ();
 b15zdnd00an1n02x5 FILLER_191_1536 ();
 b15zdnd11an1n04x5 FILLER_191_1544 ();
 b15zdnd11an1n64x5 FILLER_191_1557 ();
 b15zdnd11an1n16x5 FILLER_191_1621 ();
 b15zdnd11an1n08x5 FILLER_191_1637 ();
 b15zdnd11an1n04x5 FILLER_191_1665 ();
 b15zdnd11an1n08x5 FILLER_191_1674 ();
 b15zdnd00an1n02x5 FILLER_191_1682 ();
 b15zdnd00an1n01x5 FILLER_191_1684 ();
 b15zdnd11an1n64x5 FILLER_191_1711 ();
 b15zdnd11an1n16x5 FILLER_191_1775 ();
 b15zdnd11an1n08x5 FILLER_191_1791 ();
 b15zdnd11an1n32x5 FILLER_191_1825 ();
 b15zdnd11an1n08x5 FILLER_191_1857 ();
 b15zdnd00an1n02x5 FILLER_191_1865 ();
 b15zdnd11an1n32x5 FILLER_191_1887 ();
 b15zdnd11an1n08x5 FILLER_191_1919 ();
 b15zdnd00an1n02x5 FILLER_191_1927 ();
 b15zdnd11an1n32x5 FILLER_191_1948 ();
 b15zdnd11an1n08x5 FILLER_191_1980 ();
 b15zdnd00an1n01x5 FILLER_191_1988 ();
 b15zdnd11an1n04x5 FILLER_191_1998 ();
 b15zdnd00an1n01x5 FILLER_191_2002 ();
 b15zdnd11an1n16x5 FILLER_191_2023 ();
 b15zdnd11an1n04x5 FILLER_191_2039 ();
 b15zdnd11an1n04x5 FILLER_191_2063 ();
 b15zdnd11an1n32x5 FILLER_191_2086 ();
 b15zdnd11an1n16x5 FILLER_191_2138 ();
 b15zdnd11an1n08x5 FILLER_191_2174 ();
 b15zdnd11an1n04x5 FILLER_191_2182 ();
 b15zdnd00an1n02x5 FILLER_191_2186 ();
 b15zdnd11an1n16x5 FILLER_191_2208 ();
 b15zdnd11an1n04x5 FILLER_191_2224 ();
 b15zdnd00an1n02x5 FILLER_191_2228 ();
 b15zdnd11an1n04x5 FILLER_191_2250 ();
 b15zdnd11an1n16x5 FILLER_191_2258 ();
 b15zdnd00an1n02x5 FILLER_191_2274 ();
 b15zdnd00an1n01x5 FILLER_191_2276 ();
 b15zdnd00an1n02x5 FILLER_191_2281 ();
 b15zdnd00an1n01x5 FILLER_191_2283 ();
 b15zdnd11an1n32x5 FILLER_192_8 ();
 b15zdnd00an1n02x5 FILLER_192_40 ();
 b15zdnd11an1n08x5 FILLER_192_54 ();
 b15zdnd11an1n04x5 FILLER_192_62 ();
 b15zdnd11an1n16x5 FILLER_192_86 ();
 b15zdnd11an1n08x5 FILLER_192_102 ();
 b15zdnd00an1n02x5 FILLER_192_110 ();
 b15zdnd11an1n16x5 FILLER_192_118 ();
 b15zdnd11an1n04x5 FILLER_192_134 ();
 b15zdnd11an1n04x5 FILLER_192_147 ();
 b15zdnd00an1n01x5 FILLER_192_151 ();
 b15zdnd11an1n64x5 FILLER_192_162 ();
 b15zdnd11an1n04x5 FILLER_192_226 ();
 b15zdnd00an1n02x5 FILLER_192_230 ();
 b15zdnd11an1n08x5 FILLER_192_237 ();
 b15zdnd11an1n04x5 FILLER_192_245 ();
 b15zdnd00an1n01x5 FILLER_192_249 ();
 b15zdnd11an1n08x5 FILLER_192_268 ();
 b15zdnd00an1n01x5 FILLER_192_276 ();
 b15zdnd11an1n04x5 FILLER_192_308 ();
 b15zdnd11an1n64x5 FILLER_192_319 ();
 b15zdnd11an1n16x5 FILLER_192_383 ();
 b15zdnd11an1n64x5 FILLER_192_408 ();
 b15zdnd11an1n64x5 FILLER_192_472 ();
 b15zdnd11an1n64x5 FILLER_192_536 ();
 b15zdnd11an1n32x5 FILLER_192_600 ();
 b15zdnd11an1n16x5 FILLER_192_632 ();
 b15zdnd00an1n02x5 FILLER_192_648 ();
 b15zdnd00an1n01x5 FILLER_192_650 ();
 b15zdnd11an1n16x5 FILLER_192_657 ();
 b15zdnd11an1n08x5 FILLER_192_673 ();
 b15zdnd00an1n02x5 FILLER_192_681 ();
 b15zdnd00an1n01x5 FILLER_192_683 ();
 b15zdnd11an1n16x5 FILLER_192_689 ();
 b15zdnd11an1n08x5 FILLER_192_705 ();
 b15zdnd11an1n04x5 FILLER_192_713 ();
 b15zdnd00an1n01x5 FILLER_192_717 ();
 b15zdnd11an1n16x5 FILLER_192_726 ();
 b15zdnd00an1n01x5 FILLER_192_742 ();
 b15zdnd11an1n16x5 FILLER_192_771 ();
 b15zdnd11an1n08x5 FILLER_192_787 ();
 b15zdnd00an1n02x5 FILLER_192_795 ();
 b15zdnd11an1n16x5 FILLER_192_817 ();
 b15zdnd00an1n02x5 FILLER_192_833 ();
 b15zdnd11an1n64x5 FILLER_192_840 ();
 b15zdnd11an1n08x5 FILLER_192_904 ();
 b15zdnd00an1n01x5 FILLER_192_912 ();
 b15zdnd11an1n16x5 FILLER_192_921 ();
 b15zdnd11an1n08x5 FILLER_192_937 ();
 b15zdnd11an1n04x5 FILLER_192_945 ();
 b15zdnd00an1n02x5 FILLER_192_949 ();
 b15zdnd11an1n04x5 FILLER_192_963 ();
 b15zdnd00an1n01x5 FILLER_192_967 ();
 b15zdnd11an1n16x5 FILLER_192_974 ();
 b15zdnd11an1n08x5 FILLER_192_990 ();
 b15zdnd11an1n04x5 FILLER_192_998 ();
 b15zdnd11an1n04x5 FILLER_192_1020 ();
 b15zdnd11an1n08x5 FILLER_192_1036 ();
 b15zdnd11an1n04x5 FILLER_192_1049 ();
 b15zdnd11an1n04x5 FILLER_192_1059 ();
 b15zdnd11an1n08x5 FILLER_192_1067 ();
 b15zdnd00an1n02x5 FILLER_192_1075 ();
 b15zdnd11an1n04x5 FILLER_192_1081 ();
 b15zdnd11an1n08x5 FILLER_192_1092 ();
 b15zdnd11an1n04x5 FILLER_192_1100 ();
 b15zdnd00an1n01x5 FILLER_192_1104 ();
 b15zdnd11an1n04x5 FILLER_192_1110 ();
 b15zdnd11an1n08x5 FILLER_192_1126 ();
 b15zdnd11an1n16x5 FILLER_192_1146 ();
 b15zdnd11an1n08x5 FILLER_192_1162 ();
 b15zdnd11an1n04x5 FILLER_192_1170 ();
 b15zdnd00an1n02x5 FILLER_192_1174 ();
 b15zdnd11an1n16x5 FILLER_192_1184 ();
 b15zdnd11an1n08x5 FILLER_192_1200 ();
 b15zdnd11an1n04x5 FILLER_192_1208 ();
 b15zdnd11an1n64x5 FILLER_192_1220 ();
 b15zdnd11an1n08x5 FILLER_192_1284 ();
 b15zdnd11an1n04x5 FILLER_192_1292 ();
 b15zdnd00an1n01x5 FILLER_192_1296 ();
 b15zdnd11an1n04x5 FILLER_192_1301 ();
 b15zdnd11an1n16x5 FILLER_192_1310 ();
 b15zdnd00an1n02x5 FILLER_192_1326 ();
 b15zdnd00an1n01x5 FILLER_192_1328 ();
 b15zdnd11an1n64x5 FILLER_192_1335 ();
 b15zdnd11an1n16x5 FILLER_192_1399 ();
 b15zdnd11an1n08x5 FILLER_192_1415 ();
 b15zdnd11an1n04x5 FILLER_192_1423 ();
 b15zdnd00an1n01x5 FILLER_192_1427 ();
 b15zdnd11an1n64x5 FILLER_192_1434 ();
 b15zdnd11an1n04x5 FILLER_192_1498 ();
 b15zdnd00an1n01x5 FILLER_192_1502 ();
 b15zdnd11an1n04x5 FILLER_192_1510 ();
 b15zdnd00an1n02x5 FILLER_192_1514 ();
 b15zdnd00an1n01x5 FILLER_192_1516 ();
 b15zdnd11an1n16x5 FILLER_192_1529 ();
 b15zdnd11an1n08x5 FILLER_192_1545 ();
 b15zdnd11an1n04x5 FILLER_192_1553 ();
 b15zdnd11an1n04x5 FILLER_192_1577 ();
 b15zdnd11an1n08x5 FILLER_192_1590 ();
 b15zdnd11an1n04x5 FILLER_192_1598 ();
 b15zdnd00an1n01x5 FILLER_192_1602 ();
 b15zdnd11an1n04x5 FILLER_192_1607 ();
 b15zdnd11an1n08x5 FILLER_192_1621 ();
 b15zdnd11an1n04x5 FILLER_192_1629 ();
 b15zdnd11an1n64x5 FILLER_192_1642 ();
 b15zdnd11an1n64x5 FILLER_192_1706 ();
 b15zdnd11an1n32x5 FILLER_192_1770 ();
 b15zdnd11an1n16x5 FILLER_192_1802 ();
 b15zdnd11an1n04x5 FILLER_192_1818 ();
 b15zdnd00an1n01x5 FILLER_192_1822 ();
 b15zdnd11an1n08x5 FILLER_192_1829 ();
 b15zdnd11an1n04x5 FILLER_192_1837 ();
 b15zdnd11an1n16x5 FILLER_192_1861 ();
 b15zdnd00an1n02x5 FILLER_192_1877 ();
 b15zdnd11an1n32x5 FILLER_192_1882 ();
 b15zdnd11an1n16x5 FILLER_192_1919 ();
 b15zdnd00an1n02x5 FILLER_192_1935 ();
 b15zdnd00an1n01x5 FILLER_192_1937 ();
 b15zdnd11an1n64x5 FILLER_192_1969 ();
 b15zdnd11an1n32x5 FILLER_192_2033 ();
 b15zdnd11an1n16x5 FILLER_192_2065 ();
 b15zdnd11an1n04x5 FILLER_192_2081 ();
 b15zdnd00an1n02x5 FILLER_192_2085 ();
 b15zdnd00an1n01x5 FILLER_192_2087 ();
 b15zdnd11an1n16x5 FILLER_192_2097 ();
 b15zdnd11an1n04x5 FILLER_192_2113 ();
 b15zdnd00an1n02x5 FILLER_192_2117 ();
 b15zdnd11an1n04x5 FILLER_192_2123 ();
 b15zdnd11an1n16x5 FILLER_192_2133 ();
 b15zdnd11an1n04x5 FILLER_192_2149 ();
 b15zdnd00an1n01x5 FILLER_192_2153 ();
 b15zdnd00an1n02x5 FILLER_192_2162 ();
 b15zdnd11an1n16x5 FILLER_192_2169 ();
 b15zdnd11an1n08x5 FILLER_192_2185 ();
 b15zdnd00an1n02x5 FILLER_192_2193 ();
 b15zdnd11an1n32x5 FILLER_192_2200 ();
 b15zdnd11an1n16x5 FILLER_192_2232 ();
 b15zdnd11an1n04x5 FILLER_192_2248 ();
 b15zdnd00an1n01x5 FILLER_192_2252 ();
 b15zdnd11an1n08x5 FILLER_192_2257 ();
 b15zdnd11an1n04x5 FILLER_192_2265 ();
 b15zdnd00an1n01x5 FILLER_192_2269 ();
 b15zdnd00an1n02x5 FILLER_192_2274 ();
 b15zdnd11an1n64x5 FILLER_193_0 ();
 b15zdnd11an1n16x5 FILLER_193_64 ();
 b15zdnd11an1n04x5 FILLER_193_80 ();
 b15zdnd00an1n01x5 FILLER_193_84 ();
 b15zdnd11an1n08x5 FILLER_193_101 ();
 b15zdnd00an1n01x5 FILLER_193_109 ();
 b15zdnd11an1n08x5 FILLER_193_122 ();
 b15zdnd11an1n04x5 FILLER_193_135 ();
 b15zdnd11an1n16x5 FILLER_193_160 ();
 b15zdnd11an1n04x5 FILLER_193_176 ();
 b15zdnd11an1n64x5 FILLER_193_187 ();
 b15zdnd11an1n64x5 FILLER_193_251 ();
 b15zdnd11an1n16x5 FILLER_193_315 ();
 b15zdnd11an1n08x5 FILLER_193_331 ();
 b15zdnd00an1n02x5 FILLER_193_339 ();
 b15zdnd00an1n01x5 FILLER_193_341 ();
 b15zdnd11an1n64x5 FILLER_193_354 ();
 b15zdnd11an1n08x5 FILLER_193_418 ();
 b15zdnd00an1n01x5 FILLER_193_426 ();
 b15zdnd11an1n32x5 FILLER_193_431 ();
 b15zdnd11an1n08x5 FILLER_193_463 ();
 b15zdnd11an1n04x5 FILLER_193_471 ();
 b15zdnd00an1n02x5 FILLER_193_475 ();
 b15zdnd00an1n01x5 FILLER_193_477 ();
 b15zdnd11an1n32x5 FILLER_193_491 ();
 b15zdnd11an1n16x5 FILLER_193_523 ();
 b15zdnd11an1n04x5 FILLER_193_539 ();
 b15zdnd00an1n02x5 FILLER_193_543 ();
 b15zdnd00an1n01x5 FILLER_193_545 ();
 b15zdnd11an1n08x5 FILLER_193_553 ();
 b15zdnd11an1n04x5 FILLER_193_561 ();
 b15zdnd00an1n02x5 FILLER_193_565 ();
 b15zdnd00an1n01x5 FILLER_193_567 ();
 b15zdnd11an1n64x5 FILLER_193_579 ();
 b15zdnd11an1n08x5 FILLER_193_643 ();
 b15zdnd00an1n01x5 FILLER_193_651 ();
 b15zdnd11an1n16x5 FILLER_193_659 ();
 b15zdnd11an1n08x5 FILLER_193_675 ();
 b15zdnd00an1n01x5 FILLER_193_683 ();
 b15zdnd11an1n64x5 FILLER_193_690 ();
 b15zdnd11an1n64x5 FILLER_193_754 ();
 b15zdnd11an1n08x5 FILLER_193_818 ();
 b15zdnd00an1n02x5 FILLER_193_826 ();
 b15zdnd00an1n01x5 FILLER_193_828 ();
 b15zdnd11an1n04x5 FILLER_193_833 ();
 b15zdnd11an1n08x5 FILLER_193_846 ();
 b15zdnd11an1n08x5 FILLER_193_862 ();
 b15zdnd11an1n04x5 FILLER_193_878 ();
 b15zdnd11an1n32x5 FILLER_193_890 ();
 b15zdnd00an1n01x5 FILLER_193_922 ();
 b15zdnd11an1n64x5 FILLER_193_929 ();
 b15zdnd11an1n04x5 FILLER_193_993 ();
 b15zdnd00an1n02x5 FILLER_193_997 ();
 b15zdnd00an1n01x5 FILLER_193_999 ();
 b15zdnd11an1n16x5 FILLER_193_1006 ();
 b15zdnd11an1n08x5 FILLER_193_1022 ();
 b15zdnd00an1n02x5 FILLER_193_1030 ();
 b15zdnd00an1n01x5 FILLER_193_1032 ();
 b15zdnd11an1n04x5 FILLER_193_1053 ();
 b15zdnd11an1n04x5 FILLER_193_1070 ();
 b15zdnd11an1n04x5 FILLER_193_1088 ();
 b15zdnd11an1n16x5 FILLER_193_1101 ();
 b15zdnd11an1n04x5 FILLER_193_1117 ();
 b15zdnd00an1n02x5 FILLER_193_1121 ();
 b15zdnd00an1n01x5 FILLER_193_1123 ();
 b15zdnd11an1n32x5 FILLER_193_1128 ();
 b15zdnd11an1n16x5 FILLER_193_1160 ();
 b15zdnd11an1n04x5 FILLER_193_1176 ();
 b15zdnd00an1n02x5 FILLER_193_1180 ();
 b15zdnd11an1n04x5 FILLER_193_1207 ();
 b15zdnd11an1n64x5 FILLER_193_1222 ();
 b15zdnd11an1n64x5 FILLER_193_1286 ();
 b15zdnd11an1n08x5 FILLER_193_1350 ();
 b15zdnd11an1n04x5 FILLER_193_1358 ();
 b15zdnd11an1n32x5 FILLER_193_1368 ();
 b15zdnd00an1n02x5 FILLER_193_1400 ();
 b15zdnd11an1n16x5 FILLER_193_1408 ();
 b15zdnd11an1n08x5 FILLER_193_1424 ();
 b15zdnd11an1n04x5 FILLER_193_1432 ();
 b15zdnd00an1n02x5 FILLER_193_1436 ();
 b15zdnd11an1n16x5 FILLER_193_1452 ();
 b15zdnd11an1n04x5 FILLER_193_1468 ();
 b15zdnd11an1n08x5 FILLER_193_1483 ();
 b15zdnd00an1n02x5 FILLER_193_1491 ();
 b15zdnd00an1n01x5 FILLER_193_1493 ();
 b15zdnd11an1n16x5 FILLER_193_1501 ();
 b15zdnd11an1n04x5 FILLER_193_1523 ();
 b15zdnd11an1n04x5 FILLER_193_1532 ();
 b15zdnd11an1n04x5 FILLER_193_1542 ();
 b15zdnd00an1n02x5 FILLER_193_1546 ();
 b15zdnd11an1n32x5 FILLER_193_1560 ();
 b15zdnd11an1n08x5 FILLER_193_1592 ();
 b15zdnd11an1n04x5 FILLER_193_1600 ();
 b15zdnd00an1n02x5 FILLER_193_1604 ();
 b15zdnd11an1n08x5 FILLER_193_1614 ();
 b15zdnd00an1n02x5 FILLER_193_1622 ();
 b15zdnd11an1n04x5 FILLER_193_1629 ();
 b15zdnd11an1n08x5 FILLER_193_1644 ();
 b15zdnd00an1n02x5 FILLER_193_1652 ();
 b15zdnd00an1n01x5 FILLER_193_1654 ();
 b15zdnd11an1n04x5 FILLER_193_1668 ();
 b15zdnd11an1n32x5 FILLER_193_1677 ();
 b15zdnd11an1n08x5 FILLER_193_1709 ();
 b15zdnd11an1n04x5 FILLER_193_1717 ();
 b15zdnd11an1n32x5 FILLER_193_1745 ();
 b15zdnd11an1n08x5 FILLER_193_1777 ();
 b15zdnd11an1n04x5 FILLER_193_1785 ();
 b15zdnd00an1n01x5 FILLER_193_1789 ();
 b15zdnd11an1n16x5 FILLER_193_1800 ();
 b15zdnd11an1n08x5 FILLER_193_1816 ();
 b15zdnd00an1n01x5 FILLER_193_1824 ();
 b15zdnd11an1n64x5 FILLER_193_1840 ();
 b15zdnd11an1n08x5 FILLER_193_1904 ();
 b15zdnd00an1n02x5 FILLER_193_1912 ();
 b15zdnd00an1n01x5 FILLER_193_1914 ();
 b15zdnd11an1n64x5 FILLER_193_1935 ();
 b15zdnd11an1n32x5 FILLER_193_1999 ();
 b15zdnd11an1n16x5 FILLER_193_2031 ();
 b15zdnd11an1n32x5 FILLER_193_2056 ();
 b15zdnd00an1n02x5 FILLER_193_2088 ();
 b15zdnd11an1n16x5 FILLER_193_2099 ();
 b15zdnd11an1n08x5 FILLER_193_2115 ();
 b15zdnd00an1n02x5 FILLER_193_2123 ();
 b15zdnd11an1n32x5 FILLER_193_2130 ();
 b15zdnd11an1n16x5 FILLER_193_2162 ();
 b15zdnd11an1n08x5 FILLER_193_2178 ();
 b15zdnd11an1n04x5 FILLER_193_2186 ();
 b15zdnd00an1n01x5 FILLER_193_2190 ();
 b15zdnd11an1n16x5 FILLER_193_2197 ();
 b15zdnd00an1n02x5 FILLER_193_2213 ();
 b15zdnd11an1n04x5 FILLER_193_2220 ();
 b15zdnd11an1n04x5 FILLER_193_2228 ();
 b15zdnd11an1n16x5 FILLER_193_2236 ();
 b15zdnd11an1n08x5 FILLER_193_2252 ();
 b15zdnd11an1n04x5 FILLER_193_2260 ();
 b15zdnd00an1n02x5 FILLER_193_2264 ();
 b15zdnd11an1n04x5 FILLER_193_2269 ();
 b15zdnd00an1n02x5 FILLER_193_2273 ();
 b15zdnd00an1n01x5 FILLER_193_2275 ();
 b15zdnd00an1n02x5 FILLER_193_2281 ();
 b15zdnd00an1n01x5 FILLER_193_2283 ();
 b15zdnd11an1n04x5 FILLER_194_8 ();
 b15zdnd00an1n02x5 FILLER_194_12 ();
 b15zdnd11an1n04x5 FILLER_194_19 ();
 b15zdnd11an1n04x5 FILLER_194_31 ();
 b15zdnd11an1n64x5 FILLER_194_42 ();
 b15zdnd11an1n04x5 FILLER_194_106 ();
 b15zdnd11an1n32x5 FILLER_194_114 ();
 b15zdnd11an1n16x5 FILLER_194_146 ();
 b15zdnd11an1n04x5 FILLER_194_162 ();
 b15zdnd00an1n01x5 FILLER_194_166 ();
 b15zdnd11an1n04x5 FILLER_194_173 ();
 b15zdnd11an1n32x5 FILLER_194_188 ();
 b15zdnd11an1n04x5 FILLER_194_220 ();
 b15zdnd11an1n64x5 FILLER_194_235 ();
 b15zdnd11an1n32x5 FILLER_194_299 ();
 b15zdnd11an1n08x5 FILLER_194_331 ();
 b15zdnd00an1n02x5 FILLER_194_339 ();
 b15zdnd00an1n01x5 FILLER_194_341 ();
 b15zdnd11an1n16x5 FILLER_194_366 ();
 b15zdnd11an1n04x5 FILLER_194_391 ();
 b15zdnd00an1n02x5 FILLER_194_395 ();
 b15zdnd11an1n08x5 FILLER_194_410 ();
 b15zdnd11an1n32x5 FILLER_194_424 ();
 b15zdnd11an1n08x5 FILLER_194_456 ();
 b15zdnd11an1n04x5 FILLER_194_464 ();
 b15zdnd11an1n04x5 FILLER_194_475 ();
 b15zdnd11an1n04x5 FILLER_194_485 ();
 b15zdnd00an1n01x5 FILLER_194_489 ();
 b15zdnd11an1n04x5 FILLER_194_510 ();
 b15zdnd11an1n16x5 FILLER_194_521 ();
 b15zdnd11an1n08x5 FILLER_194_537 ();
 b15zdnd00an1n01x5 FILLER_194_545 ();
 b15zdnd11an1n04x5 FILLER_194_552 ();
 b15zdnd11an1n04x5 FILLER_194_562 ();
 b15zdnd00an1n02x5 FILLER_194_566 ();
 b15zdnd00an1n01x5 FILLER_194_568 ();
 b15zdnd11an1n04x5 FILLER_194_576 ();
 b15zdnd11an1n64x5 FILLER_194_592 ();
 b15zdnd11an1n16x5 FILLER_194_656 ();
 b15zdnd11an1n08x5 FILLER_194_672 ();
 b15zdnd11an1n04x5 FILLER_194_680 ();
 b15zdnd00an1n02x5 FILLER_194_684 ();
 b15zdnd11an1n16x5 FILLER_194_698 ();
 b15zdnd11an1n04x5 FILLER_194_714 ();
 b15zdnd11an1n64x5 FILLER_194_726 ();
 b15zdnd11an1n32x5 FILLER_194_790 ();
 b15zdnd11an1n08x5 FILLER_194_822 ();
 b15zdnd11an1n04x5 FILLER_194_830 ();
 b15zdnd00an1n02x5 FILLER_194_834 ();
 b15zdnd00an1n01x5 FILLER_194_836 ();
 b15zdnd11an1n16x5 FILLER_194_849 ();
 b15zdnd00an1n02x5 FILLER_194_865 ();
 b15zdnd11an1n08x5 FILLER_194_871 ();
 b15zdnd00an1n01x5 FILLER_194_879 ();
 b15zdnd11an1n08x5 FILLER_194_886 ();
 b15zdnd11an1n04x5 FILLER_194_894 ();
 b15zdnd00an1n01x5 FILLER_194_898 ();
 b15zdnd11an1n16x5 FILLER_194_908 ();
 b15zdnd00an1n02x5 FILLER_194_924 ();
 b15zdnd00an1n01x5 FILLER_194_926 ();
 b15zdnd11an1n16x5 FILLER_194_936 ();
 b15zdnd11an1n08x5 FILLER_194_952 ();
 b15zdnd11an1n04x5 FILLER_194_960 ();
 b15zdnd00an1n01x5 FILLER_194_964 ();
 b15zdnd11an1n64x5 FILLER_194_972 ();
 b15zdnd11an1n64x5 FILLER_194_1036 ();
 b15zdnd11an1n64x5 FILLER_194_1100 ();
 b15zdnd11an1n16x5 FILLER_194_1164 ();
 b15zdnd11an1n08x5 FILLER_194_1180 ();
 b15zdnd11an1n04x5 FILLER_194_1188 ();
 b15zdnd11an1n04x5 FILLER_194_1203 ();
 b15zdnd11an1n64x5 FILLER_194_1219 ();
 b15zdnd11an1n16x5 FILLER_194_1283 ();
 b15zdnd11an1n08x5 FILLER_194_1299 ();
 b15zdnd00an1n02x5 FILLER_194_1307 ();
 b15zdnd00an1n01x5 FILLER_194_1309 ();
 b15zdnd11an1n16x5 FILLER_194_1315 ();
 b15zdnd11an1n04x5 FILLER_194_1331 ();
 b15zdnd00an1n02x5 FILLER_194_1335 ();
 b15zdnd11an1n04x5 FILLER_194_1343 ();
 b15zdnd11an1n08x5 FILLER_194_1353 ();
 b15zdnd00an1n02x5 FILLER_194_1361 ();
 b15zdnd11an1n16x5 FILLER_194_1373 ();
 b15zdnd11an1n04x5 FILLER_194_1389 ();
 b15zdnd00an1n01x5 FILLER_194_1393 ();
 b15zdnd11an1n64x5 FILLER_194_1398 ();
 b15zdnd11an1n64x5 FILLER_194_1462 ();
 b15zdnd11an1n32x5 FILLER_194_1526 ();
 b15zdnd11an1n16x5 FILLER_194_1558 ();
 b15zdnd11an1n08x5 FILLER_194_1574 ();
 b15zdnd00an1n02x5 FILLER_194_1582 ();
 b15zdnd00an1n01x5 FILLER_194_1584 ();
 b15zdnd11an1n64x5 FILLER_194_1590 ();
 b15zdnd11an1n08x5 FILLER_194_1654 ();
 b15zdnd11an1n64x5 FILLER_194_1681 ();
 b15zdnd11an1n32x5 FILLER_194_1745 ();
 b15zdnd11an1n08x5 FILLER_194_1777 ();
 b15zdnd11an1n04x5 FILLER_194_1785 ();
 b15zdnd00an1n01x5 FILLER_194_1789 ();
 b15zdnd11an1n64x5 FILLER_194_1805 ();
 b15zdnd11an1n64x5 FILLER_194_1869 ();
 b15zdnd11an1n32x5 FILLER_194_1933 ();
 b15zdnd11an1n04x5 FILLER_194_1965 ();
 b15zdnd00an1n01x5 FILLER_194_1969 ();
 b15zdnd11an1n64x5 FILLER_194_1981 ();
 b15zdnd11an1n32x5 FILLER_194_2045 ();
 b15zdnd11an1n16x5 FILLER_194_2077 ();
 b15zdnd00an1n01x5 FILLER_194_2093 ();
 b15zdnd11an1n32x5 FILLER_194_2106 ();
 b15zdnd11an1n16x5 FILLER_194_2138 ();
 b15zdnd11an1n32x5 FILLER_194_2162 ();
 b15zdnd11an1n16x5 FILLER_194_2194 ();
 b15zdnd11an1n16x5 FILLER_194_2219 ();
 b15zdnd11an1n08x5 FILLER_194_2235 ();
 b15zdnd11an1n04x5 FILLER_194_2243 ();
 b15zdnd00an1n02x5 FILLER_194_2247 ();
 b15zdnd11an1n16x5 FILLER_194_2257 ();
 b15zdnd00an1n02x5 FILLER_194_2273 ();
 b15zdnd00an1n01x5 FILLER_194_2275 ();
 b15zdnd11an1n16x5 FILLER_195_0 ();
 b15zdnd11an1n08x5 FILLER_195_16 ();
 b15zdnd11an1n04x5 FILLER_195_24 ();
 b15zdnd00an1n02x5 FILLER_195_28 ();
 b15zdnd00an1n01x5 FILLER_195_30 ();
 b15zdnd11an1n04x5 FILLER_195_35 ();
 b15zdnd11an1n08x5 FILLER_195_50 ();
 b15zdnd11an1n04x5 FILLER_195_58 ();
 b15zdnd11an1n64x5 FILLER_195_80 ();
 b15zdnd11an1n64x5 FILLER_195_144 ();
 b15zdnd11an1n16x5 FILLER_195_208 ();
 b15zdnd11an1n08x5 FILLER_195_224 ();
 b15zdnd11an1n04x5 FILLER_195_232 ();
 b15zdnd11an1n32x5 FILLER_195_262 ();
 b15zdnd11an1n04x5 FILLER_195_294 ();
 b15zdnd00an1n02x5 FILLER_195_298 ();
 b15zdnd00an1n01x5 FILLER_195_300 ();
 b15zdnd11an1n04x5 FILLER_195_306 ();
 b15zdnd11an1n64x5 FILLER_195_336 ();
 b15zdnd11an1n16x5 FILLER_195_400 ();
 b15zdnd11an1n04x5 FILLER_195_416 ();
 b15zdnd00an1n02x5 FILLER_195_420 ();
 b15zdnd11an1n16x5 FILLER_195_428 ();
 b15zdnd11an1n08x5 FILLER_195_455 ();
 b15zdnd11an1n04x5 FILLER_195_463 ();
 b15zdnd00an1n01x5 FILLER_195_467 ();
 b15zdnd11an1n16x5 FILLER_195_479 ();
 b15zdnd11an1n08x5 FILLER_195_495 ();
 b15zdnd11an1n04x5 FILLER_195_503 ();
 b15zdnd11an1n16x5 FILLER_195_520 ();
 b15zdnd11an1n08x5 FILLER_195_536 ();
 b15zdnd11an1n04x5 FILLER_195_544 ();
 b15zdnd11an1n16x5 FILLER_195_555 ();
 b15zdnd11an1n04x5 FILLER_195_571 ();
 b15zdnd00an1n02x5 FILLER_195_575 ();
 b15zdnd00an1n01x5 FILLER_195_577 ();
 b15zdnd11an1n16x5 FILLER_195_584 ();
 b15zdnd11an1n64x5 FILLER_195_606 ();
 b15zdnd11an1n16x5 FILLER_195_670 ();
 b15zdnd11an1n04x5 FILLER_195_686 ();
 b15zdnd00an1n01x5 FILLER_195_690 ();
 b15zdnd11an1n32x5 FILLER_195_709 ();
 b15zdnd00an1n02x5 FILLER_195_741 ();
 b15zdnd11an1n64x5 FILLER_195_755 ();
 b15zdnd11an1n64x5 FILLER_195_819 ();
 b15zdnd11an1n64x5 FILLER_195_883 ();
 b15zdnd11an1n08x5 FILLER_195_947 ();
 b15zdnd00an1n02x5 FILLER_195_955 ();
 b15zdnd00an1n01x5 FILLER_195_957 ();
 b15zdnd11an1n04x5 FILLER_195_965 ();
 b15zdnd00an1n02x5 FILLER_195_969 ();
 b15zdnd00an1n01x5 FILLER_195_971 ();
 b15zdnd11an1n08x5 FILLER_195_977 ();
 b15zdnd11an1n04x5 FILLER_195_985 ();
 b15zdnd11an1n64x5 FILLER_195_995 ();
 b15zdnd11an1n32x5 FILLER_195_1059 ();
 b15zdnd11an1n16x5 FILLER_195_1091 ();
 b15zdnd11an1n08x5 FILLER_195_1107 ();
 b15zdnd11an1n04x5 FILLER_195_1115 ();
 b15zdnd00an1n02x5 FILLER_195_1119 ();
 b15zdnd00an1n01x5 FILLER_195_1121 ();
 b15zdnd11an1n64x5 FILLER_195_1132 ();
 b15zdnd11an1n08x5 FILLER_195_1196 ();
 b15zdnd11an1n04x5 FILLER_195_1204 ();
 b15zdnd11an1n64x5 FILLER_195_1213 ();
 b15zdnd11an1n04x5 FILLER_195_1277 ();
 b15zdnd00an1n01x5 FILLER_195_1281 ();
 b15zdnd11an1n16x5 FILLER_195_1289 ();
 b15zdnd11an1n08x5 FILLER_195_1305 ();
 b15zdnd11an1n32x5 FILLER_195_1323 ();
 b15zdnd11an1n08x5 FILLER_195_1355 ();
 b15zdnd11an1n04x5 FILLER_195_1363 ();
 b15zdnd11an1n16x5 FILLER_195_1376 ();
 b15zdnd00an1n02x5 FILLER_195_1392 ();
 b15zdnd11an1n08x5 FILLER_195_1403 ();
 b15zdnd11an1n04x5 FILLER_195_1411 ();
 b15zdnd00an1n02x5 FILLER_195_1415 ();
 b15zdnd00an1n01x5 FILLER_195_1417 ();
 b15zdnd11an1n64x5 FILLER_195_1424 ();
 b15zdnd11an1n08x5 FILLER_195_1488 ();
 b15zdnd00an1n02x5 FILLER_195_1496 ();
 b15zdnd00an1n01x5 FILLER_195_1498 ();
 b15zdnd11an1n32x5 FILLER_195_1510 ();
 b15zdnd00an1n02x5 FILLER_195_1542 ();
 b15zdnd00an1n01x5 FILLER_195_1544 ();
 b15zdnd11an1n64x5 FILLER_195_1561 ();
 b15zdnd11an1n08x5 FILLER_195_1625 ();
 b15zdnd00an1n02x5 FILLER_195_1633 ();
 b15zdnd11an1n16x5 FILLER_195_1640 ();
 b15zdnd11an1n08x5 FILLER_195_1656 ();
 b15zdnd00an1n02x5 FILLER_195_1664 ();
 b15zdnd00an1n01x5 FILLER_195_1666 ();
 b15zdnd11an1n16x5 FILLER_195_1678 ();
 b15zdnd11an1n08x5 FILLER_195_1694 ();
 b15zdnd11an1n04x5 FILLER_195_1702 ();
 b15zdnd00an1n02x5 FILLER_195_1706 ();
 b15zdnd11an1n04x5 FILLER_195_1739 ();
 b15zdnd11an1n04x5 FILLER_195_1764 ();
 b15zdnd11an1n16x5 FILLER_195_1777 ();
 b15zdnd00an1n02x5 FILLER_195_1793 ();
 b15zdnd11an1n64x5 FILLER_195_1805 ();
 b15zdnd11an1n64x5 FILLER_195_1869 ();
 b15zdnd11an1n16x5 FILLER_195_1933 ();
 b15zdnd11an1n08x5 FILLER_195_1949 ();
 b15zdnd11an1n04x5 FILLER_195_1957 ();
 b15zdnd00an1n02x5 FILLER_195_1961 ();
 b15zdnd11an1n32x5 FILLER_195_1983 ();
 b15zdnd11an1n08x5 FILLER_195_2015 ();
 b15zdnd11an1n04x5 FILLER_195_2023 ();
 b15zdnd00an1n02x5 FILLER_195_2027 ();
 b15zdnd11an1n64x5 FILLER_195_2032 ();
 b15zdnd11an1n64x5 FILLER_195_2096 ();
 b15zdnd11an1n64x5 FILLER_195_2160 ();
 b15zdnd11an1n16x5 FILLER_195_2224 ();
 b15zdnd11an1n04x5 FILLER_195_2240 ();
 b15zdnd00an1n01x5 FILLER_195_2244 ();
 b15zdnd11an1n08x5 FILLER_195_2251 ();
 b15zdnd00an1n02x5 FILLER_195_2259 ();
 b15zdnd11an1n04x5 FILLER_195_2269 ();
 b15zdnd00an1n01x5 FILLER_195_2273 ();
 b15zdnd00an1n02x5 FILLER_195_2282 ();
 b15zdnd11an1n16x5 FILLER_196_8 ();
 b15zdnd11an1n04x5 FILLER_196_24 ();
 b15zdnd00an1n02x5 FILLER_196_28 ();
 b15zdnd00an1n01x5 FILLER_196_30 ();
 b15zdnd11an1n08x5 FILLER_196_35 ();
 b15zdnd11an1n04x5 FILLER_196_64 ();
 b15zdnd00an1n01x5 FILLER_196_68 ();
 b15zdnd11an1n32x5 FILLER_196_73 ();
 b15zdnd11an1n16x5 FILLER_196_105 ();
 b15zdnd11an1n04x5 FILLER_196_125 ();
 b15zdnd00an1n02x5 FILLER_196_129 ();
 b15zdnd11an1n04x5 FILLER_196_136 ();
 b15zdnd11an1n04x5 FILLER_196_153 ();
 b15zdnd00an1n02x5 FILLER_196_157 ();
 b15zdnd11an1n32x5 FILLER_196_164 ();
 b15zdnd11an1n16x5 FILLER_196_196 ();
 b15zdnd11an1n04x5 FILLER_196_212 ();
 b15zdnd11an1n04x5 FILLER_196_225 ();
 b15zdnd00an1n01x5 FILLER_196_229 ();
 b15zdnd11an1n08x5 FILLER_196_234 ();
 b15zdnd00an1n02x5 FILLER_196_242 ();
 b15zdnd00an1n01x5 FILLER_196_244 ();
 b15zdnd11an1n08x5 FILLER_196_255 ();
 b15zdnd00an1n02x5 FILLER_196_263 ();
 b15zdnd11an1n04x5 FILLER_196_270 ();
 b15zdnd00an1n02x5 FILLER_196_274 ();
 b15zdnd11an1n04x5 FILLER_196_296 ();
 b15zdnd11an1n64x5 FILLER_196_314 ();
 b15zdnd11an1n04x5 FILLER_196_378 ();
 b15zdnd11an1n08x5 FILLER_196_398 ();
 b15zdnd00an1n02x5 FILLER_196_406 ();
 b15zdnd11an1n04x5 FILLER_196_418 ();
 b15zdnd11an1n08x5 FILLER_196_436 ();
 b15zdnd11an1n04x5 FILLER_196_444 ();
 b15zdnd00an1n02x5 FILLER_196_448 ();
 b15zdnd11an1n32x5 FILLER_196_456 ();
 b15zdnd11an1n04x5 FILLER_196_488 ();
 b15zdnd00an1n01x5 FILLER_196_492 ();
 b15zdnd11an1n04x5 FILLER_196_514 ();
 b15zdnd11an1n32x5 FILLER_196_523 ();
 b15zdnd11an1n16x5 FILLER_196_555 ();
 b15zdnd11an1n04x5 FILLER_196_571 ();
 b15zdnd00an1n02x5 FILLER_196_575 ();
 b15zdnd00an1n01x5 FILLER_196_577 ();
 b15zdnd11an1n16x5 FILLER_196_583 ();
 b15zdnd00an1n01x5 FILLER_196_599 ();
 b15zdnd11an1n04x5 FILLER_196_607 ();
 b15zdnd11an1n16x5 FILLER_196_619 ();
 b15zdnd00an1n02x5 FILLER_196_635 ();
 b15zdnd00an1n01x5 FILLER_196_637 ();
 b15zdnd11an1n16x5 FILLER_196_644 ();
 b15zdnd11an1n08x5 FILLER_196_660 ();
 b15zdnd11an1n04x5 FILLER_196_668 ();
 b15zdnd00an1n02x5 FILLER_196_672 ();
 b15zdnd00an1n01x5 FILLER_196_674 ();
 b15zdnd11an1n04x5 FILLER_196_680 ();
 b15zdnd11an1n08x5 FILLER_196_689 ();
 b15zdnd11an1n04x5 FILLER_196_697 ();
 b15zdnd11an1n04x5 FILLER_196_711 ();
 b15zdnd00an1n02x5 FILLER_196_715 ();
 b15zdnd00an1n01x5 FILLER_196_717 ();
 b15zdnd00an1n02x5 FILLER_196_726 ();
 b15zdnd11an1n04x5 FILLER_196_743 ();
 b15zdnd11an1n16x5 FILLER_196_752 ();
 b15zdnd11an1n04x5 FILLER_196_768 ();
 b15zdnd00an1n02x5 FILLER_196_772 ();
 b15zdnd11an1n64x5 FILLER_196_794 ();
 b15zdnd11an1n64x5 FILLER_196_877 ();
 b15zdnd11an1n16x5 FILLER_196_941 ();
 b15zdnd11an1n08x5 FILLER_196_957 ();
 b15zdnd11an1n04x5 FILLER_196_965 ();
 b15zdnd00an1n02x5 FILLER_196_969 ();
 b15zdnd11an1n32x5 FILLER_196_1007 ();
 b15zdnd11an1n08x5 FILLER_196_1039 ();
 b15zdnd11an1n04x5 FILLER_196_1047 ();
 b15zdnd11an1n32x5 FILLER_196_1057 ();
 b15zdnd11an1n16x5 FILLER_196_1089 ();
 b15zdnd11an1n04x5 FILLER_196_1105 ();
 b15zdnd11an1n16x5 FILLER_196_1126 ();
 b15zdnd11an1n08x5 FILLER_196_1142 ();
 b15zdnd00an1n02x5 FILLER_196_1150 ();
 b15zdnd11an1n64x5 FILLER_196_1172 ();
 b15zdnd11an1n32x5 FILLER_196_1236 ();
 b15zdnd11an1n08x5 FILLER_196_1268 ();
 b15zdnd11an1n08x5 FILLER_196_1286 ();
 b15zdnd11an1n04x5 FILLER_196_1294 ();
 b15zdnd00an1n01x5 FILLER_196_1298 ();
 b15zdnd11an1n16x5 FILLER_196_1308 ();
 b15zdnd11an1n08x5 FILLER_196_1324 ();
 b15zdnd11an1n04x5 FILLER_196_1332 ();
 b15zdnd11an1n64x5 FILLER_196_1341 ();
 b15zdnd11an1n32x5 FILLER_196_1405 ();
 b15zdnd11an1n16x5 FILLER_196_1437 ();
 b15zdnd00an1n01x5 FILLER_196_1453 ();
 b15zdnd11an1n08x5 FILLER_196_1460 ();
 b15zdnd00an1n02x5 FILLER_196_1468 ();
 b15zdnd00an1n01x5 FILLER_196_1470 ();
 b15zdnd11an1n04x5 FILLER_196_1481 ();
 b15zdnd11an1n04x5 FILLER_196_1494 ();
 b15zdnd00an1n02x5 FILLER_196_1498 ();
 b15zdnd00an1n01x5 FILLER_196_1500 ();
 b15zdnd11an1n04x5 FILLER_196_1505 ();
 b15zdnd11an1n04x5 FILLER_196_1514 ();
 b15zdnd00an1n01x5 FILLER_196_1518 ();
 b15zdnd11an1n04x5 FILLER_196_1535 ();
 b15zdnd00an1n01x5 FILLER_196_1539 ();
 b15zdnd11an1n04x5 FILLER_196_1561 ();
 b15zdnd00an1n01x5 FILLER_196_1565 ();
 b15zdnd11an1n64x5 FILLER_196_1570 ();
 b15zdnd00an1n01x5 FILLER_196_1634 ();
 b15zdnd11an1n64x5 FILLER_196_1645 ();
 b15zdnd11an1n64x5 FILLER_196_1709 ();
 b15zdnd11an1n64x5 FILLER_196_1773 ();
 b15zdnd11an1n64x5 FILLER_196_1837 ();
 b15zdnd11an1n32x5 FILLER_196_1901 ();
 b15zdnd00an1n01x5 FILLER_196_1933 ();
 b15zdnd11an1n16x5 FILLER_196_1949 ();
 b15zdnd00an1n01x5 FILLER_196_1965 ();
 b15zdnd11an1n08x5 FILLER_196_1990 ();
 b15zdnd11an1n16x5 FILLER_196_2018 ();
 b15zdnd00an1n02x5 FILLER_196_2034 ();
 b15zdnd11an1n16x5 FILLER_196_2053 ();
 b15zdnd11an1n04x5 FILLER_196_2069 ();
 b15zdnd00an1n02x5 FILLER_196_2073 ();
 b15zdnd11an1n32x5 FILLER_196_2095 ();
 b15zdnd11an1n16x5 FILLER_196_2127 ();
 b15zdnd11an1n08x5 FILLER_196_2143 ();
 b15zdnd00an1n02x5 FILLER_196_2151 ();
 b15zdnd00an1n01x5 FILLER_196_2153 ();
 b15zdnd11an1n08x5 FILLER_196_2162 ();
 b15zdnd00an1n02x5 FILLER_196_2170 ();
 b15zdnd00an1n01x5 FILLER_196_2172 ();
 b15zdnd11an1n32x5 FILLER_196_2179 ();
 b15zdnd11an1n04x5 FILLER_196_2211 ();
 b15zdnd11an1n32x5 FILLER_196_2224 ();
 b15zdnd11an1n16x5 FILLER_196_2256 ();
 b15zdnd11an1n04x5 FILLER_196_2272 ();
 b15zdnd11an1n32x5 FILLER_197_0 ();
 b15zdnd11an1n08x5 FILLER_197_32 ();
 b15zdnd00an1n01x5 FILLER_197_40 ();
 b15zdnd11an1n16x5 FILLER_197_57 ();
 b15zdnd00an1n02x5 FILLER_197_73 ();
 b15zdnd11an1n32x5 FILLER_197_81 ();
 b15zdnd11an1n04x5 FILLER_197_113 ();
 b15zdnd00an1n01x5 FILLER_197_117 ();
 b15zdnd11an1n32x5 FILLER_197_126 ();
 b15zdnd00an1n01x5 FILLER_197_158 ();
 b15zdnd11an1n16x5 FILLER_197_165 ();
 b15zdnd11an1n08x5 FILLER_197_195 ();
 b15zdnd00an1n02x5 FILLER_197_203 ();
 b15zdnd00an1n01x5 FILLER_197_205 ();
 b15zdnd11an1n08x5 FILLER_197_226 ();
 b15zdnd11an1n04x5 FILLER_197_234 ();
 b15zdnd00an1n02x5 FILLER_197_238 ();
 b15zdnd00an1n01x5 FILLER_197_240 ();
 b15zdnd11an1n04x5 FILLER_197_251 ();
 b15zdnd00an1n02x5 FILLER_197_255 ();
 b15zdnd11an1n16x5 FILLER_197_273 ();
 b15zdnd11an1n08x5 FILLER_197_289 ();
 b15zdnd11an1n04x5 FILLER_197_297 ();
 b15zdnd00an1n01x5 FILLER_197_301 ();
 b15zdnd11an1n04x5 FILLER_197_322 ();
 b15zdnd11an1n64x5 FILLER_197_352 ();
 b15zdnd11an1n32x5 FILLER_197_416 ();
 b15zdnd11an1n16x5 FILLER_197_448 ();
 b15zdnd00an1n01x5 FILLER_197_464 ();
 b15zdnd11an1n64x5 FILLER_197_472 ();
 b15zdnd11an1n08x5 FILLER_197_536 ();
 b15zdnd11an1n04x5 FILLER_197_544 ();
 b15zdnd00an1n02x5 FILLER_197_548 ();
 b15zdnd00an1n01x5 FILLER_197_550 ();
 b15zdnd11an1n16x5 FILLER_197_563 ();
 b15zdnd11an1n04x5 FILLER_197_579 ();
 b15zdnd00an1n02x5 FILLER_197_583 ();
 b15zdnd00an1n01x5 FILLER_197_585 ();
 b15zdnd11an1n32x5 FILLER_197_600 ();
 b15zdnd11an1n04x5 FILLER_197_632 ();
 b15zdnd00an1n02x5 FILLER_197_636 ();
 b15zdnd00an1n01x5 FILLER_197_638 ();
 b15zdnd11an1n04x5 FILLER_197_647 ();
 b15zdnd11an1n16x5 FILLER_197_656 ();
 b15zdnd11an1n08x5 FILLER_197_672 ();
 b15zdnd11an1n04x5 FILLER_197_685 ();
 b15zdnd11an1n64x5 FILLER_197_698 ();
 b15zdnd11an1n64x5 FILLER_197_762 ();
 b15zdnd11an1n64x5 FILLER_197_826 ();
 b15zdnd11an1n32x5 FILLER_197_890 ();
 b15zdnd11an1n04x5 FILLER_197_922 ();
 b15zdnd00an1n02x5 FILLER_197_926 ();
 b15zdnd11an1n04x5 FILLER_197_936 ();
 b15zdnd11an1n32x5 FILLER_197_944 ();
 b15zdnd11an1n08x5 FILLER_197_976 ();
 b15zdnd00an1n02x5 FILLER_197_984 ();
 b15zdnd00an1n01x5 FILLER_197_986 ();
 b15zdnd11an1n08x5 FILLER_197_1004 ();
 b15zdnd11an1n04x5 FILLER_197_1012 ();
 b15zdnd00an1n02x5 FILLER_197_1016 ();
 b15zdnd00an1n01x5 FILLER_197_1018 ();
 b15zdnd11an1n04x5 FILLER_197_1026 ();
 b15zdnd11an1n16x5 FILLER_197_1056 ();
 b15zdnd11an1n04x5 FILLER_197_1072 ();
 b15zdnd00an1n02x5 FILLER_197_1076 ();
 b15zdnd11an1n08x5 FILLER_197_1084 ();
 b15zdnd11an1n04x5 FILLER_197_1092 ();
 b15zdnd00an1n01x5 FILLER_197_1096 ();
 b15zdnd11an1n16x5 FILLER_197_1102 ();
 b15zdnd11an1n04x5 FILLER_197_1118 ();
 b15zdnd11an1n16x5 FILLER_197_1127 ();
 b15zdnd11an1n04x5 FILLER_197_1143 ();
 b15zdnd11an1n04x5 FILLER_197_1159 ();
 b15zdnd11an1n04x5 FILLER_197_1175 ();
 b15zdnd11an1n04x5 FILLER_197_1186 ();
 b15zdnd11an1n16x5 FILLER_197_1194 ();
 b15zdnd11an1n08x5 FILLER_197_1210 ();
 b15zdnd11an1n04x5 FILLER_197_1218 ();
 b15zdnd00an1n01x5 FILLER_197_1222 ();
 b15zdnd11an1n64x5 FILLER_197_1228 ();
 b15zdnd11an1n16x5 FILLER_197_1292 ();
 b15zdnd00an1n02x5 FILLER_197_1308 ();
 b15zdnd11an1n16x5 FILLER_197_1316 ();
 b15zdnd00an1n02x5 FILLER_197_1332 ();
 b15zdnd11an1n04x5 FILLER_197_1346 ();
 b15zdnd11an1n08x5 FILLER_197_1355 ();
 b15zdnd11an1n04x5 FILLER_197_1363 ();
 b15zdnd00an1n01x5 FILLER_197_1367 ();
 b15zdnd11an1n16x5 FILLER_197_1373 ();
 b15zdnd11an1n32x5 FILLER_197_1393 ();
 b15zdnd11an1n08x5 FILLER_197_1425 ();
 b15zdnd11an1n64x5 FILLER_197_1437 ();
 b15zdnd11an1n08x5 FILLER_197_1501 ();
 b15zdnd11an1n32x5 FILLER_197_1515 ();
 b15zdnd11an1n16x5 FILLER_197_1556 ();
 b15zdnd11an1n08x5 FILLER_197_1572 ();
 b15zdnd00an1n02x5 FILLER_197_1580 ();
 b15zdnd00an1n01x5 FILLER_197_1582 ();
 b15zdnd11an1n16x5 FILLER_197_1588 ();
 b15zdnd11an1n04x5 FILLER_197_1604 ();
 b15zdnd00an1n02x5 FILLER_197_1608 ();
 b15zdnd00an1n01x5 FILLER_197_1610 ();
 b15zdnd11an1n16x5 FILLER_197_1616 ();
 b15zdnd00an1n02x5 FILLER_197_1632 ();
 b15zdnd00an1n01x5 FILLER_197_1634 ();
 b15zdnd11an1n16x5 FILLER_197_1640 ();
 b15zdnd11an1n08x5 FILLER_197_1656 ();
 b15zdnd00an1n02x5 FILLER_197_1664 ();
 b15zdnd11an1n04x5 FILLER_197_1672 ();
 b15zdnd11an1n04x5 FILLER_197_1682 ();
 b15zdnd11an1n64x5 FILLER_197_1706 ();
 b15zdnd11an1n64x5 FILLER_197_1770 ();
 b15zdnd11an1n16x5 FILLER_197_1834 ();
 b15zdnd11an1n08x5 FILLER_197_1850 ();
 b15zdnd00an1n02x5 FILLER_197_1858 ();
 b15zdnd00an1n01x5 FILLER_197_1860 ();
 b15zdnd11an1n08x5 FILLER_197_1881 ();
 b15zdnd11an1n04x5 FILLER_197_1889 ();
 b15zdnd11an1n64x5 FILLER_197_1913 ();
 b15zdnd11an1n04x5 FILLER_197_1977 ();
 b15zdnd00an1n02x5 FILLER_197_1981 ();
 b15zdnd11an1n08x5 FILLER_197_1987 ();
 b15zdnd11an1n04x5 FILLER_197_1995 ();
 b15zdnd11an1n32x5 FILLER_197_2004 ();
 b15zdnd11an1n04x5 FILLER_197_2036 ();
 b15zdnd00an1n02x5 FILLER_197_2040 ();
 b15zdnd00an1n01x5 FILLER_197_2042 ();
 b15zdnd11an1n32x5 FILLER_197_2048 ();
 b15zdnd11an1n04x5 FILLER_197_2080 ();
 b15zdnd11an1n32x5 FILLER_197_2104 ();
 b15zdnd11an1n16x5 FILLER_197_2136 ();
 b15zdnd11an1n08x5 FILLER_197_2152 ();
 b15zdnd11an1n04x5 FILLER_197_2160 ();
 b15zdnd00an1n02x5 FILLER_197_2164 ();
 b15zdnd00an1n01x5 FILLER_197_2166 ();
 b15zdnd11an1n16x5 FILLER_197_2187 ();
 b15zdnd11an1n08x5 FILLER_197_2203 ();
 b15zdnd00an1n01x5 FILLER_197_2211 ();
 b15zdnd11an1n16x5 FILLER_197_2223 ();
 b15zdnd11an1n08x5 FILLER_197_2242 ();
 b15zdnd11an1n04x5 FILLER_197_2250 ();
 b15zdnd11an1n04x5 FILLER_197_2258 ();
 b15zdnd11an1n04x5 FILLER_197_2267 ();
 b15zdnd00an1n01x5 FILLER_197_2271 ();
 b15zdnd11an1n08x5 FILLER_197_2276 ();
 b15zdnd11an1n16x5 FILLER_198_8 ();
 b15zdnd00an1n01x5 FILLER_198_24 ();
 b15zdnd11an1n32x5 FILLER_198_33 ();
 b15zdnd00an1n02x5 FILLER_198_65 ();
 b15zdnd11an1n64x5 FILLER_198_77 ();
 b15zdnd11an1n16x5 FILLER_198_141 ();
 b15zdnd00an1n02x5 FILLER_198_157 ();
 b15zdnd11an1n16x5 FILLER_198_163 ();
 b15zdnd11an1n04x5 FILLER_198_179 ();
 b15zdnd00an1n01x5 FILLER_198_183 ();
 b15zdnd11an1n04x5 FILLER_198_189 ();
 b15zdnd11an1n04x5 FILLER_198_219 ();
 b15zdnd11an1n32x5 FILLER_198_228 ();
 b15zdnd11an1n16x5 FILLER_198_260 ();
 b15zdnd00an1n01x5 FILLER_198_276 ();
 b15zdnd11an1n08x5 FILLER_198_293 ();
 b15zdnd00an1n02x5 FILLER_198_301 ();
 b15zdnd00an1n01x5 FILLER_198_303 ();
 b15zdnd11an1n08x5 FILLER_198_330 ();
 b15zdnd00an1n01x5 FILLER_198_338 ();
 b15zdnd11an1n64x5 FILLER_198_371 ();
 b15zdnd11an1n16x5 FILLER_198_435 ();
 b15zdnd00an1n02x5 FILLER_198_451 ();
 b15zdnd11an1n08x5 FILLER_198_459 ();
 b15zdnd11an1n04x5 FILLER_198_467 ();
 b15zdnd00an1n01x5 FILLER_198_471 ();
 b15zdnd11an1n16x5 FILLER_198_480 ();
 b15zdnd11an1n32x5 FILLER_198_500 ();
 b15zdnd11an1n16x5 FILLER_198_532 ();
 b15zdnd00an1n02x5 FILLER_198_548 ();
 b15zdnd00an1n01x5 FILLER_198_550 ();
 b15zdnd11an1n32x5 FILLER_198_559 ();
 b15zdnd11an1n04x5 FILLER_198_591 ();
 b15zdnd00an1n02x5 FILLER_198_595 ();
 b15zdnd11an1n64x5 FILLER_198_603 ();
 b15zdnd11an1n16x5 FILLER_198_667 ();
 b15zdnd11an1n08x5 FILLER_198_683 ();
 b15zdnd11an1n04x5 FILLER_198_691 ();
 b15zdnd00an1n01x5 FILLER_198_695 ();
 b15zdnd00an1n02x5 FILLER_198_716 ();
 b15zdnd11an1n32x5 FILLER_198_726 ();
 b15zdnd11an1n04x5 FILLER_198_758 ();
 b15zdnd00an1n02x5 FILLER_198_762 ();
 b15zdnd11an1n64x5 FILLER_198_782 ();
 b15zdnd11an1n16x5 FILLER_198_846 ();
 b15zdnd11an1n08x5 FILLER_198_862 ();
 b15zdnd00an1n01x5 FILLER_198_870 ();
 b15zdnd11an1n16x5 FILLER_198_876 ();
 b15zdnd00an1n01x5 FILLER_198_892 ();
 b15zdnd11an1n16x5 FILLER_198_900 ();
 b15zdnd11an1n08x5 FILLER_198_916 ();
 b15zdnd11an1n04x5 FILLER_198_924 ();
 b15zdnd00an1n02x5 FILLER_198_928 ();
 b15zdnd11an1n64x5 FILLER_198_939 ();
 b15zdnd11an1n32x5 FILLER_198_1003 ();
 b15zdnd11an1n04x5 FILLER_198_1035 ();
 b15zdnd00an1n01x5 FILLER_198_1039 ();
 b15zdnd11an1n32x5 FILLER_198_1044 ();
 b15zdnd11an1n04x5 FILLER_198_1076 ();
 b15zdnd00an1n01x5 FILLER_198_1080 ();
 b15zdnd11an1n04x5 FILLER_198_1093 ();
 b15zdnd11an1n16x5 FILLER_198_1102 ();
 b15zdnd11an1n08x5 FILLER_198_1118 ();
 b15zdnd00an1n02x5 FILLER_198_1126 ();
 b15zdnd00an1n01x5 FILLER_198_1128 ();
 b15zdnd11an1n08x5 FILLER_198_1135 ();
 b15zdnd11an1n16x5 FILLER_198_1169 ();
 b15zdnd11an1n08x5 FILLER_198_1185 ();
 b15zdnd00an1n01x5 FILLER_198_1193 ();
 b15zdnd11an1n64x5 FILLER_198_1220 ();
 b15zdnd11an1n32x5 FILLER_198_1284 ();
 b15zdnd11an1n16x5 FILLER_198_1316 ();
 b15zdnd00an1n01x5 FILLER_198_1332 ();
 b15zdnd11an1n08x5 FILLER_198_1347 ();
 b15zdnd00an1n02x5 FILLER_198_1355 ();
 b15zdnd11an1n08x5 FILLER_198_1374 ();
 b15zdnd11an1n04x5 FILLER_198_1382 ();
 b15zdnd00an1n02x5 FILLER_198_1386 ();
 b15zdnd00an1n01x5 FILLER_198_1388 ();
 b15zdnd11an1n16x5 FILLER_198_1399 ();
 b15zdnd00an1n02x5 FILLER_198_1415 ();
 b15zdnd00an1n01x5 FILLER_198_1417 ();
 b15zdnd11an1n16x5 FILLER_198_1433 ();
 b15zdnd00an1n02x5 FILLER_198_1449 ();
 b15zdnd00an1n01x5 FILLER_198_1451 ();
 b15zdnd11an1n64x5 FILLER_198_1463 ();
 b15zdnd11an1n32x5 FILLER_198_1527 ();
 b15zdnd11an1n04x5 FILLER_198_1559 ();
 b15zdnd00an1n02x5 FILLER_198_1563 ();
 b15zdnd11an1n04x5 FILLER_198_1577 ();
 b15zdnd11an1n32x5 FILLER_198_1589 ();
 b15zdnd11an1n08x5 FILLER_198_1621 ();
 b15zdnd00an1n02x5 FILLER_198_1629 ();
 b15zdnd00an1n01x5 FILLER_198_1631 ();
 b15zdnd11an1n08x5 FILLER_198_1636 ();
 b15zdnd11an1n04x5 FILLER_198_1644 ();
 b15zdnd00an1n02x5 FILLER_198_1648 ();
 b15zdnd00an1n01x5 FILLER_198_1650 ();
 b15zdnd11an1n64x5 FILLER_198_1677 ();
 b15zdnd11an1n64x5 FILLER_198_1741 ();
 b15zdnd11an1n32x5 FILLER_198_1805 ();
 b15zdnd11an1n08x5 FILLER_198_1837 ();
 b15zdnd00an1n02x5 FILLER_198_1845 ();
 b15zdnd11an1n04x5 FILLER_198_1859 ();
 b15zdnd11an1n04x5 FILLER_198_1872 ();
 b15zdnd11an1n08x5 FILLER_198_1888 ();
 b15zdnd00an1n02x5 FILLER_198_1896 ();
 b15zdnd11an1n04x5 FILLER_198_1903 ();
 b15zdnd00an1n02x5 FILLER_198_1907 ();
 b15zdnd00an1n01x5 FILLER_198_1909 ();
 b15zdnd11an1n64x5 FILLER_198_1916 ();
 b15zdnd00an1n02x5 FILLER_198_1980 ();
 b15zdnd00an1n01x5 FILLER_198_1982 ();
 b15zdnd11an1n04x5 FILLER_198_1988 ();
 b15zdnd11an1n32x5 FILLER_198_2001 ();
 b15zdnd00an1n01x5 FILLER_198_2033 ();
 b15zdnd11an1n64x5 FILLER_198_2054 ();
 b15zdnd11an1n08x5 FILLER_198_2118 ();
 b15zdnd00an1n02x5 FILLER_198_2126 ();
 b15zdnd00an1n01x5 FILLER_198_2128 ();
 b15zdnd11an1n04x5 FILLER_198_2149 ();
 b15zdnd00an1n01x5 FILLER_198_2153 ();
 b15zdnd11an1n08x5 FILLER_198_2162 ();
 b15zdnd11an1n04x5 FILLER_198_2170 ();
 b15zdnd11an1n64x5 FILLER_198_2179 ();
 b15zdnd00an1n02x5 FILLER_198_2243 ();
 b15zdnd11an1n08x5 FILLER_198_2249 ();
 b15zdnd11an1n04x5 FILLER_198_2257 ();
 b15zdnd11an1n04x5 FILLER_198_2265 ();
 b15zdnd00an1n01x5 FILLER_198_2269 ();
 b15zdnd00an1n02x5 FILLER_198_2274 ();
 b15zdnd11an1n08x5 FILLER_199_0 ();
 b15zdnd11an1n04x5 FILLER_199_8 ();
 b15zdnd11an1n04x5 FILLER_199_16 ();
 b15zdnd11an1n08x5 FILLER_199_24 ();
 b15zdnd11an1n04x5 FILLER_199_32 ();
 b15zdnd00an1n02x5 FILLER_199_36 ();
 b15zdnd00an1n01x5 FILLER_199_38 ();
 b15zdnd11an1n16x5 FILLER_199_47 ();
 b15zdnd00an1n01x5 FILLER_199_63 ();
 b15zdnd11an1n04x5 FILLER_199_76 ();
 b15zdnd00an1n02x5 FILLER_199_80 ();
 b15zdnd11an1n32x5 FILLER_199_88 ();
 b15zdnd00an1n01x5 FILLER_199_120 ();
 b15zdnd11an1n32x5 FILLER_199_127 ();
 b15zdnd11an1n16x5 FILLER_199_159 ();
 b15zdnd11an1n04x5 FILLER_199_175 ();
 b15zdnd11an1n04x5 FILLER_199_189 ();
 b15zdnd11an1n64x5 FILLER_199_219 ();
 b15zdnd11an1n16x5 FILLER_199_283 ();
 b15zdnd11an1n08x5 FILLER_199_299 ();
 b15zdnd00an1n01x5 FILLER_199_307 ();
 b15zdnd11an1n32x5 FILLER_199_329 ();
 b15zdnd11an1n16x5 FILLER_199_361 ();
 b15zdnd00an1n01x5 FILLER_199_377 ();
 b15zdnd11an1n08x5 FILLER_199_399 ();
 b15zdnd00an1n02x5 FILLER_199_407 ();
 b15zdnd11an1n16x5 FILLER_199_414 ();
 b15zdnd11an1n04x5 FILLER_199_430 ();
 b15zdnd00an1n02x5 FILLER_199_434 ();
 b15zdnd11an1n08x5 FILLER_199_443 ();
 b15zdnd11an1n04x5 FILLER_199_451 ();
 b15zdnd00an1n02x5 FILLER_199_455 ();
 b15zdnd00an1n01x5 FILLER_199_457 ();
 b15zdnd11an1n04x5 FILLER_199_465 ();
 b15zdnd00an1n02x5 FILLER_199_469 ();
 b15zdnd00an1n01x5 FILLER_199_471 ();
 b15zdnd11an1n32x5 FILLER_199_477 ();
 b15zdnd11an1n04x5 FILLER_199_509 ();
 b15zdnd00an1n02x5 FILLER_199_513 ();
 b15zdnd00an1n01x5 FILLER_199_515 ();
 b15zdnd11an1n16x5 FILLER_199_520 ();
 b15zdnd11an1n08x5 FILLER_199_536 ();
 b15zdnd00an1n01x5 FILLER_199_544 ();
 b15zdnd11an1n04x5 FILLER_199_552 ();
 b15zdnd11an1n64x5 FILLER_199_566 ();
 b15zdnd11an1n32x5 FILLER_199_630 ();
 b15zdnd11an1n04x5 FILLER_199_662 ();
 b15zdnd11an1n64x5 FILLER_199_673 ();
 b15zdnd11an1n64x5 FILLER_199_737 ();
 b15zdnd11an1n64x5 FILLER_199_801 ();
 b15zdnd00an1n02x5 FILLER_199_865 ();
 b15zdnd11an1n08x5 FILLER_199_873 ();
 b15zdnd00an1n01x5 FILLER_199_881 ();
 b15zdnd11an1n16x5 FILLER_199_892 ();
 b15zdnd11an1n16x5 FILLER_199_914 ();
 b15zdnd00an1n01x5 FILLER_199_930 ();
 b15zdnd11an1n64x5 FILLER_199_935 ();
 b15zdnd11an1n04x5 FILLER_199_999 ();
 b15zdnd00an1n01x5 FILLER_199_1003 ();
 b15zdnd11an1n08x5 FILLER_199_1014 ();
 b15zdnd00an1n02x5 FILLER_199_1022 ();
 b15zdnd00an1n01x5 FILLER_199_1024 ();
 b15zdnd11an1n04x5 FILLER_199_1032 ();
 b15zdnd11an1n32x5 FILLER_199_1051 ();
 b15zdnd11an1n08x5 FILLER_199_1083 ();
 b15zdnd11an1n04x5 FILLER_199_1091 ();
 b15zdnd00an1n02x5 FILLER_199_1095 ();
 b15zdnd11an1n16x5 FILLER_199_1103 ();
 b15zdnd11an1n04x5 FILLER_199_1119 ();
 b15zdnd00an1n01x5 FILLER_199_1123 ();
 b15zdnd11an1n08x5 FILLER_199_1130 ();
 b15zdnd11an1n04x5 FILLER_199_1138 ();
 b15zdnd11an1n32x5 FILLER_199_1147 ();
 b15zdnd11an1n08x5 FILLER_199_1179 ();
 b15zdnd11an1n04x5 FILLER_199_1187 ();
 b15zdnd00an1n01x5 FILLER_199_1191 ();
 b15zdnd11an1n08x5 FILLER_199_1212 ();
 b15zdnd11an1n04x5 FILLER_199_1220 ();
 b15zdnd11an1n64x5 FILLER_199_1234 ();
 b15zdnd11an1n32x5 FILLER_199_1298 ();
 b15zdnd11an1n16x5 FILLER_199_1330 ();
 b15zdnd11an1n08x5 FILLER_199_1346 ();
 b15zdnd00an1n01x5 FILLER_199_1354 ();
 b15zdnd11an1n16x5 FILLER_199_1361 ();
 b15zdnd11an1n08x5 FILLER_199_1377 ();
 b15zdnd11an1n04x5 FILLER_199_1385 ();
 b15zdnd00an1n02x5 FILLER_199_1389 ();
 b15zdnd11an1n64x5 FILLER_199_1397 ();
 b15zdnd11an1n08x5 FILLER_199_1461 ();
 b15zdnd00an1n02x5 FILLER_199_1469 ();
 b15zdnd11an1n08x5 FILLER_199_1502 ();
 b15zdnd00an1n02x5 FILLER_199_1510 ();
 b15zdnd00an1n01x5 FILLER_199_1512 ();
 b15zdnd11an1n16x5 FILLER_199_1522 ();
 b15zdnd11an1n08x5 FILLER_199_1538 ();
 b15zdnd00an1n02x5 FILLER_199_1546 ();
 b15zdnd11an1n32x5 FILLER_199_1555 ();
 b15zdnd11an1n08x5 FILLER_199_1587 ();
 b15zdnd11an1n04x5 FILLER_199_1604 ();
 b15zdnd11an1n16x5 FILLER_199_1620 ();
 b15zdnd11an1n08x5 FILLER_199_1636 ();
 b15zdnd11an1n04x5 FILLER_199_1644 ();
 b15zdnd00an1n02x5 FILLER_199_1648 ();
 b15zdnd00an1n01x5 FILLER_199_1650 ();
 b15zdnd11an1n16x5 FILLER_199_1656 ();
 b15zdnd11an1n16x5 FILLER_199_1677 ();
 b15zdnd11an1n08x5 FILLER_199_1693 ();
 b15zdnd11an1n04x5 FILLER_199_1726 ();
 b15zdnd11an1n16x5 FILLER_199_1742 ();
 b15zdnd11an1n04x5 FILLER_199_1758 ();
 b15zdnd11an1n32x5 FILLER_199_1802 ();
 b15zdnd00an1n01x5 FILLER_199_1834 ();
 b15zdnd11an1n08x5 FILLER_199_1859 ();
 b15zdnd00an1n02x5 FILLER_199_1867 ();
 b15zdnd00an1n01x5 FILLER_199_1869 ();
 b15zdnd11an1n16x5 FILLER_199_1896 ();
 b15zdnd11an1n04x5 FILLER_199_1912 ();
 b15zdnd11an1n16x5 FILLER_199_1956 ();
 b15zdnd00an1n02x5 FILLER_199_1972 ();
 b15zdnd11an1n64x5 FILLER_199_1995 ();
 b15zdnd11an1n64x5 FILLER_199_2059 ();
 b15zdnd11an1n08x5 FILLER_199_2123 ();
 b15zdnd11an1n04x5 FILLER_199_2131 ();
 b15zdnd00an1n01x5 FILLER_199_2135 ();
 b15zdnd11an1n64x5 FILLER_199_2141 ();
 b15zdnd00an1n02x5 FILLER_199_2205 ();
 b15zdnd00an1n01x5 FILLER_199_2207 ();
 b15zdnd11an1n16x5 FILLER_199_2228 ();
 b15zdnd00an1n02x5 FILLER_199_2244 ();
 b15zdnd00an1n01x5 FILLER_199_2246 ();
 b15zdnd11an1n04x5 FILLER_199_2251 ();
 b15zdnd11an1n04x5 FILLER_199_2266 ();
 b15zdnd11an1n08x5 FILLER_199_2274 ();
 b15zdnd00an1n02x5 FILLER_199_2282 ();
 b15zdnd11an1n64x5 FILLER_200_8 ();
 b15zdnd11an1n32x5 FILLER_200_72 ();
 b15zdnd00an1n01x5 FILLER_200_104 ();
 b15zdnd11an1n16x5 FILLER_200_131 ();
 b15zdnd00an1n02x5 FILLER_200_147 ();
 b15zdnd00an1n01x5 FILLER_200_149 ();
 b15zdnd11an1n04x5 FILLER_200_156 ();
 b15zdnd00an1n02x5 FILLER_200_160 ();
 b15zdnd11an1n08x5 FILLER_200_168 ();
 b15zdnd11an1n04x5 FILLER_200_176 ();
 b15zdnd00an1n02x5 FILLER_200_180 ();
 b15zdnd11an1n32x5 FILLER_200_195 ();
 b15zdnd11an1n16x5 FILLER_200_227 ();
 b15zdnd00an1n02x5 FILLER_200_243 ();
 b15zdnd11an1n32x5 FILLER_200_251 ();
 b15zdnd11an1n08x5 FILLER_200_283 ();
 b15zdnd00an1n01x5 FILLER_200_291 ();
 b15zdnd11an1n04x5 FILLER_200_315 ();
 b15zdnd11an1n32x5 FILLER_200_343 ();
 b15zdnd11an1n08x5 FILLER_200_375 ();
 b15zdnd11an1n04x5 FILLER_200_383 ();
 b15zdnd11an1n04x5 FILLER_200_397 ();
 b15zdnd11an1n04x5 FILLER_200_407 ();
 b15zdnd11an1n64x5 FILLER_200_418 ();
 b15zdnd11an1n08x5 FILLER_200_482 ();
 b15zdnd11an1n04x5 FILLER_200_490 ();
 b15zdnd00an1n01x5 FILLER_200_494 ();
 b15zdnd11an1n32x5 FILLER_200_525 ();
 b15zdnd11an1n16x5 FILLER_200_557 ();
 b15zdnd11an1n04x5 FILLER_200_573 ();
 b15zdnd00an1n02x5 FILLER_200_577 ();
 b15zdnd00an1n01x5 FILLER_200_579 ();
 b15zdnd11an1n32x5 FILLER_200_589 ();
 b15zdnd11an1n16x5 FILLER_200_621 ();
 b15zdnd11an1n08x5 FILLER_200_637 ();
 b15zdnd11an1n04x5 FILLER_200_645 ();
 b15zdnd11an1n16x5 FILLER_200_656 ();
 b15zdnd00an1n02x5 FILLER_200_672 ();
 b15zdnd11an1n32x5 FILLER_200_683 ();
 b15zdnd00an1n02x5 FILLER_200_715 ();
 b15zdnd00an1n01x5 FILLER_200_717 ();
 b15zdnd00an1n02x5 FILLER_200_726 ();
 b15zdnd00an1n01x5 FILLER_200_728 ();
 b15zdnd11an1n64x5 FILLER_200_760 ();
 b15zdnd11an1n08x5 FILLER_200_824 ();
 b15zdnd11an1n04x5 FILLER_200_832 ();
 b15zdnd00an1n02x5 FILLER_200_836 ();
 b15zdnd11an1n64x5 FILLER_200_850 ();
 b15zdnd11an1n16x5 FILLER_200_914 ();
 b15zdnd00an1n02x5 FILLER_200_930 ();
 b15zdnd00an1n01x5 FILLER_200_932 ();
 b15zdnd11an1n16x5 FILLER_200_939 ();
 b15zdnd11an1n08x5 FILLER_200_955 ();
 b15zdnd11an1n04x5 FILLER_200_963 ();
 b15zdnd00an1n02x5 FILLER_200_967 ();
 b15zdnd11an1n04x5 FILLER_200_976 ();
 b15zdnd11an1n32x5 FILLER_200_986 ();
 b15zdnd11an1n16x5 FILLER_200_1018 ();
 b15zdnd00an1n01x5 FILLER_200_1034 ();
 b15zdnd11an1n64x5 FILLER_200_1053 ();
 b15zdnd11an1n08x5 FILLER_200_1117 ();
 b15zdnd00an1n02x5 FILLER_200_1125 ();
 b15zdnd00an1n01x5 FILLER_200_1127 ();
 b15zdnd11an1n16x5 FILLER_200_1134 ();
 b15zdnd11an1n08x5 FILLER_200_1150 ();
 b15zdnd00an1n02x5 FILLER_200_1158 ();
 b15zdnd11an1n04x5 FILLER_200_1172 ();
 b15zdnd11an1n32x5 FILLER_200_1180 ();
 b15zdnd11an1n32x5 FILLER_200_1222 ();
 b15zdnd11an1n16x5 FILLER_200_1254 ();
 b15zdnd11an1n04x5 FILLER_200_1270 ();
 b15zdnd11an1n32x5 FILLER_200_1288 ();
 b15zdnd11an1n16x5 FILLER_200_1320 ();
 b15zdnd11an1n04x5 FILLER_200_1336 ();
 b15zdnd00an1n02x5 FILLER_200_1340 ();
 b15zdnd11an1n32x5 FILLER_200_1352 ();
 b15zdnd00an1n02x5 FILLER_200_1384 ();
 b15zdnd11an1n32x5 FILLER_200_1393 ();
 b15zdnd11an1n16x5 FILLER_200_1425 ();
 b15zdnd11an1n08x5 FILLER_200_1441 ();
 b15zdnd00an1n01x5 FILLER_200_1449 ();
 b15zdnd11an1n64x5 FILLER_200_1454 ();
 b15zdnd11an1n64x5 FILLER_200_1518 ();
 b15zdnd11an1n16x5 FILLER_200_1582 ();
 b15zdnd11an1n04x5 FILLER_200_1598 ();
 b15zdnd00an1n01x5 FILLER_200_1602 ();
 b15zdnd11an1n32x5 FILLER_200_1613 ();
 b15zdnd11an1n16x5 FILLER_200_1645 ();
 b15zdnd11an1n04x5 FILLER_200_1661 ();
 b15zdnd11an1n32x5 FILLER_200_1682 ();
 b15zdnd11an1n04x5 FILLER_200_1714 ();
 b15zdnd00an1n02x5 FILLER_200_1718 ();
 b15zdnd11an1n04x5 FILLER_200_1745 ();
 b15zdnd11an1n08x5 FILLER_200_1775 ();
 b15zdnd00an1n01x5 FILLER_200_1783 ();
 b15zdnd11an1n16x5 FILLER_200_1793 ();
 b15zdnd11an1n08x5 FILLER_200_1809 ();
 b15zdnd11an1n04x5 FILLER_200_1826 ();
 b15zdnd11an1n64x5 FILLER_200_1842 ();
 b15zdnd11an1n64x5 FILLER_200_1906 ();
 b15zdnd11an1n64x5 FILLER_200_1970 ();
 b15zdnd11an1n32x5 FILLER_200_2034 ();
 b15zdnd11an1n16x5 FILLER_200_2066 ();
 b15zdnd11an1n08x5 FILLER_200_2082 ();
 b15zdnd11an1n04x5 FILLER_200_2090 ();
 b15zdnd00an1n02x5 FILLER_200_2094 ();
 b15zdnd11an1n32x5 FILLER_200_2099 ();
 b15zdnd11an1n16x5 FILLER_200_2131 ();
 b15zdnd11an1n04x5 FILLER_200_2147 ();
 b15zdnd00an1n02x5 FILLER_200_2151 ();
 b15zdnd00an1n01x5 FILLER_200_2153 ();
 b15zdnd11an1n64x5 FILLER_200_2162 ();
 b15zdnd11an1n08x5 FILLER_200_2226 ();
 b15zdnd11an1n04x5 FILLER_200_2242 ();
 b15zdnd11an1n08x5 FILLER_200_2250 ();
 b15zdnd11an1n04x5 FILLER_200_2264 ();
 b15zdnd11an1n04x5 FILLER_200_2272 ();
 b15zdnd11an1n32x5 FILLER_201_0 ();
 b15zdnd11an1n16x5 FILLER_201_32 ();
 b15zdnd11an1n08x5 FILLER_201_48 ();
 b15zdnd00an1n02x5 FILLER_201_56 ();
 b15zdnd11an1n32x5 FILLER_201_66 ();
 b15zdnd11an1n04x5 FILLER_201_98 ();
 b15zdnd00an1n02x5 FILLER_201_102 ();
 b15zdnd11an1n04x5 FILLER_201_108 ();
 b15zdnd11an1n04x5 FILLER_201_127 ();
 b15zdnd11an1n04x5 FILLER_201_136 ();
 b15zdnd00an1n02x5 FILLER_201_140 ();
 b15zdnd00an1n01x5 FILLER_201_142 ();
 b15zdnd11an1n04x5 FILLER_201_158 ();
 b15zdnd11an1n08x5 FILLER_201_166 ();
 b15zdnd11an1n04x5 FILLER_201_174 ();
 b15zdnd11an1n16x5 FILLER_201_189 ();
 b15zdnd00an1n01x5 FILLER_201_205 ();
 b15zdnd11an1n04x5 FILLER_201_229 ();
 b15zdnd11an1n08x5 FILLER_201_253 ();
 b15zdnd11an1n04x5 FILLER_201_261 ();
 b15zdnd11an1n32x5 FILLER_201_281 ();
 b15zdnd11an1n04x5 FILLER_201_313 ();
 b15zdnd00an1n02x5 FILLER_201_317 ();
 b15zdnd00an1n01x5 FILLER_201_319 ();
 b15zdnd11an1n04x5 FILLER_201_341 ();
 b15zdnd11an1n04x5 FILLER_201_371 ();
 b15zdnd00an1n02x5 FILLER_201_375 ();
 b15zdnd00an1n01x5 FILLER_201_377 ();
 b15zdnd11an1n04x5 FILLER_201_386 ();
 b15zdnd00an1n02x5 FILLER_201_390 ();
 b15zdnd11an1n16x5 FILLER_201_417 ();
 b15zdnd11an1n16x5 FILLER_201_445 ();
 b15zdnd11an1n04x5 FILLER_201_473 ();
 b15zdnd11an1n16x5 FILLER_201_490 ();
 b15zdnd11an1n08x5 FILLER_201_506 ();
 b15zdnd11an1n04x5 FILLER_201_514 ();
 b15zdnd00an1n02x5 FILLER_201_518 ();
 b15zdnd00an1n01x5 FILLER_201_520 ();
 b15zdnd11an1n08x5 FILLER_201_533 ();
 b15zdnd11an1n04x5 FILLER_201_541 ();
 b15zdnd00an1n02x5 FILLER_201_545 ();
 b15zdnd11an1n16x5 FILLER_201_553 ();
 b15zdnd11an1n08x5 FILLER_201_569 ();
 b15zdnd11an1n04x5 FILLER_201_577 ();
 b15zdnd00an1n02x5 FILLER_201_581 ();
 b15zdnd00an1n01x5 FILLER_201_583 ();
 b15zdnd11an1n04x5 FILLER_201_592 ();
 b15zdnd00an1n01x5 FILLER_201_596 ();
 b15zdnd11an1n16x5 FILLER_201_603 ();
 b15zdnd11an1n04x5 FILLER_201_619 ();
 b15zdnd00an1n01x5 FILLER_201_623 ();
 b15zdnd11an1n08x5 FILLER_201_629 ();
 b15zdnd11an1n04x5 FILLER_201_637 ();
 b15zdnd00an1n02x5 FILLER_201_641 ();
 b15zdnd00an1n01x5 FILLER_201_643 ();
 b15zdnd11an1n04x5 FILLER_201_656 ();
 b15zdnd11an1n32x5 FILLER_201_671 ();
 b15zdnd11an1n04x5 FILLER_201_703 ();
 b15zdnd00an1n02x5 FILLER_201_707 ();
 b15zdnd11an1n16x5 FILLER_201_714 ();
 b15zdnd00an1n01x5 FILLER_201_730 ();
 b15zdnd11an1n04x5 FILLER_201_747 ();
 b15zdnd00an1n01x5 FILLER_201_751 ();
 b15zdnd11an1n04x5 FILLER_201_768 ();
 b15zdnd11an1n32x5 FILLER_201_786 ();
 b15zdnd11an1n16x5 FILLER_201_818 ();
 b15zdnd11an1n08x5 FILLER_201_834 ();
 b15zdnd00an1n01x5 FILLER_201_842 ();
 b15zdnd11an1n04x5 FILLER_201_852 ();
 b15zdnd00an1n02x5 FILLER_201_856 ();
 b15zdnd11an1n04x5 FILLER_201_862 ();
 b15zdnd11an1n32x5 FILLER_201_871 ();
 b15zdnd11an1n04x5 FILLER_201_903 ();
 b15zdnd00an1n02x5 FILLER_201_907 ();
 b15zdnd00an1n01x5 FILLER_201_909 ();
 b15zdnd11an1n08x5 FILLER_201_921 ();
 b15zdnd11an1n04x5 FILLER_201_934 ();
 b15zdnd11an1n08x5 FILLER_201_944 ();
 b15zdnd11an1n04x5 FILLER_201_952 ();
 b15zdnd00an1n01x5 FILLER_201_956 ();
 b15zdnd11an1n08x5 FILLER_201_974 ();
 b15zdnd11an1n04x5 FILLER_201_982 ();
 b15zdnd11an1n64x5 FILLER_201_990 ();
 b15zdnd00an1n02x5 FILLER_201_1054 ();
 b15zdnd11an1n08x5 FILLER_201_1070 ();
 b15zdnd00an1n02x5 FILLER_201_1078 ();
 b15zdnd11an1n64x5 FILLER_201_1088 ();
 b15zdnd11an1n16x5 FILLER_201_1152 ();
 b15zdnd11an1n16x5 FILLER_201_1182 ();
 b15zdnd11an1n08x5 FILLER_201_1198 ();
 b15zdnd11an1n04x5 FILLER_201_1206 ();
 b15zdnd00an1n02x5 FILLER_201_1210 ();
 b15zdnd11an1n16x5 FILLER_201_1219 ();
 b15zdnd00an1n02x5 FILLER_201_1235 ();
 b15zdnd00an1n01x5 FILLER_201_1237 ();
 b15zdnd11an1n16x5 FILLER_201_1264 ();
 b15zdnd11an1n08x5 FILLER_201_1280 ();
 b15zdnd00an1n01x5 FILLER_201_1288 ();
 b15zdnd11an1n04x5 FILLER_201_1299 ();
 b15zdnd11an1n64x5 FILLER_201_1312 ();
 b15zdnd11an1n32x5 FILLER_201_1388 ();
 b15zdnd11an1n16x5 FILLER_201_1420 ();
 b15zdnd11an1n04x5 FILLER_201_1436 ();
 b15zdnd11an1n16x5 FILLER_201_1453 ();
 b15zdnd11an1n04x5 FILLER_201_1469 ();
 b15zdnd00an1n02x5 FILLER_201_1473 ();
 b15zdnd11an1n64x5 FILLER_201_1481 ();
 b15zdnd00an1n01x5 FILLER_201_1545 ();
 b15zdnd11an1n16x5 FILLER_201_1551 ();
 b15zdnd11an1n08x5 FILLER_201_1567 ();
 b15zdnd11an1n04x5 FILLER_201_1575 ();
 b15zdnd11an1n64x5 FILLER_201_1595 ();
 b15zdnd11an1n64x5 FILLER_201_1659 ();
 b15zdnd11an1n64x5 FILLER_201_1723 ();
 b15zdnd11an1n64x5 FILLER_201_1787 ();
 b15zdnd11an1n16x5 FILLER_201_1851 ();
 b15zdnd11an1n08x5 FILLER_201_1867 ();
 b15zdnd00an1n02x5 FILLER_201_1875 ();
 b15zdnd11an1n64x5 FILLER_201_1882 ();
 b15zdnd11an1n32x5 FILLER_201_1946 ();
 b15zdnd11an1n04x5 FILLER_201_1978 ();
 b15zdnd11an1n64x5 FILLER_201_2002 ();
 b15zdnd11an1n16x5 FILLER_201_2066 ();
 b15zdnd11an1n08x5 FILLER_201_2082 ();
 b15zdnd11an1n04x5 FILLER_201_2090 ();
 b15zdnd00an1n01x5 FILLER_201_2094 ();
 b15zdnd11an1n16x5 FILLER_201_2115 ();
 b15zdnd00an1n02x5 FILLER_201_2131 ();
 b15zdnd11an1n64x5 FILLER_201_2142 ();
 b15zdnd11an1n32x5 FILLER_201_2206 ();
 b15zdnd11an1n16x5 FILLER_201_2238 ();
 b15zdnd11an1n08x5 FILLER_201_2254 ();
 b15zdnd11an1n08x5 FILLER_201_2266 ();
 b15zdnd00an1n02x5 FILLER_201_2274 ();
 b15zdnd00an1n01x5 FILLER_201_2276 ();
 b15zdnd00an1n02x5 FILLER_201_2281 ();
 b15zdnd00an1n01x5 FILLER_201_2283 ();
 b15zdnd11an1n64x5 FILLER_202_8 ();
 b15zdnd11an1n64x5 FILLER_202_72 ();
 b15zdnd11an1n08x5 FILLER_202_136 ();
 b15zdnd11an1n16x5 FILLER_202_154 ();
 b15zdnd11an1n08x5 FILLER_202_170 ();
 b15zdnd00an1n02x5 FILLER_202_178 ();
 b15zdnd11an1n08x5 FILLER_202_198 ();
 b15zdnd11an1n04x5 FILLER_202_206 ();
 b15zdnd11an1n16x5 FILLER_202_226 ();
 b15zdnd00an1n02x5 FILLER_202_242 ();
 b15zdnd00an1n01x5 FILLER_202_244 ();
 b15zdnd11an1n32x5 FILLER_202_249 ();
 b15zdnd11an1n16x5 FILLER_202_281 ();
 b15zdnd11an1n04x5 FILLER_202_297 ();
 b15zdnd00an1n02x5 FILLER_202_301 ();
 b15zdnd11an1n32x5 FILLER_202_329 ();
 b15zdnd11an1n16x5 FILLER_202_361 ();
 b15zdnd00an1n01x5 FILLER_202_377 ();
 b15zdnd11an1n16x5 FILLER_202_390 ();
 b15zdnd11an1n08x5 FILLER_202_406 ();
 b15zdnd00an1n01x5 FILLER_202_414 ();
 b15zdnd11an1n64x5 FILLER_202_426 ();
 b15zdnd11an1n32x5 FILLER_202_490 ();
 b15zdnd11an1n16x5 FILLER_202_522 ();
 b15zdnd11an1n04x5 FILLER_202_538 ();
 b15zdnd00an1n02x5 FILLER_202_542 ();
 b15zdnd11an1n16x5 FILLER_202_550 ();
 b15zdnd11an1n08x5 FILLER_202_566 ();
 b15zdnd11an1n04x5 FILLER_202_574 ();
 b15zdnd00an1n02x5 FILLER_202_578 ();
 b15zdnd11an1n04x5 FILLER_202_587 ();
 b15zdnd11an1n16x5 FILLER_202_596 ();
 b15zdnd00an1n02x5 FILLER_202_612 ();
 b15zdnd00an1n01x5 FILLER_202_614 ();
 b15zdnd11an1n04x5 FILLER_202_621 ();
 b15zdnd11an1n16x5 FILLER_202_632 ();
 b15zdnd11an1n08x5 FILLER_202_660 ();
 b15zdnd11an1n04x5 FILLER_202_668 ();
 b15zdnd00an1n02x5 FILLER_202_672 ();
 b15zdnd11an1n16x5 FILLER_202_679 ();
 b15zdnd11an1n08x5 FILLER_202_695 ();
 b15zdnd11an1n04x5 FILLER_202_703 ();
 b15zdnd00an1n02x5 FILLER_202_716 ();
 b15zdnd11an1n64x5 FILLER_202_726 ();
 b15zdnd11an1n32x5 FILLER_202_790 ();
 b15zdnd11an1n16x5 FILLER_202_822 ();
 b15zdnd11an1n16x5 FILLER_202_846 ();
 b15zdnd11an1n04x5 FILLER_202_878 ();
 b15zdnd11an1n64x5 FILLER_202_887 ();
 b15zdnd11an1n08x5 FILLER_202_951 ();
 b15zdnd11an1n04x5 FILLER_202_959 ();
 b15zdnd11an1n16x5 FILLER_202_967 ();
 b15zdnd00an1n01x5 FILLER_202_983 ();
 b15zdnd11an1n64x5 FILLER_202_990 ();
 b15zdnd11an1n32x5 FILLER_202_1054 ();
 b15zdnd11an1n16x5 FILLER_202_1086 ();
 b15zdnd00an1n02x5 FILLER_202_1102 ();
 b15zdnd00an1n01x5 FILLER_202_1104 ();
 b15zdnd11an1n32x5 FILLER_202_1114 ();
 b15zdnd00an1n01x5 FILLER_202_1146 ();
 b15zdnd11an1n32x5 FILLER_202_1151 ();
 b15zdnd11an1n08x5 FILLER_202_1183 ();
 b15zdnd11an1n64x5 FILLER_202_1201 ();
 b15zdnd11an1n16x5 FILLER_202_1265 ();
 b15zdnd11an1n04x5 FILLER_202_1281 ();
 b15zdnd00an1n01x5 FILLER_202_1285 ();
 b15zdnd11an1n08x5 FILLER_202_1299 ();
 b15zdnd00an1n01x5 FILLER_202_1307 ();
 b15zdnd11an1n32x5 FILLER_202_1318 ();
 b15zdnd11an1n16x5 FILLER_202_1350 ();
 b15zdnd00an1n02x5 FILLER_202_1366 ();
 b15zdnd11an1n08x5 FILLER_202_1377 ();
 b15zdnd11an1n16x5 FILLER_202_1392 ();
 b15zdnd11an1n08x5 FILLER_202_1408 ();
 b15zdnd11an1n32x5 FILLER_202_1421 ();
 b15zdnd11an1n08x5 FILLER_202_1453 ();
 b15zdnd00an1n02x5 FILLER_202_1461 ();
 b15zdnd00an1n01x5 FILLER_202_1463 ();
 b15zdnd11an1n08x5 FILLER_202_1469 ();
 b15zdnd11an1n64x5 FILLER_202_1481 ();
 b15zdnd11an1n32x5 FILLER_202_1545 ();
 b15zdnd11an1n16x5 FILLER_202_1577 ();
 b15zdnd11an1n08x5 FILLER_202_1593 ();
 b15zdnd11an1n04x5 FILLER_202_1601 ();
 b15zdnd00an1n02x5 FILLER_202_1605 ();
 b15zdnd11an1n08x5 FILLER_202_1614 ();
 b15zdnd00an1n02x5 FILLER_202_1622 ();
 b15zdnd11an1n04x5 FILLER_202_1630 ();
 b15zdnd11an1n04x5 FILLER_202_1646 ();
 b15zdnd11an1n08x5 FILLER_202_1655 ();
 b15zdnd11an1n04x5 FILLER_202_1663 ();
 b15zdnd00an1n02x5 FILLER_202_1667 ();
 b15zdnd11an1n64x5 FILLER_202_1684 ();
 b15zdnd11an1n64x5 FILLER_202_1748 ();
 b15zdnd11an1n08x5 FILLER_202_1812 ();
 b15zdnd11an1n16x5 FILLER_202_1851 ();
 b15zdnd11an1n08x5 FILLER_202_1867 ();
 b15zdnd11an1n04x5 FILLER_202_1895 ();
 b15zdnd11an1n16x5 FILLER_202_1917 ();
 b15zdnd11an1n08x5 FILLER_202_1933 ();
 b15zdnd00an1n02x5 FILLER_202_1941 ();
 b15zdnd00an1n01x5 FILLER_202_1943 ();
 b15zdnd11an1n32x5 FILLER_202_1964 ();
 b15zdnd11an1n16x5 FILLER_202_1996 ();
 b15zdnd11an1n08x5 FILLER_202_2012 ();
 b15zdnd11an1n04x5 FILLER_202_2020 ();
 b15zdnd00an1n01x5 FILLER_202_2024 ();
 b15zdnd11an1n04x5 FILLER_202_2034 ();
 b15zdnd11an1n64x5 FILLER_202_2047 ();
 b15zdnd11an1n32x5 FILLER_202_2111 ();
 b15zdnd11an1n08x5 FILLER_202_2143 ();
 b15zdnd00an1n02x5 FILLER_202_2151 ();
 b15zdnd00an1n01x5 FILLER_202_2153 ();
 b15zdnd11an1n04x5 FILLER_202_2162 ();
 b15zdnd00an1n02x5 FILLER_202_2166 ();
 b15zdnd11an1n64x5 FILLER_202_2173 ();
 b15zdnd11an1n08x5 FILLER_202_2237 ();
 b15zdnd11an1n04x5 FILLER_202_2245 ();
 b15zdnd00an1n02x5 FILLER_202_2249 ();
 b15zdnd00an1n01x5 FILLER_202_2251 ();
 b15zdnd11an1n16x5 FILLER_202_2257 ();
 b15zdnd00an1n02x5 FILLER_202_2273 ();
 b15zdnd00an1n01x5 FILLER_202_2275 ();
 b15zdnd11an1n08x5 FILLER_203_0 ();
 b15zdnd00an1n01x5 FILLER_203_8 ();
 b15zdnd11an1n64x5 FILLER_203_17 ();
 b15zdnd11an1n64x5 FILLER_203_81 ();
 b15zdnd11an1n64x5 FILLER_203_145 ();
 b15zdnd11an1n16x5 FILLER_203_209 ();
 b15zdnd11an1n08x5 FILLER_203_225 ();
 b15zdnd11an1n04x5 FILLER_203_233 ();
 b15zdnd00an1n01x5 FILLER_203_237 ();
 b15zdnd11an1n04x5 FILLER_203_243 ();
 b15zdnd11an1n64x5 FILLER_203_257 ();
 b15zdnd11an1n08x5 FILLER_203_321 ();
 b15zdnd00an1n02x5 FILLER_203_329 ();
 b15zdnd00an1n01x5 FILLER_203_331 ();
 b15zdnd11an1n64x5 FILLER_203_358 ();
 b15zdnd11an1n64x5 FILLER_203_422 ();
 b15zdnd11an1n32x5 FILLER_203_486 ();
 b15zdnd11an1n16x5 FILLER_203_518 ();
 b15zdnd11an1n08x5 FILLER_203_534 ();
 b15zdnd11an1n04x5 FILLER_203_542 ();
 b15zdnd11an1n32x5 FILLER_203_555 ();
 b15zdnd11an1n04x5 FILLER_203_587 ();
 b15zdnd11an1n64x5 FILLER_203_598 ();
 b15zdnd11an1n08x5 FILLER_203_662 ();
 b15zdnd00an1n02x5 FILLER_203_670 ();
 b15zdnd00an1n01x5 FILLER_203_672 ();
 b15zdnd11an1n16x5 FILLER_203_678 ();
 b15zdnd00an1n01x5 FILLER_203_694 ();
 b15zdnd11an1n64x5 FILLER_203_709 ();
 b15zdnd11an1n16x5 FILLER_203_773 ();
 b15zdnd11an1n08x5 FILLER_203_789 ();
 b15zdnd00an1n02x5 FILLER_203_797 ();
 b15zdnd11an1n16x5 FILLER_203_819 ();
 b15zdnd00an1n01x5 FILLER_203_835 ();
 b15zdnd11an1n08x5 FILLER_203_846 ();
 b15zdnd11an1n04x5 FILLER_203_854 ();
 b15zdnd00an1n01x5 FILLER_203_858 ();
 b15zdnd11an1n08x5 FILLER_203_865 ();
 b15zdnd11an1n04x5 FILLER_203_873 ();
 b15zdnd11an1n64x5 FILLER_203_883 ();
 b15zdnd11an1n32x5 FILLER_203_947 ();
 b15zdnd11an1n08x5 FILLER_203_979 ();
 b15zdnd00an1n02x5 FILLER_203_987 ();
 b15zdnd00an1n01x5 FILLER_203_989 ();
 b15zdnd11an1n64x5 FILLER_203_996 ();
 b15zdnd11an1n32x5 FILLER_203_1060 ();
 b15zdnd11an1n16x5 FILLER_203_1092 ();
 b15zdnd00an1n01x5 FILLER_203_1108 ();
 b15zdnd11an1n04x5 FILLER_203_1122 ();
 b15zdnd11an1n04x5 FILLER_203_1138 ();
 b15zdnd11an1n64x5 FILLER_203_1149 ();
 b15zdnd11an1n64x5 FILLER_203_1213 ();
 b15zdnd11an1n16x5 FILLER_203_1277 ();
 b15zdnd11an1n04x5 FILLER_203_1293 ();
 b15zdnd11an1n04x5 FILLER_203_1323 ();
 b15zdnd11an1n08x5 FILLER_203_1339 ();
 b15zdnd00an1n02x5 FILLER_203_1347 ();
 b15zdnd11an1n16x5 FILLER_203_1354 ();
 b15zdnd11an1n08x5 FILLER_203_1370 ();
 b15zdnd11an1n04x5 FILLER_203_1378 ();
 b15zdnd00an1n01x5 FILLER_203_1382 ();
 b15zdnd11an1n16x5 FILLER_203_1399 ();
 b15zdnd11an1n08x5 FILLER_203_1415 ();
 b15zdnd11an1n32x5 FILLER_203_1428 ();
 b15zdnd11an1n16x5 FILLER_203_1460 ();
 b15zdnd00an1n02x5 FILLER_203_1476 ();
 b15zdnd11an1n08x5 FILLER_203_1489 ();
 b15zdnd11an1n04x5 FILLER_203_1497 ();
 b15zdnd00an1n01x5 FILLER_203_1501 ();
 b15zdnd11an1n04x5 FILLER_203_1509 ();
 b15zdnd00an1n02x5 FILLER_203_1513 ();
 b15zdnd11an1n04x5 FILLER_203_1521 ();
 b15zdnd11an1n16x5 FILLER_203_1530 ();
 b15zdnd11an1n04x5 FILLER_203_1546 ();
 b15zdnd00an1n02x5 FILLER_203_1550 ();
 b15zdnd00an1n01x5 FILLER_203_1552 ();
 b15zdnd11an1n16x5 FILLER_203_1559 ();
 b15zdnd11an1n08x5 FILLER_203_1575 ();
 b15zdnd11an1n16x5 FILLER_203_1590 ();
 b15zdnd11an1n04x5 FILLER_203_1606 ();
 b15zdnd00an1n02x5 FILLER_203_1610 ();
 b15zdnd11an1n08x5 FILLER_203_1633 ();
 b15zdnd11an1n04x5 FILLER_203_1641 ();
 b15zdnd00an1n02x5 FILLER_203_1645 ();
 b15zdnd11an1n16x5 FILLER_203_1651 ();
 b15zdnd00an1n01x5 FILLER_203_1667 ();
 b15zdnd11an1n16x5 FILLER_203_1677 ();
 b15zdnd11an1n08x5 FILLER_203_1693 ();
 b15zdnd11an1n04x5 FILLER_203_1701 ();
 b15zdnd00an1n01x5 FILLER_203_1705 ();
 b15zdnd11an1n64x5 FILLER_203_1716 ();
 b15zdnd11an1n16x5 FILLER_203_1780 ();
 b15zdnd11an1n08x5 FILLER_203_1796 ();
 b15zdnd11an1n04x5 FILLER_203_1804 ();
 b15zdnd11an1n64x5 FILLER_203_1839 ();
 b15zdnd11an1n32x5 FILLER_203_1903 ();
 b15zdnd00an1n01x5 FILLER_203_1935 ();
 b15zdnd11an1n16x5 FILLER_203_1945 ();
 b15zdnd11an1n08x5 FILLER_203_1961 ();
 b15zdnd11an1n04x5 FILLER_203_1969 ();
 b15zdnd00an1n02x5 FILLER_203_1973 ();
 b15zdnd00an1n01x5 FILLER_203_1975 ();
 b15zdnd11an1n16x5 FILLER_203_1981 ();
 b15zdnd11an1n08x5 FILLER_203_1997 ();
 b15zdnd11an1n04x5 FILLER_203_2005 ();
 b15zdnd00an1n02x5 FILLER_203_2009 ();
 b15zdnd00an1n01x5 FILLER_203_2011 ();
 b15zdnd11an1n08x5 FILLER_203_2032 ();
 b15zdnd00an1n02x5 FILLER_203_2040 ();
 b15zdnd11an1n64x5 FILLER_203_2047 ();
 b15zdnd11an1n16x5 FILLER_203_2111 ();
 b15zdnd11an1n16x5 FILLER_203_2147 ();
 b15zdnd11an1n04x5 FILLER_203_2163 ();
 b15zdnd11an1n32x5 FILLER_203_2173 ();
 b15zdnd11an1n08x5 FILLER_203_2205 ();
 b15zdnd11an1n04x5 FILLER_203_2213 ();
 b15zdnd00an1n01x5 FILLER_203_2217 ();
 b15zdnd11an1n04x5 FILLER_203_2238 ();
 b15zdnd11an1n08x5 FILLER_203_2246 ();
 b15zdnd11an1n04x5 FILLER_203_2254 ();
 b15zdnd00an1n01x5 FILLER_203_2258 ();
 b15zdnd11an1n04x5 FILLER_203_2263 ();
 b15zdnd11an1n04x5 FILLER_203_2271 ();
 b15zdnd00an1n02x5 FILLER_203_2275 ();
 b15zdnd00an1n01x5 FILLER_203_2277 ();
 b15zdnd00an1n02x5 FILLER_203_2282 ();
 b15zdnd11an1n64x5 FILLER_204_8 ();
 b15zdnd11an1n64x5 FILLER_204_72 ();
 b15zdnd11an1n64x5 FILLER_204_136 ();
 b15zdnd11an1n32x5 FILLER_204_200 ();
 b15zdnd11an1n16x5 FILLER_204_232 ();
 b15zdnd11an1n04x5 FILLER_204_248 ();
 b15zdnd00an1n01x5 FILLER_204_252 ();
 b15zdnd11an1n64x5 FILLER_204_258 ();
 b15zdnd11an1n64x5 FILLER_204_322 ();
 b15zdnd11an1n64x5 FILLER_204_386 ();
 b15zdnd11an1n16x5 FILLER_204_450 ();
 b15zdnd11an1n08x5 FILLER_204_466 ();
 b15zdnd11an1n04x5 FILLER_204_474 ();
 b15zdnd11an1n16x5 FILLER_204_487 ();
 b15zdnd11an1n04x5 FILLER_204_503 ();
 b15zdnd00an1n02x5 FILLER_204_507 ();
 b15zdnd00an1n01x5 FILLER_204_509 ();
 b15zdnd11an1n08x5 FILLER_204_521 ();
 b15zdnd11an1n04x5 FILLER_204_529 ();
 b15zdnd00an1n02x5 FILLER_204_533 ();
 b15zdnd00an1n01x5 FILLER_204_535 ();
 b15zdnd11an1n64x5 FILLER_204_545 ();
 b15zdnd11an1n64x5 FILLER_204_609 ();
 b15zdnd11an1n16x5 FILLER_204_673 ();
 b15zdnd00an1n02x5 FILLER_204_689 ();
 b15zdnd11an1n16x5 FILLER_204_696 ();
 b15zdnd11an1n04x5 FILLER_204_712 ();
 b15zdnd00an1n02x5 FILLER_204_716 ();
 b15zdnd11an1n08x5 FILLER_204_726 ();
 b15zdnd11an1n04x5 FILLER_204_734 ();
 b15zdnd00an1n02x5 FILLER_204_738 ();
 b15zdnd00an1n01x5 FILLER_204_740 ();
 b15zdnd11an1n64x5 FILLER_204_755 ();
 b15zdnd11an1n16x5 FILLER_204_819 ();
 b15zdnd11an1n32x5 FILLER_204_840 ();
 b15zdnd11an1n08x5 FILLER_204_872 ();
 b15zdnd11an1n32x5 FILLER_204_887 ();
 b15zdnd11an1n16x5 FILLER_204_919 ();
 b15zdnd00an1n01x5 FILLER_204_935 ();
 b15zdnd11an1n16x5 FILLER_204_940 ();
 b15zdnd00an1n01x5 FILLER_204_956 ();
 b15zdnd11an1n32x5 FILLER_204_969 ();
 b15zdnd11an1n04x5 FILLER_204_1001 ();
 b15zdnd00an1n02x5 FILLER_204_1005 ();
 b15zdnd11an1n04x5 FILLER_204_1012 ();
 b15zdnd11an1n16x5 FILLER_204_1026 ();
 b15zdnd11an1n08x5 FILLER_204_1042 ();
 b15zdnd11an1n04x5 FILLER_204_1057 ();
 b15zdnd11an1n04x5 FILLER_204_1071 ();
 b15zdnd11an1n04x5 FILLER_204_1087 ();
 b15zdnd11an1n08x5 FILLER_204_1098 ();
 b15zdnd00an1n02x5 FILLER_204_1106 ();
 b15zdnd00an1n01x5 FILLER_204_1108 ();
 b15zdnd11an1n16x5 FILLER_204_1118 ();
 b15zdnd00an1n02x5 FILLER_204_1134 ();
 b15zdnd00an1n01x5 FILLER_204_1136 ();
 b15zdnd11an1n16x5 FILLER_204_1145 ();
 b15zdnd11an1n08x5 FILLER_204_1161 ();
 b15zdnd11an1n04x5 FILLER_204_1169 ();
 b15zdnd00an1n02x5 FILLER_204_1173 ();
 b15zdnd00an1n01x5 FILLER_204_1175 ();
 b15zdnd11an1n64x5 FILLER_204_1187 ();
 b15zdnd11an1n64x5 FILLER_204_1251 ();
 b15zdnd11an1n32x5 FILLER_204_1315 ();
 b15zdnd11an1n16x5 FILLER_204_1347 ();
 b15zdnd11an1n08x5 FILLER_204_1363 ();
 b15zdnd11an1n04x5 FILLER_204_1371 ();
 b15zdnd00an1n02x5 FILLER_204_1375 ();
 b15zdnd00an1n01x5 FILLER_204_1377 ();
 b15zdnd11an1n04x5 FILLER_204_1391 ();
 b15zdnd11an1n16x5 FILLER_204_1400 ();
 b15zdnd00an1n01x5 FILLER_204_1416 ();
 b15zdnd11an1n16x5 FILLER_204_1433 ();
 b15zdnd00an1n02x5 FILLER_204_1449 ();
 b15zdnd00an1n01x5 FILLER_204_1451 ();
 b15zdnd11an1n16x5 FILLER_204_1459 ();
 b15zdnd11an1n08x5 FILLER_204_1475 ();
 b15zdnd00an1n01x5 FILLER_204_1483 ();
 b15zdnd11an1n32x5 FILLER_204_1490 ();
 b15zdnd11an1n16x5 FILLER_204_1522 ();
 b15zdnd11an1n08x5 FILLER_204_1538 ();
 b15zdnd11an1n04x5 FILLER_204_1546 ();
 b15zdnd00an1n02x5 FILLER_204_1550 ();
 b15zdnd00an1n01x5 FILLER_204_1552 ();
 b15zdnd11an1n16x5 FILLER_204_1562 ();
 b15zdnd11an1n08x5 FILLER_204_1578 ();
 b15zdnd00an1n01x5 FILLER_204_1586 ();
 b15zdnd11an1n04x5 FILLER_204_1594 ();
 b15zdnd11an1n04x5 FILLER_204_1605 ();
 b15zdnd00an1n02x5 FILLER_204_1609 ();
 b15zdnd00an1n01x5 FILLER_204_1611 ();
 b15zdnd11an1n08x5 FILLER_204_1638 ();
 b15zdnd00an1n01x5 FILLER_204_1646 ();
 b15zdnd11an1n04x5 FILLER_204_1660 ();
 b15zdnd11an1n32x5 FILLER_204_1684 ();
 b15zdnd11an1n16x5 FILLER_204_1716 ();
 b15zdnd11an1n04x5 FILLER_204_1732 ();
 b15zdnd00an1n01x5 FILLER_204_1736 ();
 b15zdnd11an1n04x5 FILLER_204_1768 ();
 b15zdnd11an1n64x5 FILLER_204_1803 ();
 b15zdnd11an1n64x5 FILLER_204_1867 ();
 b15zdnd11an1n16x5 FILLER_204_1931 ();
 b15zdnd11an1n08x5 FILLER_204_1947 ();
 b15zdnd11an1n04x5 FILLER_204_1955 ();
 b15zdnd00an1n02x5 FILLER_204_1959 ();
 b15zdnd00an1n01x5 FILLER_204_1961 ();
 b15zdnd11an1n64x5 FILLER_204_1982 ();
 b15zdnd11an1n64x5 FILLER_204_2046 ();
 b15zdnd11an1n16x5 FILLER_204_2110 ();
 b15zdnd11an1n08x5 FILLER_204_2126 ();
 b15zdnd11an1n08x5 FILLER_204_2139 ();
 b15zdnd11an1n04x5 FILLER_204_2147 ();
 b15zdnd00an1n02x5 FILLER_204_2151 ();
 b15zdnd00an1n01x5 FILLER_204_2153 ();
 b15zdnd00an1n02x5 FILLER_204_2162 ();
 b15zdnd11an1n04x5 FILLER_204_2184 ();
 b15zdnd00an1n02x5 FILLER_204_2188 ();
 b15zdnd11an1n04x5 FILLER_204_2201 ();
 b15zdnd11an1n32x5 FILLER_204_2216 ();
 b15zdnd11an1n04x5 FILLER_204_2248 ();
 b15zdnd11an1n04x5 FILLER_204_2256 ();
 b15zdnd00an1n02x5 FILLER_204_2260 ();
 b15zdnd11an1n04x5 FILLER_204_2265 ();
 b15zdnd00an1n01x5 FILLER_204_2269 ();
 b15zdnd00an1n02x5 FILLER_204_2274 ();
 b15zdnd00an1n02x5 FILLER_205_0 ();
 b15zdnd11an1n64x5 FILLER_205_6 ();
 b15zdnd11an1n64x5 FILLER_205_70 ();
 b15zdnd11an1n64x5 FILLER_205_134 ();
 b15zdnd11an1n64x5 FILLER_205_198 ();
 b15zdnd11an1n64x5 FILLER_205_262 ();
 b15zdnd11an1n32x5 FILLER_205_326 ();
 b15zdnd11an1n08x5 FILLER_205_358 ();
 b15zdnd11an1n04x5 FILLER_205_366 ();
 b15zdnd00an1n02x5 FILLER_205_370 ();
 b15zdnd00an1n01x5 FILLER_205_372 ();
 b15zdnd11an1n64x5 FILLER_205_405 ();
 b15zdnd00an1n01x5 FILLER_205_469 ();
 b15zdnd11an1n04x5 FILLER_205_475 ();
 b15zdnd11an1n04x5 FILLER_205_493 ();
 b15zdnd11an1n08x5 FILLER_205_505 ();
 b15zdnd11an1n04x5 FILLER_205_513 ();
 b15zdnd11an1n08x5 FILLER_205_524 ();
 b15zdnd11an1n04x5 FILLER_205_532 ();
 b15zdnd11an1n64x5 FILLER_205_552 ();
 b15zdnd11an1n64x5 FILLER_205_616 ();
 b15zdnd11an1n16x5 FILLER_205_680 ();
 b15zdnd11an1n08x5 FILLER_205_696 ();
 b15zdnd00an1n02x5 FILLER_205_704 ();
 b15zdnd00an1n01x5 FILLER_205_706 ();
 b15zdnd11an1n08x5 FILLER_205_712 ();
 b15zdnd11an1n04x5 FILLER_205_720 ();
 b15zdnd00an1n01x5 FILLER_205_724 ();
 b15zdnd11an1n64x5 FILLER_205_744 ();
 b15zdnd11an1n16x5 FILLER_205_808 ();
 b15zdnd11an1n04x5 FILLER_205_824 ();
 b15zdnd00an1n02x5 FILLER_205_828 ();
 b15zdnd11an1n16x5 FILLER_205_850 ();
 b15zdnd11an1n04x5 FILLER_205_866 ();
 b15zdnd00an1n02x5 FILLER_205_870 ();
 b15zdnd11an1n04x5 FILLER_205_877 ();
 b15zdnd11an1n08x5 FILLER_205_890 ();
 b15zdnd00an1n01x5 FILLER_205_898 ();
 b15zdnd11an1n08x5 FILLER_205_903 ();
 b15zdnd11an1n04x5 FILLER_205_911 ();
 b15zdnd00an1n02x5 FILLER_205_915 ();
 b15zdnd00an1n01x5 FILLER_205_917 ();
 b15zdnd11an1n08x5 FILLER_205_922 ();
 b15zdnd00an1n02x5 FILLER_205_930 ();
 b15zdnd00an1n01x5 FILLER_205_932 ();
 b15zdnd11an1n32x5 FILLER_205_938 ();
 b15zdnd11an1n08x5 FILLER_205_970 ();
 b15zdnd11an1n16x5 FILLER_205_985 ();
 b15zdnd11an1n08x5 FILLER_205_1001 ();
 b15zdnd11an1n04x5 FILLER_205_1009 ();
 b15zdnd00an1n02x5 FILLER_205_1013 ();
 b15zdnd11an1n08x5 FILLER_205_1031 ();
 b15zdnd00an1n02x5 FILLER_205_1039 ();
 b15zdnd11an1n32x5 FILLER_205_1054 ();
 b15zdnd11an1n16x5 FILLER_205_1086 ();
 b15zdnd11an1n04x5 FILLER_205_1102 ();
 b15zdnd00an1n02x5 FILLER_205_1106 ();
 b15zdnd11an1n32x5 FILLER_205_1114 ();
 b15zdnd11an1n16x5 FILLER_205_1146 ();
 b15zdnd00an1n02x5 FILLER_205_1162 ();
 b15zdnd11an1n64x5 FILLER_205_1174 ();
 b15zdnd11an1n64x5 FILLER_205_1238 ();
 b15zdnd11an1n08x5 FILLER_205_1302 ();
 b15zdnd11an1n04x5 FILLER_205_1310 ();
 b15zdnd11an1n16x5 FILLER_205_1323 ();
 b15zdnd11an1n16x5 FILLER_205_1351 ();
 b15zdnd11an1n08x5 FILLER_205_1367 ();
 b15zdnd11an1n04x5 FILLER_205_1375 ();
 b15zdnd11an1n64x5 FILLER_205_1391 ();
 b15zdnd11an1n32x5 FILLER_205_1455 ();
 b15zdnd00an1n01x5 FILLER_205_1487 ();
 b15zdnd11an1n08x5 FILLER_205_1494 ();
 b15zdnd00an1n01x5 FILLER_205_1502 ();
 b15zdnd11an1n08x5 FILLER_205_1508 ();
 b15zdnd11an1n16x5 FILLER_205_1521 ();
 b15zdnd11an1n08x5 FILLER_205_1537 ();
 b15zdnd11an1n04x5 FILLER_205_1545 ();
 b15zdnd00an1n01x5 FILLER_205_1549 ();
 b15zdnd11an1n16x5 FILLER_205_1555 ();
 b15zdnd11an1n08x5 FILLER_205_1571 ();
 b15zdnd11an1n04x5 FILLER_205_1579 ();
 b15zdnd00an1n02x5 FILLER_205_1583 ();
 b15zdnd11an1n64x5 FILLER_205_1593 ();
 b15zdnd11an1n08x5 FILLER_205_1657 ();
 b15zdnd00an1n02x5 FILLER_205_1665 ();
 b15zdnd11an1n32x5 FILLER_205_1683 ();
 b15zdnd11an1n08x5 FILLER_205_1715 ();
 b15zdnd00an1n01x5 FILLER_205_1723 ();
 b15zdnd11an1n04x5 FILLER_205_1742 ();
 b15zdnd11an1n64x5 FILLER_205_1758 ();
 b15zdnd11an1n32x5 FILLER_205_1822 ();
 b15zdnd11an1n04x5 FILLER_205_1854 ();
 b15zdnd00an1n02x5 FILLER_205_1858 ();
 b15zdnd11an1n64x5 FILLER_205_1875 ();
 b15zdnd11an1n32x5 FILLER_205_1939 ();
 b15zdnd00an1n02x5 FILLER_205_1971 ();
 b15zdnd11an1n64x5 FILLER_205_1982 ();
 b15zdnd11an1n08x5 FILLER_205_2046 ();
 b15zdnd11an1n04x5 FILLER_205_2054 ();
 b15zdnd00an1n02x5 FILLER_205_2058 ();
 b15zdnd11an1n08x5 FILLER_205_2080 ();
 b15zdnd11an1n04x5 FILLER_205_2088 ();
 b15zdnd00an1n02x5 FILLER_205_2092 ();
 b15zdnd00an1n01x5 FILLER_205_2094 ();
 b15zdnd11an1n16x5 FILLER_205_2100 ();
 b15zdnd11an1n08x5 FILLER_205_2116 ();
 b15zdnd11an1n04x5 FILLER_205_2124 ();
 b15zdnd00an1n01x5 FILLER_205_2128 ();
 b15zdnd11an1n64x5 FILLER_205_2138 ();
 b15zdnd00an1n02x5 FILLER_205_2202 ();
 b15zdnd00an1n01x5 FILLER_205_2204 ();
 b15zdnd11an1n16x5 FILLER_205_2225 ();
 b15zdnd11an1n08x5 FILLER_205_2241 ();
 b15zdnd11an1n04x5 FILLER_205_2249 ();
 b15zdnd00an1n02x5 FILLER_205_2253 ();
 b15zdnd00an1n01x5 FILLER_205_2255 ();
 b15zdnd11an1n04x5 FILLER_205_2261 ();
 b15zdnd11an1n08x5 FILLER_205_2269 ();
 b15zdnd00an1n02x5 FILLER_205_2282 ();
 b15zdnd11an1n16x5 FILLER_206_8 ();
 b15zdnd11an1n08x5 FILLER_206_24 ();
 b15zdnd11an1n04x5 FILLER_206_32 ();
 b15zdnd00an1n02x5 FILLER_206_36 ();
 b15zdnd11an1n64x5 FILLER_206_45 ();
 b15zdnd11an1n64x5 FILLER_206_109 ();
 b15zdnd11an1n64x5 FILLER_206_173 ();
 b15zdnd11an1n64x5 FILLER_206_237 ();
 b15zdnd11an1n64x5 FILLER_206_301 ();
 b15zdnd11an1n08x5 FILLER_206_365 ();
 b15zdnd11an1n08x5 FILLER_206_383 ();
 b15zdnd11an1n04x5 FILLER_206_391 ();
 b15zdnd00an1n01x5 FILLER_206_395 ();
 b15zdnd11an1n04x5 FILLER_206_403 ();
 b15zdnd11an1n08x5 FILLER_206_411 ();
 b15zdnd11an1n04x5 FILLER_206_419 ();
 b15zdnd11an1n04x5 FILLER_206_428 ();
 b15zdnd11an1n16x5 FILLER_206_438 ();
 b15zdnd11an1n08x5 FILLER_206_454 ();
 b15zdnd11an1n04x5 FILLER_206_462 ();
 b15zdnd00an1n02x5 FILLER_206_466 ();
 b15zdnd00an1n01x5 FILLER_206_468 ();
 b15zdnd11an1n04x5 FILLER_206_475 ();
 b15zdnd00an1n01x5 FILLER_206_479 ();
 b15zdnd11an1n32x5 FILLER_206_488 ();
 b15zdnd11an1n16x5 FILLER_206_520 ();
 b15zdnd11an1n08x5 FILLER_206_536 ();
 b15zdnd00an1n02x5 FILLER_206_544 ();
 b15zdnd00an1n01x5 FILLER_206_546 ();
 b15zdnd11an1n04x5 FILLER_206_553 ();
 b15zdnd00an1n02x5 FILLER_206_557 ();
 b15zdnd00an1n01x5 FILLER_206_559 ();
 b15zdnd11an1n04x5 FILLER_206_572 ();
 b15zdnd11an1n08x5 FILLER_206_588 ();
 b15zdnd11an1n04x5 FILLER_206_596 ();
 b15zdnd11an1n08x5 FILLER_206_605 ();
 b15zdnd11an1n32x5 FILLER_206_630 ();
 b15zdnd00an1n01x5 FILLER_206_662 ();
 b15zdnd11an1n04x5 FILLER_206_671 ();
 b15zdnd11an1n04x5 FILLER_206_679 ();
 b15zdnd00an1n02x5 FILLER_206_683 ();
 b15zdnd00an1n01x5 FILLER_206_685 ();
 b15zdnd11an1n16x5 FILLER_206_700 ();
 b15zdnd00an1n02x5 FILLER_206_716 ();
 b15zdnd11an1n08x5 FILLER_206_726 ();
 b15zdnd11an1n04x5 FILLER_206_734 ();
 b15zdnd11an1n64x5 FILLER_206_748 ();
 b15zdnd11an1n32x5 FILLER_206_812 ();
 b15zdnd00an1n02x5 FILLER_206_844 ();
 b15zdnd11an1n04x5 FILLER_206_852 ();
 b15zdnd11an1n32x5 FILLER_206_868 ();
 b15zdnd11an1n16x5 FILLER_206_900 ();
 b15zdnd11an1n32x5 FILLER_206_928 ();
 b15zdnd11an1n16x5 FILLER_206_960 ();
 b15zdnd11an1n04x5 FILLER_206_976 ();
 b15zdnd11an1n04x5 FILLER_206_985 ();
 b15zdnd11an1n08x5 FILLER_206_998 ();
 b15zdnd11an1n16x5 FILLER_206_1012 ();
 b15zdnd11an1n04x5 FILLER_206_1028 ();
 b15zdnd00an1n02x5 FILLER_206_1032 ();
 b15zdnd11an1n64x5 FILLER_206_1048 ();
 b15zdnd11an1n32x5 FILLER_206_1112 ();
 b15zdnd11an1n08x5 FILLER_206_1144 ();
 b15zdnd11an1n04x5 FILLER_206_1159 ();
 b15zdnd11an1n08x5 FILLER_206_1187 ();
 b15zdnd00an1n02x5 FILLER_206_1195 ();
 b15zdnd00an1n01x5 FILLER_206_1197 ();
 b15zdnd11an1n64x5 FILLER_206_1207 ();
 b15zdnd11an1n16x5 FILLER_206_1271 ();
 b15zdnd00an1n01x5 FILLER_206_1287 ();
 b15zdnd11an1n16x5 FILLER_206_1298 ();
 b15zdnd11an1n04x5 FILLER_206_1314 ();
 b15zdnd00an1n01x5 FILLER_206_1318 ();
 b15zdnd11an1n04x5 FILLER_206_1323 ();
 b15zdnd00an1n01x5 FILLER_206_1327 ();
 b15zdnd11an1n04x5 FILLER_206_1339 ();
 b15zdnd11an1n64x5 FILLER_206_1352 ();
 b15zdnd11an1n32x5 FILLER_206_1430 ();
 b15zdnd11an1n16x5 FILLER_206_1466 ();
 b15zdnd00an1n02x5 FILLER_206_1482 ();
 b15zdnd00an1n01x5 FILLER_206_1484 ();
 b15zdnd11an1n32x5 FILLER_206_1492 ();
 b15zdnd11an1n16x5 FILLER_206_1524 ();
 b15zdnd11an1n08x5 FILLER_206_1540 ();
 b15zdnd00an1n02x5 FILLER_206_1548 ();
 b15zdnd00an1n01x5 FILLER_206_1550 ();
 b15zdnd11an1n16x5 FILLER_206_1557 ();
 b15zdnd11an1n04x5 FILLER_206_1573 ();
 b15zdnd00an1n01x5 FILLER_206_1577 ();
 b15zdnd11an1n64x5 FILLER_206_1585 ();
 b15zdnd11an1n16x5 FILLER_206_1649 ();
 b15zdnd11an1n08x5 FILLER_206_1665 ();
 b15zdnd11an1n04x5 FILLER_206_1673 ();
 b15zdnd11an1n64x5 FILLER_206_1686 ();
 b15zdnd11an1n32x5 FILLER_206_1750 ();
 b15zdnd11an1n16x5 FILLER_206_1782 ();
 b15zdnd11an1n08x5 FILLER_206_1798 ();
 b15zdnd00an1n02x5 FILLER_206_1806 ();
 b15zdnd00an1n01x5 FILLER_206_1808 ();
 b15zdnd11an1n16x5 FILLER_206_1833 ();
 b15zdnd11an1n08x5 FILLER_206_1849 ();
 b15zdnd00an1n02x5 FILLER_206_1857 ();
 b15zdnd00an1n01x5 FILLER_206_1859 ();
 b15zdnd11an1n64x5 FILLER_206_1871 ();
 b15zdnd11an1n64x5 FILLER_206_1935 ();
 b15zdnd11an1n64x5 FILLER_206_1999 ();
 b15zdnd11an1n32x5 FILLER_206_2063 ();
 b15zdnd00an1n01x5 FILLER_206_2095 ();
 b15zdnd11an1n32x5 FILLER_206_2100 ();
 b15zdnd11an1n16x5 FILLER_206_2132 ();
 b15zdnd11an1n04x5 FILLER_206_2148 ();
 b15zdnd00an1n02x5 FILLER_206_2152 ();
 b15zdnd11an1n64x5 FILLER_206_2162 ();
 b15zdnd11an1n32x5 FILLER_206_2226 ();
 b15zdnd11an1n16x5 FILLER_206_2258 ();
 b15zdnd00an1n02x5 FILLER_206_2274 ();
 b15zdnd11an1n16x5 FILLER_207_0 ();
 b15zdnd00an1n02x5 FILLER_207_16 ();
 b15zdnd00an1n01x5 FILLER_207_18 ();
 b15zdnd11an1n64x5 FILLER_207_23 ();
 b15zdnd11an1n64x5 FILLER_207_87 ();
 b15zdnd11an1n64x5 FILLER_207_151 ();
 b15zdnd11an1n64x5 FILLER_207_215 ();
 b15zdnd11an1n64x5 FILLER_207_279 ();
 b15zdnd11an1n32x5 FILLER_207_343 ();
 b15zdnd11an1n16x5 FILLER_207_375 ();
 b15zdnd11an1n08x5 FILLER_207_391 ();
 b15zdnd00an1n02x5 FILLER_207_399 ();
 b15zdnd11an1n16x5 FILLER_207_408 ();
 b15zdnd11an1n16x5 FILLER_207_439 ();
 b15zdnd00an1n02x5 FILLER_207_455 ();
 b15zdnd11an1n64x5 FILLER_207_469 ();
 b15zdnd11an1n08x5 FILLER_207_533 ();
 b15zdnd11an1n04x5 FILLER_207_541 ();
 b15zdnd00an1n02x5 FILLER_207_545 ();
 b15zdnd11an1n08x5 FILLER_207_553 ();
 b15zdnd11an1n04x5 FILLER_207_561 ();
 b15zdnd00an1n02x5 FILLER_207_565 ();
 b15zdnd11an1n16x5 FILLER_207_572 ();
 b15zdnd11an1n04x5 FILLER_207_588 ();
 b15zdnd11an1n04x5 FILLER_207_600 ();
 b15zdnd11an1n32x5 FILLER_207_616 ();
 b15zdnd11an1n16x5 FILLER_207_648 ();
 b15zdnd11an1n04x5 FILLER_207_664 ();
 b15zdnd00an1n02x5 FILLER_207_668 ();
 b15zdnd11an1n32x5 FILLER_207_682 ();
 b15zdnd11an1n16x5 FILLER_207_714 ();
 b15zdnd11an1n08x5 FILLER_207_730 ();
 b15zdnd11an1n04x5 FILLER_207_738 ();
 b15zdnd11an1n32x5 FILLER_207_746 ();
 b15zdnd11an1n16x5 FILLER_207_778 ();
 b15zdnd11an1n08x5 FILLER_207_794 ();
 b15zdnd00an1n01x5 FILLER_207_802 ();
 b15zdnd11an1n32x5 FILLER_207_823 ();
 b15zdnd11an1n08x5 FILLER_207_855 ();
 b15zdnd00an1n02x5 FILLER_207_863 ();
 b15zdnd00an1n01x5 FILLER_207_865 ();
 b15zdnd11an1n32x5 FILLER_207_882 ();
 b15zdnd11an1n04x5 FILLER_207_914 ();
 b15zdnd00an1n02x5 FILLER_207_918 ();
 b15zdnd00an1n01x5 FILLER_207_920 ();
 b15zdnd11an1n04x5 FILLER_207_928 ();
 b15zdnd00an1n02x5 FILLER_207_932 ();
 b15zdnd00an1n01x5 FILLER_207_934 ();
 b15zdnd11an1n16x5 FILLER_207_951 ();
 b15zdnd11an1n08x5 FILLER_207_967 ();
 b15zdnd11an1n08x5 FILLER_207_985 ();
 b15zdnd11an1n04x5 FILLER_207_993 ();
 b15zdnd00an1n02x5 FILLER_207_997 ();
 b15zdnd11an1n08x5 FILLER_207_1005 ();
 b15zdnd11an1n04x5 FILLER_207_1013 ();
 b15zdnd00an1n01x5 FILLER_207_1017 ();
 b15zdnd11an1n64x5 FILLER_207_1023 ();
 b15zdnd11an1n32x5 FILLER_207_1087 ();
 b15zdnd00an1n01x5 FILLER_207_1119 ();
 b15zdnd11an1n04x5 FILLER_207_1126 ();
 b15zdnd00an1n02x5 FILLER_207_1130 ();
 b15zdnd11an1n08x5 FILLER_207_1138 ();
 b15zdnd11an1n04x5 FILLER_207_1146 ();
 b15zdnd00an1n02x5 FILLER_207_1150 ();
 b15zdnd11an1n32x5 FILLER_207_1160 ();
 b15zdnd11an1n04x5 FILLER_207_1192 ();
 b15zdnd00an1n02x5 FILLER_207_1196 ();
 b15zdnd00an1n01x5 FILLER_207_1198 ();
 b15zdnd11an1n04x5 FILLER_207_1204 ();
 b15zdnd11an1n64x5 FILLER_207_1214 ();
 b15zdnd11an1n08x5 FILLER_207_1278 ();
 b15zdnd00an1n02x5 FILLER_207_1286 ();
 b15zdnd11an1n64x5 FILLER_207_1295 ();
 b15zdnd11an1n04x5 FILLER_207_1359 ();
 b15zdnd00an1n01x5 FILLER_207_1363 ();
 b15zdnd11an1n04x5 FILLER_207_1374 ();
 b15zdnd11an1n04x5 FILLER_207_1398 ();
 b15zdnd11an1n64x5 FILLER_207_1414 ();
 b15zdnd11an1n64x5 FILLER_207_1478 ();
 b15zdnd11an1n08x5 FILLER_207_1542 ();
 b15zdnd11an1n04x5 FILLER_207_1550 ();
 b15zdnd00an1n02x5 FILLER_207_1554 ();
 b15zdnd00an1n01x5 FILLER_207_1556 ();
 b15zdnd11an1n16x5 FILLER_207_1567 ();
 b15zdnd11an1n08x5 FILLER_207_1583 ();
 b15zdnd11an1n64x5 FILLER_207_1596 ();
 b15zdnd00an1n02x5 FILLER_207_1660 ();
 b15zdnd00an1n01x5 FILLER_207_1662 ();
 b15zdnd11an1n64x5 FILLER_207_1669 ();
 b15zdnd11an1n32x5 FILLER_207_1733 ();
 b15zdnd11an1n08x5 FILLER_207_1765 ();
 b15zdnd00an1n02x5 FILLER_207_1773 ();
 b15zdnd11an1n08x5 FILLER_207_1785 ();
 b15zdnd00an1n01x5 FILLER_207_1793 ();
 b15zdnd11an1n64x5 FILLER_207_1812 ();
 b15zdnd11an1n64x5 FILLER_207_1876 ();
 b15zdnd11an1n32x5 FILLER_207_1940 ();
 b15zdnd11an1n16x5 FILLER_207_1972 ();
 b15zdnd00an1n01x5 FILLER_207_1988 ();
 b15zdnd11an1n64x5 FILLER_207_1993 ();
 b15zdnd11an1n32x5 FILLER_207_2057 ();
 b15zdnd11an1n08x5 FILLER_207_2089 ();
 b15zdnd11an1n04x5 FILLER_207_2097 ();
 b15zdnd11an1n16x5 FILLER_207_2105 ();
 b15zdnd11an1n04x5 FILLER_207_2121 ();
 b15zdnd11an1n64x5 FILLER_207_2129 ();
 b15zdnd11an1n64x5 FILLER_207_2193 ();
 b15zdnd11an1n16x5 FILLER_207_2257 ();
 b15zdnd11an1n08x5 FILLER_207_2273 ();
 b15zdnd00an1n02x5 FILLER_207_2281 ();
 b15zdnd00an1n01x5 FILLER_207_2283 ();
 b15zdnd11an1n64x5 FILLER_208_8 ();
 b15zdnd11an1n64x5 FILLER_208_72 ();
 b15zdnd11an1n64x5 FILLER_208_136 ();
 b15zdnd11an1n64x5 FILLER_208_200 ();
 b15zdnd11an1n64x5 FILLER_208_264 ();
 b15zdnd11an1n32x5 FILLER_208_328 ();
 b15zdnd11an1n08x5 FILLER_208_360 ();
 b15zdnd11an1n04x5 FILLER_208_368 ();
 b15zdnd00an1n01x5 FILLER_208_372 ();
 b15zdnd11an1n16x5 FILLER_208_385 ();
 b15zdnd11an1n08x5 FILLER_208_411 ();
 b15zdnd00an1n02x5 FILLER_208_419 ();
 b15zdnd11an1n32x5 FILLER_208_428 ();
 b15zdnd11an1n08x5 FILLER_208_460 ();
 b15zdnd11an1n04x5 FILLER_208_468 ();
 b15zdnd11an1n04x5 FILLER_208_484 ();
 b15zdnd11an1n04x5 FILLER_208_495 ();
 b15zdnd11an1n64x5 FILLER_208_504 ();
 b15zdnd11an1n16x5 FILLER_208_568 ();
 b15zdnd11an1n08x5 FILLER_208_584 ();
 b15zdnd00an1n02x5 FILLER_208_592 ();
 b15zdnd00an1n01x5 FILLER_208_594 ();
 b15zdnd11an1n16x5 FILLER_208_603 ();
 b15zdnd11an1n04x5 FILLER_208_619 ();
 b15zdnd00an1n02x5 FILLER_208_623 ();
 b15zdnd11an1n04x5 FILLER_208_641 ();
 b15zdnd11an1n04x5 FILLER_208_676 ();
 b15zdnd11an1n32x5 FILLER_208_684 ();
 b15zdnd00an1n02x5 FILLER_208_716 ();
 b15zdnd11an1n64x5 FILLER_208_726 ();
 b15zdnd11an1n32x5 FILLER_208_790 ();
 b15zdnd11an1n16x5 FILLER_208_822 ();
 b15zdnd11an1n08x5 FILLER_208_838 ();
 b15zdnd00an1n01x5 FILLER_208_846 ();
 b15zdnd11an1n16x5 FILLER_208_857 ();
 b15zdnd11an1n04x5 FILLER_208_873 ();
 b15zdnd11an1n32x5 FILLER_208_889 ();
 b15zdnd00an1n01x5 FILLER_208_921 ();
 b15zdnd11an1n64x5 FILLER_208_930 ();
 b15zdnd11an1n32x5 FILLER_208_994 ();
 b15zdnd11an1n16x5 FILLER_208_1026 ();
 b15zdnd11an1n08x5 FILLER_208_1042 ();
 b15zdnd11an1n64x5 FILLER_208_1066 ();
 b15zdnd11an1n64x5 FILLER_208_1130 ();
 b15zdnd11an1n64x5 FILLER_208_1194 ();
 b15zdnd11an1n64x5 FILLER_208_1258 ();
 b15zdnd00an1n01x5 FILLER_208_1322 ();
 b15zdnd11an1n04x5 FILLER_208_1336 ();
 b15zdnd11an1n16x5 FILLER_208_1357 ();
 b15zdnd11an1n04x5 FILLER_208_1373 ();
 b15zdnd00an1n02x5 FILLER_208_1377 ();
 b15zdnd11an1n32x5 FILLER_208_1387 ();
 b15zdnd11an1n04x5 FILLER_208_1419 ();
 b15zdnd00an1n02x5 FILLER_208_1423 ();
 b15zdnd00an1n01x5 FILLER_208_1425 ();
 b15zdnd11an1n04x5 FILLER_208_1440 ();
 b15zdnd11an1n32x5 FILLER_208_1449 ();
 b15zdnd00an1n02x5 FILLER_208_1481 ();
 b15zdnd00an1n01x5 FILLER_208_1483 ();
 b15zdnd11an1n64x5 FILLER_208_1495 ();
 b15zdnd11an1n16x5 FILLER_208_1559 ();
 b15zdnd11an1n08x5 FILLER_208_1575 ();
 b15zdnd00an1n02x5 FILLER_208_1583 ();
 b15zdnd11an1n32x5 FILLER_208_1594 ();
 b15zdnd11an1n04x5 FILLER_208_1631 ();
 b15zdnd11an1n08x5 FILLER_208_1647 ();
 b15zdnd11an1n04x5 FILLER_208_1655 ();
 b15zdnd00an1n02x5 FILLER_208_1659 ();
 b15zdnd00an1n01x5 FILLER_208_1661 ();
 b15zdnd11an1n64x5 FILLER_208_1672 ();
 b15zdnd00an1n02x5 FILLER_208_1736 ();
 b15zdnd11an1n04x5 FILLER_208_1769 ();
 b15zdnd11an1n08x5 FILLER_208_1798 ();
 b15zdnd11an1n04x5 FILLER_208_1806 ();
 b15zdnd00an1n01x5 FILLER_208_1810 ();
 b15zdnd11an1n32x5 FILLER_208_1850 ();
 b15zdnd11an1n08x5 FILLER_208_1882 ();
 b15zdnd00an1n01x5 FILLER_208_1890 ();
 b15zdnd11an1n08x5 FILLER_208_1900 ();
 b15zdnd11an1n04x5 FILLER_208_1908 ();
 b15zdnd00an1n02x5 FILLER_208_1912 ();
 b15zdnd00an1n01x5 FILLER_208_1914 ();
 b15zdnd11an1n64x5 FILLER_208_1935 ();
 b15zdnd11an1n32x5 FILLER_208_1999 ();
 b15zdnd11an1n08x5 FILLER_208_2031 ();
 b15zdnd11an1n04x5 FILLER_208_2039 ();
 b15zdnd11an1n64x5 FILLER_208_2063 ();
 b15zdnd11an1n16x5 FILLER_208_2127 ();
 b15zdnd11an1n08x5 FILLER_208_2143 ();
 b15zdnd00an1n02x5 FILLER_208_2151 ();
 b15zdnd00an1n01x5 FILLER_208_2153 ();
 b15zdnd11an1n64x5 FILLER_208_2162 ();
 b15zdnd00an1n02x5 FILLER_208_2226 ();
 b15zdnd00an1n01x5 FILLER_208_2228 ();
 b15zdnd11an1n04x5 FILLER_208_2249 ();
 b15zdnd11an1n04x5 FILLER_208_2257 ();
 b15zdnd11an1n08x5 FILLER_208_2265 ();
 b15zdnd00an1n02x5 FILLER_208_2273 ();
 b15zdnd00an1n01x5 FILLER_208_2275 ();
 b15zdnd11an1n64x5 FILLER_209_0 ();
 b15zdnd11an1n64x5 FILLER_209_64 ();
 b15zdnd11an1n64x5 FILLER_209_128 ();
 b15zdnd11an1n64x5 FILLER_209_192 ();
 b15zdnd11an1n64x5 FILLER_209_256 ();
 b15zdnd11an1n32x5 FILLER_209_320 ();
 b15zdnd11an1n16x5 FILLER_209_352 ();
 b15zdnd11an1n04x5 FILLER_209_368 ();
 b15zdnd11an1n64x5 FILLER_209_378 ();
 b15zdnd11an1n32x5 FILLER_209_442 ();
 b15zdnd11an1n08x5 FILLER_209_474 ();
 b15zdnd11an1n04x5 FILLER_209_482 ();
 b15zdnd00an1n02x5 FILLER_209_486 ();
 b15zdnd00an1n01x5 FILLER_209_488 ();
 b15zdnd11an1n64x5 FILLER_209_501 ();
 b15zdnd11an1n16x5 FILLER_209_565 ();
 b15zdnd11an1n08x5 FILLER_209_581 ();
 b15zdnd00an1n02x5 FILLER_209_589 ();
 b15zdnd00an1n01x5 FILLER_209_591 ();
 b15zdnd11an1n04x5 FILLER_209_601 ();
 b15zdnd11an1n32x5 FILLER_209_619 ();
 b15zdnd11an1n16x5 FILLER_209_651 ();
 b15zdnd00an1n02x5 FILLER_209_667 ();
 b15zdnd00an1n01x5 FILLER_209_669 ();
 b15zdnd11an1n16x5 FILLER_209_675 ();
 b15zdnd00an1n02x5 FILLER_209_691 ();
 b15zdnd00an1n01x5 FILLER_209_693 ();
 b15zdnd11an1n16x5 FILLER_209_699 ();
 b15zdnd11an1n04x5 FILLER_209_715 ();
 b15zdnd11an1n64x5 FILLER_209_750 ();
 b15zdnd11an1n16x5 FILLER_209_814 ();
 b15zdnd11an1n08x5 FILLER_209_830 ();
 b15zdnd00an1n02x5 FILLER_209_838 ();
 b15zdnd00an1n01x5 FILLER_209_840 ();
 b15zdnd11an1n32x5 FILLER_209_853 ();
 b15zdnd11an1n16x5 FILLER_209_885 ();
 b15zdnd11an1n08x5 FILLER_209_901 ();
 b15zdnd00an1n02x5 FILLER_209_909 ();
 b15zdnd00an1n01x5 FILLER_209_911 ();
 b15zdnd11an1n32x5 FILLER_209_918 ();
 b15zdnd11an1n16x5 FILLER_209_950 ();
 b15zdnd00an1n02x5 FILLER_209_966 ();
 b15zdnd00an1n01x5 FILLER_209_968 ();
 b15zdnd11an1n16x5 FILLER_209_978 ();
 b15zdnd11an1n04x5 FILLER_209_994 ();
 b15zdnd00an1n01x5 FILLER_209_998 ();
 b15zdnd11an1n32x5 FILLER_209_1015 ();
 b15zdnd11an1n04x5 FILLER_209_1047 ();
 b15zdnd00an1n02x5 FILLER_209_1051 ();
 b15zdnd11an1n04x5 FILLER_209_1062 ();
 b15zdnd11an1n08x5 FILLER_209_1071 ();
 b15zdnd11an1n04x5 FILLER_209_1079 ();
 b15zdnd00an1n01x5 FILLER_209_1083 ();
 b15zdnd11an1n16x5 FILLER_209_1090 ();
 b15zdnd11an1n08x5 FILLER_209_1106 ();
 b15zdnd00an1n02x5 FILLER_209_1114 ();
 b15zdnd11an1n04x5 FILLER_209_1128 ();
 b15zdnd11an1n64x5 FILLER_209_1136 ();
 b15zdnd11an1n32x5 FILLER_209_1200 ();
 b15zdnd11an1n16x5 FILLER_209_1232 ();
 b15zdnd11an1n08x5 FILLER_209_1248 ();
 b15zdnd11an1n04x5 FILLER_209_1256 ();
 b15zdnd11an1n08x5 FILLER_209_1280 ();
 b15zdnd11an1n04x5 FILLER_209_1288 ();
 b15zdnd11an1n64x5 FILLER_209_1297 ();
 b15zdnd11an1n08x5 FILLER_209_1361 ();
 b15zdnd11an1n04x5 FILLER_209_1375 ();
 b15zdnd11an1n08x5 FILLER_209_1383 ();
 b15zdnd11an1n04x5 FILLER_209_1391 ();
 b15zdnd00an1n01x5 FILLER_209_1395 ();
 b15zdnd11an1n08x5 FILLER_209_1408 ();
 b15zdnd11an1n04x5 FILLER_209_1416 ();
 b15zdnd00an1n01x5 FILLER_209_1420 ();
 b15zdnd11an1n16x5 FILLER_209_1430 ();
 b15zdnd11an1n04x5 FILLER_209_1446 ();
 b15zdnd00an1n02x5 FILLER_209_1450 ();
 b15zdnd11an1n04x5 FILLER_209_1472 ();
 b15zdnd11an1n08x5 FILLER_209_1493 ();
 b15zdnd11an1n04x5 FILLER_209_1501 ();
 b15zdnd00an1n01x5 FILLER_209_1505 ();
 b15zdnd11an1n16x5 FILLER_209_1511 ();
 b15zdnd00an1n01x5 FILLER_209_1527 ();
 b15zdnd11an1n16x5 FILLER_209_1533 ();
 b15zdnd11an1n04x5 FILLER_209_1549 ();
 b15zdnd00an1n02x5 FILLER_209_1553 ();
 b15zdnd00an1n01x5 FILLER_209_1555 ();
 b15zdnd11an1n32x5 FILLER_209_1560 ();
 b15zdnd11an1n08x5 FILLER_209_1592 ();
 b15zdnd11an1n04x5 FILLER_209_1600 ();
 b15zdnd00an1n02x5 FILLER_209_1604 ();
 b15zdnd00an1n01x5 FILLER_209_1606 ();
 b15zdnd11an1n04x5 FILLER_209_1612 ();
 b15zdnd00an1n02x5 FILLER_209_1616 ();
 b15zdnd11an1n32x5 FILLER_209_1623 ();
 b15zdnd11an1n16x5 FILLER_209_1662 ();
 b15zdnd11an1n08x5 FILLER_209_1678 ();
 b15zdnd00an1n01x5 FILLER_209_1686 ();
 b15zdnd11an1n16x5 FILLER_209_1699 ();
 b15zdnd11an1n04x5 FILLER_209_1715 ();
 b15zdnd11an1n64x5 FILLER_209_1744 ();
 b15zdnd11an1n32x5 FILLER_209_1808 ();
 b15zdnd11an1n16x5 FILLER_209_1840 ();
 b15zdnd11an1n08x5 FILLER_209_1856 ();
 b15zdnd11an1n04x5 FILLER_209_1864 ();
 b15zdnd00an1n02x5 FILLER_209_1868 ();
 b15zdnd00an1n01x5 FILLER_209_1870 ();
 b15zdnd11an1n16x5 FILLER_209_1896 ();
 b15zdnd11an1n04x5 FILLER_209_1940 ();
 b15zdnd11an1n04x5 FILLER_209_1964 ();
 b15zdnd11an1n16x5 FILLER_209_1973 ();
 b15zdnd11an1n04x5 FILLER_209_2004 ();
 b15zdnd11an1n16x5 FILLER_209_2013 ();
 b15zdnd11an1n08x5 FILLER_209_2029 ();
 b15zdnd00an1n02x5 FILLER_209_2037 ();
 b15zdnd00an1n01x5 FILLER_209_2039 ();
 b15zdnd11an1n16x5 FILLER_209_2049 ();
 b15zdnd11an1n04x5 FILLER_209_2065 ();
 b15zdnd00an1n02x5 FILLER_209_2069 ();
 b15zdnd00an1n01x5 FILLER_209_2071 ();
 b15zdnd11an1n32x5 FILLER_209_2091 ();
 b15zdnd11an1n16x5 FILLER_209_2123 ();
 b15zdnd11an1n08x5 FILLER_209_2139 ();
 b15zdnd11an1n04x5 FILLER_209_2147 ();
 b15zdnd11an1n16x5 FILLER_209_2172 ();
 b15zdnd11an1n08x5 FILLER_209_2188 ();
 b15zdnd11an1n04x5 FILLER_209_2196 ();
 b15zdnd00an1n02x5 FILLER_209_2200 ();
 b15zdnd00an1n01x5 FILLER_209_2202 ();
 b15zdnd11an1n16x5 FILLER_209_2212 ();
 b15zdnd11an1n08x5 FILLER_209_2228 ();
 b15zdnd00an1n01x5 FILLER_209_2236 ();
 b15zdnd11an1n04x5 FILLER_209_2257 ();
 b15zdnd11an1n08x5 FILLER_209_2265 ();
 b15zdnd11an1n04x5 FILLER_209_2277 ();
 b15zdnd00an1n02x5 FILLER_209_2281 ();
 b15zdnd00an1n01x5 FILLER_209_2283 ();
 b15zdnd11an1n64x5 FILLER_210_8 ();
 b15zdnd11an1n64x5 FILLER_210_72 ();
 b15zdnd11an1n64x5 FILLER_210_136 ();
 b15zdnd11an1n64x5 FILLER_210_200 ();
 b15zdnd11an1n64x5 FILLER_210_264 ();
 b15zdnd11an1n64x5 FILLER_210_328 ();
 b15zdnd11an1n32x5 FILLER_210_392 ();
 b15zdnd11an1n16x5 FILLER_210_424 ();
 b15zdnd11an1n08x5 FILLER_210_440 ();
 b15zdnd11an1n04x5 FILLER_210_448 ();
 b15zdnd00an1n02x5 FILLER_210_452 ();
 b15zdnd11an1n04x5 FILLER_210_458 ();
 b15zdnd11an1n32x5 FILLER_210_469 ();
 b15zdnd11an1n16x5 FILLER_210_501 ();
 b15zdnd11an1n08x5 FILLER_210_517 ();
 b15zdnd11an1n04x5 FILLER_210_525 ();
 b15zdnd00an1n02x5 FILLER_210_529 ();
 b15zdnd11an1n64x5 FILLER_210_536 ();
 b15zdnd11an1n64x5 FILLER_210_600 ();
 b15zdnd11an1n32x5 FILLER_210_664 ();
 b15zdnd11an1n16x5 FILLER_210_696 ();
 b15zdnd11an1n04x5 FILLER_210_712 ();
 b15zdnd00an1n02x5 FILLER_210_716 ();
 b15zdnd11an1n64x5 FILLER_210_726 ();
 b15zdnd11an1n64x5 FILLER_210_790 ();
 b15zdnd11an1n16x5 FILLER_210_854 ();
 b15zdnd11an1n08x5 FILLER_210_870 ();
 b15zdnd11an1n64x5 FILLER_210_890 ();
 b15zdnd11an1n16x5 FILLER_210_954 ();
 b15zdnd00an1n02x5 FILLER_210_970 ();
 b15zdnd11an1n16x5 FILLER_210_979 ();
 b15zdnd11an1n04x5 FILLER_210_995 ();
 b15zdnd00an1n02x5 FILLER_210_999 ();
 b15zdnd00an1n01x5 FILLER_210_1001 ();
 b15zdnd11an1n16x5 FILLER_210_1034 ();
 b15zdnd11an1n08x5 FILLER_210_1050 ();
 b15zdnd11an1n08x5 FILLER_210_1063 ();
 b15zdnd11an1n04x5 FILLER_210_1071 ();
 b15zdnd00an1n01x5 FILLER_210_1075 ();
 b15zdnd11an1n04x5 FILLER_210_1084 ();
 b15zdnd11an1n16x5 FILLER_210_1100 ();
 b15zdnd00an1n02x5 FILLER_210_1116 ();
 b15zdnd11an1n04x5 FILLER_210_1124 ();
 b15zdnd11an1n64x5 FILLER_210_1134 ();
 b15zdnd11an1n64x5 FILLER_210_1198 ();
 b15zdnd11an1n64x5 FILLER_210_1262 ();
 b15zdnd11an1n64x5 FILLER_210_1326 ();
 b15zdnd11an1n64x5 FILLER_210_1390 ();
 b15zdnd11an1n04x5 FILLER_210_1466 ();
 b15zdnd00an1n02x5 FILLER_210_1470 ();
 b15zdnd11an1n16x5 FILLER_210_1478 ();
 b15zdnd11an1n08x5 FILLER_210_1494 ();
 b15zdnd00an1n01x5 FILLER_210_1502 ();
 b15zdnd11an1n08x5 FILLER_210_1509 ();
 b15zdnd11an1n04x5 FILLER_210_1527 ();
 b15zdnd11an1n64x5 FILLER_210_1538 ();
 b15zdnd11an1n08x5 FILLER_210_1602 ();
 b15zdnd00an1n02x5 FILLER_210_1610 ();
 b15zdnd00an1n01x5 FILLER_210_1612 ();
 b15zdnd11an1n08x5 FILLER_210_1619 ();
 b15zdnd11an1n04x5 FILLER_210_1627 ();
 b15zdnd00an1n02x5 FILLER_210_1631 ();
 b15zdnd00an1n01x5 FILLER_210_1633 ();
 b15zdnd11an1n32x5 FILLER_210_1640 ();
 b15zdnd11an1n04x5 FILLER_210_1672 ();
 b15zdnd00an1n02x5 FILLER_210_1676 ();
 b15zdnd00an1n01x5 FILLER_210_1678 ();
 b15zdnd11an1n08x5 FILLER_210_1705 ();
 b15zdnd11an1n04x5 FILLER_210_1713 ();
 b15zdnd11an1n64x5 FILLER_210_1739 ();
 b15zdnd11an1n32x5 FILLER_210_1803 ();
 b15zdnd11an1n16x5 FILLER_210_1835 ();
 b15zdnd11an1n08x5 FILLER_210_1851 ();
 b15zdnd11an1n32x5 FILLER_210_1879 ();
 b15zdnd11an1n16x5 FILLER_210_1911 ();
 b15zdnd11an1n04x5 FILLER_210_1958 ();
 b15zdnd11an1n04x5 FILLER_210_1965 ();
 b15zdnd00an1n02x5 FILLER_210_1969 ();
 b15zdnd11an1n08x5 FILLER_210_1997 ();
 b15zdnd11an1n04x5 FILLER_210_2005 ();
 b15zdnd11an1n32x5 FILLER_210_2029 ();
 b15zdnd11an1n16x5 FILLER_210_2061 ();
 b15zdnd11an1n08x5 FILLER_210_2077 ();
 b15zdnd00an1n01x5 FILLER_210_2085 ();
 b15zdnd11an1n08x5 FILLER_210_2090 ();
 b15zdnd11an1n04x5 FILLER_210_2098 ();
 b15zdnd00an1n02x5 FILLER_210_2102 ();
 b15zdnd00an1n01x5 FILLER_210_2104 ();
 b15zdnd11an1n16x5 FILLER_210_2125 ();
 b15zdnd00an1n02x5 FILLER_210_2152 ();
 b15zdnd00an1n02x5 FILLER_210_2162 ();
 b15zdnd11an1n08x5 FILLER_210_2195 ();
 b15zdnd00an1n01x5 FILLER_210_2203 ();
 b15zdnd11an1n04x5 FILLER_210_2214 ();
 b15zdnd00an1n02x5 FILLER_210_2218 ();
 b15zdnd11an1n08x5 FILLER_210_2225 ();
 b15zdnd11an1n04x5 FILLER_210_2233 ();
 b15zdnd00an1n02x5 FILLER_210_2237 ();
 b15zdnd00an1n01x5 FILLER_210_2239 ();
 b15zdnd11an1n08x5 FILLER_210_2244 ();
 b15zdnd11an1n04x5 FILLER_210_2252 ();
 b15zdnd11an1n04x5 FILLER_210_2260 ();
 b15zdnd11an1n08x5 FILLER_210_2268 ();
 b15zdnd11an1n32x5 FILLER_211_0 ();
 b15zdnd00an1n01x5 FILLER_211_32 ();
 b15zdnd11an1n64x5 FILLER_211_37 ();
 b15zdnd11an1n64x5 FILLER_211_101 ();
 b15zdnd11an1n16x5 FILLER_211_165 ();
 b15zdnd11an1n32x5 FILLER_211_190 ();
 b15zdnd11an1n16x5 FILLER_211_222 ();
 b15zdnd11an1n04x5 FILLER_211_238 ();
 b15zdnd00an1n02x5 FILLER_211_242 ();
 b15zdnd11an1n64x5 FILLER_211_249 ();
 b15zdnd11an1n32x5 FILLER_211_313 ();
 b15zdnd11an1n16x5 FILLER_211_345 ();
 b15zdnd11an1n08x5 FILLER_211_361 ();
 b15zdnd11an1n04x5 FILLER_211_376 ();
 b15zdnd11an1n04x5 FILLER_211_385 ();
 b15zdnd00an1n02x5 FILLER_211_389 ();
 b15zdnd00an1n01x5 FILLER_211_391 ();
 b15zdnd11an1n32x5 FILLER_211_424 ();
 b15zdnd11an1n04x5 FILLER_211_456 ();
 b15zdnd00an1n02x5 FILLER_211_460 ();
 b15zdnd11an1n64x5 FILLER_211_468 ();
 b15zdnd11an1n32x5 FILLER_211_532 ();
 b15zdnd11an1n16x5 FILLER_211_564 ();
 b15zdnd11an1n08x5 FILLER_211_580 ();
 b15zdnd11an1n04x5 FILLER_211_588 ();
 b15zdnd00an1n02x5 FILLER_211_592 ();
 b15zdnd00an1n01x5 FILLER_211_594 ();
 b15zdnd11an1n64x5 FILLER_211_600 ();
 b15zdnd11an1n16x5 FILLER_211_664 ();
 b15zdnd11an1n08x5 FILLER_211_680 ();
 b15zdnd11an1n04x5 FILLER_211_688 ();
 b15zdnd00an1n02x5 FILLER_211_692 ();
 b15zdnd11an1n64x5 FILLER_211_699 ();
 b15zdnd11an1n64x5 FILLER_211_763 ();
 b15zdnd11an1n08x5 FILLER_211_827 ();
 b15zdnd11an1n04x5 FILLER_211_835 ();
 b15zdnd00an1n02x5 FILLER_211_839 ();
 b15zdnd00an1n01x5 FILLER_211_841 ();
 b15zdnd11an1n32x5 FILLER_211_847 ();
 b15zdnd00an1n02x5 FILLER_211_879 ();
 b15zdnd11an1n08x5 FILLER_211_891 ();
 b15zdnd11an1n32x5 FILLER_211_903 ();
 b15zdnd11an1n16x5 FILLER_211_935 ();
 b15zdnd11an1n08x5 FILLER_211_951 ();
 b15zdnd11an1n04x5 FILLER_211_959 ();
 b15zdnd00an1n01x5 FILLER_211_963 ();
 b15zdnd11an1n16x5 FILLER_211_969 ();
 b15zdnd11an1n04x5 FILLER_211_985 ();
 b15zdnd00an1n01x5 FILLER_211_989 ();
 b15zdnd11an1n16x5 FILLER_211_1004 ();
 b15zdnd00an1n02x5 FILLER_211_1020 ();
 b15zdnd11an1n32x5 FILLER_211_1027 ();
 b15zdnd11an1n16x5 FILLER_211_1059 ();
 b15zdnd11an1n08x5 FILLER_211_1075 ();
 b15zdnd00an1n01x5 FILLER_211_1083 ();
 b15zdnd11an1n32x5 FILLER_211_1089 ();
 b15zdnd00an1n02x5 FILLER_211_1121 ();
 b15zdnd11an1n32x5 FILLER_211_1134 ();
 b15zdnd11an1n08x5 FILLER_211_1166 ();
 b15zdnd11an1n04x5 FILLER_211_1174 ();
 b15zdnd00an1n02x5 FILLER_211_1178 ();
 b15zdnd00an1n01x5 FILLER_211_1180 ();
 b15zdnd11an1n16x5 FILLER_211_1186 ();
 b15zdnd11an1n08x5 FILLER_211_1202 ();
 b15zdnd11an1n04x5 FILLER_211_1210 ();
 b15zdnd00an1n02x5 FILLER_211_1214 ();
 b15zdnd11an1n64x5 FILLER_211_1226 ();
 b15zdnd11an1n04x5 FILLER_211_1290 ();
 b15zdnd00an1n02x5 FILLER_211_1294 ();
 b15zdnd11an1n08x5 FILLER_211_1302 ();
 b15zdnd11an1n04x5 FILLER_211_1310 ();
 b15zdnd11an1n08x5 FILLER_211_1318 ();
 b15zdnd11an1n04x5 FILLER_211_1326 ();
 b15zdnd11an1n16x5 FILLER_211_1348 ();
 b15zdnd11an1n04x5 FILLER_211_1364 ();
 b15zdnd00an1n02x5 FILLER_211_1368 ();
 b15zdnd11an1n04x5 FILLER_211_1376 ();
 b15zdnd00an1n02x5 FILLER_211_1380 ();
 b15zdnd00an1n01x5 FILLER_211_1382 ();
 b15zdnd11an1n64x5 FILLER_211_1388 ();
 b15zdnd11an1n04x5 FILLER_211_1452 ();
 b15zdnd00an1n02x5 FILLER_211_1456 ();
 b15zdnd00an1n01x5 FILLER_211_1458 ();
 b15zdnd11an1n64x5 FILLER_211_1468 ();
 b15zdnd11an1n08x5 FILLER_211_1532 ();
 b15zdnd11an1n04x5 FILLER_211_1540 ();
 b15zdnd00an1n02x5 FILLER_211_1544 ();
 b15zdnd00an1n01x5 FILLER_211_1546 ();
 b15zdnd11an1n08x5 FILLER_211_1554 ();
 b15zdnd00an1n01x5 FILLER_211_1562 ();
 b15zdnd11an1n16x5 FILLER_211_1568 ();
 b15zdnd11an1n08x5 FILLER_211_1584 ();
 b15zdnd00an1n02x5 FILLER_211_1592 ();
 b15zdnd00an1n01x5 FILLER_211_1594 ();
 b15zdnd11an1n32x5 FILLER_211_1601 ();
 b15zdnd11an1n04x5 FILLER_211_1633 ();
 b15zdnd11an1n64x5 FILLER_211_1653 ();
 b15zdnd11an1n16x5 FILLER_211_1717 ();
 b15zdnd11an1n08x5 FILLER_211_1733 ();
 b15zdnd11an1n64x5 FILLER_211_1750 ();
 b15zdnd11an1n64x5 FILLER_211_1814 ();
 b15zdnd11an1n64x5 FILLER_211_1878 ();
 b15zdnd00an1n02x5 FILLER_211_1942 ();
 b15zdnd00an1n01x5 FILLER_211_1944 ();
 b15zdnd11an1n64x5 FILLER_211_1954 ();
 b15zdnd11an1n64x5 FILLER_211_2018 ();
 b15zdnd11an1n32x5 FILLER_211_2082 ();
 b15zdnd11an1n08x5 FILLER_211_2114 ();
 b15zdnd00an1n02x5 FILLER_211_2122 ();
 b15zdnd11an1n08x5 FILLER_211_2142 ();
 b15zdnd11an1n04x5 FILLER_211_2150 ();
 b15zdnd11an1n08x5 FILLER_211_2182 ();
 b15zdnd00an1n02x5 FILLER_211_2190 ();
 b15zdnd00an1n01x5 FILLER_211_2192 ();
 b15zdnd11an1n16x5 FILLER_211_2196 ();
 b15zdnd00an1n02x5 FILLER_211_2212 ();
 b15zdnd11an1n04x5 FILLER_211_2217 ();
 b15zdnd11an1n08x5 FILLER_211_2241 ();
 b15zdnd11an1n04x5 FILLER_211_2249 ();
 b15zdnd11an1n04x5 FILLER_211_2257 ();
 b15zdnd11an1n04x5 FILLER_211_2265 ();
 b15zdnd11an1n04x5 FILLER_211_2273 ();
 b15zdnd00an1n01x5 FILLER_211_2277 ();
 b15zdnd00an1n02x5 FILLER_211_2282 ();
 b15zdnd11an1n64x5 FILLER_212_8 ();
 b15zdnd11an1n08x5 FILLER_212_72 ();
 b15zdnd00an1n02x5 FILLER_212_80 ();
 b15zdnd00an1n01x5 FILLER_212_82 ();
 b15zdnd11an1n64x5 FILLER_212_99 ();
 b15zdnd11an1n08x5 FILLER_212_163 ();
 b15zdnd11an1n08x5 FILLER_212_180 ();
 b15zdnd11an1n16x5 FILLER_212_197 ();
 b15zdnd00an1n02x5 FILLER_212_213 ();
 b15zdnd11an1n16x5 FILLER_212_220 ();
 b15zdnd11an1n08x5 FILLER_212_236 ();
 b15zdnd00an1n02x5 FILLER_212_244 ();
 b15zdnd11an1n16x5 FILLER_212_255 ();
 b15zdnd11an1n08x5 FILLER_212_271 ();
 b15zdnd00an1n02x5 FILLER_212_279 ();
 b15zdnd11an1n08x5 FILLER_212_285 ();
 b15zdnd11an1n32x5 FILLER_212_313 ();
 b15zdnd11an1n16x5 FILLER_212_345 ();
 b15zdnd11an1n08x5 FILLER_212_361 ();
 b15zdnd11an1n04x5 FILLER_212_369 ();
 b15zdnd00an1n02x5 FILLER_212_373 ();
 b15zdnd00an1n01x5 FILLER_212_375 ();
 b15zdnd11an1n04x5 FILLER_212_382 ();
 b15zdnd11an1n16x5 FILLER_212_392 ();
 b15zdnd11an1n08x5 FILLER_212_408 ();
 b15zdnd11an1n04x5 FILLER_212_416 ();
 b15zdnd00an1n02x5 FILLER_212_420 ();
 b15zdnd11an1n32x5 FILLER_212_428 ();
 b15zdnd11an1n16x5 FILLER_212_460 ();
 b15zdnd11an1n04x5 FILLER_212_476 ();
 b15zdnd11an1n16x5 FILLER_212_490 ();
 b15zdnd11an1n08x5 FILLER_212_506 ();
 b15zdnd11an1n04x5 FILLER_212_514 ();
 b15zdnd00an1n01x5 FILLER_212_518 ();
 b15zdnd11an1n16x5 FILLER_212_526 ();
 b15zdnd11an1n04x5 FILLER_212_552 ();
 b15zdnd11an1n08x5 FILLER_212_562 ();
 b15zdnd00an1n01x5 FILLER_212_570 ();
 b15zdnd11an1n04x5 FILLER_212_576 ();
 b15zdnd00an1n01x5 FILLER_212_580 ();
 b15zdnd11an1n08x5 FILLER_212_586 ();
 b15zdnd00an1n02x5 FILLER_212_594 ();
 b15zdnd00an1n01x5 FILLER_212_596 ();
 b15zdnd11an1n16x5 FILLER_212_602 ();
 b15zdnd11an1n04x5 FILLER_212_618 ();
 b15zdnd00an1n02x5 FILLER_212_622 ();
 b15zdnd11an1n16x5 FILLER_212_631 ();
 b15zdnd00an1n02x5 FILLER_212_647 ();
 b15zdnd00an1n01x5 FILLER_212_649 ();
 b15zdnd11an1n16x5 FILLER_212_659 ();
 b15zdnd11an1n04x5 FILLER_212_675 ();
 b15zdnd00an1n02x5 FILLER_212_679 ();
 b15zdnd00an1n01x5 FILLER_212_681 ();
 b15zdnd11an1n08x5 FILLER_212_708 ();
 b15zdnd00an1n02x5 FILLER_212_716 ();
 b15zdnd00an1n02x5 FILLER_212_726 ();
 b15zdnd11an1n64x5 FILLER_212_760 ();
 b15zdnd11an1n32x5 FILLER_212_824 ();
 b15zdnd11an1n04x5 FILLER_212_864 ();
 b15zdnd11an1n16x5 FILLER_212_896 ();
 b15zdnd11an1n04x5 FILLER_212_912 ();
 b15zdnd11an1n04x5 FILLER_212_922 ();
 b15zdnd11an1n16x5 FILLER_212_936 ();
 b15zdnd11an1n08x5 FILLER_212_952 ();
 b15zdnd00an1n02x5 FILLER_212_960 ();
 b15zdnd00an1n01x5 FILLER_212_962 ();
 b15zdnd11an1n32x5 FILLER_212_977 ();
 b15zdnd11an1n16x5 FILLER_212_1009 ();
 b15zdnd00an1n02x5 FILLER_212_1025 ();
 b15zdnd11an1n16x5 FILLER_212_1031 ();
 b15zdnd11an1n08x5 FILLER_212_1047 ();
 b15zdnd11an1n04x5 FILLER_212_1055 ();
 b15zdnd00an1n02x5 FILLER_212_1059 ();
 b15zdnd11an1n64x5 FILLER_212_1077 ();
 b15zdnd11an1n08x5 FILLER_212_1141 ();
 b15zdnd11an1n04x5 FILLER_212_1149 ();
 b15zdnd00an1n02x5 FILLER_212_1153 ();
 b15zdnd00an1n01x5 FILLER_212_1155 ();
 b15zdnd11an1n08x5 FILLER_212_1160 ();
 b15zdnd11an1n04x5 FILLER_212_1168 ();
 b15zdnd00an1n02x5 FILLER_212_1172 ();
 b15zdnd11an1n08x5 FILLER_212_1180 ();
 b15zdnd11an1n08x5 FILLER_212_1194 ();
 b15zdnd11an1n04x5 FILLER_212_1208 ();
 b15zdnd00an1n02x5 FILLER_212_1212 ();
 b15zdnd00an1n01x5 FILLER_212_1214 ();
 b15zdnd11an1n32x5 FILLER_212_1246 ();
 b15zdnd11an1n08x5 FILLER_212_1278 ();
 b15zdnd11an1n04x5 FILLER_212_1286 ();
 b15zdnd00an1n02x5 FILLER_212_1290 ();
 b15zdnd11an1n04x5 FILLER_212_1299 ();
 b15zdnd11an1n16x5 FILLER_212_1307 ();
 b15zdnd11an1n08x5 FILLER_212_1323 ();
 b15zdnd00an1n02x5 FILLER_212_1331 ();
 b15zdnd11an1n04x5 FILLER_212_1347 ();
 b15zdnd11an1n04x5 FILLER_212_1374 ();
 b15zdnd00an1n01x5 FILLER_212_1378 ();
 b15zdnd11an1n64x5 FILLER_212_1387 ();
 b15zdnd11an1n64x5 FILLER_212_1451 ();
 b15zdnd11an1n16x5 FILLER_212_1515 ();
 b15zdnd00an1n02x5 FILLER_212_1531 ();
 b15zdnd11an1n08x5 FILLER_212_1541 ();
 b15zdnd00an1n02x5 FILLER_212_1549 ();
 b15zdnd00an1n01x5 FILLER_212_1551 ();
 b15zdnd11an1n08x5 FILLER_212_1564 ();
 b15zdnd11an1n04x5 FILLER_212_1572 ();
 b15zdnd11an1n64x5 FILLER_212_1588 ();
 b15zdnd11an1n04x5 FILLER_212_1652 ();
 b15zdnd11an1n64x5 FILLER_212_1671 ();
 b15zdnd11an1n32x5 FILLER_212_1735 ();
 b15zdnd11an1n08x5 FILLER_212_1767 ();
 b15zdnd00an1n01x5 FILLER_212_1775 ();
 b15zdnd11an1n04x5 FILLER_212_1802 ();
 b15zdnd11an1n64x5 FILLER_212_1831 ();
 b15zdnd00an1n01x5 FILLER_212_1895 ();
 b15zdnd11an1n64x5 FILLER_212_1900 ();
 b15zdnd11an1n04x5 FILLER_212_1964 ();
 b15zdnd00an1n02x5 FILLER_212_1968 ();
 b15zdnd11an1n64x5 FILLER_212_1988 ();
 b15zdnd11an1n32x5 FILLER_212_2052 ();
 b15zdnd11an1n08x5 FILLER_212_2084 ();
 b15zdnd11an1n04x5 FILLER_212_2092 ();
 b15zdnd00an1n02x5 FILLER_212_2096 ();
 b15zdnd00an1n01x5 FILLER_212_2098 ();
 b15zdnd11an1n32x5 FILLER_212_2110 ();
 b15zdnd11an1n08x5 FILLER_212_2142 ();
 b15zdnd11an1n04x5 FILLER_212_2150 ();
 b15zdnd11an1n64x5 FILLER_212_2162 ();
 b15zdnd11an1n16x5 FILLER_212_2226 ();
 b15zdnd11an1n08x5 FILLER_212_2242 ();
 b15zdnd00an1n01x5 FILLER_212_2250 ();
 b15zdnd11an1n16x5 FILLER_212_2255 ();
 b15zdnd11an1n04x5 FILLER_212_2271 ();
 b15zdnd00an1n01x5 FILLER_212_2275 ();
 b15zdnd11an1n64x5 FILLER_213_0 ();
 b15zdnd11an1n64x5 FILLER_213_64 ();
 b15zdnd11an1n08x5 FILLER_213_128 ();
 b15zdnd11an1n04x5 FILLER_213_136 ();
 b15zdnd11an1n32x5 FILLER_213_145 ();
 b15zdnd11an1n04x5 FILLER_213_177 ();
 b15zdnd00an1n02x5 FILLER_213_181 ();
 b15zdnd00an1n01x5 FILLER_213_183 ();
 b15zdnd11an1n16x5 FILLER_213_193 ();
 b15zdnd11an1n32x5 FILLER_213_215 ();
 b15zdnd11an1n04x5 FILLER_213_247 ();
 b15zdnd00an1n01x5 FILLER_213_251 ();
 b15zdnd11an1n16x5 FILLER_213_259 ();
 b15zdnd11an1n04x5 FILLER_213_275 ();
 b15zdnd00an1n02x5 FILLER_213_279 ();
 b15zdnd11an1n04x5 FILLER_213_296 ();
 b15zdnd00an1n02x5 FILLER_213_300 ();
 b15zdnd11an1n04x5 FILLER_213_314 ();
 b15zdnd11an1n32x5 FILLER_213_334 ();
 b15zdnd11an1n04x5 FILLER_213_366 ();
 b15zdnd00an1n02x5 FILLER_213_370 ();
 b15zdnd11an1n08x5 FILLER_213_379 ();
 b15zdnd11an1n04x5 FILLER_213_387 ();
 b15zdnd00an1n01x5 FILLER_213_391 ();
 b15zdnd11an1n04x5 FILLER_213_408 ();
 b15zdnd00an1n02x5 FILLER_213_412 ();
 b15zdnd11an1n08x5 FILLER_213_425 ();
 b15zdnd11an1n08x5 FILLER_213_443 ();
 b15zdnd11an1n04x5 FILLER_213_467 ();
 b15zdnd00an1n02x5 FILLER_213_471 ();
 b15zdnd00an1n01x5 FILLER_213_473 ();
 b15zdnd11an1n16x5 FILLER_213_478 ();
 b15zdnd00an1n02x5 FILLER_213_494 ();
 b15zdnd11an1n16x5 FILLER_213_505 ();
 b15zdnd11an1n08x5 FILLER_213_521 ();
 b15zdnd00an1n01x5 FILLER_213_529 ();
 b15zdnd11an1n04x5 FILLER_213_540 ();
 b15zdnd11an1n04x5 FILLER_213_553 ();
 b15zdnd11an1n16x5 FILLER_213_561 ();
 b15zdnd11an1n08x5 FILLER_213_577 ();
 b15zdnd00an1n02x5 FILLER_213_585 ();
 b15zdnd00an1n01x5 FILLER_213_587 ();
 b15zdnd11an1n16x5 FILLER_213_597 ();
 b15zdnd11an1n04x5 FILLER_213_613 ();
 b15zdnd00an1n02x5 FILLER_213_617 ();
 b15zdnd00an1n01x5 FILLER_213_619 ();
 b15zdnd11an1n16x5 FILLER_213_625 ();
 b15zdnd11an1n04x5 FILLER_213_641 ();
 b15zdnd00an1n02x5 FILLER_213_645 ();
 b15zdnd00an1n01x5 FILLER_213_647 ();
 b15zdnd11an1n08x5 FILLER_213_656 ();
 b15zdnd00an1n02x5 FILLER_213_664 ();
 b15zdnd11an1n04x5 FILLER_213_687 ();
 b15zdnd11an1n08x5 FILLER_213_698 ();
 b15zdnd11an1n04x5 FILLER_213_706 ();
 b15zdnd00an1n02x5 FILLER_213_710 ();
 b15zdnd00an1n01x5 FILLER_213_712 ();
 b15zdnd11an1n04x5 FILLER_213_717 ();
 b15zdnd00an1n02x5 FILLER_213_721 ();
 b15zdnd00an1n01x5 FILLER_213_723 ();
 b15zdnd11an1n04x5 FILLER_213_756 ();
 b15zdnd11an1n04x5 FILLER_213_774 ();
 b15zdnd11an1n04x5 FILLER_213_804 ();
 b15zdnd00an1n01x5 FILLER_213_808 ();
 b15zdnd11an1n16x5 FILLER_213_829 ();
 b15zdnd11an1n08x5 FILLER_213_845 ();
 b15zdnd11an1n04x5 FILLER_213_860 ();
 b15zdnd11an1n64x5 FILLER_213_875 ();
 b15zdnd11an1n32x5 FILLER_213_939 ();
 b15zdnd11an1n16x5 FILLER_213_971 ();
 b15zdnd00an1n02x5 FILLER_213_987 ();
 b15zdnd11an1n04x5 FILLER_213_998 ();
 b15zdnd11an1n04x5 FILLER_213_1008 ();
 b15zdnd00an1n01x5 FILLER_213_1012 ();
 b15zdnd11an1n64x5 FILLER_213_1024 ();
 b15zdnd11an1n64x5 FILLER_213_1088 ();
 b15zdnd11an1n08x5 FILLER_213_1152 ();
 b15zdnd11an1n08x5 FILLER_213_1172 ();
 b15zdnd11an1n04x5 FILLER_213_1180 ();
 b15zdnd00an1n01x5 FILLER_213_1184 ();
 b15zdnd11an1n08x5 FILLER_213_1189 ();
 b15zdnd11an1n04x5 FILLER_213_1197 ();
 b15zdnd00an1n01x5 FILLER_213_1201 ();
 b15zdnd11an1n04x5 FILLER_213_1207 ();
 b15zdnd00an1n02x5 FILLER_213_1211 ();
 b15zdnd11an1n64x5 FILLER_213_1222 ();
 b15zdnd00an1n01x5 FILLER_213_1286 ();
 b15zdnd11an1n64x5 FILLER_213_1292 ();
 b15zdnd11an1n16x5 FILLER_213_1356 ();
 b15zdnd11an1n04x5 FILLER_213_1372 ();
 b15zdnd00an1n02x5 FILLER_213_1376 ();
 b15zdnd11an1n04x5 FILLER_213_1385 ();
 b15zdnd11an1n16x5 FILLER_213_1404 ();
 b15zdnd11an1n64x5 FILLER_213_1440 ();
 b15zdnd11an1n04x5 FILLER_213_1509 ();
 b15zdnd00an1n02x5 FILLER_213_1513 ();
 b15zdnd11an1n64x5 FILLER_213_1532 ();
 b15zdnd11an1n16x5 FILLER_213_1596 ();
 b15zdnd00an1n02x5 FILLER_213_1612 ();
 b15zdnd11an1n08x5 FILLER_213_1623 ();
 b15zdnd11an1n04x5 FILLER_213_1631 ();
 b15zdnd00an1n01x5 FILLER_213_1635 ();
 b15zdnd11an1n32x5 FILLER_213_1641 ();
 b15zdnd11an1n04x5 FILLER_213_1673 ();
 b15zdnd00an1n02x5 FILLER_213_1677 ();
 b15zdnd11an1n32x5 FILLER_213_1696 ();
 b15zdnd11an1n16x5 FILLER_213_1728 ();
 b15zdnd00an1n02x5 FILLER_213_1744 ();
 b15zdnd00an1n01x5 FILLER_213_1746 ();
 b15zdnd11an1n64x5 FILLER_213_1756 ();
 b15zdnd11an1n64x5 FILLER_213_1820 ();
 b15zdnd11an1n64x5 FILLER_213_1884 ();
 b15zdnd11an1n64x5 FILLER_213_1948 ();
 b15zdnd11an1n64x5 FILLER_213_2012 ();
 b15zdnd11an1n64x5 FILLER_213_2076 ();
 b15zdnd11an1n04x5 FILLER_213_2140 ();
 b15zdnd00an1n01x5 FILLER_213_2144 ();
 b15zdnd11an1n64x5 FILLER_213_2165 ();
 b15zdnd00an1n02x5 FILLER_213_2229 ();
 b15zdnd00an1n01x5 FILLER_213_2231 ();
 b15zdnd11an1n16x5 FILLER_213_2236 ();
 b15zdnd00an1n02x5 FILLER_213_2252 ();
 b15zdnd00an1n01x5 FILLER_213_2254 ();
 b15zdnd11an1n04x5 FILLER_213_2260 ();
 b15zdnd11an1n04x5 FILLER_213_2268 ();
 b15zdnd00an1n01x5 FILLER_213_2272 ();
 b15zdnd11an1n04x5 FILLER_213_2277 ();
 b15zdnd00an1n02x5 FILLER_213_2281 ();
 b15zdnd00an1n01x5 FILLER_213_2283 ();
 b15zdnd11an1n16x5 FILLER_214_8 ();
 b15zdnd11an1n04x5 FILLER_214_24 ();
 b15zdnd00an1n01x5 FILLER_214_28 ();
 b15zdnd11an1n32x5 FILLER_214_33 ();
 b15zdnd11an1n08x5 FILLER_214_65 ();
 b15zdnd11an1n04x5 FILLER_214_73 ();
 b15zdnd00an1n02x5 FILLER_214_77 ();
 b15zdnd11an1n04x5 FILLER_214_97 ();
 b15zdnd00an1n02x5 FILLER_214_101 ();
 b15zdnd00an1n01x5 FILLER_214_103 ();
 b15zdnd11an1n08x5 FILLER_214_116 ();
 b15zdnd00an1n01x5 FILLER_214_124 ();
 b15zdnd11an1n04x5 FILLER_214_131 ();
 b15zdnd00an1n02x5 FILLER_214_135 ();
 b15zdnd00an1n01x5 FILLER_214_137 ();
 b15zdnd11an1n08x5 FILLER_214_144 ();
 b15zdnd11an1n04x5 FILLER_214_152 ();
 b15zdnd00an1n02x5 FILLER_214_156 ();
 b15zdnd00an1n01x5 FILLER_214_158 ();
 b15zdnd11an1n04x5 FILLER_214_169 ();
 b15zdnd11an1n08x5 FILLER_214_180 ();
 b15zdnd11an1n16x5 FILLER_214_197 ();
 b15zdnd11an1n04x5 FILLER_214_213 ();
 b15zdnd00an1n01x5 FILLER_214_217 ();
 b15zdnd11an1n32x5 FILLER_214_244 ();
 b15zdnd11an1n16x5 FILLER_214_276 ();
 b15zdnd11an1n08x5 FILLER_214_292 ();
 b15zdnd11an1n04x5 FILLER_214_300 ();
 b15zdnd11an1n64x5 FILLER_214_330 ();
 b15zdnd11an1n32x5 FILLER_214_394 ();
 b15zdnd11an1n08x5 FILLER_214_426 ();
 b15zdnd11an1n04x5 FILLER_214_434 ();
 b15zdnd11an1n16x5 FILLER_214_454 ();
 b15zdnd11an1n04x5 FILLER_214_470 ();
 b15zdnd11an1n04x5 FILLER_214_480 ();
 b15zdnd11an1n04x5 FILLER_214_496 ();
 b15zdnd11an1n04x5 FILLER_214_504 ();
 b15zdnd11an1n16x5 FILLER_214_524 ();
 b15zdnd11an1n04x5 FILLER_214_540 ();
 b15zdnd00an1n02x5 FILLER_214_544 ();
 b15zdnd00an1n01x5 FILLER_214_546 ();
 b15zdnd11an1n64x5 FILLER_214_552 ();
 b15zdnd11an1n16x5 FILLER_214_616 ();
 b15zdnd00an1n02x5 FILLER_214_632 ();
 b15zdnd00an1n01x5 FILLER_214_634 ();
 b15zdnd11an1n04x5 FILLER_214_643 ();
 b15zdnd11an1n64x5 FILLER_214_654 ();
 b15zdnd00an1n02x5 FILLER_214_726 ();
 b15zdnd00an1n01x5 FILLER_214_728 ();
 b15zdnd11an1n32x5 FILLER_214_746 ();
 b15zdnd11an1n08x5 FILLER_214_778 ();
 b15zdnd11an1n08x5 FILLER_214_806 ();
 b15zdnd00an1n02x5 FILLER_214_814 ();
 b15zdnd11an1n64x5 FILLER_214_842 ();
 b15zdnd11an1n04x5 FILLER_214_906 ();
 b15zdnd11an1n32x5 FILLER_214_917 ();
 b15zdnd11an1n16x5 FILLER_214_949 ();
 b15zdnd11an1n04x5 FILLER_214_965 ();
 b15zdnd00an1n02x5 FILLER_214_969 ();
 b15zdnd11an1n32x5 FILLER_214_977 ();
 b15zdnd11an1n16x5 FILLER_214_1009 ();
 b15zdnd11an1n08x5 FILLER_214_1025 ();
 b15zdnd11an1n04x5 FILLER_214_1033 ();
 b15zdnd00an1n01x5 FILLER_214_1037 ();
 b15zdnd11an1n08x5 FILLER_214_1043 ();
 b15zdnd11an1n04x5 FILLER_214_1051 ();
 b15zdnd11an1n64x5 FILLER_214_1059 ();
 b15zdnd11an1n16x5 FILLER_214_1123 ();
 b15zdnd11an1n04x5 FILLER_214_1139 ();
 b15zdnd00an1n01x5 FILLER_214_1143 ();
 b15zdnd11an1n64x5 FILLER_214_1148 ();
 b15zdnd11an1n64x5 FILLER_214_1212 ();
 b15zdnd11an1n08x5 FILLER_214_1276 ();
 b15zdnd00an1n02x5 FILLER_214_1284 ();
 b15zdnd11an1n04x5 FILLER_214_1296 ();
 b15zdnd00an1n02x5 FILLER_214_1300 ();
 b15zdnd00an1n01x5 FILLER_214_1302 ();
 b15zdnd11an1n04x5 FILLER_214_1323 ();
 b15zdnd00an1n01x5 FILLER_214_1327 ();
 b15zdnd11an1n04x5 FILLER_214_1348 ();
 b15zdnd11an1n04x5 FILLER_214_1366 ();
 b15zdnd11an1n04x5 FILLER_214_1387 ();
 b15zdnd11an1n16x5 FILLER_214_1411 ();
 b15zdnd11an1n16x5 FILLER_214_1441 ();
 b15zdnd11an1n08x5 FILLER_214_1457 ();
 b15zdnd00an1n01x5 FILLER_214_1465 ();
 b15zdnd11an1n16x5 FILLER_214_1472 ();
 b15zdnd11an1n04x5 FILLER_214_1488 ();
 b15zdnd00an1n01x5 FILLER_214_1492 ();
 b15zdnd11an1n64x5 FILLER_214_1499 ();
 b15zdnd11an1n08x5 FILLER_214_1563 ();
 b15zdnd00an1n01x5 FILLER_214_1571 ();
 b15zdnd11an1n04x5 FILLER_214_1598 ();
 b15zdnd11an1n04x5 FILLER_214_1618 ();
 b15zdnd11an1n32x5 FILLER_214_1628 ();
 b15zdnd11an1n08x5 FILLER_214_1660 ();
 b15zdnd00an1n01x5 FILLER_214_1668 ();
 b15zdnd11an1n04x5 FILLER_214_1675 ();
 b15zdnd11an1n16x5 FILLER_214_1689 ();
 b15zdnd00an1n01x5 FILLER_214_1705 ();
 b15zdnd11an1n64x5 FILLER_214_1716 ();
 b15zdnd11an1n64x5 FILLER_214_1780 ();
 b15zdnd11an1n08x5 FILLER_214_1844 ();
 b15zdnd00an1n02x5 FILLER_214_1852 ();
 b15zdnd11an1n64x5 FILLER_214_1859 ();
 b15zdnd11an1n16x5 FILLER_214_1923 ();
 b15zdnd00an1n02x5 FILLER_214_1939 ();
 b15zdnd11an1n64x5 FILLER_214_1961 ();
 b15zdnd11an1n32x5 FILLER_214_2025 ();
 b15zdnd11an1n16x5 FILLER_214_2057 ();
 b15zdnd11an1n08x5 FILLER_214_2073 ();
 b15zdnd11an1n04x5 FILLER_214_2081 ();
 b15zdnd11an1n08x5 FILLER_214_2103 ();
 b15zdnd00an1n02x5 FILLER_214_2111 ();
 b15zdnd00an1n01x5 FILLER_214_2113 ();
 b15zdnd11an1n32x5 FILLER_214_2119 ();
 b15zdnd00an1n02x5 FILLER_214_2151 ();
 b15zdnd00an1n01x5 FILLER_214_2153 ();
 b15zdnd11an1n64x5 FILLER_214_2162 ();
 b15zdnd11an1n16x5 FILLER_214_2226 ();
 b15zdnd11an1n08x5 FILLER_214_2242 ();
 b15zdnd00an1n02x5 FILLER_214_2250 ();
 b15zdnd00an1n01x5 FILLER_214_2252 ();
 b15zdnd11an1n16x5 FILLER_214_2257 ();
 b15zdnd00an1n02x5 FILLER_214_2273 ();
 b15zdnd00an1n01x5 FILLER_214_2275 ();
 b15zdnd11an1n64x5 FILLER_215_0 ();
 b15zdnd11an1n32x5 FILLER_215_64 ();
 b15zdnd00an1n02x5 FILLER_215_96 ();
 b15zdnd00an1n01x5 FILLER_215_98 ();
 b15zdnd11an1n32x5 FILLER_215_120 ();
 b15zdnd00an1n01x5 FILLER_215_152 ();
 b15zdnd11an1n04x5 FILLER_215_161 ();
 b15zdnd11an1n08x5 FILLER_215_179 ();
 b15zdnd11an1n08x5 FILLER_215_194 ();
 b15zdnd00an1n01x5 FILLER_215_202 ();
 b15zdnd11an1n64x5 FILLER_215_207 ();
 b15zdnd11an1n16x5 FILLER_215_271 ();
 b15zdnd11an1n08x5 FILLER_215_287 ();
 b15zdnd11an1n64x5 FILLER_215_321 ();
 b15zdnd11an1n64x5 FILLER_215_385 ();
 b15zdnd11an1n64x5 FILLER_215_449 ();
 b15zdnd11an1n32x5 FILLER_215_513 ();
 b15zdnd11an1n16x5 FILLER_215_545 ();
 b15zdnd11an1n64x5 FILLER_215_568 ();
 b15zdnd11an1n64x5 FILLER_215_632 ();
 b15zdnd11an1n64x5 FILLER_215_696 ();
 b15zdnd11an1n16x5 FILLER_215_760 ();
 b15zdnd00an1n02x5 FILLER_215_776 ();
 b15zdnd00an1n01x5 FILLER_215_778 ();
 b15zdnd11an1n32x5 FILLER_215_799 ();
 b15zdnd11an1n08x5 FILLER_215_831 ();
 b15zdnd11an1n04x5 FILLER_215_839 ();
 b15zdnd00an1n02x5 FILLER_215_843 ();
 b15zdnd00an1n01x5 FILLER_215_845 ();
 b15zdnd11an1n16x5 FILLER_215_862 ();
 b15zdnd11an1n04x5 FILLER_215_878 ();
 b15zdnd00an1n01x5 FILLER_215_882 ();
 b15zdnd11an1n16x5 FILLER_215_887 ();
 b15zdnd00an1n02x5 FILLER_215_903 ();
 b15zdnd00an1n01x5 FILLER_215_905 ();
 b15zdnd11an1n04x5 FILLER_215_912 ();
 b15zdnd11an1n08x5 FILLER_215_925 ();
 b15zdnd11an1n04x5 FILLER_215_933 ();
 b15zdnd00an1n01x5 FILLER_215_937 ();
 b15zdnd11an1n32x5 FILLER_215_943 ();
 b15zdnd00an1n02x5 FILLER_215_975 ();
 b15zdnd11an1n16x5 FILLER_215_984 ();
 b15zdnd11an1n08x5 FILLER_215_1000 ();
 b15zdnd11an1n04x5 FILLER_215_1008 ();
 b15zdnd00an1n01x5 FILLER_215_1012 ();
 b15zdnd11an1n08x5 FILLER_215_1027 ();
 b15zdnd11an1n04x5 FILLER_215_1035 ();
 b15zdnd00an1n02x5 FILLER_215_1039 ();
 b15zdnd11an1n04x5 FILLER_215_1046 ();
 b15zdnd00an1n01x5 FILLER_215_1050 ();
 b15zdnd11an1n16x5 FILLER_215_1061 ();
 b15zdnd11an1n08x5 FILLER_215_1077 ();
 b15zdnd11an1n04x5 FILLER_215_1085 ();
 b15zdnd00an1n02x5 FILLER_215_1089 ();
 b15zdnd11an1n08x5 FILLER_215_1101 ();
 b15zdnd00an1n02x5 FILLER_215_1109 ();
 b15zdnd11an1n04x5 FILLER_215_1117 ();
 b15zdnd00an1n01x5 FILLER_215_1121 ();
 b15zdnd11an1n04x5 FILLER_215_1135 ();
 b15zdnd00an1n01x5 FILLER_215_1139 ();
 b15zdnd11an1n08x5 FILLER_215_1147 ();
 b15zdnd00an1n01x5 FILLER_215_1155 ();
 b15zdnd11an1n08x5 FILLER_215_1176 ();
 b15zdnd11an1n04x5 FILLER_215_1184 ();
 b15zdnd11an1n08x5 FILLER_215_1212 ();
 b15zdnd11an1n04x5 FILLER_215_1220 ();
 b15zdnd00an1n01x5 FILLER_215_1224 ();
 b15zdnd11an1n64x5 FILLER_215_1251 ();
 b15zdnd11an1n16x5 FILLER_215_1315 ();
 b15zdnd11an1n08x5 FILLER_215_1331 ();
 b15zdnd11an1n04x5 FILLER_215_1339 ();
 b15zdnd11an1n64x5 FILLER_215_1359 ();
 b15zdnd11an1n08x5 FILLER_215_1423 ();
 b15zdnd11an1n04x5 FILLER_215_1431 ();
 b15zdnd00an1n02x5 FILLER_215_1435 ();
 b15zdnd00an1n01x5 FILLER_215_1437 ();
 b15zdnd11an1n16x5 FILLER_215_1442 ();
 b15zdnd11an1n04x5 FILLER_215_1458 ();
 b15zdnd11an1n16x5 FILLER_215_1467 ();
 b15zdnd11an1n08x5 FILLER_215_1483 ();
 b15zdnd00an1n02x5 FILLER_215_1491 ();
 b15zdnd00an1n01x5 FILLER_215_1493 ();
 b15zdnd11an1n32x5 FILLER_215_1500 ();
 b15zdnd11an1n08x5 FILLER_215_1532 ();
 b15zdnd11an1n16x5 FILLER_215_1552 ();
 b15zdnd11an1n08x5 FILLER_215_1568 ();
 b15zdnd11an1n04x5 FILLER_215_1576 ();
 b15zdnd11an1n04x5 FILLER_215_1585 ();
 b15zdnd11an1n32x5 FILLER_215_1594 ();
 b15zdnd11an1n16x5 FILLER_215_1626 ();
 b15zdnd11an1n04x5 FILLER_215_1652 ();
 b15zdnd11an1n64x5 FILLER_215_1661 ();
 b15zdnd11an1n64x5 FILLER_215_1725 ();
 b15zdnd11an1n32x5 FILLER_215_1789 ();
 b15zdnd11an1n16x5 FILLER_215_1821 ();
 b15zdnd11an1n04x5 FILLER_215_1848 ();
 b15zdnd11an1n32x5 FILLER_215_1872 ();
 b15zdnd11an1n16x5 FILLER_215_1904 ();
 b15zdnd00an1n02x5 FILLER_215_1920 ();
 b15zdnd11an1n64x5 FILLER_215_1928 ();
 b15zdnd11an1n08x5 FILLER_215_1992 ();
 b15zdnd11an1n04x5 FILLER_215_2000 ();
 b15zdnd00an1n02x5 FILLER_215_2004 ();
 b15zdnd00an1n01x5 FILLER_215_2006 ();
 b15zdnd11an1n08x5 FILLER_215_2027 ();
 b15zdnd11an1n04x5 FILLER_215_2035 ();
 b15zdnd00an1n02x5 FILLER_215_2039 ();
 b15zdnd11an1n04x5 FILLER_215_2052 ();
 b15zdnd11an1n16x5 FILLER_215_2061 ();
 b15zdnd11an1n04x5 FILLER_215_2077 ();
 b15zdnd11an1n04x5 FILLER_215_2099 ();
 b15zdnd11an1n64x5 FILLER_215_2123 ();
 b15zdnd00an1n02x5 FILLER_215_2187 ();
 b15zdnd00an1n01x5 FILLER_215_2189 ();
 b15zdnd11an1n32x5 FILLER_215_2196 ();
 b15zdnd11an1n08x5 FILLER_215_2228 ();
 b15zdnd00an1n02x5 FILLER_215_2236 ();
 b15zdnd11an1n04x5 FILLER_215_2246 ();
 b15zdnd11an1n16x5 FILLER_215_2266 ();
 b15zdnd00an1n02x5 FILLER_215_2282 ();
 b15zdnd11an1n32x5 FILLER_216_8 ();
 b15zdnd11an1n08x5 FILLER_216_40 ();
 b15zdnd11an1n04x5 FILLER_216_48 ();
 b15zdnd00an1n02x5 FILLER_216_52 ();
 b15zdnd11an1n32x5 FILLER_216_77 ();
 b15zdnd11an1n16x5 FILLER_216_109 ();
 b15zdnd00an1n02x5 FILLER_216_125 ();
 b15zdnd00an1n01x5 FILLER_216_127 ();
 b15zdnd11an1n08x5 FILLER_216_149 ();
 b15zdnd00an1n01x5 FILLER_216_157 ();
 b15zdnd11an1n04x5 FILLER_216_178 ();
 b15zdnd00an1n01x5 FILLER_216_182 ();
 b15zdnd11an1n32x5 FILLER_216_199 ();
 b15zdnd11an1n16x5 FILLER_216_231 ();
 b15zdnd11an1n08x5 FILLER_216_247 ();
 b15zdnd00an1n02x5 FILLER_216_255 ();
 b15zdnd00an1n01x5 FILLER_216_257 ();
 b15zdnd11an1n32x5 FILLER_216_269 ();
 b15zdnd11an1n16x5 FILLER_216_301 ();
 b15zdnd11an1n04x5 FILLER_216_317 ();
 b15zdnd11an1n32x5 FILLER_216_347 ();
 b15zdnd11an1n16x5 FILLER_216_379 ();
 b15zdnd11an1n04x5 FILLER_216_395 ();
 b15zdnd11an1n64x5 FILLER_216_403 ();
 b15zdnd11an1n64x5 FILLER_216_467 ();
 b15zdnd11an1n16x5 FILLER_216_531 ();
 b15zdnd11an1n08x5 FILLER_216_547 ();
 b15zdnd11an1n64x5 FILLER_216_567 ();
 b15zdnd11an1n64x5 FILLER_216_631 ();
 b15zdnd11an1n16x5 FILLER_216_695 ();
 b15zdnd11an1n04x5 FILLER_216_711 ();
 b15zdnd00an1n02x5 FILLER_216_715 ();
 b15zdnd00an1n01x5 FILLER_216_717 ();
 b15zdnd11an1n64x5 FILLER_216_726 ();
 b15zdnd00an1n02x5 FILLER_216_790 ();
 b15zdnd00an1n01x5 FILLER_216_792 ();
 b15zdnd11an1n32x5 FILLER_216_819 ();
 b15zdnd11an1n04x5 FILLER_216_851 ();
 b15zdnd00an1n02x5 FILLER_216_855 ();
 b15zdnd11an1n04x5 FILLER_216_875 ();
 b15zdnd11an1n16x5 FILLER_216_891 ();
 b15zdnd11an1n04x5 FILLER_216_913 ();
 b15zdnd00an1n02x5 FILLER_216_917 ();
 b15zdnd00an1n01x5 FILLER_216_919 ();
 b15zdnd11an1n08x5 FILLER_216_924 ();
 b15zdnd11an1n32x5 FILLER_216_937 ();
 b15zdnd00an1n01x5 FILLER_216_969 ();
 b15zdnd11an1n32x5 FILLER_216_979 ();
 b15zdnd11an1n16x5 FILLER_216_1011 ();
 b15zdnd11an1n08x5 FILLER_216_1027 ();
 b15zdnd00an1n02x5 FILLER_216_1035 ();
 b15zdnd00an1n01x5 FILLER_216_1037 ();
 b15zdnd11an1n16x5 FILLER_216_1043 ();
 b15zdnd00an1n01x5 FILLER_216_1059 ();
 b15zdnd11an1n08x5 FILLER_216_1064 ();
 b15zdnd00an1n02x5 FILLER_216_1072 ();
 b15zdnd00an1n01x5 FILLER_216_1074 ();
 b15zdnd11an1n16x5 FILLER_216_1086 ();
 b15zdnd11an1n04x5 FILLER_216_1102 ();
 b15zdnd00an1n01x5 FILLER_216_1106 ();
 b15zdnd11an1n16x5 FILLER_216_1117 ();
 b15zdnd11an1n08x5 FILLER_216_1133 ();
 b15zdnd00an1n02x5 FILLER_216_1141 ();
 b15zdnd11an1n08x5 FILLER_216_1155 ();
 b15zdnd00an1n01x5 FILLER_216_1163 ();
 b15zdnd11an1n16x5 FILLER_216_1169 ();
 b15zdnd11an1n08x5 FILLER_216_1185 ();
 b15zdnd00an1n01x5 FILLER_216_1193 ();
 b15zdnd11an1n64x5 FILLER_216_1220 ();
 b15zdnd00an1n02x5 FILLER_216_1284 ();
 b15zdnd00an1n01x5 FILLER_216_1286 ();
 b15zdnd11an1n32x5 FILLER_216_1293 ();
 b15zdnd11an1n08x5 FILLER_216_1325 ();
 b15zdnd00an1n01x5 FILLER_216_1333 ();
 b15zdnd11an1n08x5 FILLER_216_1345 ();
 b15zdnd00an1n01x5 FILLER_216_1353 ();
 b15zdnd11an1n16x5 FILLER_216_1374 ();
 b15zdnd11an1n32x5 FILLER_216_1394 ();
 b15zdnd00an1n01x5 FILLER_216_1426 ();
 b15zdnd11an1n04x5 FILLER_216_1431 ();
 b15zdnd11an1n32x5 FILLER_216_1440 ();
 b15zdnd11an1n16x5 FILLER_216_1472 ();
 b15zdnd11an1n16x5 FILLER_216_1496 ();
 b15zdnd11an1n08x5 FILLER_216_1512 ();
 b15zdnd11an1n04x5 FILLER_216_1520 ();
 b15zdnd00an1n02x5 FILLER_216_1524 ();
 b15zdnd11an1n04x5 FILLER_216_1542 ();
 b15zdnd11an1n16x5 FILLER_216_1558 ();
 b15zdnd11an1n08x5 FILLER_216_1574 ();
 b15zdnd11an1n04x5 FILLER_216_1582 ();
 b15zdnd00an1n01x5 FILLER_216_1586 ();
 b15zdnd11an1n64x5 FILLER_216_1593 ();
 b15zdnd11an1n04x5 FILLER_216_1662 ();
 b15zdnd00an1n02x5 FILLER_216_1666 ();
 b15zdnd11an1n32x5 FILLER_216_1675 ();
 b15zdnd11an1n16x5 FILLER_216_1707 ();
 b15zdnd00an1n02x5 FILLER_216_1723 ();
 b15zdnd00an1n01x5 FILLER_216_1725 ();
 b15zdnd11an1n16x5 FILLER_216_1736 ();
 b15zdnd11an1n08x5 FILLER_216_1752 ();
 b15zdnd11an1n04x5 FILLER_216_1760 ();
 b15zdnd00an1n01x5 FILLER_216_1764 ();
 b15zdnd11an1n08x5 FILLER_216_1777 ();
 b15zdnd00an1n02x5 FILLER_216_1785 ();
 b15zdnd11an1n04x5 FILLER_216_1802 ();
 b15zdnd11an1n04x5 FILLER_216_1837 ();
 b15zdnd11an1n08x5 FILLER_216_1860 ();
 b15zdnd11an1n04x5 FILLER_216_1868 ();
 b15zdnd11an1n16x5 FILLER_216_1892 ();
 b15zdnd00an1n02x5 FILLER_216_1908 ();
 b15zdnd00an1n01x5 FILLER_216_1910 ();
 b15zdnd11an1n32x5 FILLER_216_1931 ();
 b15zdnd11an1n16x5 FILLER_216_1963 ();
 b15zdnd00an1n02x5 FILLER_216_1979 ();
 b15zdnd11an1n04x5 FILLER_216_2002 ();
 b15zdnd11an1n04x5 FILLER_216_2012 ();
 b15zdnd11an1n16x5 FILLER_216_2021 ();
 b15zdnd11an1n08x5 FILLER_216_2037 ();
 b15zdnd00an1n02x5 FILLER_216_2045 ();
 b15zdnd11an1n32x5 FILLER_216_2067 ();
 b15zdnd00an1n01x5 FILLER_216_2099 ();
 b15zdnd11an1n16x5 FILLER_216_2104 ();
 b15zdnd11an1n08x5 FILLER_216_2120 ();
 b15zdnd00an1n02x5 FILLER_216_2128 ();
 b15zdnd00an1n02x5 FILLER_216_2152 ();
 b15zdnd11an1n16x5 FILLER_216_2162 ();
 b15zdnd11an1n04x5 FILLER_216_2178 ();
 b15zdnd00an1n01x5 FILLER_216_2182 ();
 b15zdnd11an1n04x5 FILLER_216_2203 ();
 b15zdnd11an1n08x5 FILLER_216_2227 ();
 b15zdnd00an1n02x5 FILLER_216_2235 ();
 b15zdnd00an1n01x5 FILLER_216_2237 ();
 b15zdnd11an1n04x5 FILLER_216_2242 ();
 b15zdnd11an1n04x5 FILLER_216_2250 ();
 b15zdnd11an1n04x5 FILLER_216_2262 ();
 b15zdnd11an1n04x5 FILLER_216_2270 ();
 b15zdnd00an1n02x5 FILLER_216_2274 ();
 b15zdnd11an1n32x5 FILLER_217_0 ();
 b15zdnd11an1n08x5 FILLER_217_32 ();
 b15zdnd11an1n04x5 FILLER_217_40 ();
 b15zdnd11an1n64x5 FILLER_217_62 ();
 b15zdnd11an1n64x5 FILLER_217_126 ();
 b15zdnd11an1n16x5 FILLER_217_190 ();
 b15zdnd11an1n08x5 FILLER_217_206 ();
 b15zdnd11an1n04x5 FILLER_217_214 ();
 b15zdnd00an1n02x5 FILLER_217_218 ();
 b15zdnd11an1n04x5 FILLER_217_225 ();
 b15zdnd11an1n04x5 FILLER_217_255 ();
 b15zdnd11an1n08x5 FILLER_217_264 ();
 b15zdnd00an1n02x5 FILLER_217_272 ();
 b15zdnd11an1n16x5 FILLER_217_286 ();
 b15zdnd11an1n08x5 FILLER_217_302 ();
 b15zdnd11an1n04x5 FILLER_217_310 ();
 b15zdnd00an1n01x5 FILLER_217_314 ();
 b15zdnd11an1n04x5 FILLER_217_346 ();
 b15zdnd11an1n16x5 FILLER_217_376 ();
 b15zdnd11an1n08x5 FILLER_217_392 ();
 b15zdnd00an1n02x5 FILLER_217_400 ();
 b15zdnd00an1n01x5 FILLER_217_402 ();
 b15zdnd11an1n04x5 FILLER_217_413 ();
 b15zdnd00an1n02x5 FILLER_217_417 ();
 b15zdnd11an1n08x5 FILLER_217_427 ();
 b15zdnd11an1n04x5 FILLER_217_435 ();
 b15zdnd00an1n01x5 FILLER_217_439 ();
 b15zdnd11an1n32x5 FILLER_217_456 ();
 b15zdnd00an1n02x5 FILLER_217_488 ();
 b15zdnd00an1n01x5 FILLER_217_490 ();
 b15zdnd11an1n16x5 FILLER_217_513 ();
 b15zdnd00an1n02x5 FILLER_217_529 ();
 b15zdnd00an1n01x5 FILLER_217_531 ();
 b15zdnd11an1n08x5 FILLER_217_537 ();
 b15zdnd00an1n02x5 FILLER_217_545 ();
 b15zdnd00an1n01x5 FILLER_217_547 ();
 b15zdnd11an1n04x5 FILLER_217_574 ();
 b15zdnd11an1n32x5 FILLER_217_588 ();
 b15zdnd11an1n08x5 FILLER_217_620 ();
 b15zdnd11an1n04x5 FILLER_217_628 ();
 b15zdnd00an1n01x5 FILLER_217_632 ();
 b15zdnd11an1n08x5 FILLER_217_637 ();
 b15zdnd00an1n02x5 FILLER_217_645 ();
 b15zdnd00an1n01x5 FILLER_217_647 ();
 b15zdnd11an1n08x5 FILLER_217_660 ();
 b15zdnd00an1n02x5 FILLER_217_668 ();
 b15zdnd11an1n04x5 FILLER_217_678 ();
 b15zdnd11an1n32x5 FILLER_217_688 ();
 b15zdnd11an1n16x5 FILLER_217_720 ();
 b15zdnd00an1n01x5 FILLER_217_736 ();
 b15zdnd11an1n04x5 FILLER_217_749 ();
 b15zdnd11an1n04x5 FILLER_217_765 ();
 b15zdnd11an1n64x5 FILLER_217_789 ();
 b15zdnd11an1n08x5 FILLER_217_853 ();
 b15zdnd11an1n04x5 FILLER_217_861 ();
 b15zdnd00an1n02x5 FILLER_217_865 ();
 b15zdnd00an1n01x5 FILLER_217_867 ();
 b15zdnd11an1n16x5 FILLER_217_878 ();
 b15zdnd11an1n64x5 FILLER_217_900 ();
 b15zdnd11an1n16x5 FILLER_217_964 ();
 b15zdnd00an1n02x5 FILLER_217_980 ();
 b15zdnd00an1n01x5 FILLER_217_982 ();
 b15zdnd11an1n16x5 FILLER_217_988 ();
 b15zdnd00an1n02x5 FILLER_217_1004 ();
 b15zdnd00an1n01x5 FILLER_217_1006 ();
 b15zdnd11an1n08x5 FILLER_217_1025 ();
 b15zdnd00an1n02x5 FILLER_217_1033 ();
 b15zdnd11an1n32x5 FILLER_217_1040 ();
 b15zdnd11an1n16x5 FILLER_217_1072 ();
 b15zdnd11an1n04x5 FILLER_217_1088 ();
 b15zdnd00an1n02x5 FILLER_217_1092 ();
 b15zdnd00an1n01x5 FILLER_217_1094 ();
 b15zdnd11an1n32x5 FILLER_217_1101 ();
 b15zdnd00an1n02x5 FILLER_217_1133 ();
 b15zdnd00an1n01x5 FILLER_217_1135 ();
 b15zdnd11an1n16x5 FILLER_217_1141 ();
 b15zdnd00an1n02x5 FILLER_217_1157 ();
 b15zdnd11an1n08x5 FILLER_217_1177 ();
 b15zdnd11an1n04x5 FILLER_217_1185 ();
 b15zdnd00an1n01x5 FILLER_217_1189 ();
 b15zdnd11an1n64x5 FILLER_217_1198 ();
 b15zdnd11an1n16x5 FILLER_217_1262 ();
 b15zdnd00an1n01x5 FILLER_217_1278 ();
 b15zdnd11an1n04x5 FILLER_217_1286 ();
 b15zdnd11an1n16x5 FILLER_217_1294 ();
 b15zdnd00an1n01x5 FILLER_217_1310 ();
 b15zdnd11an1n04x5 FILLER_217_1320 ();
 b15zdnd11an1n16x5 FILLER_217_1337 ();
 b15zdnd11an1n04x5 FILLER_217_1369 ();
 b15zdnd11an1n04x5 FILLER_217_1383 ();
 b15zdnd11an1n16x5 FILLER_217_1399 ();
 b15zdnd11an1n08x5 FILLER_217_1415 ();
 b15zdnd11an1n04x5 FILLER_217_1423 ();
 b15zdnd00an1n01x5 FILLER_217_1427 ();
 b15zdnd11an1n64x5 FILLER_217_1435 ();
 b15zdnd11an1n32x5 FILLER_217_1499 ();
 b15zdnd11an1n08x5 FILLER_217_1531 ();
 b15zdnd11an1n04x5 FILLER_217_1539 ();
 b15zdnd11an1n04x5 FILLER_217_1550 ();
 b15zdnd00an1n02x5 FILLER_217_1554 ();
 b15zdnd00an1n01x5 FILLER_217_1556 ();
 b15zdnd11an1n64x5 FILLER_217_1569 ();
 b15zdnd11an1n32x5 FILLER_217_1633 ();
 b15zdnd11an1n08x5 FILLER_217_1665 ();
 b15zdnd00an1n01x5 FILLER_217_1673 ();
 b15zdnd11an1n64x5 FILLER_217_1681 ();
 b15zdnd11an1n16x5 FILLER_217_1745 ();
 b15zdnd11an1n04x5 FILLER_217_1761 ();
 b15zdnd11an1n32x5 FILLER_217_1774 ();
 b15zdnd11an1n16x5 FILLER_217_1806 ();
 b15zdnd11an1n08x5 FILLER_217_1822 ();
 b15zdnd11an1n04x5 FILLER_217_1830 ();
 b15zdnd00an1n02x5 FILLER_217_1834 ();
 b15zdnd00an1n01x5 FILLER_217_1836 ();
 b15zdnd11an1n04x5 FILLER_217_1868 ();
 b15zdnd11an1n16x5 FILLER_217_1883 ();
 b15zdnd00an1n01x5 FILLER_217_1899 ();
 b15zdnd11an1n08x5 FILLER_217_1912 ();
 b15zdnd11an1n04x5 FILLER_217_1920 ();
 b15zdnd11an1n64x5 FILLER_217_1929 ();
 b15zdnd11an1n08x5 FILLER_217_1993 ();
 b15zdnd11an1n04x5 FILLER_217_2001 ();
 b15zdnd11an1n32x5 FILLER_217_2012 ();
 b15zdnd11an1n16x5 FILLER_217_2044 ();
 b15zdnd11an1n04x5 FILLER_217_2060 ();
 b15zdnd00an1n01x5 FILLER_217_2064 ();
 b15zdnd11an1n64x5 FILLER_217_2068 ();
 b15zdnd11an1n08x5 FILLER_217_2132 ();
 b15zdnd00an1n01x5 FILLER_217_2140 ();
 b15zdnd11an1n16x5 FILLER_217_2166 ();
 b15zdnd11an1n08x5 FILLER_217_2182 ();
 b15zdnd00an1n01x5 FILLER_217_2190 ();
 b15zdnd11an1n08x5 FILLER_217_2196 ();
 b15zdnd00an1n02x5 FILLER_217_2204 ();
 b15zdnd11an1n08x5 FILLER_217_2211 ();
 b15zdnd00an1n01x5 FILLER_217_2219 ();
 b15zdnd11an1n08x5 FILLER_217_2223 ();
 b15zdnd00an1n01x5 FILLER_217_2231 ();
 b15zdnd11an1n08x5 FILLER_217_2236 ();
 b15zdnd11an1n04x5 FILLER_217_2244 ();
 b15zdnd11an1n04x5 FILLER_217_2253 ();
 b15zdnd11an1n08x5 FILLER_217_2261 ();
 b15zdnd11an1n04x5 FILLER_217_2269 ();
 b15zdnd00an1n02x5 FILLER_217_2273 ();
 b15zdnd11an1n04x5 FILLER_217_2279 ();
 b15zdnd00an1n01x5 FILLER_217_2283 ();
 b15zdnd11an1n32x5 FILLER_218_8 ();
 b15zdnd11an1n16x5 FILLER_218_40 ();
 b15zdnd00an1n01x5 FILLER_218_56 ();
 b15zdnd11an1n32x5 FILLER_218_61 ();
 b15zdnd11an1n08x5 FILLER_218_93 ();
 b15zdnd00an1n01x5 FILLER_218_101 ();
 b15zdnd11an1n64x5 FILLER_218_118 ();
 b15zdnd11an1n08x5 FILLER_218_182 ();
 b15zdnd11an1n04x5 FILLER_218_190 ();
 b15zdnd11an1n16x5 FILLER_218_198 ();
 b15zdnd11an1n04x5 FILLER_218_214 ();
 b15zdnd00an1n02x5 FILLER_218_218 ();
 b15zdnd11an1n16x5 FILLER_218_229 ();
 b15zdnd11an1n04x5 FILLER_218_245 ();
 b15zdnd00an1n01x5 FILLER_218_249 ();
 b15zdnd11an1n08x5 FILLER_218_256 ();
 b15zdnd11an1n04x5 FILLER_218_264 ();
 b15zdnd00an1n02x5 FILLER_218_268 ();
 b15zdnd00an1n01x5 FILLER_218_270 ();
 b15zdnd11an1n16x5 FILLER_218_276 ();
 b15zdnd11an1n16x5 FILLER_218_301 ();
 b15zdnd11an1n08x5 FILLER_218_317 ();
 b15zdnd00an1n02x5 FILLER_218_325 ();
 b15zdnd00an1n01x5 FILLER_218_327 ();
 b15zdnd11an1n32x5 FILLER_218_354 ();
 b15zdnd11an1n08x5 FILLER_218_386 ();
 b15zdnd11an1n04x5 FILLER_218_394 ();
 b15zdnd00an1n01x5 FILLER_218_398 ();
 b15zdnd11an1n16x5 FILLER_218_406 ();
 b15zdnd11an1n08x5 FILLER_218_422 ();
 b15zdnd11an1n04x5 FILLER_218_451 ();
 b15zdnd11an1n04x5 FILLER_218_486 ();
 b15zdnd00an1n01x5 FILLER_218_490 ();
 b15zdnd11an1n08x5 FILLER_218_507 ();
 b15zdnd00an1n01x5 FILLER_218_515 ();
 b15zdnd11an1n08x5 FILLER_218_526 ();
 b15zdnd11an1n04x5 FILLER_218_534 ();
 b15zdnd00an1n02x5 FILLER_218_538 ();
 b15zdnd00an1n01x5 FILLER_218_540 ();
 b15zdnd11an1n32x5 FILLER_218_545 ();
 b15zdnd11an1n04x5 FILLER_218_577 ();
 b15zdnd00an1n01x5 FILLER_218_581 ();
 b15zdnd11an1n16x5 FILLER_218_597 ();
 b15zdnd11an1n08x5 FILLER_218_613 ();
 b15zdnd11an1n04x5 FILLER_218_625 ();
 b15zdnd00an1n02x5 FILLER_218_629 ();
 b15zdnd00an1n01x5 FILLER_218_631 ();
 b15zdnd11an1n08x5 FILLER_218_640 ();
 b15zdnd00an1n02x5 FILLER_218_648 ();
 b15zdnd11an1n08x5 FILLER_218_662 ();
 b15zdnd11an1n04x5 FILLER_218_670 ();
 b15zdnd11an1n04x5 FILLER_218_683 ();
 b15zdnd11an1n08x5 FILLER_218_707 ();
 b15zdnd00an1n02x5 FILLER_218_715 ();
 b15zdnd00an1n01x5 FILLER_218_717 ();
 b15zdnd00an1n02x5 FILLER_218_726 ();
 b15zdnd11an1n64x5 FILLER_218_748 ();
 b15zdnd11an1n64x5 FILLER_218_812 ();
 b15zdnd11an1n08x5 FILLER_218_876 ();
 b15zdnd00an1n02x5 FILLER_218_884 ();
 b15zdnd11an1n64x5 FILLER_218_892 ();
 b15zdnd00an1n02x5 FILLER_218_956 ();
 b15zdnd00an1n01x5 FILLER_218_958 ();
 b15zdnd11an1n08x5 FILLER_218_968 ();
 b15zdnd11an1n04x5 FILLER_218_976 ();
 b15zdnd11an1n16x5 FILLER_218_992 ();
 b15zdnd11an1n64x5 FILLER_218_1024 ();
 b15zdnd11an1n32x5 FILLER_218_1088 ();
 b15zdnd11an1n16x5 FILLER_218_1120 ();
 b15zdnd11an1n08x5 FILLER_218_1152 ();
 b15zdnd00an1n02x5 FILLER_218_1160 ();
 b15zdnd11an1n08x5 FILLER_218_1166 ();
 b15zdnd11an1n04x5 FILLER_218_1174 ();
 b15zdnd00an1n02x5 FILLER_218_1178 ();
 b15zdnd00an1n01x5 FILLER_218_1180 ();
 b15zdnd11an1n08x5 FILLER_218_1213 ();
 b15zdnd00an1n01x5 FILLER_218_1221 ();
 b15zdnd11an1n32x5 FILLER_218_1242 ();
 b15zdnd11an1n08x5 FILLER_218_1274 ();
 b15zdnd00an1n02x5 FILLER_218_1282 ();
 b15zdnd11an1n04x5 FILLER_218_1289 ();
 b15zdnd11an1n64x5 FILLER_218_1312 ();
 b15zdnd11an1n08x5 FILLER_218_1376 ();
 b15zdnd11an1n16x5 FILLER_218_1390 ();
 b15zdnd00an1n02x5 FILLER_218_1406 ();
 b15zdnd11an1n16x5 FILLER_218_1426 ();
 b15zdnd11an1n04x5 FILLER_218_1442 ();
 b15zdnd00an1n02x5 FILLER_218_1446 ();
 b15zdnd00an1n01x5 FILLER_218_1448 ();
 b15zdnd11an1n04x5 FILLER_218_1456 ();
 b15zdnd11an1n08x5 FILLER_218_1466 ();
 b15zdnd00an1n01x5 FILLER_218_1474 ();
 b15zdnd11an1n64x5 FILLER_218_1481 ();
 b15zdnd11an1n16x5 FILLER_218_1545 ();
 b15zdnd00an1n02x5 FILLER_218_1561 ();
 b15zdnd11an1n16x5 FILLER_218_1577 ();
 b15zdnd11an1n08x5 FILLER_218_1593 ();
 b15zdnd11an1n04x5 FILLER_218_1601 ();
 b15zdnd00an1n02x5 FILLER_218_1605 ();
 b15zdnd11an1n04x5 FILLER_218_1612 ();
 b15zdnd11an1n32x5 FILLER_218_1628 ();
 b15zdnd11an1n16x5 FILLER_218_1660 ();
 b15zdnd11an1n08x5 FILLER_218_1676 ();
 b15zdnd00an1n01x5 FILLER_218_1684 ();
 b15zdnd11an1n32x5 FILLER_218_1694 ();
 b15zdnd11an1n08x5 FILLER_218_1726 ();
 b15zdnd00an1n02x5 FILLER_218_1734 ();
 b15zdnd11an1n64x5 FILLER_218_1751 ();
 b15zdnd11an1n32x5 FILLER_218_1815 ();
 b15zdnd11an1n16x5 FILLER_218_1847 ();
 b15zdnd11an1n32x5 FILLER_218_1894 ();
 b15zdnd11an1n16x5 FILLER_218_1926 ();
 b15zdnd11an1n04x5 FILLER_218_1942 ();
 b15zdnd00an1n02x5 FILLER_218_1946 ();
 b15zdnd00an1n01x5 FILLER_218_1948 ();
 b15zdnd11an1n64x5 FILLER_218_1954 ();
 b15zdnd11an1n64x5 FILLER_218_2018 ();
 b15zdnd11an1n64x5 FILLER_218_2082 ();
 b15zdnd11an1n08x5 FILLER_218_2146 ();
 b15zdnd11an1n64x5 FILLER_218_2162 ();
 b15zdnd11an1n16x5 FILLER_218_2226 ();
 b15zdnd11an1n08x5 FILLER_218_2242 ();
 b15zdnd11an1n04x5 FILLER_218_2250 ();
 b15zdnd11an1n04x5 FILLER_218_2258 ();
 b15zdnd11an1n08x5 FILLER_218_2267 ();
 b15zdnd00an1n01x5 FILLER_218_2275 ();
 b15zdnd11an1n32x5 FILLER_219_0 ();
 b15zdnd11an1n16x5 FILLER_219_32 ();
 b15zdnd11an1n04x5 FILLER_219_48 ();
 b15zdnd00an1n02x5 FILLER_219_52 ();
 b15zdnd00an1n01x5 FILLER_219_54 ();
 b15zdnd11an1n04x5 FILLER_219_73 ();
 b15zdnd00an1n01x5 FILLER_219_77 ();
 b15zdnd11an1n04x5 FILLER_219_83 ();
 b15zdnd11an1n08x5 FILLER_219_95 ();
 b15zdnd11an1n04x5 FILLER_219_103 ();
 b15zdnd00an1n02x5 FILLER_219_107 ();
 b15zdnd11an1n08x5 FILLER_219_125 ();
 b15zdnd11an1n04x5 FILLER_219_133 ();
 b15zdnd00an1n02x5 FILLER_219_137 ();
 b15zdnd11an1n32x5 FILLER_219_144 ();
 b15zdnd11an1n08x5 FILLER_219_176 ();
 b15zdnd00an1n02x5 FILLER_219_184 ();
 b15zdnd00an1n01x5 FILLER_219_186 ();
 b15zdnd11an1n32x5 FILLER_219_193 ();
 b15zdnd11an1n16x5 FILLER_219_225 ();
 b15zdnd11an1n08x5 FILLER_219_241 ();
 b15zdnd11an1n04x5 FILLER_219_249 ();
 b15zdnd11an1n64x5 FILLER_219_263 ();
 b15zdnd11an1n16x5 FILLER_219_327 ();
 b15zdnd11an1n08x5 FILLER_219_343 ();
 b15zdnd11an1n04x5 FILLER_219_351 ();
 b15zdnd11an1n16x5 FILLER_219_371 ();
 b15zdnd00an1n01x5 FILLER_219_387 ();
 b15zdnd11an1n32x5 FILLER_219_411 ();
 b15zdnd11an1n16x5 FILLER_219_443 ();
 b15zdnd11an1n04x5 FILLER_219_459 ();
 b15zdnd00an1n02x5 FILLER_219_463 ();
 b15zdnd11an1n08x5 FILLER_219_481 ();
 b15zdnd11an1n04x5 FILLER_219_489 ();
 b15zdnd00an1n01x5 FILLER_219_493 ();
 b15zdnd11an1n04x5 FILLER_219_504 ();
 b15zdnd11an1n08x5 FILLER_219_519 ();
 b15zdnd11an1n04x5 FILLER_219_527 ();
 b15zdnd00an1n01x5 FILLER_219_531 ();
 b15zdnd11an1n32x5 FILLER_219_537 ();
 b15zdnd11an1n08x5 FILLER_219_569 ();
 b15zdnd00an1n02x5 FILLER_219_577 ();
 b15zdnd00an1n01x5 FILLER_219_579 ();
 b15zdnd11an1n32x5 FILLER_219_587 ();
 b15zdnd11an1n16x5 FILLER_219_619 ();
 b15zdnd00an1n02x5 FILLER_219_635 ();
 b15zdnd11an1n04x5 FILLER_219_646 ();
 b15zdnd00an1n02x5 FILLER_219_650 ();
 b15zdnd00an1n01x5 FILLER_219_652 ();
 b15zdnd11an1n64x5 FILLER_219_659 ();
 b15zdnd11an1n04x5 FILLER_219_723 ();
 b15zdnd00an1n02x5 FILLER_219_727 ();
 b15zdnd11an1n64x5 FILLER_219_755 ();
 b15zdnd11an1n08x5 FILLER_219_819 ();
 b15zdnd11an1n04x5 FILLER_219_827 ();
 b15zdnd00an1n02x5 FILLER_219_831 ();
 b15zdnd00an1n01x5 FILLER_219_833 ();
 b15zdnd11an1n08x5 FILLER_219_843 ();
 b15zdnd11an1n04x5 FILLER_219_851 ();
 b15zdnd00an1n01x5 FILLER_219_855 ();
 b15zdnd11an1n64x5 FILLER_219_870 ();
 b15zdnd00an1n01x5 FILLER_219_934 ();
 b15zdnd11an1n32x5 FILLER_219_941 ();
 b15zdnd11an1n04x5 FILLER_219_973 ();
 b15zdnd00an1n02x5 FILLER_219_977 ();
 b15zdnd00an1n01x5 FILLER_219_979 ();
 b15zdnd11an1n16x5 FILLER_219_985 ();
 b15zdnd11an1n08x5 FILLER_219_1001 ();
 b15zdnd11an1n04x5 FILLER_219_1009 ();
 b15zdnd11an1n04x5 FILLER_219_1033 ();
 b15zdnd11an1n64x5 FILLER_219_1053 ();
 b15zdnd11an1n64x5 FILLER_219_1117 ();
 b15zdnd00an1n02x5 FILLER_219_1181 ();
 b15zdnd11an1n04x5 FILLER_219_1199 ();
 b15zdnd11an1n64x5 FILLER_219_1221 ();
 b15zdnd11an1n16x5 FILLER_219_1285 ();
 b15zdnd11an1n04x5 FILLER_219_1301 ();
 b15zdnd00an1n02x5 FILLER_219_1305 ();
 b15zdnd11an1n64x5 FILLER_219_1327 ();
 b15zdnd11an1n32x5 FILLER_219_1391 ();
 b15zdnd11an1n16x5 FILLER_219_1423 ();
 b15zdnd11an1n04x5 FILLER_219_1439 ();
 b15zdnd00an1n02x5 FILLER_219_1443 ();
 b15zdnd00an1n01x5 FILLER_219_1445 ();
 b15zdnd11an1n08x5 FILLER_219_1453 ();
 b15zdnd11an1n04x5 FILLER_219_1461 ();
 b15zdnd00an1n01x5 FILLER_219_1465 ();
 b15zdnd11an1n16x5 FILLER_219_1472 ();
 b15zdnd11an1n08x5 FILLER_219_1488 ();
 b15zdnd11an1n04x5 FILLER_219_1496 ();
 b15zdnd00an1n01x5 FILLER_219_1500 ();
 b15zdnd11an1n16x5 FILLER_219_1512 ();
 b15zdnd11an1n08x5 FILLER_219_1528 ();
 b15zdnd11an1n04x5 FILLER_219_1536 ();
 b15zdnd11an1n08x5 FILLER_219_1546 ();
 b15zdnd00an1n02x5 FILLER_219_1554 ();
 b15zdnd00an1n01x5 FILLER_219_1556 ();
 b15zdnd11an1n32x5 FILLER_219_1563 ();
 b15zdnd11an1n16x5 FILLER_219_1595 ();
 b15zdnd00an1n02x5 FILLER_219_1611 ();
 b15zdnd00an1n01x5 FILLER_219_1613 ();
 b15zdnd11an1n32x5 FILLER_219_1620 ();
 b15zdnd11an1n16x5 FILLER_219_1652 ();
 b15zdnd11an1n04x5 FILLER_219_1668 ();
 b15zdnd00an1n02x5 FILLER_219_1672 ();
 b15zdnd11an1n64x5 FILLER_219_1681 ();
 b15zdnd11an1n16x5 FILLER_219_1745 ();
 b15zdnd11an1n04x5 FILLER_219_1761 ();
 b15zdnd00an1n01x5 FILLER_219_1765 ();
 b15zdnd11an1n64x5 FILLER_219_1786 ();
 b15zdnd11an1n64x5 FILLER_219_1850 ();
 b15zdnd11an1n32x5 FILLER_219_1914 ();
 b15zdnd11an1n04x5 FILLER_219_1946 ();
 b15zdnd11an1n64x5 FILLER_219_1970 ();
 b15zdnd11an1n32x5 FILLER_219_2034 ();
 b15zdnd11an1n08x5 FILLER_219_2066 ();
 b15zdnd11an1n32x5 FILLER_219_2079 ();
 b15zdnd00an1n02x5 FILLER_219_2111 ();
 b15zdnd00an1n01x5 FILLER_219_2113 ();
 b15zdnd11an1n64x5 FILLER_219_2134 ();
 b15zdnd11an1n32x5 FILLER_219_2198 ();
 b15zdnd11an1n16x5 FILLER_219_2230 ();
 b15zdnd11an1n08x5 FILLER_219_2246 ();
 b15zdnd00an1n02x5 FILLER_219_2254 ();
 b15zdnd11an1n16x5 FILLER_219_2260 ();
 b15zdnd00an1n01x5 FILLER_219_2276 ();
 b15zdnd00an1n02x5 FILLER_219_2282 ();
 b15zdnd11an1n32x5 FILLER_220_8 ();
 b15zdnd11an1n04x5 FILLER_220_40 ();
 b15zdnd00an1n02x5 FILLER_220_44 ();
 b15zdnd00an1n01x5 FILLER_220_46 ();
 b15zdnd11an1n04x5 FILLER_220_54 ();
 b15zdnd11an1n16x5 FILLER_220_74 ();
 b15zdnd11an1n08x5 FILLER_220_90 ();
 b15zdnd11an1n04x5 FILLER_220_98 ();
 b15zdnd11an1n16x5 FILLER_220_107 ();
 b15zdnd00an1n02x5 FILLER_220_123 ();
 b15zdnd00an1n01x5 FILLER_220_125 ();
 b15zdnd11an1n04x5 FILLER_220_131 ();
 b15zdnd11an1n04x5 FILLER_220_145 ();
 b15zdnd11an1n04x5 FILLER_220_153 ();
 b15zdnd00an1n02x5 FILLER_220_157 ();
 b15zdnd00an1n01x5 FILLER_220_159 ();
 b15zdnd11an1n08x5 FILLER_220_165 ();
 b15zdnd00an1n01x5 FILLER_220_173 ();
 b15zdnd11an1n64x5 FILLER_220_186 ();
 b15zdnd11an1n32x5 FILLER_220_250 ();
 b15zdnd11an1n16x5 FILLER_220_282 ();
 b15zdnd11an1n08x5 FILLER_220_305 ();
 b15zdnd11an1n04x5 FILLER_220_313 ();
 b15zdnd00an1n01x5 FILLER_220_317 ();
 b15zdnd11an1n64x5 FILLER_220_326 ();
 b15zdnd11an1n64x5 FILLER_220_390 ();
 b15zdnd11an1n32x5 FILLER_220_454 ();
 b15zdnd11an1n16x5 FILLER_220_486 ();
 b15zdnd00an1n02x5 FILLER_220_502 ();
 b15zdnd00an1n01x5 FILLER_220_504 ();
 b15zdnd11an1n64x5 FILLER_220_515 ();
 b15zdnd11an1n64x5 FILLER_220_579 ();
 b15zdnd11an1n64x5 FILLER_220_643 ();
 b15zdnd11an1n08x5 FILLER_220_707 ();
 b15zdnd00an1n02x5 FILLER_220_715 ();
 b15zdnd00an1n01x5 FILLER_220_717 ();
 b15zdnd11an1n16x5 FILLER_220_726 ();
 b15zdnd11an1n08x5 FILLER_220_742 ();
 b15zdnd00an1n01x5 FILLER_220_750 ();
 b15zdnd11an1n64x5 FILLER_220_777 ();
 b15zdnd11an1n08x5 FILLER_220_841 ();
 b15zdnd00an1n02x5 FILLER_220_849 ();
 b15zdnd11an1n32x5 FILLER_220_869 ();
 b15zdnd11an1n16x5 FILLER_220_901 ();
 b15zdnd11an1n16x5 FILLER_220_923 ();
 b15zdnd11an1n08x5 FILLER_220_939 ();
 b15zdnd11an1n16x5 FILLER_220_961 ();
 b15zdnd11an1n04x5 FILLER_220_977 ();
 b15zdnd00an1n01x5 FILLER_220_981 ();
 b15zdnd11an1n64x5 FILLER_220_986 ();
 b15zdnd11an1n16x5 FILLER_220_1050 ();
 b15zdnd11an1n04x5 FILLER_220_1066 ();
 b15zdnd00an1n02x5 FILLER_220_1070 ();
 b15zdnd11an1n64x5 FILLER_220_1082 ();
 b15zdnd11an1n64x5 FILLER_220_1146 ();
 b15zdnd11an1n64x5 FILLER_220_1210 ();
 b15zdnd11an1n04x5 FILLER_220_1274 ();
 b15zdnd00an1n02x5 FILLER_220_1278 ();
 b15zdnd11an1n04x5 FILLER_220_1300 ();
 b15zdnd11an1n08x5 FILLER_220_1319 ();
 b15zdnd00an1n02x5 FILLER_220_1327 ();
 b15zdnd11an1n08x5 FILLER_220_1342 ();
 b15zdnd11an1n04x5 FILLER_220_1350 ();
 b15zdnd00an1n02x5 FILLER_220_1354 ();
 b15zdnd11an1n08x5 FILLER_220_1370 ();
 b15zdnd11an1n04x5 FILLER_220_1378 ();
 b15zdnd00an1n02x5 FILLER_220_1382 ();
 b15zdnd00an1n01x5 FILLER_220_1384 ();
 b15zdnd11an1n32x5 FILLER_220_1394 ();
 b15zdnd11an1n16x5 FILLER_220_1426 ();
 b15zdnd11an1n04x5 FILLER_220_1442 ();
 b15zdnd00an1n02x5 FILLER_220_1446 ();
 b15zdnd11an1n04x5 FILLER_220_1452 ();
 b15zdnd00an1n01x5 FILLER_220_1456 ();
 b15zdnd11an1n32x5 FILLER_220_1461 ();
 b15zdnd11an1n08x5 FILLER_220_1493 ();
 b15zdnd11an1n04x5 FILLER_220_1501 ();
 b15zdnd00an1n01x5 FILLER_220_1505 ();
 b15zdnd11an1n08x5 FILLER_220_1522 ();
 b15zdnd11an1n04x5 FILLER_220_1530 ();
 b15zdnd11an1n32x5 FILLER_220_1552 ();
 b15zdnd11an1n08x5 FILLER_220_1584 ();
 b15zdnd11an1n64x5 FILLER_220_1604 ();
 b15zdnd11an1n08x5 FILLER_220_1668 ();
 b15zdnd00an1n02x5 FILLER_220_1676 ();
 b15zdnd00an1n01x5 FILLER_220_1678 ();
 b15zdnd11an1n64x5 FILLER_220_1688 ();
 b15zdnd11an1n32x5 FILLER_220_1752 ();
 b15zdnd11an1n16x5 FILLER_220_1784 ();
 b15zdnd11an1n04x5 FILLER_220_1800 ();
 b15zdnd11an1n64x5 FILLER_220_1825 ();
 b15zdnd11an1n32x5 FILLER_220_1889 ();
 b15zdnd11an1n16x5 FILLER_220_1921 ();
 b15zdnd11an1n08x5 FILLER_220_1937 ();
 b15zdnd00an1n02x5 FILLER_220_1945 ();
 b15zdnd11an1n64x5 FILLER_220_1967 ();
 b15zdnd11an1n08x5 FILLER_220_2031 ();
 b15zdnd00an1n02x5 FILLER_220_2039 ();
 b15zdnd00an1n01x5 FILLER_220_2041 ();
 b15zdnd11an1n16x5 FILLER_220_2046 ();
 b15zdnd11an1n08x5 FILLER_220_2062 ();
 b15zdnd11an1n04x5 FILLER_220_2070 ();
 b15zdnd00an1n01x5 FILLER_220_2074 ();
 b15zdnd11an1n32x5 FILLER_220_2095 ();
 b15zdnd11an1n16x5 FILLER_220_2127 ();
 b15zdnd11an1n08x5 FILLER_220_2143 ();
 b15zdnd00an1n02x5 FILLER_220_2151 ();
 b15zdnd00an1n01x5 FILLER_220_2153 ();
 b15zdnd11an1n16x5 FILLER_220_2162 ();
 b15zdnd11an1n08x5 FILLER_220_2178 ();
 b15zdnd11an1n04x5 FILLER_220_2186 ();
 b15zdnd00an1n02x5 FILLER_220_2190 ();
 b15zdnd00an1n01x5 FILLER_220_2192 ();
 b15zdnd11an1n32x5 FILLER_220_2197 ();
 b15zdnd11an1n08x5 FILLER_220_2229 ();
 b15zdnd11an1n04x5 FILLER_220_2237 ();
 b15zdnd00an1n01x5 FILLER_220_2241 ();
 b15zdnd11an1n04x5 FILLER_220_2246 ();
 b15zdnd11an1n04x5 FILLER_220_2256 ();
 b15zdnd11an1n04x5 FILLER_220_2266 ();
 b15zdnd00an1n02x5 FILLER_220_2274 ();
 b15zdnd11an1n32x5 FILLER_221_0 ();
 b15zdnd11an1n16x5 FILLER_221_32 ();
 b15zdnd11an1n08x5 FILLER_221_48 ();
 b15zdnd11an1n04x5 FILLER_221_56 ();
 b15zdnd11an1n08x5 FILLER_221_74 ();
 b15zdnd11an1n04x5 FILLER_221_82 ();
 b15zdnd00an1n02x5 FILLER_221_86 ();
 b15zdnd00an1n01x5 FILLER_221_88 ();
 b15zdnd11an1n08x5 FILLER_221_102 ();
 b15zdnd00an1n02x5 FILLER_221_110 ();
 b15zdnd11an1n08x5 FILLER_221_117 ();
 b15zdnd00an1n02x5 FILLER_221_125 ();
 b15zdnd11an1n04x5 FILLER_221_153 ();
 b15zdnd11an1n32x5 FILLER_221_164 ();
 b15zdnd11an1n08x5 FILLER_221_196 ();
 b15zdnd00an1n01x5 FILLER_221_204 ();
 b15zdnd11an1n64x5 FILLER_221_214 ();
 b15zdnd11an1n16x5 FILLER_221_278 ();
 b15zdnd00an1n02x5 FILLER_221_294 ();
 b15zdnd00an1n01x5 FILLER_221_296 ();
 b15zdnd11an1n08x5 FILLER_221_312 ();
 b15zdnd11an1n04x5 FILLER_221_320 ();
 b15zdnd11an1n04x5 FILLER_221_329 ();
 b15zdnd11an1n64x5 FILLER_221_359 ();
 b15zdnd11an1n64x5 FILLER_221_423 ();
 b15zdnd11an1n64x5 FILLER_221_487 ();
 b15zdnd11an1n64x5 FILLER_221_551 ();
 b15zdnd11an1n64x5 FILLER_221_615 ();
 b15zdnd11an1n32x5 FILLER_221_679 ();
 b15zdnd11an1n16x5 FILLER_221_711 ();
 b15zdnd11an1n04x5 FILLER_221_727 ();
 b15zdnd11an1n16x5 FILLER_221_751 ();
 b15zdnd11an1n08x5 FILLER_221_767 ();
 b15zdnd11an1n04x5 FILLER_221_775 ();
 b15zdnd00an1n02x5 FILLER_221_779 ();
 b15zdnd00an1n01x5 FILLER_221_781 ();
 b15zdnd11an1n64x5 FILLER_221_802 ();
 b15zdnd11an1n16x5 FILLER_221_866 ();
 b15zdnd00an1n01x5 FILLER_221_882 ();
 b15zdnd11an1n08x5 FILLER_221_891 ();
 b15zdnd11an1n04x5 FILLER_221_899 ();
 b15zdnd00an1n01x5 FILLER_221_903 ();
 b15zdnd11an1n04x5 FILLER_221_915 ();
 b15zdnd11an1n08x5 FILLER_221_926 ();
 b15zdnd11an1n64x5 FILLER_221_940 ();
 b15zdnd11an1n16x5 FILLER_221_1004 ();
 b15zdnd11an1n08x5 FILLER_221_1020 ();
 b15zdnd11an1n04x5 FILLER_221_1028 ();
 b15zdnd00an1n02x5 FILLER_221_1032 ();
 b15zdnd00an1n01x5 FILLER_221_1034 ();
 b15zdnd11an1n16x5 FILLER_221_1041 ();
 b15zdnd11an1n08x5 FILLER_221_1057 ();
 b15zdnd11an1n32x5 FILLER_221_1073 ();
 b15zdnd11an1n08x5 FILLER_221_1105 ();
 b15zdnd00an1n02x5 FILLER_221_1113 ();
 b15zdnd11an1n04x5 FILLER_221_1131 ();
 b15zdnd11an1n16x5 FILLER_221_1139 ();
 b15zdnd11an1n64x5 FILLER_221_1186 ();
 b15zdnd11an1n32x5 FILLER_221_1250 ();
 b15zdnd11an1n16x5 FILLER_221_1282 ();
 b15zdnd11an1n04x5 FILLER_221_1298 ();
 b15zdnd00an1n02x5 FILLER_221_1302 ();
 b15zdnd11an1n04x5 FILLER_221_1317 ();
 b15zdnd11an1n16x5 FILLER_221_1334 ();
 b15zdnd11an1n04x5 FILLER_221_1350 ();
 b15zdnd00an1n02x5 FILLER_221_1354 ();
 b15zdnd11an1n08x5 FILLER_221_1372 ();
 b15zdnd00an1n02x5 FILLER_221_1380 ();
 b15zdnd11an1n04x5 FILLER_221_1388 ();
 b15zdnd11an1n32x5 FILLER_221_1398 ();
 b15zdnd11an1n16x5 FILLER_221_1430 ();
 b15zdnd00an1n02x5 FILLER_221_1446 ();
 b15zdnd00an1n01x5 FILLER_221_1448 ();
 b15zdnd11an1n32x5 FILLER_221_1455 ();
 b15zdnd00an1n01x5 FILLER_221_1487 ();
 b15zdnd11an1n64x5 FILLER_221_1498 ();
 b15zdnd11an1n08x5 FILLER_221_1562 ();
 b15zdnd11an1n32x5 FILLER_221_1576 ();
 b15zdnd11an1n08x5 FILLER_221_1608 ();
 b15zdnd11an1n04x5 FILLER_221_1616 ();
 b15zdnd11an1n04x5 FILLER_221_1625 ();
 b15zdnd11an1n04x5 FILLER_221_1639 ();
 b15zdnd11an1n16x5 FILLER_221_1650 ();
 b15zdnd11an1n08x5 FILLER_221_1666 ();
 b15zdnd11an1n04x5 FILLER_221_1674 ();
 b15zdnd11an1n32x5 FILLER_221_1682 ();
 b15zdnd11an1n08x5 FILLER_221_1714 ();
 b15zdnd00an1n02x5 FILLER_221_1722 ();
 b15zdnd00an1n01x5 FILLER_221_1724 ();
 b15zdnd11an1n32x5 FILLER_221_1734 ();
 b15zdnd11an1n08x5 FILLER_221_1766 ();
 b15zdnd11an1n04x5 FILLER_221_1774 ();
 b15zdnd11an1n04x5 FILLER_221_1810 ();
 b15zdnd11an1n04x5 FILLER_221_1834 ();
 b15zdnd00an1n01x5 FILLER_221_1838 ();
 b15zdnd11an1n08x5 FILLER_221_1859 ();
 b15zdnd11an1n64x5 FILLER_221_1893 ();
 b15zdnd11an1n16x5 FILLER_221_1957 ();
 b15zdnd00an1n02x5 FILLER_221_1973 ();
 b15zdnd11an1n04x5 FILLER_221_1995 ();
 b15zdnd11an1n04x5 FILLER_221_2004 ();
 b15zdnd11an1n08x5 FILLER_221_2029 ();
 b15zdnd11an1n04x5 FILLER_221_2037 ();
 b15zdnd00an1n01x5 FILLER_221_2041 ();
 b15zdnd11an1n16x5 FILLER_221_2067 ();
 b15zdnd00an1n02x5 FILLER_221_2083 ();
 b15zdnd11an1n64x5 FILLER_221_2095 ();
 b15zdnd11an1n08x5 FILLER_221_2159 ();
 b15zdnd11an1n04x5 FILLER_221_2167 ();
 b15zdnd00an1n01x5 FILLER_221_2171 ();
 b15zdnd11an1n04x5 FILLER_221_2181 ();
 b15zdnd11an1n04x5 FILLER_221_2190 ();
 b15zdnd00an1n02x5 FILLER_221_2194 ();
 b15zdnd11an1n64x5 FILLER_221_2201 ();
 b15zdnd11an1n04x5 FILLER_221_2269 ();
 b15zdnd11an1n04x5 FILLER_221_2277 ();
 b15zdnd00an1n02x5 FILLER_221_2281 ();
 b15zdnd00an1n01x5 FILLER_221_2283 ();
 b15zdnd11an1n32x5 FILLER_222_8 ();
 b15zdnd11an1n08x5 FILLER_222_40 ();
 b15zdnd11an1n04x5 FILLER_222_48 ();
 b15zdnd00an1n01x5 FILLER_222_52 ();
 b15zdnd11an1n32x5 FILLER_222_73 ();
 b15zdnd11an1n08x5 FILLER_222_105 ();
 b15zdnd00an1n02x5 FILLER_222_113 ();
 b15zdnd00an1n01x5 FILLER_222_115 ();
 b15zdnd11an1n32x5 FILLER_222_123 ();
 b15zdnd11an1n16x5 FILLER_222_155 ();
 b15zdnd11an1n08x5 FILLER_222_171 ();
 b15zdnd11an1n04x5 FILLER_222_179 ();
 b15zdnd00an1n02x5 FILLER_222_183 ();
 b15zdnd11an1n04x5 FILLER_222_191 ();
 b15zdnd11an1n04x5 FILLER_222_205 ();
 b15zdnd00an1n02x5 FILLER_222_209 ();
 b15zdnd11an1n32x5 FILLER_222_219 ();
 b15zdnd00an1n02x5 FILLER_222_251 ();
 b15zdnd11an1n04x5 FILLER_222_262 ();
 b15zdnd11an1n04x5 FILLER_222_270 ();
 b15zdnd11an1n16x5 FILLER_222_300 ();
 b15zdnd11an1n04x5 FILLER_222_316 ();
 b15zdnd00an1n02x5 FILLER_222_320 ();
 b15zdnd11an1n16x5 FILLER_222_329 ();
 b15zdnd11an1n08x5 FILLER_222_345 ();
 b15zdnd11an1n04x5 FILLER_222_353 ();
 b15zdnd00an1n01x5 FILLER_222_357 ();
 b15zdnd11an1n64x5 FILLER_222_384 ();
 b15zdnd11an1n64x5 FILLER_222_448 ();
 b15zdnd11an1n64x5 FILLER_222_512 ();
 b15zdnd11an1n64x5 FILLER_222_576 ();
 b15zdnd11an1n64x5 FILLER_222_640 ();
 b15zdnd11an1n08x5 FILLER_222_704 ();
 b15zdnd11an1n04x5 FILLER_222_712 ();
 b15zdnd00an1n02x5 FILLER_222_716 ();
 b15zdnd11an1n64x5 FILLER_222_726 ();
 b15zdnd11an1n64x5 FILLER_222_790 ();
 b15zdnd11an1n16x5 FILLER_222_854 ();
 b15zdnd11an1n04x5 FILLER_222_870 ();
 b15zdnd00an1n02x5 FILLER_222_874 ();
 b15zdnd11an1n04x5 FILLER_222_883 ();
 b15zdnd11an1n32x5 FILLER_222_913 ();
 b15zdnd11an1n16x5 FILLER_222_945 ();
 b15zdnd11an1n04x5 FILLER_222_968 ();
 b15zdnd11an1n16x5 FILLER_222_982 ();
 b15zdnd11an1n04x5 FILLER_222_998 ();
 b15zdnd00an1n02x5 FILLER_222_1002 ();
 b15zdnd11an1n16x5 FILLER_222_1013 ();
 b15zdnd00an1n02x5 FILLER_222_1029 ();
 b15zdnd00an1n01x5 FILLER_222_1031 ();
 b15zdnd11an1n16x5 FILLER_222_1039 ();
 b15zdnd11an1n08x5 FILLER_222_1055 ();
 b15zdnd11an1n04x5 FILLER_222_1063 ();
 b15zdnd11an1n08x5 FILLER_222_1071 ();
 b15zdnd11an1n04x5 FILLER_222_1079 ();
 b15zdnd00an1n01x5 FILLER_222_1083 ();
 b15zdnd11an1n04x5 FILLER_222_1097 ();
 b15zdnd11an1n04x5 FILLER_222_1105 ();
 b15zdnd00an1n02x5 FILLER_222_1109 ();
 b15zdnd11an1n08x5 FILLER_222_1117 ();
 b15zdnd11an1n04x5 FILLER_222_1125 ();
 b15zdnd00an1n02x5 FILLER_222_1129 ();
 b15zdnd00an1n01x5 FILLER_222_1131 ();
 b15zdnd11an1n04x5 FILLER_222_1141 ();
 b15zdnd00an1n01x5 FILLER_222_1145 ();
 b15zdnd11an1n64x5 FILLER_222_1156 ();
 b15zdnd11an1n64x5 FILLER_222_1220 ();
 b15zdnd11an1n04x5 FILLER_222_1284 ();
 b15zdnd11an1n16x5 FILLER_222_1300 ();
 b15zdnd11an1n16x5 FILLER_222_1335 ();
 b15zdnd11an1n08x5 FILLER_222_1351 ();
 b15zdnd00an1n02x5 FILLER_222_1359 ();
 b15zdnd00an1n01x5 FILLER_222_1361 ();
 b15zdnd11an1n16x5 FILLER_222_1367 ();
 b15zdnd00an1n02x5 FILLER_222_1383 ();
 b15zdnd00an1n01x5 FILLER_222_1385 ();
 b15zdnd11an1n16x5 FILLER_222_1401 ();
 b15zdnd11an1n04x5 FILLER_222_1417 ();
 b15zdnd00an1n02x5 FILLER_222_1421 ();
 b15zdnd11an1n32x5 FILLER_222_1428 ();
 b15zdnd11an1n16x5 FILLER_222_1460 ();
 b15zdnd00an1n01x5 FILLER_222_1476 ();
 b15zdnd11an1n32x5 FILLER_222_1497 ();
 b15zdnd11an1n08x5 FILLER_222_1529 ();
 b15zdnd11an1n04x5 FILLER_222_1537 ();
 b15zdnd11an1n08x5 FILLER_222_1568 ();
 b15zdnd00an1n01x5 FILLER_222_1576 ();
 b15zdnd11an1n32x5 FILLER_222_1589 ();
 b15zdnd11an1n16x5 FILLER_222_1621 ();
 b15zdnd00an1n02x5 FILLER_222_1637 ();
 b15zdnd11an1n04x5 FILLER_222_1643 ();
 b15zdnd11an1n16x5 FILLER_222_1653 ();
 b15zdnd11an1n04x5 FILLER_222_1669 ();
 b15zdnd00an1n02x5 FILLER_222_1673 ();
 b15zdnd00an1n01x5 FILLER_222_1675 ();
 b15zdnd11an1n64x5 FILLER_222_1686 ();
 b15zdnd11an1n64x5 FILLER_222_1750 ();
 b15zdnd11an1n64x5 FILLER_222_1814 ();
 b15zdnd11an1n16x5 FILLER_222_1878 ();
 b15zdnd11an1n04x5 FILLER_222_1894 ();
 b15zdnd00an1n01x5 FILLER_222_1898 ();
 b15zdnd11an1n04x5 FILLER_222_1904 ();
 b15zdnd11an1n32x5 FILLER_222_1929 ();
 b15zdnd11an1n16x5 FILLER_222_1961 ();
 b15zdnd11an1n08x5 FILLER_222_1977 ();
 b15zdnd00an1n02x5 FILLER_222_1985 ();
 b15zdnd11an1n16x5 FILLER_222_1991 ();
 b15zdnd11an1n08x5 FILLER_222_2007 ();
 b15zdnd00an1n02x5 FILLER_222_2015 ();
 b15zdnd00an1n01x5 FILLER_222_2017 ();
 b15zdnd11an1n16x5 FILLER_222_2023 ();
 b15zdnd11an1n04x5 FILLER_222_2039 ();
 b15zdnd11an1n04x5 FILLER_222_2052 ();
 b15zdnd00an1n01x5 FILLER_222_2056 ();
 b15zdnd11an1n64x5 FILLER_222_2061 ();
 b15zdnd11an1n16x5 FILLER_222_2125 ();
 b15zdnd11an1n08x5 FILLER_222_2141 ();
 b15zdnd11an1n04x5 FILLER_222_2149 ();
 b15zdnd00an1n01x5 FILLER_222_2153 ();
 b15zdnd11an1n16x5 FILLER_222_2162 ();
 b15zdnd11an1n08x5 FILLER_222_2178 ();
 b15zdnd00an1n02x5 FILLER_222_2186 ();
 b15zdnd00an1n01x5 FILLER_222_2188 ();
 b15zdnd11an1n08x5 FILLER_222_2209 ();
 b15zdnd00an1n02x5 FILLER_222_2217 ();
 b15zdnd00an1n01x5 FILLER_222_2219 ();
 b15zdnd11an1n04x5 FILLER_222_2240 ();
 b15zdnd11an1n08x5 FILLER_222_2252 ();
 b15zdnd11an1n04x5 FILLER_222_2260 ();
 b15zdnd11an1n08x5 FILLER_222_2268 ();
 b15zdnd11an1n64x5 FILLER_223_0 ();
 b15zdnd11an1n64x5 FILLER_223_64 ();
 b15zdnd11an1n32x5 FILLER_223_128 ();
 b15zdnd11an1n16x5 FILLER_223_160 ();
 b15zdnd11an1n08x5 FILLER_223_176 ();
 b15zdnd00an1n01x5 FILLER_223_184 ();
 b15zdnd11an1n16x5 FILLER_223_195 ();
 b15zdnd00an1n01x5 FILLER_223_211 ();
 b15zdnd11an1n64x5 FILLER_223_225 ();
 b15zdnd11an1n32x5 FILLER_223_289 ();
 b15zdnd11an1n16x5 FILLER_223_321 ();
 b15zdnd00an1n01x5 FILLER_223_337 ();
 b15zdnd11an1n08x5 FILLER_223_355 ();
 b15zdnd11an1n04x5 FILLER_223_373 ();
 b15zdnd11an1n64x5 FILLER_223_403 ();
 b15zdnd11an1n64x5 FILLER_223_467 ();
 b15zdnd11an1n64x5 FILLER_223_531 ();
 b15zdnd11an1n64x5 FILLER_223_595 ();
 b15zdnd11an1n64x5 FILLER_223_659 ();
 b15zdnd11an1n32x5 FILLER_223_723 ();
 b15zdnd11an1n16x5 FILLER_223_755 ();
 b15zdnd00an1n02x5 FILLER_223_771 ();
 b15zdnd11an1n08x5 FILLER_223_793 ();
 b15zdnd00an1n02x5 FILLER_223_801 ();
 b15zdnd11an1n04x5 FILLER_223_823 ();
 b15zdnd11an1n16x5 FILLER_223_847 ();
 b15zdnd11an1n08x5 FILLER_223_863 ();
 b15zdnd00an1n01x5 FILLER_223_871 ();
 b15zdnd11an1n32x5 FILLER_223_878 ();
 b15zdnd11an1n16x5 FILLER_223_910 ();
 b15zdnd11an1n08x5 FILLER_223_926 ();
 b15zdnd11an1n04x5 FILLER_223_934 ();
 b15zdnd00an1n02x5 FILLER_223_938 ();
 b15zdnd11an1n16x5 FILLER_223_950 ();
 b15zdnd11an1n08x5 FILLER_223_966 ();
 b15zdnd00an1n01x5 FILLER_223_974 ();
 b15zdnd11an1n16x5 FILLER_223_979 ();
 b15zdnd11an1n04x5 FILLER_223_995 ();
 b15zdnd11an1n16x5 FILLER_223_1006 ();
 b15zdnd11an1n08x5 FILLER_223_1022 ();
 b15zdnd11an1n04x5 FILLER_223_1030 ();
 b15zdnd00an1n01x5 FILLER_223_1034 ();
 b15zdnd11an1n32x5 FILLER_223_1041 ();
 b15zdnd11an1n04x5 FILLER_223_1073 ();
 b15zdnd11an1n32x5 FILLER_223_1093 ();
 b15zdnd11an1n16x5 FILLER_223_1125 ();
 b15zdnd00an1n02x5 FILLER_223_1141 ();
 b15zdnd00an1n01x5 FILLER_223_1143 ();
 b15zdnd11an1n04x5 FILLER_223_1155 ();
 b15zdnd00an1n02x5 FILLER_223_1159 ();
 b15zdnd11an1n04x5 FILLER_223_1177 ();
 b15zdnd11an1n04x5 FILLER_223_1197 ();
 b15zdnd11an1n64x5 FILLER_223_1217 ();
 b15zdnd11an1n32x5 FILLER_223_1281 ();
 b15zdnd00an1n02x5 FILLER_223_1313 ();
 b15zdnd00an1n01x5 FILLER_223_1315 ();
 b15zdnd11an1n64x5 FILLER_223_1322 ();
 b15zdnd11an1n16x5 FILLER_223_1386 ();
 b15zdnd00an1n02x5 FILLER_223_1402 ();
 b15zdnd00an1n01x5 FILLER_223_1404 ();
 b15zdnd11an1n32x5 FILLER_223_1411 ();
 b15zdnd11an1n08x5 FILLER_223_1443 ();
 b15zdnd11an1n64x5 FILLER_223_1460 ();
 b15zdnd11an1n04x5 FILLER_223_1524 ();
 b15zdnd00an1n02x5 FILLER_223_1528 ();
 b15zdnd11an1n16x5 FILLER_223_1546 ();
 b15zdnd11an1n08x5 FILLER_223_1562 ();
 b15zdnd11an1n04x5 FILLER_223_1570 ();
 b15zdnd00an1n02x5 FILLER_223_1574 ();
 b15zdnd00an1n01x5 FILLER_223_1576 ();
 b15zdnd11an1n32x5 FILLER_223_1582 ();
 b15zdnd11an1n32x5 FILLER_223_1626 ();
 b15zdnd11an1n08x5 FILLER_223_1658 ();
 b15zdnd11an1n64x5 FILLER_223_1685 ();
 b15zdnd11an1n32x5 FILLER_223_1749 ();
 b15zdnd00an1n02x5 FILLER_223_1781 ();
 b15zdnd00an1n01x5 FILLER_223_1783 ();
 b15zdnd11an1n64x5 FILLER_223_1788 ();
 b15zdnd11an1n08x5 FILLER_223_1852 ();
 b15zdnd11an1n04x5 FILLER_223_1860 ();
 b15zdnd11an1n16x5 FILLER_223_1875 ();
 b15zdnd11an1n08x5 FILLER_223_1891 ();
 b15zdnd00an1n01x5 FILLER_223_1899 ();
 b15zdnd11an1n64x5 FILLER_223_1920 ();
 b15zdnd11an1n64x5 FILLER_223_1984 ();
 b15zdnd11an1n16x5 FILLER_223_2048 ();
 b15zdnd11an1n08x5 FILLER_223_2064 ();
 b15zdnd00an1n01x5 FILLER_223_2072 ();
 b15zdnd11an1n64x5 FILLER_223_2078 ();
 b15zdnd11an1n32x5 FILLER_223_2142 ();
 b15zdnd11an1n16x5 FILLER_223_2174 ();
 b15zdnd11an1n08x5 FILLER_223_2190 ();
 b15zdnd00an1n02x5 FILLER_223_2198 ();
 b15zdnd00an1n01x5 FILLER_223_2200 ();
 b15zdnd11an1n32x5 FILLER_223_2204 ();
 b15zdnd11an1n04x5 FILLER_223_2236 ();
 b15zdnd11an1n04x5 FILLER_223_2244 ();
 b15zdnd11an1n08x5 FILLER_223_2252 ();
 b15zdnd11an1n04x5 FILLER_223_2260 ();
 b15zdnd11an1n04x5 FILLER_223_2268 ();
 b15zdnd11an1n08x5 FILLER_223_2276 ();
 b15zdnd11an1n16x5 FILLER_224_8 ();
 b15zdnd11an1n04x5 FILLER_224_24 ();
 b15zdnd00an1n02x5 FILLER_224_28 ();
 b15zdnd00an1n01x5 FILLER_224_30 ();
 b15zdnd11an1n16x5 FILLER_224_47 ();
 b15zdnd11an1n04x5 FILLER_224_63 ();
 b15zdnd11an1n16x5 FILLER_224_80 ();
 b15zdnd00an1n01x5 FILLER_224_96 ();
 b15zdnd11an1n04x5 FILLER_224_101 ();
 b15zdnd11an1n64x5 FILLER_224_121 ();
 b15zdnd00an1n01x5 FILLER_224_185 ();
 b15zdnd11an1n16x5 FILLER_224_197 ();
 b15zdnd11an1n08x5 FILLER_224_213 ();
 b15zdnd11an1n04x5 FILLER_224_227 ();
 b15zdnd11an1n08x5 FILLER_224_236 ();
 b15zdnd00an1n02x5 FILLER_224_244 ();
 b15zdnd00an1n01x5 FILLER_224_246 ();
 b15zdnd11an1n08x5 FILLER_224_253 ();
 b15zdnd11an1n04x5 FILLER_224_261 ();
 b15zdnd11an1n16x5 FILLER_224_275 ();
 b15zdnd11an1n08x5 FILLER_224_291 ();
 b15zdnd00an1n01x5 FILLER_224_299 ();
 b15zdnd11an1n16x5 FILLER_224_316 ();
 b15zdnd11an1n08x5 FILLER_224_332 ();
 b15zdnd11an1n04x5 FILLER_224_347 ();
 b15zdnd11an1n04x5 FILLER_224_377 ();
 b15zdnd11an1n64x5 FILLER_224_388 ();
 b15zdnd11an1n64x5 FILLER_224_452 ();
 b15zdnd11an1n32x5 FILLER_224_516 ();
 b15zdnd11an1n08x5 FILLER_224_548 ();
 b15zdnd11an1n04x5 FILLER_224_556 ();
 b15zdnd00an1n02x5 FILLER_224_560 ();
 b15zdnd11an1n04x5 FILLER_224_571 ();
 b15zdnd00an1n02x5 FILLER_224_575 ();
 b15zdnd00an1n01x5 FILLER_224_577 ();
 b15zdnd11an1n32x5 FILLER_224_582 ();
 b15zdnd11an1n16x5 FILLER_224_614 ();
 b15zdnd00an1n02x5 FILLER_224_630 ();
 b15zdnd00an1n01x5 FILLER_224_632 ();
 b15zdnd11an1n32x5 FILLER_224_641 ();
 b15zdnd11an1n16x5 FILLER_224_673 ();
 b15zdnd00an1n01x5 FILLER_224_689 ();
 b15zdnd00an1n02x5 FILLER_224_716 ();
 b15zdnd11an1n64x5 FILLER_224_726 ();
 b15zdnd11an1n16x5 FILLER_224_790 ();
 b15zdnd11an1n08x5 FILLER_224_806 ();
 b15zdnd00an1n02x5 FILLER_224_814 ();
 b15zdnd00an1n01x5 FILLER_224_816 ();
 b15zdnd11an1n04x5 FILLER_224_826 ();
 b15zdnd11an1n32x5 FILLER_224_839 ();
 b15zdnd11an1n08x5 FILLER_224_871 ();
 b15zdnd11an1n04x5 FILLER_224_884 ();
 b15zdnd11an1n32x5 FILLER_224_892 ();
 b15zdnd11an1n16x5 FILLER_224_924 ();
 b15zdnd11an1n08x5 FILLER_224_940 ();
 b15zdnd11an1n04x5 FILLER_224_948 ();
 b15zdnd00an1n02x5 FILLER_224_952 ();
 b15zdnd00an1n01x5 FILLER_224_954 ();
 b15zdnd11an1n08x5 FILLER_224_967 ();
 b15zdnd00an1n01x5 FILLER_224_975 ();
 b15zdnd11an1n64x5 FILLER_224_980 ();
 b15zdnd11an1n64x5 FILLER_224_1044 ();
 b15zdnd11an1n32x5 FILLER_224_1108 ();
 b15zdnd00an1n02x5 FILLER_224_1140 ();
 b15zdnd11an1n32x5 FILLER_224_1158 ();
 b15zdnd11an1n16x5 FILLER_224_1190 ();
 b15zdnd00an1n01x5 FILLER_224_1206 ();
 b15zdnd11an1n04x5 FILLER_224_1223 ();
 b15zdnd00an1n01x5 FILLER_224_1227 ();
 b15zdnd11an1n64x5 FILLER_224_1248 ();
 b15zdnd11an1n64x5 FILLER_224_1312 ();
 b15zdnd11an1n16x5 FILLER_224_1376 ();
 b15zdnd11an1n08x5 FILLER_224_1392 ();
 b15zdnd11an1n04x5 FILLER_224_1400 ();
 b15zdnd11an1n04x5 FILLER_224_1412 ();
 b15zdnd11an1n16x5 FILLER_224_1422 ();
 b15zdnd11an1n08x5 FILLER_224_1438 ();
 b15zdnd11an1n04x5 FILLER_224_1446 ();
 b15zdnd00an1n02x5 FILLER_224_1450 ();
 b15zdnd00an1n01x5 FILLER_224_1452 ();
 b15zdnd11an1n64x5 FILLER_224_1464 ();
 b15zdnd11an1n64x5 FILLER_224_1528 ();
 b15zdnd11an1n64x5 FILLER_224_1592 ();
 b15zdnd11an1n32x5 FILLER_224_1656 ();
 b15zdnd11an1n08x5 FILLER_224_1688 ();
 b15zdnd00an1n01x5 FILLER_224_1696 ();
 b15zdnd11an1n04x5 FILLER_224_1722 ();
 b15zdnd11an1n32x5 FILLER_224_1748 ();
 b15zdnd11an1n04x5 FILLER_224_1811 ();
 b15zdnd00an1n01x5 FILLER_224_1815 ();
 b15zdnd11an1n04x5 FILLER_224_1847 ();
 b15zdnd11an1n64x5 FILLER_224_1877 ();
 b15zdnd11an1n64x5 FILLER_224_1941 ();
 b15zdnd11an1n64x5 FILLER_224_2005 ();
 b15zdnd11an1n32x5 FILLER_224_2069 ();
 b15zdnd11an1n08x5 FILLER_224_2101 ();
 b15zdnd11an1n04x5 FILLER_224_2109 ();
 b15zdnd11an1n32x5 FILLER_224_2118 ();
 b15zdnd11an1n04x5 FILLER_224_2150 ();
 b15zdnd11an1n64x5 FILLER_224_2162 ();
 b15zdnd11an1n16x5 FILLER_224_2226 ();
 b15zdnd11an1n08x5 FILLER_224_2242 ();
 b15zdnd11an1n08x5 FILLER_224_2254 ();
 b15zdnd11an1n08x5 FILLER_224_2266 ();
 b15zdnd00an1n02x5 FILLER_224_2274 ();
 b15zdnd11an1n16x5 FILLER_225_0 ();
 b15zdnd11an1n08x5 FILLER_225_16 ();
 b15zdnd11an1n04x5 FILLER_225_24 ();
 b15zdnd11an1n16x5 FILLER_225_59 ();
 b15zdnd11an1n08x5 FILLER_225_75 ();
 b15zdnd11an1n32x5 FILLER_225_90 ();
 b15zdnd11an1n04x5 FILLER_225_122 ();
 b15zdnd00an1n01x5 FILLER_225_126 ();
 b15zdnd11an1n04x5 FILLER_225_132 ();
 b15zdnd11an1n64x5 FILLER_225_142 ();
 b15zdnd11an1n64x5 FILLER_225_206 ();
 b15zdnd11an1n08x5 FILLER_225_287 ();
 b15zdnd00an1n02x5 FILLER_225_295 ();
 b15zdnd00an1n01x5 FILLER_225_297 ();
 b15zdnd11an1n04x5 FILLER_225_324 ();
 b15zdnd00an1n01x5 FILLER_225_328 ();
 b15zdnd11an1n08x5 FILLER_225_342 ();
 b15zdnd11an1n04x5 FILLER_225_350 ();
 b15zdnd11an1n64x5 FILLER_225_361 ();
 b15zdnd11an1n64x5 FILLER_225_425 ();
 b15zdnd11an1n08x5 FILLER_225_489 ();
 b15zdnd00an1n02x5 FILLER_225_497 ();
 b15zdnd00an1n01x5 FILLER_225_499 ();
 b15zdnd11an1n16x5 FILLER_225_532 ();
 b15zdnd11an1n08x5 FILLER_225_548 ();
 b15zdnd11an1n08x5 FILLER_225_565 ();
 b15zdnd00an1n02x5 FILLER_225_573 ();
 b15zdnd00an1n01x5 FILLER_225_575 ();
 b15zdnd11an1n08x5 FILLER_225_590 ();
 b15zdnd11an1n04x5 FILLER_225_598 ();
 b15zdnd00an1n01x5 FILLER_225_602 ();
 b15zdnd11an1n16x5 FILLER_225_607 ();
 b15zdnd11an1n08x5 FILLER_225_623 ();
 b15zdnd00an1n01x5 FILLER_225_631 ();
 b15zdnd11an1n04x5 FILLER_225_644 ();
 b15zdnd11an1n32x5 FILLER_225_656 ();
 b15zdnd11an1n08x5 FILLER_225_688 ();
 b15zdnd00an1n02x5 FILLER_225_696 ();
 b15zdnd11an1n64x5 FILLER_225_718 ();
 b15zdnd11an1n64x5 FILLER_225_782 ();
 b15zdnd11an1n32x5 FILLER_225_846 ();
 b15zdnd11an1n16x5 FILLER_225_878 ();
 b15zdnd11an1n08x5 FILLER_225_894 ();
 b15zdnd00an1n02x5 FILLER_225_902 ();
 b15zdnd00an1n01x5 FILLER_225_904 ();
 b15zdnd11an1n64x5 FILLER_225_913 ();
 b15zdnd11an1n08x5 FILLER_225_977 ();
 b15zdnd11an1n04x5 FILLER_225_985 ();
 b15zdnd11an1n32x5 FILLER_225_993 ();
 b15zdnd11an1n08x5 FILLER_225_1025 ();
 b15zdnd00an1n01x5 FILLER_225_1033 ();
 b15zdnd11an1n64x5 FILLER_225_1041 ();
 b15zdnd11an1n32x5 FILLER_225_1105 ();
 b15zdnd11an1n16x5 FILLER_225_1137 ();
 b15zdnd11an1n04x5 FILLER_225_1153 ();
 b15zdnd11an1n08x5 FILLER_225_1177 ();
 b15zdnd11an1n04x5 FILLER_225_1185 ();
 b15zdnd00an1n01x5 FILLER_225_1189 ();
 b15zdnd11an1n32x5 FILLER_225_1196 ();
 b15zdnd11an1n16x5 FILLER_225_1228 ();
 b15zdnd11an1n08x5 FILLER_225_1244 ();
 b15zdnd00an1n02x5 FILLER_225_1252 ();
 b15zdnd00an1n01x5 FILLER_225_1254 ();
 b15zdnd11an1n04x5 FILLER_225_1275 ();
 b15zdnd11an1n04x5 FILLER_225_1295 ();
 b15zdnd11an1n08x5 FILLER_225_1322 ();
 b15zdnd11an1n04x5 FILLER_225_1336 ();
 b15zdnd00an1n02x5 FILLER_225_1340 ();
 b15zdnd11an1n08x5 FILLER_225_1349 ();
 b15zdnd11an1n08x5 FILLER_225_1362 ();
 b15zdnd11an1n64x5 FILLER_225_1386 ();
 b15zdnd11an1n16x5 FILLER_225_1450 ();
 b15zdnd11an1n08x5 FILLER_225_1466 ();
 b15zdnd11an1n04x5 FILLER_225_1474 ();
 b15zdnd00an1n02x5 FILLER_225_1478 ();
 b15zdnd11an1n04x5 FILLER_225_1486 ();
 b15zdnd11an1n08x5 FILLER_225_1502 ();
 b15zdnd11an1n04x5 FILLER_225_1519 ();
 b15zdnd11an1n04x5 FILLER_225_1527 ();
 b15zdnd11an1n32x5 FILLER_225_1541 ();
 b15zdnd11an1n04x5 FILLER_225_1573 ();
 b15zdnd00an1n02x5 FILLER_225_1577 ();
 b15zdnd11an1n16x5 FILLER_225_1589 ();
 b15zdnd11an1n08x5 FILLER_225_1605 ();
 b15zdnd11an1n04x5 FILLER_225_1613 ();
 b15zdnd00an1n02x5 FILLER_225_1617 ();
 b15zdnd00an1n01x5 FILLER_225_1619 ();
 b15zdnd11an1n32x5 FILLER_225_1629 ();
 b15zdnd11an1n04x5 FILLER_225_1672 ();
 b15zdnd11an1n32x5 FILLER_225_1689 ();
 b15zdnd11an1n16x5 FILLER_225_1721 ();
 b15zdnd11an1n08x5 FILLER_225_1737 ();
 b15zdnd11an1n04x5 FILLER_225_1745 ();
 b15zdnd11an1n08x5 FILLER_225_1769 ();
 b15zdnd11an1n04x5 FILLER_225_1777 ();
 b15zdnd00an1n02x5 FILLER_225_1781 ();
 b15zdnd11an1n64x5 FILLER_225_1792 ();
 b15zdnd11an1n08x5 FILLER_225_1856 ();
 b15zdnd11an1n04x5 FILLER_225_1864 ();
 b15zdnd00an1n01x5 FILLER_225_1868 ();
 b15zdnd11an1n04x5 FILLER_225_1879 ();
 b15zdnd11an1n32x5 FILLER_225_1888 ();
 b15zdnd11an1n16x5 FILLER_225_1920 ();
 b15zdnd11an1n08x5 FILLER_225_1936 ();
 b15zdnd11an1n04x5 FILLER_225_1944 ();
 b15zdnd00an1n02x5 FILLER_225_1948 ();
 b15zdnd00an1n01x5 FILLER_225_1950 ();
 b15zdnd11an1n04x5 FILLER_225_1966 ();
 b15zdnd11an1n32x5 FILLER_225_1975 ();
 b15zdnd11an1n04x5 FILLER_225_2007 ();
 b15zdnd00an1n02x5 FILLER_225_2011 ();
 b15zdnd11an1n64x5 FILLER_225_2033 ();
 b15zdnd11an1n16x5 FILLER_225_2097 ();
 b15zdnd11an1n32x5 FILLER_225_2133 ();
 b15zdnd11an1n16x5 FILLER_225_2165 ();
 b15zdnd00an1n02x5 FILLER_225_2181 ();
 b15zdnd11an1n04x5 FILLER_225_2203 ();
 b15zdnd11an1n04x5 FILLER_225_2227 ();
 b15zdnd00an1n01x5 FILLER_225_2231 ();
 b15zdnd11an1n04x5 FILLER_225_2236 ();
 b15zdnd11an1n08x5 FILLER_225_2248 ();
 b15zdnd00an1n02x5 FILLER_225_2256 ();
 b15zdnd00an1n01x5 FILLER_225_2258 ();
 b15zdnd11an1n16x5 FILLER_225_2263 ();
 b15zdnd11an1n04x5 FILLER_225_2279 ();
 b15zdnd00an1n01x5 FILLER_225_2283 ();
 b15zdnd11an1n32x5 FILLER_226_8 ();
 b15zdnd11an1n16x5 FILLER_226_40 ();
 b15zdnd00an1n01x5 FILLER_226_56 ();
 b15zdnd11an1n08x5 FILLER_226_71 ();
 b15zdnd00an1n02x5 FILLER_226_79 ();
 b15zdnd00an1n01x5 FILLER_226_81 ();
 b15zdnd11an1n32x5 FILLER_226_94 ();
 b15zdnd11an1n08x5 FILLER_226_126 ();
 b15zdnd11an1n04x5 FILLER_226_134 ();
 b15zdnd00an1n02x5 FILLER_226_138 ();
 b15zdnd00an1n01x5 FILLER_226_140 ();
 b15zdnd11an1n04x5 FILLER_226_157 ();
 b15zdnd11an1n04x5 FILLER_226_176 ();
 b15zdnd11an1n04x5 FILLER_226_193 ();
 b15zdnd11an1n08x5 FILLER_226_201 ();
 b15zdnd00an1n02x5 FILLER_226_209 ();
 b15zdnd11an1n16x5 FILLER_226_223 ();
 b15zdnd11an1n08x5 FILLER_226_239 ();
 b15zdnd00an1n02x5 FILLER_226_247 ();
 b15zdnd11an1n08x5 FILLER_226_258 ();
 b15zdnd11an1n16x5 FILLER_226_281 ();
 b15zdnd11an1n04x5 FILLER_226_297 ();
 b15zdnd00an1n02x5 FILLER_226_301 ();
 b15zdnd00an1n01x5 FILLER_226_303 ();
 b15zdnd11an1n16x5 FILLER_226_324 ();
 b15zdnd11an1n04x5 FILLER_226_340 ();
 b15zdnd00an1n02x5 FILLER_226_344 ();
 b15zdnd00an1n01x5 FILLER_226_346 ();
 b15zdnd11an1n08x5 FILLER_226_361 ();
 b15zdnd11an1n64x5 FILLER_226_382 ();
 b15zdnd00an1n01x5 FILLER_226_446 ();
 b15zdnd11an1n04x5 FILLER_226_454 ();
 b15zdnd00an1n01x5 FILLER_226_458 ();
 b15zdnd11an1n08x5 FILLER_226_465 ();
 b15zdnd00an1n02x5 FILLER_226_473 ();
 b15zdnd00an1n01x5 FILLER_226_475 ();
 b15zdnd11an1n08x5 FILLER_226_486 ();
 b15zdnd11an1n04x5 FILLER_226_502 ();
 b15zdnd11an1n04x5 FILLER_226_524 ();
 b15zdnd00an1n01x5 FILLER_226_528 ();
 b15zdnd11an1n32x5 FILLER_226_538 ();
 b15zdnd11an1n16x5 FILLER_226_570 ();
 b15zdnd11an1n08x5 FILLER_226_586 ();
 b15zdnd00an1n01x5 FILLER_226_594 ();
 b15zdnd11an1n04x5 FILLER_226_625 ();
 b15zdnd11an1n04x5 FILLER_226_639 ();
 b15zdnd11an1n32x5 FILLER_226_675 ();
 b15zdnd11an1n08x5 FILLER_226_707 ();
 b15zdnd00an1n02x5 FILLER_226_715 ();
 b15zdnd00an1n01x5 FILLER_226_717 ();
 b15zdnd11an1n32x5 FILLER_226_726 ();
 b15zdnd11an1n16x5 FILLER_226_758 ();
 b15zdnd00an1n01x5 FILLER_226_774 ();
 b15zdnd11an1n04x5 FILLER_226_795 ();
 b15zdnd11an1n32x5 FILLER_226_809 ();
 b15zdnd11an1n08x5 FILLER_226_841 ();
 b15zdnd00an1n02x5 FILLER_226_849 ();
 b15zdnd00an1n01x5 FILLER_226_851 ();
 b15zdnd11an1n08x5 FILLER_226_870 ();
 b15zdnd11an1n04x5 FILLER_226_878 ();
 b15zdnd00an1n02x5 FILLER_226_882 ();
 b15zdnd11an1n08x5 FILLER_226_896 ();
 b15zdnd11an1n04x5 FILLER_226_904 ();
 b15zdnd00an1n02x5 FILLER_226_908 ();
 b15zdnd11an1n04x5 FILLER_226_915 ();
 b15zdnd11an1n32x5 FILLER_226_937 ();
 b15zdnd11an1n08x5 FILLER_226_969 ();
 b15zdnd11an1n04x5 FILLER_226_977 ();
 b15zdnd11an1n32x5 FILLER_226_988 ();
 b15zdnd11an1n08x5 FILLER_226_1020 ();
 b15zdnd00an1n02x5 FILLER_226_1028 ();
 b15zdnd00an1n01x5 FILLER_226_1030 ();
 b15zdnd11an1n16x5 FILLER_226_1037 ();
 b15zdnd11an1n08x5 FILLER_226_1053 ();
 b15zdnd11an1n04x5 FILLER_226_1061 ();
 b15zdnd00an1n02x5 FILLER_226_1065 ();
 b15zdnd11an1n32x5 FILLER_226_1072 ();
 b15zdnd11an1n04x5 FILLER_226_1104 ();
 b15zdnd00an1n02x5 FILLER_226_1108 ();
 b15zdnd00an1n01x5 FILLER_226_1110 ();
 b15zdnd11an1n08x5 FILLER_226_1127 ();
 b15zdnd11an1n04x5 FILLER_226_1135 ();
 b15zdnd00an1n02x5 FILLER_226_1139 ();
 b15zdnd11an1n08x5 FILLER_226_1161 ();
 b15zdnd11an1n04x5 FILLER_226_1169 ();
 b15zdnd11an1n64x5 FILLER_226_1204 ();
 b15zdnd11an1n08x5 FILLER_226_1268 ();
 b15zdnd11an1n04x5 FILLER_226_1276 ();
 b15zdnd11an1n04x5 FILLER_226_1293 ();
 b15zdnd11an1n16x5 FILLER_226_1315 ();
 b15zdnd11an1n08x5 FILLER_226_1331 ();
 b15zdnd00an1n02x5 FILLER_226_1339 ();
 b15zdnd00an1n01x5 FILLER_226_1341 ();
 b15zdnd11an1n04x5 FILLER_226_1355 ();
 b15zdnd11an1n16x5 FILLER_226_1371 ();
 b15zdnd11an1n04x5 FILLER_226_1387 ();
 b15zdnd00an1n02x5 FILLER_226_1391 ();
 b15zdnd00an1n01x5 FILLER_226_1393 ();
 b15zdnd11an1n64x5 FILLER_226_1400 ();
 b15zdnd11an1n16x5 FILLER_226_1464 ();
 b15zdnd11an1n08x5 FILLER_226_1480 ();
 b15zdnd11an1n04x5 FILLER_226_1488 ();
 b15zdnd00an1n02x5 FILLER_226_1492 ();
 b15zdnd00an1n01x5 FILLER_226_1494 ();
 b15zdnd11an1n04x5 FILLER_226_1519 ();
 b15zdnd11an1n08x5 FILLER_226_1533 ();
 b15zdnd00an1n01x5 FILLER_226_1541 ();
 b15zdnd11an1n16x5 FILLER_226_1551 ();
 b15zdnd11an1n08x5 FILLER_226_1567 ();
 b15zdnd11an1n32x5 FILLER_226_1586 ();
 b15zdnd11an1n08x5 FILLER_226_1618 ();
 b15zdnd11an1n04x5 FILLER_226_1626 ();
 b15zdnd00an1n02x5 FILLER_226_1630 ();
 b15zdnd11an1n32x5 FILLER_226_1636 ();
 b15zdnd00an1n02x5 FILLER_226_1668 ();
 b15zdnd11an1n08x5 FILLER_226_1675 ();
 b15zdnd11an1n04x5 FILLER_226_1683 ();
 b15zdnd11an1n64x5 FILLER_226_1705 ();
 b15zdnd11an1n08x5 FILLER_226_1769 ();
 b15zdnd00an1n02x5 FILLER_226_1777 ();
 b15zdnd00an1n01x5 FILLER_226_1779 ();
 b15zdnd11an1n32x5 FILLER_226_1785 ();
 b15zdnd11an1n04x5 FILLER_226_1817 ();
 b15zdnd00an1n02x5 FILLER_226_1821 ();
 b15zdnd11an1n32x5 FILLER_226_1828 ();
 b15zdnd11an1n16x5 FILLER_226_1860 ();
 b15zdnd11an1n08x5 FILLER_226_1876 ();
 b15zdnd11an1n64x5 FILLER_226_1904 ();
 b15zdnd11an1n08x5 FILLER_226_1968 ();
 b15zdnd11an1n04x5 FILLER_226_1976 ();
 b15zdnd11an1n16x5 FILLER_226_2001 ();
 b15zdnd11an1n08x5 FILLER_226_2017 ();
 b15zdnd00an1n02x5 FILLER_226_2025 ();
 b15zdnd00an1n01x5 FILLER_226_2027 ();
 b15zdnd11an1n16x5 FILLER_226_2048 ();
 b15zdnd11an1n08x5 FILLER_226_2064 ();
 b15zdnd11an1n04x5 FILLER_226_2072 ();
 b15zdnd11an1n16x5 FILLER_226_2085 ();
 b15zdnd11an1n08x5 FILLER_226_2101 ();
 b15zdnd11an1n04x5 FILLER_226_2109 ();
 b15zdnd11an1n08x5 FILLER_226_2124 ();
 b15zdnd00an1n02x5 FILLER_226_2152 ();
 b15zdnd11an1n64x5 FILLER_226_2162 ();
 b15zdnd11an1n16x5 FILLER_226_2226 ();
 b15zdnd11an1n08x5 FILLER_226_2242 ();
 b15zdnd11an1n08x5 FILLER_226_2261 ();
 b15zdnd11an1n04x5 FILLER_226_2269 ();
 b15zdnd00an1n02x5 FILLER_226_2273 ();
 b15zdnd00an1n01x5 FILLER_226_2275 ();
 b15zdnd11an1n64x5 FILLER_227_0 ();
 b15zdnd11an1n16x5 FILLER_227_64 ();
 b15zdnd00an1n02x5 FILLER_227_80 ();
 b15zdnd11an1n64x5 FILLER_227_93 ();
 b15zdnd11an1n16x5 FILLER_227_157 ();
 b15zdnd11an1n08x5 FILLER_227_173 ();
 b15zdnd11an1n04x5 FILLER_227_181 ();
 b15zdnd11an1n08x5 FILLER_227_201 ();
 b15zdnd00an1n02x5 FILLER_227_209 ();
 b15zdnd11an1n16x5 FILLER_227_226 ();
 b15zdnd11an1n04x5 FILLER_227_242 ();
 b15zdnd00an1n02x5 FILLER_227_246 ();
 b15zdnd11an1n16x5 FILLER_227_252 ();
 b15zdnd11an1n08x5 FILLER_227_268 ();
 b15zdnd11an1n04x5 FILLER_227_276 ();
 b15zdnd00an1n02x5 FILLER_227_280 ();
 b15zdnd00an1n01x5 FILLER_227_282 ();
 b15zdnd11an1n32x5 FILLER_227_309 ();
 b15zdnd11an1n08x5 FILLER_227_341 ();
 b15zdnd11an1n64x5 FILLER_227_369 ();
 b15zdnd11an1n16x5 FILLER_227_433 ();
 b15zdnd11an1n08x5 FILLER_227_449 ();
 b15zdnd00an1n02x5 FILLER_227_457 ();
 b15zdnd11an1n04x5 FILLER_227_466 ();
 b15zdnd00an1n02x5 FILLER_227_470 ();
 b15zdnd00an1n01x5 FILLER_227_472 ();
 b15zdnd11an1n32x5 FILLER_227_483 ();
 b15zdnd11an1n08x5 FILLER_227_515 ();
 b15zdnd11an1n08x5 FILLER_227_532 ();
 b15zdnd11an1n04x5 FILLER_227_540 ();
 b15zdnd11an1n08x5 FILLER_227_551 ();
 b15zdnd11an1n32x5 FILLER_227_563 ();
 b15zdnd11an1n04x5 FILLER_227_595 ();
 b15zdnd00an1n02x5 FILLER_227_599 ();
 b15zdnd11an1n64x5 FILLER_227_618 ();
 b15zdnd00an1n01x5 FILLER_227_682 ();
 b15zdnd11an1n32x5 FILLER_227_700 ();
 b15zdnd11an1n04x5 FILLER_227_732 ();
 b15zdnd00an1n02x5 FILLER_227_736 ();
 b15zdnd00an1n01x5 FILLER_227_738 ();
 b15zdnd11an1n64x5 FILLER_227_765 ();
 b15zdnd11an1n32x5 FILLER_227_829 ();
 b15zdnd11an1n16x5 FILLER_227_861 ();
 b15zdnd00an1n02x5 FILLER_227_877 ();
 b15zdnd00an1n01x5 FILLER_227_879 ();
 b15zdnd11an1n32x5 FILLER_227_900 ();
 b15zdnd11an1n08x5 FILLER_227_932 ();
 b15zdnd00an1n01x5 FILLER_227_940 ();
 b15zdnd11an1n08x5 FILLER_227_959 ();
 b15zdnd00an1n02x5 FILLER_227_967 ();
 b15zdnd11an1n32x5 FILLER_227_984 ();
 b15zdnd11an1n08x5 FILLER_227_1016 ();
 b15zdnd00an1n02x5 FILLER_227_1024 ();
 b15zdnd11an1n16x5 FILLER_227_1031 ();
 b15zdnd11an1n04x5 FILLER_227_1047 ();
 b15zdnd00an1n01x5 FILLER_227_1051 ();
 b15zdnd11an1n08x5 FILLER_227_1062 ();
 b15zdnd11an1n04x5 FILLER_227_1070 ();
 b15zdnd00an1n01x5 FILLER_227_1074 ();
 b15zdnd11an1n64x5 FILLER_227_1083 ();
 b15zdnd11an1n64x5 FILLER_227_1147 ();
 b15zdnd11an1n64x5 FILLER_227_1211 ();
 b15zdnd00an1n02x5 FILLER_227_1275 ();
 b15zdnd00an1n01x5 FILLER_227_1277 ();
 b15zdnd11an1n32x5 FILLER_227_1296 ();
 b15zdnd00an1n02x5 FILLER_227_1328 ();
 b15zdnd11an1n32x5 FILLER_227_1350 ();
 b15zdnd11an1n08x5 FILLER_227_1382 ();
 b15zdnd11an1n04x5 FILLER_227_1390 ();
 b15zdnd00an1n01x5 FILLER_227_1394 ();
 b15zdnd11an1n08x5 FILLER_227_1405 ();
 b15zdnd11an1n04x5 FILLER_227_1413 ();
 b15zdnd00an1n02x5 FILLER_227_1417 ();
 b15zdnd00an1n01x5 FILLER_227_1419 ();
 b15zdnd11an1n08x5 FILLER_227_1433 ();
 b15zdnd11an1n64x5 FILLER_227_1455 ();
 b15zdnd11an1n64x5 FILLER_227_1519 ();
 b15zdnd00an1n01x5 FILLER_227_1583 ();
 b15zdnd11an1n16x5 FILLER_227_1589 ();
 b15zdnd11an1n08x5 FILLER_227_1605 ();
 b15zdnd11an1n04x5 FILLER_227_1613 ();
 b15zdnd00an1n02x5 FILLER_227_1617 ();
 b15zdnd11an1n04x5 FILLER_227_1627 ();
 b15zdnd11an1n04x5 FILLER_227_1636 ();
 b15zdnd00an1n01x5 FILLER_227_1640 ();
 b15zdnd11an1n64x5 FILLER_227_1647 ();
 b15zdnd11an1n64x5 FILLER_227_1711 ();
 b15zdnd11an1n64x5 FILLER_227_1775 ();
 b15zdnd11an1n16x5 FILLER_227_1839 ();
 b15zdnd11an1n16x5 FILLER_227_1870 ();
 b15zdnd00an1n02x5 FILLER_227_1886 ();
 b15zdnd11an1n32x5 FILLER_227_1898 ();
 b15zdnd11an1n04x5 FILLER_227_1930 ();
 b15zdnd00an1n02x5 FILLER_227_1934 ();
 b15zdnd11an1n04x5 FILLER_227_1956 ();
 b15zdnd11an1n64x5 FILLER_227_1980 ();
 b15zdnd11an1n16x5 FILLER_227_2064 ();
 b15zdnd11an1n08x5 FILLER_227_2080 ();
 b15zdnd11an1n04x5 FILLER_227_2088 ();
 b15zdnd11an1n64x5 FILLER_227_2113 ();
 b15zdnd11an1n16x5 FILLER_227_2177 ();
 b15zdnd11an1n08x5 FILLER_227_2193 ();
 b15zdnd00an1n02x5 FILLER_227_2201 ();
 b15zdnd00an1n01x5 FILLER_227_2203 ();
 b15zdnd11an1n64x5 FILLER_227_2209 ();
 b15zdnd11an1n08x5 FILLER_227_2273 ();
 b15zdnd00an1n02x5 FILLER_227_2281 ();
 b15zdnd00an1n01x5 FILLER_227_2283 ();
 b15zdnd00an1n02x5 FILLER_228_8 ();
 b15zdnd11an1n08x5 FILLER_228_17 ();
 b15zdnd11an1n04x5 FILLER_228_25 ();
 b15zdnd11an1n32x5 FILLER_228_52 ();
 b15zdnd11an1n16x5 FILLER_228_84 ();
 b15zdnd11an1n04x5 FILLER_228_100 ();
 b15zdnd11an1n16x5 FILLER_228_109 ();
 b15zdnd11an1n08x5 FILLER_228_125 ();
 b15zdnd00an1n02x5 FILLER_228_133 ();
 b15zdnd00an1n01x5 FILLER_228_135 ();
 b15zdnd11an1n64x5 FILLER_228_155 ();
 b15zdnd11an1n16x5 FILLER_228_219 ();
 b15zdnd11an1n08x5 FILLER_228_235 ();
 b15zdnd11an1n04x5 FILLER_228_243 ();
 b15zdnd11an1n32x5 FILLER_228_263 ();
 b15zdnd11an1n08x5 FILLER_228_295 ();
 b15zdnd11an1n04x5 FILLER_228_303 ();
 b15zdnd00an1n02x5 FILLER_228_307 ();
 b15zdnd11an1n32x5 FILLER_228_314 ();
 b15zdnd11an1n08x5 FILLER_228_346 ();
 b15zdnd11an1n04x5 FILLER_228_354 ();
 b15zdnd00an1n02x5 FILLER_228_358 ();
 b15zdnd00an1n01x5 FILLER_228_360 ();
 b15zdnd11an1n64x5 FILLER_228_380 ();
 b15zdnd11an1n32x5 FILLER_228_444 ();
 b15zdnd00an1n02x5 FILLER_228_476 ();
 b15zdnd11an1n32x5 FILLER_228_502 ();
 b15zdnd11an1n08x5 FILLER_228_534 ();
 b15zdnd00an1n02x5 FILLER_228_542 ();
 b15zdnd00an1n01x5 FILLER_228_544 ();
 b15zdnd11an1n08x5 FILLER_228_550 ();
 b15zdnd11an1n32x5 FILLER_228_565 ();
 b15zdnd11an1n08x5 FILLER_228_597 ();
 b15zdnd00an1n02x5 FILLER_228_605 ();
 b15zdnd00an1n01x5 FILLER_228_607 ();
 b15zdnd11an1n32x5 FILLER_228_616 ();
 b15zdnd11an1n16x5 FILLER_228_648 ();
 b15zdnd00an1n02x5 FILLER_228_664 ();
 b15zdnd00an1n01x5 FILLER_228_666 ();
 b15zdnd11an1n32x5 FILLER_228_672 ();
 b15zdnd11an1n08x5 FILLER_228_704 ();
 b15zdnd11an1n04x5 FILLER_228_712 ();
 b15zdnd00an1n02x5 FILLER_228_716 ();
 b15zdnd11an1n08x5 FILLER_228_726 ();
 b15zdnd11an1n04x5 FILLER_228_734 ();
 b15zdnd11an1n64x5 FILLER_228_748 ();
 b15zdnd11an1n64x5 FILLER_228_812 ();
 b15zdnd11an1n16x5 FILLER_228_876 ();
 b15zdnd11an1n04x5 FILLER_228_892 ();
 b15zdnd00an1n02x5 FILLER_228_896 ();
 b15zdnd00an1n01x5 FILLER_228_898 ();
 b15zdnd11an1n08x5 FILLER_228_917 ();
 b15zdnd11an1n04x5 FILLER_228_925 ();
 b15zdnd00an1n02x5 FILLER_228_929 ();
 b15zdnd11an1n08x5 FILLER_228_950 ();
 b15zdnd11an1n04x5 FILLER_228_958 ();
 b15zdnd00an1n01x5 FILLER_228_962 ();
 b15zdnd11an1n16x5 FILLER_228_968 ();
 b15zdnd11an1n08x5 FILLER_228_984 ();
 b15zdnd11an1n04x5 FILLER_228_1006 ();
 b15zdnd11an1n32x5 FILLER_228_1017 ();
 b15zdnd11an1n16x5 FILLER_228_1049 ();
 b15zdnd00an1n01x5 FILLER_228_1065 ();
 b15zdnd11an1n04x5 FILLER_228_1070 ();
 b15zdnd11an1n64x5 FILLER_228_1086 ();
 b15zdnd00an1n01x5 FILLER_228_1150 ();
 b15zdnd11an1n04x5 FILLER_228_1171 ();
 b15zdnd00an1n02x5 FILLER_228_1175 ();
 b15zdnd00an1n01x5 FILLER_228_1177 ();
 b15zdnd11an1n64x5 FILLER_228_1196 ();
 b15zdnd11an1n64x5 FILLER_228_1260 ();
 b15zdnd11an1n64x5 FILLER_228_1324 ();
 b15zdnd11an1n08x5 FILLER_228_1388 ();
 b15zdnd11an1n04x5 FILLER_228_1396 ();
 b15zdnd11an1n04x5 FILLER_228_1404 ();
 b15zdnd11an1n08x5 FILLER_228_1424 ();
 b15zdnd11an1n04x5 FILLER_228_1432 ();
 b15zdnd00an1n02x5 FILLER_228_1436 ();
 b15zdnd11an1n64x5 FILLER_228_1444 ();
 b15zdnd11an1n32x5 FILLER_228_1508 ();
 b15zdnd11an1n16x5 FILLER_228_1540 ();
 b15zdnd11an1n04x5 FILLER_228_1556 ();
 b15zdnd00an1n02x5 FILLER_228_1560 ();
 b15zdnd00an1n01x5 FILLER_228_1562 ();
 b15zdnd11an1n04x5 FILLER_228_1575 ();
 b15zdnd11an1n16x5 FILLER_228_1595 ();
 b15zdnd11an1n08x5 FILLER_228_1611 ();
 b15zdnd00an1n01x5 FILLER_228_1619 ();
 b15zdnd11an1n04x5 FILLER_228_1626 ();
 b15zdnd00an1n01x5 FILLER_228_1630 ();
 b15zdnd11an1n64x5 FILLER_228_1639 ();
 b15zdnd11an1n16x5 FILLER_228_1703 ();
 b15zdnd11an1n08x5 FILLER_228_1719 ();
 b15zdnd00an1n01x5 FILLER_228_1727 ();
 b15zdnd11an1n16x5 FILLER_228_1733 ();
 b15zdnd11an1n08x5 FILLER_228_1749 ();
 b15zdnd11an1n04x5 FILLER_228_1757 ();
 b15zdnd00an1n02x5 FILLER_228_1761 ();
 b15zdnd00an1n01x5 FILLER_228_1763 ();
 b15zdnd11an1n32x5 FILLER_228_1789 ();
 b15zdnd00an1n02x5 FILLER_228_1821 ();
 b15zdnd00an1n01x5 FILLER_228_1823 ();
 b15zdnd11an1n32x5 FILLER_228_1844 ();
 b15zdnd11an1n32x5 FILLER_228_1888 ();
 b15zdnd11an1n16x5 FILLER_228_1920 ();
 b15zdnd11an1n08x5 FILLER_228_1936 ();
 b15zdnd00an1n02x5 FILLER_228_1944 ();
 b15zdnd00an1n01x5 FILLER_228_1946 ();
 b15zdnd11an1n04x5 FILLER_228_1973 ();
 b15zdnd11an1n64x5 FILLER_228_1980 ();
 b15zdnd11an1n64x5 FILLER_228_2044 ();
 b15zdnd11an1n32x5 FILLER_228_2108 ();
 b15zdnd11an1n08x5 FILLER_228_2140 ();
 b15zdnd11an1n04x5 FILLER_228_2148 ();
 b15zdnd00an1n02x5 FILLER_228_2152 ();
 b15zdnd11an1n32x5 FILLER_228_2162 ();
 b15zdnd11an1n08x5 FILLER_228_2194 ();
 b15zdnd00an1n01x5 FILLER_228_2202 ();
 b15zdnd11an1n32x5 FILLER_228_2212 ();
 b15zdnd11an1n04x5 FILLER_228_2244 ();
 b15zdnd00an1n02x5 FILLER_228_2248 ();
 b15zdnd11an1n16x5 FILLER_228_2254 ();
 b15zdnd11an1n04x5 FILLER_228_2270 ();
 b15zdnd00an1n02x5 FILLER_228_2274 ();
 b15zdnd11an1n32x5 FILLER_229_0 ();
 b15zdnd11an1n16x5 FILLER_229_32 ();
 b15zdnd11an1n04x5 FILLER_229_48 ();
 b15zdnd00an1n01x5 FILLER_229_52 ();
 b15zdnd11an1n32x5 FILLER_229_57 ();
 b15zdnd11an1n08x5 FILLER_229_89 ();
 b15zdnd11an1n04x5 FILLER_229_97 ();
 b15zdnd00an1n02x5 FILLER_229_101 ();
 b15zdnd00an1n01x5 FILLER_229_103 ();
 b15zdnd11an1n64x5 FILLER_229_112 ();
 b15zdnd11an1n08x5 FILLER_229_176 ();
 b15zdnd00an1n02x5 FILLER_229_184 ();
 b15zdnd00an1n01x5 FILLER_229_186 ();
 b15zdnd11an1n64x5 FILLER_229_191 ();
 b15zdnd00an1n02x5 FILLER_229_255 ();
 b15zdnd11an1n08x5 FILLER_229_263 ();
 b15zdnd11an1n04x5 FILLER_229_271 ();
 b15zdnd00an1n02x5 FILLER_229_275 ();
 b15zdnd11an1n32x5 FILLER_229_283 ();
 b15zdnd00an1n02x5 FILLER_229_315 ();
 b15zdnd00an1n01x5 FILLER_229_317 ();
 b15zdnd11an1n16x5 FILLER_229_335 ();
 b15zdnd00an1n02x5 FILLER_229_351 ();
 b15zdnd11an1n64x5 FILLER_229_367 ();
 b15zdnd11an1n04x5 FILLER_229_431 ();
 b15zdnd00an1n02x5 FILLER_229_435 ();
 b15zdnd11an1n32x5 FILLER_229_447 ();
 b15zdnd11an1n16x5 FILLER_229_479 ();
 b15zdnd11an1n08x5 FILLER_229_507 ();
 b15zdnd11an1n04x5 FILLER_229_528 ();
 b15zdnd00an1n02x5 FILLER_229_532 ();
 b15zdnd11an1n08x5 FILLER_229_540 ();
 b15zdnd11an1n04x5 FILLER_229_548 ();
 b15zdnd00an1n01x5 FILLER_229_552 ();
 b15zdnd11an1n64x5 FILLER_229_564 ();
 b15zdnd11an1n32x5 FILLER_229_628 ();
 b15zdnd11an1n04x5 FILLER_229_660 ();
 b15zdnd00an1n02x5 FILLER_229_664 ();
 b15zdnd11an1n16x5 FILLER_229_673 ();
 b15zdnd11an1n04x5 FILLER_229_689 ();
 b15zdnd00an1n02x5 FILLER_229_693 ();
 b15zdnd00an1n01x5 FILLER_229_695 ();
 b15zdnd11an1n16x5 FILLER_229_706 ();
 b15zdnd11an1n04x5 FILLER_229_722 ();
 b15zdnd00an1n02x5 FILLER_229_726 ();
 b15zdnd00an1n01x5 FILLER_229_728 ();
 b15zdnd11an1n04x5 FILLER_229_736 ();
 b15zdnd11an1n08x5 FILLER_229_756 ();
 b15zdnd00an1n02x5 FILLER_229_764 ();
 b15zdnd00an1n01x5 FILLER_229_766 ();
 b15zdnd11an1n16x5 FILLER_229_781 ();
 b15zdnd11an1n08x5 FILLER_229_797 ();
 b15zdnd11an1n04x5 FILLER_229_805 ();
 b15zdnd00an1n02x5 FILLER_229_809 ();
 b15zdnd11an1n64x5 FILLER_229_831 ();
 b15zdnd11an1n08x5 FILLER_229_895 ();
 b15zdnd00an1n02x5 FILLER_229_903 ();
 b15zdnd00an1n01x5 FILLER_229_905 ();
 b15zdnd11an1n16x5 FILLER_229_927 ();
 b15zdnd11an1n08x5 FILLER_229_943 ();
 b15zdnd00an1n02x5 FILLER_229_951 ();
 b15zdnd00an1n01x5 FILLER_229_953 ();
 b15zdnd11an1n04x5 FILLER_229_957 ();
 b15zdnd00an1n01x5 FILLER_229_961 ();
 b15zdnd11an1n04x5 FILLER_229_969 ();
 b15zdnd00an1n01x5 FILLER_229_973 ();
 b15zdnd11an1n32x5 FILLER_229_978 ();
 b15zdnd00an1n01x5 FILLER_229_1010 ();
 b15zdnd11an1n64x5 FILLER_229_1015 ();
 b15zdnd11an1n32x5 FILLER_229_1079 ();
 b15zdnd11an1n16x5 FILLER_229_1111 ();
 b15zdnd11an1n04x5 FILLER_229_1127 ();
 b15zdnd00an1n01x5 FILLER_229_1131 ();
 b15zdnd11an1n64x5 FILLER_229_1139 ();
 b15zdnd11an1n64x5 FILLER_229_1203 ();
 b15zdnd11an1n64x5 FILLER_229_1267 ();
 b15zdnd11an1n08x5 FILLER_229_1331 ();
 b15zdnd11an1n04x5 FILLER_229_1339 ();
 b15zdnd11an1n16x5 FILLER_229_1348 ();
 b15zdnd11an1n04x5 FILLER_229_1364 ();
 b15zdnd00an1n02x5 FILLER_229_1368 ();
 b15zdnd00an1n01x5 FILLER_229_1370 ();
 b15zdnd11an1n32x5 FILLER_229_1381 ();
 b15zdnd11an1n08x5 FILLER_229_1413 ();
 b15zdnd11an1n04x5 FILLER_229_1421 ();
 b15zdnd00an1n02x5 FILLER_229_1425 ();
 b15zdnd00an1n01x5 FILLER_229_1427 ();
 b15zdnd11an1n32x5 FILLER_229_1436 ();
 b15zdnd11an1n04x5 FILLER_229_1468 ();
 b15zdnd00an1n02x5 FILLER_229_1472 ();
 b15zdnd00an1n01x5 FILLER_229_1474 ();
 b15zdnd11an1n32x5 FILLER_229_1483 ();
 b15zdnd11an1n08x5 FILLER_229_1515 ();
 b15zdnd11an1n04x5 FILLER_229_1523 ();
 b15zdnd00an1n02x5 FILLER_229_1527 ();
 b15zdnd11an1n64x5 FILLER_229_1535 ();
 b15zdnd11an1n16x5 FILLER_229_1599 ();
 b15zdnd11an1n04x5 FILLER_229_1615 ();
 b15zdnd11an1n32x5 FILLER_229_1625 ();
 b15zdnd11an1n04x5 FILLER_229_1657 ();
 b15zdnd11an1n04x5 FILLER_229_1679 ();
 b15zdnd11an1n16x5 FILLER_229_1699 ();
 b15zdnd11an1n04x5 FILLER_229_1735 ();
 b15zdnd11an1n64x5 FILLER_229_1770 ();
 b15zdnd11an1n64x5 FILLER_229_1834 ();
 b15zdnd11an1n08x5 FILLER_229_1898 ();
 b15zdnd11an1n04x5 FILLER_229_1906 ();
 b15zdnd11an1n64x5 FILLER_229_1941 ();
 b15zdnd11an1n64x5 FILLER_229_2005 ();
 b15zdnd11an1n64x5 FILLER_229_2069 ();
 b15zdnd11an1n32x5 FILLER_229_2133 ();
 b15zdnd11an1n16x5 FILLER_229_2165 ();
 b15zdnd11an1n04x5 FILLER_229_2181 ();
 b15zdnd11an1n16x5 FILLER_229_2205 ();
 b15zdnd11an1n08x5 FILLER_229_2221 ();
 b15zdnd11an1n04x5 FILLER_229_2229 ();
 b15zdnd11an1n16x5 FILLER_229_2253 ();
 b15zdnd00an1n01x5 FILLER_229_2269 ();
 b15zdnd11an1n08x5 FILLER_229_2274 ();
 b15zdnd00an1n02x5 FILLER_229_2282 ();
 b15zdnd11an1n16x5 FILLER_230_8 ();
 b15zdnd11an1n04x5 FILLER_230_24 ();
 b15zdnd00an1n02x5 FILLER_230_28 ();
 b15zdnd00an1n01x5 FILLER_230_30 ();
 b15zdnd11an1n04x5 FILLER_230_48 ();
 b15zdnd11an1n04x5 FILLER_230_58 ();
 b15zdnd00an1n02x5 FILLER_230_62 ();
 b15zdnd00an1n01x5 FILLER_230_64 ();
 b15zdnd11an1n08x5 FILLER_230_88 ();
 b15zdnd11an1n04x5 FILLER_230_96 ();
 b15zdnd11an1n04x5 FILLER_230_104 ();
 b15zdnd11an1n64x5 FILLER_230_114 ();
 b15zdnd11an1n32x5 FILLER_230_178 ();
 b15zdnd11an1n08x5 FILLER_230_210 ();
 b15zdnd00an1n01x5 FILLER_230_218 ();
 b15zdnd11an1n04x5 FILLER_230_225 ();
 b15zdnd11an1n32x5 FILLER_230_235 ();
 b15zdnd11an1n08x5 FILLER_230_267 ();
 b15zdnd00an1n01x5 FILLER_230_275 ();
 b15zdnd11an1n08x5 FILLER_230_288 ();
 b15zdnd00an1n02x5 FILLER_230_296 ();
 b15zdnd11an1n04x5 FILLER_230_312 ();
 b15zdnd11an1n04x5 FILLER_230_337 ();
 b15zdnd11an1n64x5 FILLER_230_361 ();
 b15zdnd11an1n32x5 FILLER_230_425 ();
 b15zdnd11an1n08x5 FILLER_230_457 ();
 b15zdnd00an1n02x5 FILLER_230_465 ();
 b15zdnd00an1n01x5 FILLER_230_467 ();
 b15zdnd11an1n04x5 FILLER_230_478 ();
 b15zdnd11an1n16x5 FILLER_230_496 ();
 b15zdnd11an1n04x5 FILLER_230_512 ();
 b15zdnd00an1n01x5 FILLER_230_516 ();
 b15zdnd11an1n32x5 FILLER_230_530 ();
 b15zdnd00an1n01x5 FILLER_230_562 ();
 b15zdnd11an1n32x5 FILLER_230_568 ();
 b15zdnd11an1n04x5 FILLER_230_600 ();
 b15zdnd00an1n02x5 FILLER_230_604 ();
 b15zdnd00an1n01x5 FILLER_230_606 ();
 b15zdnd11an1n04x5 FILLER_230_617 ();
 b15zdnd11an1n08x5 FILLER_230_633 ();
 b15zdnd11an1n04x5 FILLER_230_641 ();
 b15zdnd00an1n02x5 FILLER_230_645 ();
 b15zdnd00an1n01x5 FILLER_230_647 ();
 b15zdnd11an1n04x5 FILLER_230_658 ();
 b15zdnd11an1n16x5 FILLER_230_672 ();
 b15zdnd11an1n08x5 FILLER_230_688 ();
 b15zdnd00an1n01x5 FILLER_230_696 ();
 b15zdnd11an1n08x5 FILLER_230_706 ();
 b15zdnd11an1n04x5 FILLER_230_714 ();
 b15zdnd11an1n08x5 FILLER_230_726 ();
 b15zdnd11an1n04x5 FILLER_230_734 ();
 b15zdnd00an1n02x5 FILLER_230_738 ();
 b15zdnd11an1n64x5 FILLER_230_766 ();
 b15zdnd11an1n16x5 FILLER_230_830 ();
 b15zdnd00an1n02x5 FILLER_230_846 ();
 b15zdnd00an1n01x5 FILLER_230_848 ();
 b15zdnd11an1n32x5 FILLER_230_869 ();
 b15zdnd11an1n16x5 FILLER_230_901 ();
 b15zdnd00an1n02x5 FILLER_230_917 ();
 b15zdnd11an1n04x5 FILLER_230_950 ();
 b15zdnd00an1n02x5 FILLER_230_954 ();
 b15zdnd11an1n64x5 FILLER_230_988 ();
 b15zdnd11an1n64x5 FILLER_230_1052 ();
 b15zdnd11an1n08x5 FILLER_230_1116 ();
 b15zdnd11an1n04x5 FILLER_230_1124 ();
 b15zdnd00an1n02x5 FILLER_230_1128 ();
 b15zdnd00an1n01x5 FILLER_230_1130 ();
 b15zdnd11an1n08x5 FILLER_230_1141 ();
 b15zdnd11an1n04x5 FILLER_230_1149 ();
 b15zdnd00an1n02x5 FILLER_230_1153 ();
 b15zdnd11an1n16x5 FILLER_230_1180 ();
 b15zdnd00an1n01x5 FILLER_230_1196 ();
 b15zdnd11an1n16x5 FILLER_230_1202 ();
 b15zdnd11an1n04x5 FILLER_230_1218 ();
 b15zdnd11an1n64x5 FILLER_230_1238 ();
 b15zdnd11an1n04x5 FILLER_230_1302 ();
 b15zdnd00an1n02x5 FILLER_230_1306 ();
 b15zdnd00an1n01x5 FILLER_230_1308 ();
 b15zdnd11an1n16x5 FILLER_230_1325 ();
 b15zdnd11an1n04x5 FILLER_230_1341 ();
 b15zdnd00an1n01x5 FILLER_230_1345 ();
 b15zdnd11an1n04x5 FILLER_230_1355 ();
 b15zdnd11an1n32x5 FILLER_230_1391 ();
 b15zdnd00an1n01x5 FILLER_230_1423 ();
 b15zdnd11an1n16x5 FILLER_230_1432 ();
 b15zdnd00an1n02x5 FILLER_230_1448 ();
 b15zdnd11an1n04x5 FILLER_230_1465 ();
 b15zdnd00an1n02x5 FILLER_230_1469 ();
 b15zdnd11an1n04x5 FILLER_230_1478 ();
 b15zdnd11an1n04x5 FILLER_230_1508 ();
 b15zdnd00an1n02x5 FILLER_230_1512 ();
 b15zdnd11an1n04x5 FILLER_230_1522 ();
 b15zdnd00an1n02x5 FILLER_230_1526 ();
 b15zdnd11an1n08x5 FILLER_230_1540 ();
 b15zdnd00an1n01x5 FILLER_230_1548 ();
 b15zdnd11an1n08x5 FILLER_230_1556 ();
 b15zdnd11an1n04x5 FILLER_230_1564 ();
 b15zdnd00an1n02x5 FILLER_230_1568 ();
 b15zdnd00an1n01x5 FILLER_230_1570 ();
 b15zdnd11an1n32x5 FILLER_230_1580 ();
 b15zdnd11an1n04x5 FILLER_230_1612 ();
 b15zdnd00an1n01x5 FILLER_230_1616 ();
 b15zdnd11an1n16x5 FILLER_230_1627 ();
 b15zdnd11an1n08x5 FILLER_230_1643 ();
 b15zdnd00an1n02x5 FILLER_230_1651 ();
 b15zdnd00an1n01x5 FILLER_230_1653 ();
 b15zdnd11an1n32x5 FILLER_230_1674 ();
 b15zdnd00an1n01x5 FILLER_230_1706 ();
 b15zdnd11an1n08x5 FILLER_230_1721 ();
 b15zdnd11an1n04x5 FILLER_230_1729 ();
 b15zdnd11an1n64x5 FILLER_230_1736 ();
 b15zdnd11an1n64x5 FILLER_230_1800 ();
 b15zdnd11an1n64x5 FILLER_230_1864 ();
 b15zdnd11an1n64x5 FILLER_230_1928 ();
 b15zdnd11an1n64x5 FILLER_230_1992 ();
 b15zdnd11an1n64x5 FILLER_230_2056 ();
 b15zdnd11an1n32x5 FILLER_230_2120 ();
 b15zdnd00an1n02x5 FILLER_230_2152 ();
 b15zdnd11an1n32x5 FILLER_230_2162 ();
 b15zdnd11an1n04x5 FILLER_230_2194 ();
 b15zdnd00an1n02x5 FILLER_230_2198 ();
 b15zdnd11an1n16x5 FILLER_230_2226 ();
 b15zdnd11an1n08x5 FILLER_230_2242 ();
 b15zdnd00an1n02x5 FILLER_230_2250 ();
 b15zdnd11an1n04x5 FILLER_230_2263 ();
 b15zdnd00an1n02x5 FILLER_230_2267 ();
 b15zdnd00an1n01x5 FILLER_230_2269 ();
 b15zdnd00an1n02x5 FILLER_230_2274 ();
 b15zdnd11an1n16x5 FILLER_231_0 ();
 b15zdnd11an1n08x5 FILLER_231_16 ();
 b15zdnd11an1n04x5 FILLER_231_24 ();
 b15zdnd11an1n08x5 FILLER_231_50 ();
 b15zdnd11an1n04x5 FILLER_231_58 ();
 b15zdnd11an1n16x5 FILLER_231_76 ();
 b15zdnd11an1n08x5 FILLER_231_92 ();
 b15zdnd00an1n02x5 FILLER_231_100 ();
 b15zdnd00an1n01x5 FILLER_231_102 ();
 b15zdnd11an1n08x5 FILLER_231_110 ();
 b15zdnd11an1n04x5 FILLER_231_118 ();
 b15zdnd00an1n02x5 FILLER_231_122 ();
 b15zdnd11an1n08x5 FILLER_231_130 ();
 b15zdnd11an1n04x5 FILLER_231_138 ();
 b15zdnd00an1n02x5 FILLER_231_142 ();
 b15zdnd11an1n04x5 FILLER_231_154 ();
 b15zdnd11an1n16x5 FILLER_231_164 ();
 b15zdnd00an1n02x5 FILLER_231_180 ();
 b15zdnd11an1n16x5 FILLER_231_187 ();
 b15zdnd11an1n08x5 FILLER_231_203 ();
 b15zdnd11an1n04x5 FILLER_231_211 ();
 b15zdnd00an1n02x5 FILLER_231_215 ();
 b15zdnd00an1n01x5 FILLER_231_217 ();
 b15zdnd11an1n04x5 FILLER_231_223 ();
 b15zdnd00an1n02x5 FILLER_231_227 ();
 b15zdnd11an1n32x5 FILLER_231_239 ();
 b15zdnd11an1n04x5 FILLER_231_271 ();
 b15zdnd00an1n02x5 FILLER_231_275 ();
 b15zdnd11an1n08x5 FILLER_231_281 ();
 b15zdnd11an1n04x5 FILLER_231_289 ();
 b15zdnd00an1n02x5 FILLER_231_293 ();
 b15zdnd11an1n08x5 FILLER_231_321 ();
 b15zdnd11an1n04x5 FILLER_231_329 ();
 b15zdnd00an1n02x5 FILLER_231_333 ();
 b15zdnd11an1n04x5 FILLER_231_341 ();
 b15zdnd11an1n08x5 FILLER_231_349 ();
 b15zdnd11an1n04x5 FILLER_231_357 ();
 b15zdnd00an1n02x5 FILLER_231_361 ();
 b15zdnd11an1n64x5 FILLER_231_371 ();
 b15zdnd11an1n64x5 FILLER_231_435 ();
 b15zdnd11an1n16x5 FILLER_231_499 ();
 b15zdnd11an1n08x5 FILLER_231_515 ();
 b15zdnd11an1n04x5 FILLER_231_523 ();
 b15zdnd00an1n01x5 FILLER_231_527 ();
 b15zdnd11an1n04x5 FILLER_231_535 ();
 b15zdnd11an1n64x5 FILLER_231_565 ();
 b15zdnd11an1n64x5 FILLER_231_629 ();
 b15zdnd11an1n04x5 FILLER_231_693 ();
 b15zdnd00an1n01x5 FILLER_231_697 ();
 b15zdnd11an1n32x5 FILLER_231_707 ();
 b15zdnd11an1n16x5 FILLER_231_739 ();
 b15zdnd11an1n08x5 FILLER_231_755 ();
 b15zdnd11an1n04x5 FILLER_231_763 ();
 b15zdnd00an1n02x5 FILLER_231_767 ();
 b15zdnd00an1n01x5 FILLER_231_769 ();
 b15zdnd11an1n16x5 FILLER_231_786 ();
 b15zdnd00an1n01x5 FILLER_231_802 ();
 b15zdnd11an1n16x5 FILLER_231_829 ();
 b15zdnd11an1n08x5 FILLER_231_845 ();
 b15zdnd00an1n02x5 FILLER_231_853 ();
 b15zdnd11an1n08x5 FILLER_231_859 ();
 b15zdnd11an1n04x5 FILLER_231_867 ();
 b15zdnd00an1n01x5 FILLER_231_871 ();
 b15zdnd11an1n64x5 FILLER_231_884 ();
 b15zdnd11an1n64x5 FILLER_231_948 ();
 b15zdnd11an1n64x5 FILLER_231_1012 ();
 b15zdnd11an1n32x5 FILLER_231_1076 ();
 b15zdnd11an1n08x5 FILLER_231_1108 ();
 b15zdnd00an1n01x5 FILLER_231_1116 ();
 b15zdnd11an1n08x5 FILLER_231_1122 ();
 b15zdnd00an1n02x5 FILLER_231_1130 ();
 b15zdnd11an1n08x5 FILLER_231_1146 ();
 b15zdnd00an1n01x5 FILLER_231_1154 ();
 b15zdnd11an1n04x5 FILLER_231_1161 ();
 b15zdnd00an1n02x5 FILLER_231_1165 ();
 b15zdnd11an1n16x5 FILLER_231_1186 ();
 b15zdnd11an1n04x5 FILLER_231_1202 ();
 b15zdnd11an1n16x5 FILLER_231_1214 ();
 b15zdnd11an1n08x5 FILLER_231_1230 ();
 b15zdnd00an1n02x5 FILLER_231_1238 ();
 b15zdnd11an1n32x5 FILLER_231_1258 ();
 b15zdnd11an1n08x5 FILLER_231_1290 ();
 b15zdnd11an1n16x5 FILLER_231_1320 ();
 b15zdnd00an1n02x5 FILLER_231_1336 ();
 b15zdnd11an1n04x5 FILLER_231_1353 ();
 b15zdnd00an1n02x5 FILLER_231_1357 ();
 b15zdnd00an1n01x5 FILLER_231_1359 ();
 b15zdnd11an1n32x5 FILLER_231_1381 ();
 b15zdnd11an1n16x5 FILLER_231_1413 ();
 b15zdnd11an1n16x5 FILLER_231_1435 ();
 b15zdnd11an1n08x5 FILLER_231_1451 ();
 b15zdnd00an1n02x5 FILLER_231_1459 ();
 b15zdnd11an1n16x5 FILLER_231_1472 ();
 b15zdnd11an1n08x5 FILLER_231_1488 ();
 b15zdnd11an1n04x5 FILLER_231_1496 ();
 b15zdnd00an1n02x5 FILLER_231_1500 ();
 b15zdnd11an1n04x5 FILLER_231_1518 ();
 b15zdnd11an1n32x5 FILLER_231_1528 ();
 b15zdnd11an1n16x5 FILLER_231_1560 ();
 b15zdnd11an1n04x5 FILLER_231_1576 ();
 b15zdnd11an1n04x5 FILLER_231_1594 ();
 b15zdnd11an1n04x5 FILLER_231_1610 ();
 b15zdnd00an1n01x5 FILLER_231_1614 ();
 b15zdnd11an1n04x5 FILLER_231_1626 ();
 b15zdnd00an1n01x5 FILLER_231_1630 ();
 b15zdnd11an1n04x5 FILLER_231_1639 ();
 b15zdnd00an1n02x5 FILLER_231_1643 ();
 b15zdnd11an1n16x5 FILLER_231_1660 ();
 b15zdnd11an1n04x5 FILLER_231_1676 ();
 b15zdnd00an1n02x5 FILLER_231_1680 ();
 b15zdnd00an1n01x5 FILLER_231_1682 ();
 b15zdnd11an1n64x5 FILLER_231_1699 ();
 b15zdnd11an1n16x5 FILLER_231_1763 ();
 b15zdnd11an1n04x5 FILLER_231_1779 ();
 b15zdnd00an1n02x5 FILLER_231_1783 ();
 b15zdnd11an1n16x5 FILLER_231_1794 ();
 b15zdnd11an1n04x5 FILLER_231_1810 ();
 b15zdnd11an1n64x5 FILLER_231_1820 ();
 b15zdnd11an1n64x5 FILLER_231_1884 ();
 b15zdnd11an1n64x5 FILLER_231_1948 ();
 b15zdnd11an1n64x5 FILLER_231_2012 ();
 b15zdnd11an1n64x5 FILLER_231_2076 ();
 b15zdnd11an1n64x5 FILLER_231_2140 ();
 b15zdnd11an1n16x5 FILLER_231_2204 ();
 b15zdnd11an1n08x5 FILLER_231_2220 ();
 b15zdnd00an1n02x5 FILLER_231_2228 ();
 b15zdnd11an1n32x5 FILLER_231_2250 ();
 b15zdnd00an1n02x5 FILLER_231_2282 ();
 b15zdnd11an1n32x5 FILLER_232_8 ();
 b15zdnd11an1n04x5 FILLER_232_40 ();
 b15zdnd00an1n02x5 FILLER_232_44 ();
 b15zdnd00an1n01x5 FILLER_232_46 ();
 b15zdnd11an1n32x5 FILLER_232_57 ();
 b15zdnd11an1n16x5 FILLER_232_89 ();
 b15zdnd00an1n02x5 FILLER_232_105 ();
 b15zdnd11an1n04x5 FILLER_232_112 ();
 b15zdnd11an1n04x5 FILLER_232_123 ();
 b15zdnd00an1n01x5 FILLER_232_127 ();
 b15zdnd11an1n16x5 FILLER_232_140 ();
 b15zdnd11an1n08x5 FILLER_232_156 ();
 b15zdnd11an1n04x5 FILLER_232_164 ();
 b15zdnd00an1n02x5 FILLER_232_168 ();
 b15zdnd11an1n04x5 FILLER_232_175 ();
 b15zdnd11an1n04x5 FILLER_232_185 ();
 b15zdnd00an1n02x5 FILLER_232_189 ();
 b15zdnd11an1n04x5 FILLER_232_212 ();
 b15zdnd11an1n64x5 FILLER_232_224 ();
 b15zdnd11an1n04x5 FILLER_232_288 ();
 b15zdnd00an1n02x5 FILLER_232_292 ();
 b15zdnd00an1n01x5 FILLER_232_294 ();
 b15zdnd11an1n08x5 FILLER_232_309 ();
 b15zdnd11an1n04x5 FILLER_232_317 ();
 b15zdnd11an1n16x5 FILLER_232_325 ();
 b15zdnd11an1n04x5 FILLER_232_347 ();
 b15zdnd11an1n64x5 FILLER_232_368 ();
 b15zdnd11an1n64x5 FILLER_232_432 ();
 b15zdnd11an1n16x5 FILLER_232_496 ();
 b15zdnd11an1n08x5 FILLER_232_512 ();
 b15zdnd11an1n64x5 FILLER_232_525 ();
 b15zdnd11an1n08x5 FILLER_232_589 ();
 b15zdnd00an1n02x5 FILLER_232_597 ();
 b15zdnd00an1n01x5 FILLER_232_599 ();
 b15zdnd11an1n08x5 FILLER_232_606 ();
 b15zdnd00an1n02x5 FILLER_232_614 ();
 b15zdnd11an1n08x5 FILLER_232_632 ();
 b15zdnd00an1n02x5 FILLER_232_640 ();
 b15zdnd11an1n04x5 FILLER_232_656 ();
 b15zdnd11an1n16x5 FILLER_232_665 ();
 b15zdnd11an1n04x5 FILLER_232_681 ();
 b15zdnd00an1n02x5 FILLER_232_685 ();
 b15zdnd00an1n01x5 FILLER_232_687 ();
 b15zdnd11an1n16x5 FILLER_232_700 ();
 b15zdnd00an1n02x5 FILLER_232_716 ();
 b15zdnd11an1n16x5 FILLER_232_726 ();
 b15zdnd11an1n08x5 FILLER_232_742 ();
 b15zdnd00an1n02x5 FILLER_232_750 ();
 b15zdnd11an1n04x5 FILLER_232_773 ();
 b15zdnd11an1n32x5 FILLER_232_803 ();
 b15zdnd11an1n16x5 FILLER_232_835 ();
 b15zdnd11an1n04x5 FILLER_232_851 ();
 b15zdnd00an1n02x5 FILLER_232_855 ();
 b15zdnd11an1n32x5 FILLER_232_862 ();
 b15zdnd11an1n16x5 FILLER_232_894 ();
 b15zdnd11an1n08x5 FILLER_232_910 ();
 b15zdnd11an1n64x5 FILLER_232_927 ();
 b15zdnd11an1n64x5 FILLER_232_991 ();
 b15zdnd11an1n64x5 FILLER_232_1055 ();
 b15zdnd11an1n64x5 FILLER_232_1119 ();
 b15zdnd11an1n16x5 FILLER_232_1183 ();
 b15zdnd11an1n08x5 FILLER_232_1199 ();
 b15zdnd00an1n02x5 FILLER_232_1207 ();
 b15zdnd11an1n64x5 FILLER_232_1217 ();
 b15zdnd11an1n32x5 FILLER_232_1281 ();
 b15zdnd11an1n16x5 FILLER_232_1313 ();
 b15zdnd11an1n08x5 FILLER_232_1329 ();
 b15zdnd11an1n16x5 FILLER_232_1345 ();
 b15zdnd11an1n08x5 FILLER_232_1361 ();
 b15zdnd00an1n02x5 FILLER_232_1369 ();
 b15zdnd00an1n01x5 FILLER_232_1371 ();
 b15zdnd11an1n16x5 FILLER_232_1385 ();
 b15zdnd11an1n08x5 FILLER_232_1401 ();
 b15zdnd00an1n02x5 FILLER_232_1409 ();
 b15zdnd00an1n01x5 FILLER_232_1411 ();
 b15zdnd11an1n04x5 FILLER_232_1416 ();
 b15zdnd11an1n64x5 FILLER_232_1427 ();
 b15zdnd11an1n08x5 FILLER_232_1491 ();
 b15zdnd00an1n02x5 FILLER_232_1499 ();
 b15zdnd00an1n01x5 FILLER_232_1501 ();
 b15zdnd11an1n32x5 FILLER_232_1507 ();
 b15zdnd11an1n08x5 FILLER_232_1539 ();
 b15zdnd00an1n02x5 FILLER_232_1547 ();
 b15zdnd11an1n04x5 FILLER_232_1554 ();
 b15zdnd11an1n04x5 FILLER_232_1565 ();
 b15zdnd11an1n16x5 FILLER_232_1574 ();
 b15zdnd11an1n08x5 FILLER_232_1590 ();
 b15zdnd00an1n02x5 FILLER_232_1598 ();
 b15zdnd11an1n08x5 FILLER_232_1606 ();
 b15zdnd00an1n02x5 FILLER_232_1614 ();
 b15zdnd00an1n01x5 FILLER_232_1616 ();
 b15zdnd11an1n64x5 FILLER_232_1622 ();
 b15zdnd11an1n64x5 FILLER_232_1686 ();
 b15zdnd11an1n32x5 FILLER_232_1750 ();
 b15zdnd00an1n02x5 FILLER_232_1782 ();
 b15zdnd00an1n01x5 FILLER_232_1784 ();
 b15zdnd11an1n08x5 FILLER_232_1790 ();
 b15zdnd11an1n04x5 FILLER_232_1798 ();
 b15zdnd00an1n02x5 FILLER_232_1802 ();
 b15zdnd00an1n01x5 FILLER_232_1804 ();
 b15zdnd11an1n64x5 FILLER_232_1825 ();
 b15zdnd11an1n16x5 FILLER_232_1889 ();
 b15zdnd11an1n64x5 FILLER_232_1937 ();
 b15zdnd11an1n08x5 FILLER_232_2001 ();
 b15zdnd11an1n04x5 FILLER_232_2009 ();
 b15zdnd00an1n02x5 FILLER_232_2013 ();
 b15zdnd00an1n01x5 FILLER_232_2015 ();
 b15zdnd11an1n32x5 FILLER_232_2033 ();
 b15zdnd11an1n16x5 FILLER_232_2065 ();
 b15zdnd11an1n08x5 FILLER_232_2081 ();
 b15zdnd11an1n04x5 FILLER_232_2089 ();
 b15zdnd00an1n01x5 FILLER_232_2093 ();
 b15zdnd11an1n32x5 FILLER_232_2106 ();
 b15zdnd11an1n16x5 FILLER_232_2138 ();
 b15zdnd11an1n64x5 FILLER_232_2162 ();
 b15zdnd11an1n32x5 FILLER_232_2226 ();
 b15zdnd11an1n16x5 FILLER_232_2258 ();
 b15zdnd00an1n02x5 FILLER_232_2274 ();
 b15zdnd11an1n16x5 FILLER_233_0 ();
 b15zdnd00an1n02x5 FILLER_233_16 ();
 b15zdnd11an1n64x5 FILLER_233_22 ();
 b15zdnd11an1n04x5 FILLER_233_86 ();
 b15zdnd00an1n01x5 FILLER_233_90 ();
 b15zdnd11an1n64x5 FILLER_233_97 ();
 b15zdnd11an1n64x5 FILLER_233_161 ();
 b15zdnd11an1n64x5 FILLER_233_225 ();
 b15zdnd11an1n16x5 FILLER_233_289 ();
 b15zdnd11an1n08x5 FILLER_233_305 ();
 b15zdnd11an1n04x5 FILLER_233_313 ();
 b15zdnd00an1n02x5 FILLER_233_317 ();
 b15zdnd11an1n32x5 FILLER_233_325 ();
 b15zdnd00an1n02x5 FILLER_233_357 ();
 b15zdnd11an1n64x5 FILLER_233_366 ();
 b15zdnd11an1n04x5 FILLER_233_430 ();
 b15zdnd00an1n01x5 FILLER_233_434 ();
 b15zdnd11an1n08x5 FILLER_233_441 ();
 b15zdnd11an1n04x5 FILLER_233_449 ();
 b15zdnd00an1n02x5 FILLER_233_453 ();
 b15zdnd00an1n01x5 FILLER_233_455 ();
 b15zdnd11an1n04x5 FILLER_233_462 ();
 b15zdnd11an1n16x5 FILLER_233_472 ();
 b15zdnd11an1n08x5 FILLER_233_488 ();
 b15zdnd00an1n01x5 FILLER_233_496 ();
 b15zdnd11an1n08x5 FILLER_233_505 ();
 b15zdnd11an1n04x5 FILLER_233_513 ();
 b15zdnd00an1n02x5 FILLER_233_517 ();
 b15zdnd00an1n01x5 FILLER_233_519 ();
 b15zdnd11an1n04x5 FILLER_233_526 ();
 b15zdnd11an1n32x5 FILLER_233_536 ();
 b15zdnd11an1n16x5 FILLER_233_568 ();
 b15zdnd11an1n08x5 FILLER_233_584 ();
 b15zdnd00an1n01x5 FILLER_233_592 ();
 b15zdnd11an1n04x5 FILLER_233_619 ();
 b15zdnd11an1n64x5 FILLER_233_632 ();
 b15zdnd11an1n16x5 FILLER_233_696 ();
 b15zdnd11an1n16x5 FILLER_233_719 ();
 b15zdnd11an1n04x5 FILLER_233_753 ();
 b15zdnd11an1n16x5 FILLER_233_775 ();
 b15zdnd11an1n08x5 FILLER_233_791 ();
 b15zdnd11an1n04x5 FILLER_233_799 ();
 b15zdnd11an1n16x5 FILLER_233_829 ();
 b15zdnd11an1n08x5 FILLER_233_845 ();
 b15zdnd11an1n04x5 FILLER_233_853 ();
 b15zdnd00an1n02x5 FILLER_233_857 ();
 b15zdnd11an1n64x5 FILLER_233_879 ();
 b15zdnd11an1n64x5 FILLER_233_943 ();
 b15zdnd11an1n32x5 FILLER_233_1007 ();
 b15zdnd11an1n16x5 FILLER_233_1039 ();
 b15zdnd11an1n04x5 FILLER_233_1073 ();
 b15zdnd11an1n64x5 FILLER_233_1083 ();
 b15zdnd11an1n16x5 FILLER_233_1147 ();
 b15zdnd11an1n08x5 FILLER_233_1163 ();
 b15zdnd00an1n02x5 FILLER_233_1171 ();
 b15zdnd00an1n01x5 FILLER_233_1173 ();
 b15zdnd11an1n16x5 FILLER_233_1179 ();
 b15zdnd11an1n08x5 FILLER_233_1195 ();
 b15zdnd11an1n04x5 FILLER_233_1203 ();
 b15zdnd00an1n01x5 FILLER_233_1207 ();
 b15zdnd11an1n04x5 FILLER_233_1213 ();
 b15zdnd00an1n01x5 FILLER_233_1217 ();
 b15zdnd11an1n32x5 FILLER_233_1234 ();
 b15zdnd11an1n16x5 FILLER_233_1266 ();
 b15zdnd11an1n16x5 FILLER_233_1298 ();
 b15zdnd11an1n08x5 FILLER_233_1314 ();
 b15zdnd11an1n04x5 FILLER_233_1322 ();
 b15zdnd11an1n32x5 FILLER_233_1336 ();
 b15zdnd11an1n16x5 FILLER_233_1368 ();
 b15zdnd00an1n01x5 FILLER_233_1384 ();
 b15zdnd11an1n08x5 FILLER_233_1395 ();
 b15zdnd00an1n01x5 FILLER_233_1403 ();
 b15zdnd11an1n08x5 FILLER_233_1410 ();
 b15zdnd11an1n04x5 FILLER_233_1418 ();
 b15zdnd11an1n16x5 FILLER_233_1436 ();
 b15zdnd00an1n01x5 FILLER_233_1452 ();
 b15zdnd11an1n64x5 FILLER_233_1459 ();
 b15zdnd11an1n64x5 FILLER_233_1523 ();
 b15zdnd11an1n32x5 FILLER_233_1587 ();
 b15zdnd11an1n16x5 FILLER_233_1619 ();
 b15zdnd11an1n08x5 FILLER_233_1635 ();
 b15zdnd11an1n04x5 FILLER_233_1643 ();
 b15zdnd11an1n64x5 FILLER_233_1654 ();
 b15zdnd11an1n64x5 FILLER_233_1718 ();
 b15zdnd11an1n04x5 FILLER_233_1782 ();
 b15zdnd11an1n08x5 FILLER_233_1806 ();
 b15zdnd00an1n01x5 FILLER_233_1814 ();
 b15zdnd11an1n16x5 FILLER_233_1820 ();
 b15zdnd11an1n08x5 FILLER_233_1836 ();
 b15zdnd11an1n04x5 FILLER_233_1844 ();
 b15zdnd00an1n02x5 FILLER_233_1848 ();
 b15zdnd11an1n32x5 FILLER_233_1870 ();
 b15zdnd11an1n08x5 FILLER_233_1902 ();
 b15zdnd00an1n02x5 FILLER_233_1910 ();
 b15zdnd00an1n01x5 FILLER_233_1912 ();
 b15zdnd11an1n08x5 FILLER_233_1945 ();
 b15zdnd11an1n04x5 FILLER_233_1953 ();
 b15zdnd00an1n01x5 FILLER_233_1957 ();
 b15zdnd11an1n08x5 FILLER_233_1963 ();
 b15zdnd11an1n04x5 FILLER_233_1971 ();
 b15zdnd00an1n01x5 FILLER_233_1975 ();
 b15zdnd11an1n04x5 FILLER_233_1982 ();
 b15zdnd00an1n01x5 FILLER_233_1986 ();
 b15zdnd11an1n08x5 FILLER_233_1991 ();
 b15zdnd00an1n01x5 FILLER_233_1999 ();
 b15zdnd11an1n04x5 FILLER_233_2005 ();
 b15zdnd11an1n04x5 FILLER_233_2020 ();
 b15zdnd11an1n04x5 FILLER_233_2031 ();
 b15zdnd00an1n01x5 FILLER_233_2035 ();
 b15zdnd11an1n16x5 FILLER_233_2042 ();
 b15zdnd11an1n16x5 FILLER_233_2065 ();
 b15zdnd11an1n04x5 FILLER_233_2081 ();
 b15zdnd11an1n04x5 FILLER_233_2094 ();
 b15zdnd00an1n02x5 FILLER_233_2098 ();
 b15zdnd11an1n16x5 FILLER_233_2106 ();
 b15zdnd00an1n02x5 FILLER_233_2122 ();
 b15zdnd11an1n08x5 FILLER_233_2136 ();
 b15zdnd11an1n04x5 FILLER_233_2144 ();
 b15zdnd00an1n02x5 FILLER_233_2148 ();
 b15zdnd11an1n64x5 FILLER_233_2161 ();
 b15zdnd11an1n32x5 FILLER_233_2225 ();
 b15zdnd11an1n04x5 FILLER_233_2257 ();
 b15zdnd11an1n16x5 FILLER_233_2265 ();
 b15zdnd00an1n02x5 FILLER_233_2281 ();
 b15zdnd00an1n01x5 FILLER_233_2283 ();
 b15zdnd11an1n64x5 FILLER_234_8 ();
 b15zdnd11an1n32x5 FILLER_234_72 ();
 b15zdnd11an1n04x5 FILLER_234_104 ();
 b15zdnd00an1n02x5 FILLER_234_108 ();
 b15zdnd11an1n64x5 FILLER_234_116 ();
 b15zdnd11an1n16x5 FILLER_234_180 ();
 b15zdnd00an1n01x5 FILLER_234_196 ();
 b15zdnd11an1n16x5 FILLER_234_206 ();
 b15zdnd00an1n02x5 FILLER_234_222 ();
 b15zdnd00an1n01x5 FILLER_234_224 ();
 b15zdnd11an1n64x5 FILLER_234_236 ();
 b15zdnd11an1n08x5 FILLER_234_300 ();
 b15zdnd11an1n04x5 FILLER_234_308 ();
 b15zdnd00an1n02x5 FILLER_234_312 ();
 b15zdnd00an1n01x5 FILLER_234_314 ();
 b15zdnd11an1n32x5 FILLER_234_327 ();
 b15zdnd11an1n16x5 FILLER_234_359 ();
 b15zdnd11an1n04x5 FILLER_234_375 ();
 b15zdnd00an1n02x5 FILLER_234_379 ();
 b15zdnd11an1n16x5 FILLER_234_413 ();
 b15zdnd00an1n02x5 FILLER_234_429 ();
 b15zdnd11an1n16x5 FILLER_234_447 ();
 b15zdnd11an1n04x5 FILLER_234_476 ();
 b15zdnd11an1n32x5 FILLER_234_484 ();
 b15zdnd11an1n16x5 FILLER_234_516 ();
 b15zdnd11an1n04x5 FILLER_234_532 ();
 b15zdnd00an1n02x5 FILLER_234_536 ();
 b15zdnd11an1n04x5 FILLER_234_548 ();
 b15zdnd11an1n08x5 FILLER_234_560 ();
 b15zdnd11an1n04x5 FILLER_234_568 ();
 b15zdnd00an1n02x5 FILLER_234_572 ();
 b15zdnd00an1n01x5 FILLER_234_574 ();
 b15zdnd11an1n16x5 FILLER_234_583 ();
 b15zdnd11an1n08x5 FILLER_234_599 ();
 b15zdnd00an1n02x5 FILLER_234_607 ();
 b15zdnd11an1n16x5 FILLER_234_616 ();
 b15zdnd11an1n08x5 FILLER_234_632 ();
 b15zdnd11an1n32x5 FILLER_234_660 ();
 b15zdnd11an1n04x5 FILLER_234_692 ();
 b15zdnd00an1n02x5 FILLER_234_696 ();
 b15zdnd11an1n08x5 FILLER_234_708 ();
 b15zdnd00an1n02x5 FILLER_234_716 ();
 b15zdnd11an1n08x5 FILLER_234_726 ();
 b15zdnd11an1n04x5 FILLER_234_734 ();
 b15zdnd00an1n01x5 FILLER_234_738 ();
 b15zdnd11an1n08x5 FILLER_234_755 ();
 b15zdnd11an1n04x5 FILLER_234_763 ();
 b15zdnd00an1n01x5 FILLER_234_767 ();
 b15zdnd11an1n16x5 FILLER_234_788 ();
 b15zdnd11an1n08x5 FILLER_234_804 ();
 b15zdnd11an1n04x5 FILLER_234_812 ();
 b15zdnd11an1n32x5 FILLER_234_836 ();
 b15zdnd11an1n08x5 FILLER_234_868 ();
 b15zdnd00an1n01x5 FILLER_234_876 ();
 b15zdnd11an1n64x5 FILLER_234_881 ();
 b15zdnd00an1n02x5 FILLER_234_945 ();
 b15zdnd00an1n01x5 FILLER_234_947 ();
 b15zdnd11an1n32x5 FILLER_234_960 ();
 b15zdnd11an1n16x5 FILLER_234_992 ();
 b15zdnd11an1n08x5 FILLER_234_1008 ();
 b15zdnd00an1n02x5 FILLER_234_1016 ();
 b15zdnd00an1n01x5 FILLER_234_1018 ();
 b15zdnd11an1n16x5 FILLER_234_1035 ();
 b15zdnd11an1n08x5 FILLER_234_1051 ();
 b15zdnd11an1n04x5 FILLER_234_1069 ();
 b15zdnd11an1n16x5 FILLER_234_1080 ();
 b15zdnd11an1n04x5 FILLER_234_1096 ();
 b15zdnd00an1n01x5 FILLER_234_1100 ();
 b15zdnd11an1n04x5 FILLER_234_1106 ();
 b15zdnd11an1n32x5 FILLER_234_1115 ();
 b15zdnd11an1n16x5 FILLER_234_1147 ();
 b15zdnd11an1n08x5 FILLER_234_1163 ();
 b15zdnd00an1n02x5 FILLER_234_1171 ();
 b15zdnd00an1n01x5 FILLER_234_1173 ();
 b15zdnd11an1n04x5 FILLER_234_1179 ();
 b15zdnd11an1n32x5 FILLER_234_1188 ();
 b15zdnd11an1n04x5 FILLER_234_1220 ();
 b15zdnd11an1n16x5 FILLER_234_1237 ();
 b15zdnd11an1n04x5 FILLER_234_1253 ();
 b15zdnd11an1n04x5 FILLER_234_1262 ();
 b15zdnd11an1n16x5 FILLER_234_1278 ();
 b15zdnd11an1n08x5 FILLER_234_1294 ();
 b15zdnd11an1n04x5 FILLER_234_1302 ();
 b15zdnd00an1n02x5 FILLER_234_1306 ();
 b15zdnd11an1n64x5 FILLER_234_1334 ();
 b15zdnd11an1n16x5 FILLER_234_1407 ();
 b15zdnd11an1n08x5 FILLER_234_1423 ();
 b15zdnd00an1n02x5 FILLER_234_1431 ();
 b15zdnd11an1n64x5 FILLER_234_1439 ();
 b15zdnd11an1n32x5 FILLER_234_1503 ();
 b15zdnd11an1n08x5 FILLER_234_1535 ();
 b15zdnd11an1n16x5 FILLER_234_1552 ();
 b15zdnd11an1n08x5 FILLER_234_1568 ();
 b15zdnd11an1n04x5 FILLER_234_1576 ();
 b15zdnd00an1n02x5 FILLER_234_1580 ();
 b15zdnd11an1n64x5 FILLER_234_1594 ();
 b15zdnd11an1n64x5 FILLER_234_1658 ();
 b15zdnd11an1n64x5 FILLER_234_1722 ();
 b15zdnd11an1n64x5 FILLER_234_1786 ();
 b15zdnd11an1n32x5 FILLER_234_1850 ();
 b15zdnd11an1n08x5 FILLER_234_1882 ();
 b15zdnd00an1n02x5 FILLER_234_1890 ();
 b15zdnd00an1n01x5 FILLER_234_1892 ();
 b15zdnd11an1n08x5 FILLER_234_1919 ();
 b15zdnd11an1n04x5 FILLER_234_1927 ();
 b15zdnd00an1n01x5 FILLER_234_1931 ();
 b15zdnd11an1n04x5 FILLER_234_1939 ();
 b15zdnd11an1n16x5 FILLER_234_1951 ();
 b15zdnd00an1n02x5 FILLER_234_1967 ();
 b15zdnd11an1n04x5 FILLER_234_2000 ();
 b15zdnd11an1n32x5 FILLER_234_2009 ();
 b15zdnd11an1n16x5 FILLER_234_2041 ();
 b15zdnd00an1n01x5 FILLER_234_2057 ();
 b15zdnd11an1n04x5 FILLER_234_2068 ();
 b15zdnd11an1n16x5 FILLER_234_2076 ();
 b15zdnd11an1n04x5 FILLER_234_2092 ();
 b15zdnd11an1n04x5 FILLER_234_2109 ();
 b15zdnd11an1n16x5 FILLER_234_2126 ();
 b15zdnd11an1n04x5 FILLER_234_2142 ();
 b15zdnd00an1n02x5 FILLER_234_2152 ();
 b15zdnd11an1n04x5 FILLER_234_2162 ();
 b15zdnd00an1n02x5 FILLER_234_2166 ();
 b15zdnd00an1n01x5 FILLER_234_2168 ();
 b15zdnd11an1n64x5 FILLER_234_2185 ();
 b15zdnd11an1n04x5 FILLER_234_2249 ();
 b15zdnd11an1n16x5 FILLER_234_2258 ();
 b15zdnd00an1n02x5 FILLER_234_2274 ();
 b15zdnd11an1n16x5 FILLER_235_0 ();
 b15zdnd00an1n01x5 FILLER_235_16 ();
 b15zdnd11an1n08x5 FILLER_235_21 ();
 b15zdnd11an1n04x5 FILLER_235_29 ();
 b15zdnd00an1n02x5 FILLER_235_33 ();
 b15zdnd00an1n01x5 FILLER_235_35 ();
 b15zdnd11an1n32x5 FILLER_235_54 ();
 b15zdnd11an1n16x5 FILLER_235_86 ();
 b15zdnd11an1n08x5 FILLER_235_102 ();
 b15zdnd11an1n04x5 FILLER_235_110 ();
 b15zdnd00an1n01x5 FILLER_235_114 ();
 b15zdnd11an1n32x5 FILLER_235_122 ();
 b15zdnd11an1n64x5 FILLER_235_159 ();
 b15zdnd11an1n08x5 FILLER_235_223 ();
 b15zdnd00an1n02x5 FILLER_235_231 ();
 b15zdnd11an1n08x5 FILLER_235_240 ();
 b15zdnd11an1n04x5 FILLER_235_248 ();
 b15zdnd00an1n01x5 FILLER_235_252 ();
 b15zdnd11an1n04x5 FILLER_235_258 ();
 b15zdnd11an1n08x5 FILLER_235_268 ();
 b15zdnd00an1n02x5 FILLER_235_276 ();
 b15zdnd00an1n01x5 FILLER_235_278 ();
 b15zdnd11an1n32x5 FILLER_235_284 ();
 b15zdnd00an1n02x5 FILLER_235_316 ();
 b15zdnd00an1n01x5 FILLER_235_318 ();
 b15zdnd11an1n16x5 FILLER_235_323 ();
 b15zdnd11an1n08x5 FILLER_235_339 ();
 b15zdnd11an1n04x5 FILLER_235_347 ();
 b15zdnd11an1n64x5 FILLER_235_369 ();
 b15zdnd11an1n16x5 FILLER_235_433 ();
 b15zdnd11an1n08x5 FILLER_235_449 ();
 b15zdnd00an1n02x5 FILLER_235_457 ();
 b15zdnd00an1n01x5 FILLER_235_459 ();
 b15zdnd11an1n04x5 FILLER_235_472 ();
 b15zdnd00an1n02x5 FILLER_235_476 ();
 b15zdnd11an1n08x5 FILLER_235_484 ();
 b15zdnd11an1n04x5 FILLER_235_492 ();
 b15zdnd00an1n02x5 FILLER_235_496 ();
 b15zdnd00an1n01x5 FILLER_235_498 ();
 b15zdnd11an1n32x5 FILLER_235_504 ();
 b15zdnd11an1n08x5 FILLER_235_536 ();
 b15zdnd11an1n04x5 FILLER_235_544 ();
 b15zdnd00an1n02x5 FILLER_235_548 ();
 b15zdnd11an1n04x5 FILLER_235_557 ();
 b15zdnd11an1n04x5 FILLER_235_571 ();
 b15zdnd00an1n01x5 FILLER_235_575 ();
 b15zdnd11an1n64x5 FILLER_235_592 ();
 b15zdnd11an1n08x5 FILLER_235_656 ();
 b15zdnd11an1n04x5 FILLER_235_664 ();
 b15zdnd00an1n02x5 FILLER_235_668 ();
 b15zdnd00an1n01x5 FILLER_235_670 ();
 b15zdnd11an1n32x5 FILLER_235_691 ();
 b15zdnd00an1n02x5 FILLER_235_723 ();
 b15zdnd00an1n01x5 FILLER_235_725 ();
 b15zdnd11an1n32x5 FILLER_235_736 ();
 b15zdnd11an1n08x5 FILLER_235_768 ();
 b15zdnd11an1n04x5 FILLER_235_776 ();
 b15zdnd00an1n02x5 FILLER_235_780 ();
 b15zdnd11an1n08x5 FILLER_235_802 ();
 b15zdnd11an1n04x5 FILLER_235_810 ();
 b15zdnd00an1n01x5 FILLER_235_814 ();
 b15zdnd11an1n64x5 FILLER_235_824 ();
 b15zdnd11an1n08x5 FILLER_235_888 ();
 b15zdnd00an1n02x5 FILLER_235_896 ();
 b15zdnd11an1n16x5 FILLER_235_923 ();
 b15zdnd11an1n08x5 FILLER_235_939 ();
 b15zdnd11an1n04x5 FILLER_235_947 ();
 b15zdnd11an1n16x5 FILLER_235_971 ();
 b15zdnd11an1n08x5 FILLER_235_987 ();
 b15zdnd11an1n04x5 FILLER_235_995 ();
 b15zdnd11an1n16x5 FILLER_235_1017 ();
 b15zdnd00an1n02x5 FILLER_235_1033 ();
 b15zdnd11an1n04x5 FILLER_235_1047 ();
 b15zdnd00an1n01x5 FILLER_235_1051 ();
 b15zdnd11an1n08x5 FILLER_235_1068 ();
 b15zdnd00an1n02x5 FILLER_235_1076 ();
 b15zdnd00an1n01x5 FILLER_235_1078 ();
 b15zdnd11an1n08x5 FILLER_235_1085 ();
 b15zdnd11an1n04x5 FILLER_235_1093 ();
 b15zdnd00an1n01x5 FILLER_235_1097 ();
 b15zdnd11an1n08x5 FILLER_235_1108 ();
 b15zdnd11an1n04x5 FILLER_235_1116 ();
 b15zdnd11an1n08x5 FILLER_235_1135 ();
 b15zdnd11an1n04x5 FILLER_235_1143 ();
 b15zdnd00an1n02x5 FILLER_235_1147 ();
 b15zdnd00an1n01x5 FILLER_235_1149 ();
 b15zdnd11an1n16x5 FILLER_235_1157 ();
 b15zdnd11an1n08x5 FILLER_235_1173 ();
 b15zdnd11an1n04x5 FILLER_235_1181 ();
 b15zdnd00an1n01x5 FILLER_235_1185 ();
 b15zdnd11an1n16x5 FILLER_235_1192 ();
 b15zdnd11an1n04x5 FILLER_235_1208 ();
 b15zdnd00an1n01x5 FILLER_235_1212 ();
 b15zdnd11an1n32x5 FILLER_235_1222 ();
 b15zdnd11an1n08x5 FILLER_235_1254 ();
 b15zdnd00an1n01x5 FILLER_235_1262 ();
 b15zdnd11an1n16x5 FILLER_235_1295 ();
 b15zdnd11an1n04x5 FILLER_235_1311 ();
 b15zdnd00an1n01x5 FILLER_235_1315 ();
 b15zdnd11an1n32x5 FILLER_235_1329 ();
 b15zdnd00an1n02x5 FILLER_235_1361 ();
 b15zdnd00an1n01x5 FILLER_235_1363 ();
 b15zdnd11an1n16x5 FILLER_235_1375 ();
 b15zdnd11an1n08x5 FILLER_235_1391 ();
 b15zdnd11an1n64x5 FILLER_235_1404 ();
 b15zdnd11an1n08x5 FILLER_235_1468 ();
 b15zdnd11an1n04x5 FILLER_235_1476 ();
 b15zdnd11an1n04x5 FILLER_235_1485 ();
 b15zdnd11an1n16x5 FILLER_235_1496 ();
 b15zdnd11an1n04x5 FILLER_235_1512 ();
 b15zdnd11an1n08x5 FILLER_235_1522 ();
 b15zdnd11an1n08x5 FILLER_235_1534 ();
 b15zdnd11an1n64x5 FILLER_235_1567 ();
 b15zdnd11an1n64x5 FILLER_235_1631 ();
 b15zdnd11an1n64x5 FILLER_235_1695 ();
 b15zdnd11an1n16x5 FILLER_235_1759 ();
 b15zdnd11an1n04x5 FILLER_235_1775 ();
 b15zdnd00an1n02x5 FILLER_235_1779 ();
 b15zdnd11an1n16x5 FILLER_235_1807 ();
 b15zdnd11an1n04x5 FILLER_235_1823 ();
 b15zdnd00an1n01x5 FILLER_235_1827 ();
 b15zdnd11an1n32x5 FILLER_235_1854 ();
 b15zdnd00an1n02x5 FILLER_235_1886 ();
 b15zdnd11an1n16x5 FILLER_235_1909 ();
 b15zdnd11an1n08x5 FILLER_235_1925 ();
 b15zdnd11an1n32x5 FILLER_235_1949 ();
 b15zdnd00an1n02x5 FILLER_235_1981 ();
 b15zdnd00an1n01x5 FILLER_235_1983 ();
 b15zdnd11an1n16x5 FILLER_235_1997 ();
 b15zdnd00an1n01x5 FILLER_235_2013 ();
 b15zdnd11an1n04x5 FILLER_235_2034 ();
 b15zdnd11an1n64x5 FILLER_235_2046 ();
 b15zdnd11an1n16x5 FILLER_235_2110 ();
 b15zdnd11an1n08x5 FILLER_235_2126 ();
 b15zdnd11an1n04x5 FILLER_235_2134 ();
 b15zdnd00an1n02x5 FILLER_235_2138 ();
 b15zdnd00an1n01x5 FILLER_235_2140 ();
 b15zdnd11an1n16x5 FILLER_235_2147 ();
 b15zdnd11an1n04x5 FILLER_235_2163 ();
 b15zdnd00an1n02x5 FILLER_235_2167 ();
 b15zdnd11an1n04x5 FILLER_235_2187 ();
 b15zdnd11an1n04x5 FILLER_235_2202 ();
 b15zdnd11an1n16x5 FILLER_235_2222 ();
 b15zdnd11an1n08x5 FILLER_235_2238 ();
 b15zdnd11an1n08x5 FILLER_235_2266 ();
 b15zdnd11an1n04x5 FILLER_235_2274 ();
 b15zdnd00an1n02x5 FILLER_235_2282 ();
 b15zdnd11an1n64x5 FILLER_236_8 ();
 b15zdnd11an1n32x5 FILLER_236_77 ();
 b15zdnd11an1n16x5 FILLER_236_109 ();
 b15zdnd11an1n08x5 FILLER_236_125 ();
 b15zdnd11an1n04x5 FILLER_236_133 ();
 b15zdnd00an1n02x5 FILLER_236_137 ();
 b15zdnd00an1n01x5 FILLER_236_139 ();
 b15zdnd11an1n04x5 FILLER_236_150 ();
 b15zdnd11an1n08x5 FILLER_236_160 ();
 b15zdnd11an1n04x5 FILLER_236_168 ();
 b15zdnd00an1n01x5 FILLER_236_172 ();
 b15zdnd11an1n32x5 FILLER_236_178 ();
 b15zdnd11an1n16x5 FILLER_236_210 ();
 b15zdnd11an1n08x5 FILLER_236_226 ();
 b15zdnd00an1n02x5 FILLER_236_234 ();
 b15zdnd00an1n01x5 FILLER_236_236 ();
 b15zdnd11an1n04x5 FILLER_236_250 ();
 b15zdnd11an1n08x5 FILLER_236_259 ();
 b15zdnd00an1n02x5 FILLER_236_267 ();
 b15zdnd11an1n32x5 FILLER_236_281 ();
 b15zdnd11an1n16x5 FILLER_236_313 ();
 b15zdnd00an1n02x5 FILLER_236_329 ();
 b15zdnd11an1n64x5 FILLER_236_347 ();
 b15zdnd11an1n08x5 FILLER_236_411 ();
 b15zdnd11an1n64x5 FILLER_236_430 ();
 b15zdnd11an1n04x5 FILLER_236_494 ();
 b15zdnd00an1n01x5 FILLER_236_498 ();
 b15zdnd11an1n04x5 FILLER_236_508 ();
 b15zdnd11an1n04x5 FILLER_236_519 ();
 b15zdnd00an1n02x5 FILLER_236_523 ();
 b15zdnd11an1n64x5 FILLER_236_537 ();
 b15zdnd00an1n01x5 FILLER_236_601 ();
 b15zdnd11an1n16x5 FILLER_236_628 ();
 b15zdnd11an1n04x5 FILLER_236_644 ();
 b15zdnd00an1n01x5 FILLER_236_648 ();
 b15zdnd11an1n08x5 FILLER_236_654 ();
 b15zdnd11an1n04x5 FILLER_236_662 ();
 b15zdnd00an1n01x5 FILLER_236_666 ();
 b15zdnd11an1n08x5 FILLER_236_671 ();
 b15zdnd00an1n02x5 FILLER_236_679 ();
 b15zdnd00an1n01x5 FILLER_236_681 ();
 b15zdnd11an1n04x5 FILLER_236_694 ();
 b15zdnd11an1n04x5 FILLER_236_712 ();
 b15zdnd00an1n02x5 FILLER_236_716 ();
 b15zdnd11an1n08x5 FILLER_236_726 ();
 b15zdnd11an1n64x5 FILLER_236_743 ();
 b15zdnd11an1n64x5 FILLER_236_807 ();
 b15zdnd11an1n32x5 FILLER_236_871 ();
 b15zdnd11an1n08x5 FILLER_236_903 ();
 b15zdnd00an1n01x5 FILLER_236_911 ();
 b15zdnd11an1n16x5 FILLER_236_932 ();
 b15zdnd11an1n08x5 FILLER_236_948 ();
 b15zdnd00an1n01x5 FILLER_236_956 ();
 b15zdnd11an1n32x5 FILLER_236_977 ();
 b15zdnd11an1n08x5 FILLER_236_1009 ();
 b15zdnd00an1n02x5 FILLER_236_1017 ();
 b15zdnd00an1n01x5 FILLER_236_1019 ();
 b15zdnd11an1n08x5 FILLER_236_1032 ();
 b15zdnd11an1n16x5 FILLER_236_1051 ();
 b15zdnd00an1n02x5 FILLER_236_1067 ();
 b15zdnd11an1n16x5 FILLER_236_1079 ();
 b15zdnd11an1n08x5 FILLER_236_1095 ();
 b15zdnd11an1n04x5 FILLER_236_1109 ();
 b15zdnd11an1n16x5 FILLER_236_1125 ();
 b15zdnd11an1n08x5 FILLER_236_1141 ();
 b15zdnd00an1n02x5 FILLER_236_1149 ();
 b15zdnd11an1n04x5 FILLER_236_1163 ();
 b15zdnd00an1n02x5 FILLER_236_1167 ();
 b15zdnd11an1n04x5 FILLER_236_1184 ();
 b15zdnd11an1n16x5 FILLER_236_1196 ();
 b15zdnd11an1n04x5 FILLER_236_1212 ();
 b15zdnd00an1n01x5 FILLER_236_1216 ();
 b15zdnd11an1n32x5 FILLER_236_1223 ();
 b15zdnd11an1n04x5 FILLER_236_1255 ();
 b15zdnd00an1n02x5 FILLER_236_1259 ();
 b15zdnd00an1n01x5 FILLER_236_1261 ();
 b15zdnd11an1n32x5 FILLER_236_1272 ();
 b15zdnd00an1n02x5 FILLER_236_1304 ();
 b15zdnd11an1n16x5 FILLER_236_1320 ();
 b15zdnd11an1n04x5 FILLER_236_1336 ();
 b15zdnd00an1n02x5 FILLER_236_1340 ();
 b15zdnd11an1n32x5 FILLER_236_1373 ();
 b15zdnd11an1n16x5 FILLER_236_1405 ();
 b15zdnd00an1n02x5 FILLER_236_1421 ();
 b15zdnd00an1n01x5 FILLER_236_1423 ();
 b15zdnd11an1n08x5 FILLER_236_1434 ();
 b15zdnd00an1n02x5 FILLER_236_1442 ();
 b15zdnd00an1n01x5 FILLER_236_1444 ();
 b15zdnd11an1n04x5 FILLER_236_1455 ();
 b15zdnd11an1n08x5 FILLER_236_1467 ();
 b15zdnd11an1n04x5 FILLER_236_1475 ();
 b15zdnd11an1n04x5 FILLER_236_1487 ();
 b15zdnd11an1n08x5 FILLER_236_1496 ();
 b15zdnd11an1n64x5 FILLER_236_1513 ();
 b15zdnd11an1n64x5 FILLER_236_1577 ();
 b15zdnd11an1n32x5 FILLER_236_1641 ();
 b15zdnd11an1n08x5 FILLER_236_1673 ();
 b15zdnd00an1n02x5 FILLER_236_1681 ();
 b15zdnd11an1n64x5 FILLER_236_1695 ();
 b15zdnd11an1n08x5 FILLER_236_1759 ();
 b15zdnd11an1n64x5 FILLER_236_1787 ();
 b15zdnd11an1n16x5 FILLER_236_1851 ();
 b15zdnd11an1n08x5 FILLER_236_1867 ();
 b15zdnd11an1n16x5 FILLER_236_1907 ();
 b15zdnd11an1n08x5 FILLER_236_1923 ();
 b15zdnd11an1n04x5 FILLER_236_1931 ();
 b15zdnd00an1n02x5 FILLER_236_1935 ();
 b15zdnd11an1n08x5 FILLER_236_1969 ();
 b15zdnd11an1n04x5 FILLER_236_1977 ();
 b15zdnd00an1n02x5 FILLER_236_1981 ();
 b15zdnd11an1n32x5 FILLER_236_2003 ();
 b15zdnd11an1n04x5 FILLER_236_2035 ();
 b15zdnd00an1n02x5 FILLER_236_2039 ();
 b15zdnd00an1n01x5 FILLER_236_2041 ();
 b15zdnd11an1n32x5 FILLER_236_2048 ();
 b15zdnd11an1n16x5 FILLER_236_2080 ();
 b15zdnd11an1n08x5 FILLER_236_2096 ();
 b15zdnd11an1n04x5 FILLER_236_2104 ();
 b15zdnd11an1n04x5 FILLER_236_2114 ();
 b15zdnd11an1n08x5 FILLER_236_2124 ();
 b15zdnd11an1n04x5 FILLER_236_2132 ();
 b15zdnd00an1n02x5 FILLER_236_2136 ();
 b15zdnd11an1n04x5 FILLER_236_2150 ();
 b15zdnd11an1n16x5 FILLER_236_2162 ();
 b15zdnd11an1n04x5 FILLER_236_2178 ();
 b15zdnd00an1n02x5 FILLER_236_2182 ();
 b15zdnd00an1n01x5 FILLER_236_2184 ();
 b15zdnd11an1n32x5 FILLER_236_2201 ();
 b15zdnd11an1n16x5 FILLER_236_2233 ();
 b15zdnd11an1n08x5 FILLER_236_2249 ();
 b15zdnd00an1n02x5 FILLER_236_2257 ();
 b15zdnd11an1n08x5 FILLER_236_2264 ();
 b15zdnd11an1n04x5 FILLER_236_2272 ();
 b15zdnd11an1n32x5 FILLER_237_0 ();
 b15zdnd11an1n16x5 FILLER_237_32 ();
 b15zdnd11an1n04x5 FILLER_237_48 ();
 b15zdnd00an1n01x5 FILLER_237_52 ();
 b15zdnd11an1n16x5 FILLER_237_59 ();
 b15zdnd00an1n01x5 FILLER_237_75 ();
 b15zdnd11an1n08x5 FILLER_237_91 ();
 b15zdnd00an1n01x5 FILLER_237_99 ();
 b15zdnd11an1n16x5 FILLER_237_105 ();
 b15zdnd11an1n04x5 FILLER_237_121 ();
 b15zdnd11an1n16x5 FILLER_237_140 ();
 b15zdnd00an1n01x5 FILLER_237_156 ();
 b15zdnd11an1n04x5 FILLER_237_173 ();
 b15zdnd11an1n64x5 FILLER_237_186 ();
 b15zdnd11an1n16x5 FILLER_237_250 ();
 b15zdnd11an1n04x5 FILLER_237_266 ();
 b15zdnd11an1n32x5 FILLER_237_274 ();
 b15zdnd11an1n08x5 FILLER_237_306 ();
 b15zdnd11an1n08x5 FILLER_237_330 ();
 b15zdnd00an1n01x5 FILLER_237_338 ();
 b15zdnd11an1n64x5 FILLER_237_355 ();
 b15zdnd11an1n08x5 FILLER_237_419 ();
 b15zdnd11an1n04x5 FILLER_237_427 ();
 b15zdnd00an1n02x5 FILLER_237_431 ();
 b15zdnd11an1n32x5 FILLER_237_449 ();
 b15zdnd11an1n16x5 FILLER_237_481 ();
 b15zdnd11an1n04x5 FILLER_237_497 ();
 b15zdnd11an1n04x5 FILLER_237_507 ();
 b15zdnd11an1n04x5 FILLER_237_527 ();
 b15zdnd11an1n16x5 FILLER_237_541 ();
 b15zdnd11an1n04x5 FILLER_237_557 ();
 b15zdnd00an1n01x5 FILLER_237_561 ();
 b15zdnd11an1n32x5 FILLER_237_573 ();
 b15zdnd11an1n08x5 FILLER_237_605 ();
 b15zdnd11an1n04x5 FILLER_237_613 ();
 b15zdnd11an1n04x5 FILLER_237_626 ();
 b15zdnd00an1n01x5 FILLER_237_630 ();
 b15zdnd11an1n04x5 FILLER_237_641 ();
 b15zdnd00an1n02x5 FILLER_237_645 ();
 b15zdnd00an1n01x5 FILLER_237_647 ();
 b15zdnd11an1n04x5 FILLER_237_658 ();
 b15zdnd11an1n16x5 FILLER_237_676 ();
 b15zdnd11an1n08x5 FILLER_237_692 ();
 b15zdnd11an1n16x5 FILLER_237_706 ();
 b15zdnd11an1n08x5 FILLER_237_722 ();
 b15zdnd11an1n04x5 FILLER_237_730 ();
 b15zdnd00an1n02x5 FILLER_237_734 ();
 b15zdnd11an1n32x5 FILLER_237_742 ();
 b15zdnd11an1n16x5 FILLER_237_774 ();
 b15zdnd11an1n08x5 FILLER_237_790 ();
 b15zdnd11an1n04x5 FILLER_237_798 ();
 b15zdnd11an1n32x5 FILLER_237_811 ();
 b15zdnd11an1n16x5 FILLER_237_843 ();
 b15zdnd11an1n08x5 FILLER_237_859 ();
 b15zdnd00an1n01x5 FILLER_237_867 ();
 b15zdnd11an1n64x5 FILLER_237_872 ();
 b15zdnd11an1n64x5 FILLER_237_936 ();
 b15zdnd11an1n64x5 FILLER_237_1000 ();
 b15zdnd11an1n64x5 FILLER_237_1064 ();
 b15zdnd11an1n16x5 FILLER_237_1128 ();
 b15zdnd11an1n08x5 FILLER_237_1144 ();
 b15zdnd00an1n02x5 FILLER_237_1152 ();
 b15zdnd11an1n32x5 FILLER_237_1160 ();
 b15zdnd11an1n16x5 FILLER_237_1192 ();
 b15zdnd11an1n08x5 FILLER_237_1208 ();
 b15zdnd00an1n02x5 FILLER_237_1216 ();
 b15zdnd00an1n01x5 FILLER_237_1218 ();
 b15zdnd11an1n32x5 FILLER_237_1229 ();
 b15zdnd11an1n16x5 FILLER_237_1261 ();
 b15zdnd11an1n04x5 FILLER_237_1277 ();
 b15zdnd00an1n02x5 FILLER_237_1281 ();
 b15zdnd00an1n01x5 FILLER_237_1283 ();
 b15zdnd11an1n64x5 FILLER_237_1315 ();
 b15zdnd11an1n16x5 FILLER_237_1379 ();
 b15zdnd11an1n04x5 FILLER_237_1395 ();
 b15zdnd11an1n08x5 FILLER_237_1430 ();
 b15zdnd11an1n04x5 FILLER_237_1438 ();
 b15zdnd11an1n64x5 FILLER_237_1461 ();
 b15zdnd00an1n02x5 FILLER_237_1525 ();
 b15zdnd00an1n01x5 FILLER_237_1527 ();
 b15zdnd11an1n64x5 FILLER_237_1536 ();
 b15zdnd11an1n32x5 FILLER_237_1600 ();
 b15zdnd11an1n16x5 FILLER_237_1632 ();
 b15zdnd11an1n04x5 FILLER_237_1648 ();
 b15zdnd11an1n04x5 FILLER_237_1661 ();
 b15zdnd00an1n02x5 FILLER_237_1665 ();
 b15zdnd00an1n01x5 FILLER_237_1667 ();
 b15zdnd11an1n32x5 FILLER_237_1672 ();
 b15zdnd11an1n16x5 FILLER_237_1704 ();
 b15zdnd00an1n01x5 FILLER_237_1720 ();
 b15zdnd11an1n32x5 FILLER_237_1726 ();
 b15zdnd00an1n01x5 FILLER_237_1758 ();
 b15zdnd11an1n32x5 FILLER_237_1791 ();
 b15zdnd11an1n08x5 FILLER_237_1823 ();
 b15zdnd00an1n01x5 FILLER_237_1831 ();
 b15zdnd11an1n64x5 FILLER_237_1852 ();
 b15zdnd11an1n16x5 FILLER_237_1916 ();
 b15zdnd11an1n08x5 FILLER_237_1932 ();
 b15zdnd11an1n04x5 FILLER_237_1940 ();
 b15zdnd11an1n32x5 FILLER_237_1948 ();
 b15zdnd11an1n08x5 FILLER_237_1980 ();
 b15zdnd11an1n04x5 FILLER_237_1988 ();
 b15zdnd00an1n01x5 FILLER_237_1992 ();
 b15zdnd11an1n64x5 FILLER_237_2019 ();
 b15zdnd11an1n64x5 FILLER_237_2083 ();
 b15zdnd11an1n64x5 FILLER_237_2147 ();
 b15zdnd11an1n64x5 FILLER_237_2211 ();
 b15zdnd11an1n08x5 FILLER_237_2275 ();
 b15zdnd00an1n01x5 FILLER_237_2283 ();
 b15zdnd11an1n32x5 FILLER_238_8 ();
 b15zdnd11an1n08x5 FILLER_238_40 ();
 b15zdnd11an1n04x5 FILLER_238_48 ();
 b15zdnd00an1n02x5 FILLER_238_52 ();
 b15zdnd11an1n16x5 FILLER_238_60 ();
 b15zdnd11an1n08x5 FILLER_238_76 ();
 b15zdnd00an1n02x5 FILLER_238_84 ();
 b15zdnd11an1n08x5 FILLER_238_95 ();
 b15zdnd00an1n01x5 FILLER_238_103 ();
 b15zdnd11an1n04x5 FILLER_238_110 ();
 b15zdnd11an1n32x5 FILLER_238_119 ();
 b15zdnd11an1n16x5 FILLER_238_161 ();
 b15zdnd11an1n08x5 FILLER_238_177 ();
 b15zdnd11an1n04x5 FILLER_238_185 ();
 b15zdnd00an1n02x5 FILLER_238_189 ();
 b15zdnd00an1n01x5 FILLER_238_191 ();
 b15zdnd11an1n04x5 FILLER_238_199 ();
 b15zdnd11an1n32x5 FILLER_238_209 ();
 b15zdnd11an1n16x5 FILLER_238_241 ();
 b15zdnd11an1n08x5 FILLER_238_257 ();
 b15zdnd11an1n04x5 FILLER_238_265 ();
 b15zdnd11an1n08x5 FILLER_238_275 ();
 b15zdnd11an1n04x5 FILLER_238_283 ();
 b15zdnd00an1n01x5 FILLER_238_287 ();
 b15zdnd11an1n16x5 FILLER_238_308 ();
 b15zdnd00an1n01x5 FILLER_238_324 ();
 b15zdnd11an1n08x5 FILLER_238_351 ();
 b15zdnd11an1n04x5 FILLER_238_359 ();
 b15zdnd11an1n08x5 FILLER_238_370 ();
 b15zdnd11an1n64x5 FILLER_238_382 ();
 b15zdnd11an1n08x5 FILLER_238_446 ();
 b15zdnd11an1n04x5 FILLER_238_454 ();
 b15zdnd00an1n01x5 FILLER_238_458 ();
 b15zdnd11an1n64x5 FILLER_238_464 ();
 b15zdnd11an1n32x5 FILLER_238_528 ();
 b15zdnd11an1n16x5 FILLER_238_560 ();
 b15zdnd11an1n08x5 FILLER_238_576 ();
 b15zdnd11an1n16x5 FILLER_238_594 ();
 b15zdnd11an1n64x5 FILLER_238_620 ();
 b15zdnd11an1n16x5 FILLER_238_684 ();
 b15zdnd00an1n02x5 FILLER_238_700 ();
 b15zdnd00an1n01x5 FILLER_238_702 ();
 b15zdnd11an1n08x5 FILLER_238_709 ();
 b15zdnd00an1n01x5 FILLER_238_717 ();
 b15zdnd11an1n08x5 FILLER_238_726 ();
 b15zdnd11an1n04x5 FILLER_238_734 ();
 b15zdnd11an1n16x5 FILLER_238_743 ();
 b15zdnd11an1n04x5 FILLER_238_759 ();
 b15zdnd00an1n02x5 FILLER_238_763 ();
 b15zdnd11an1n64x5 FILLER_238_775 ();
 b15zdnd11an1n04x5 FILLER_238_839 ();
 b15zdnd11an1n64x5 FILLER_238_863 ();
 b15zdnd11an1n64x5 FILLER_238_927 ();
 b15zdnd11an1n16x5 FILLER_238_991 ();
 b15zdnd11an1n08x5 FILLER_238_1007 ();
 b15zdnd00an1n02x5 FILLER_238_1015 ();
 b15zdnd00an1n01x5 FILLER_238_1017 ();
 b15zdnd11an1n64x5 FILLER_238_1025 ();
 b15zdnd11an1n64x5 FILLER_238_1089 ();
 b15zdnd11an1n64x5 FILLER_238_1153 ();
 b15zdnd00an1n02x5 FILLER_238_1217 ();
 b15zdnd11an1n16x5 FILLER_238_1224 ();
 b15zdnd11an1n04x5 FILLER_238_1240 ();
 b15zdnd11an1n64x5 FILLER_238_1248 ();
 b15zdnd11an1n16x5 FILLER_238_1312 ();
 b15zdnd00an1n02x5 FILLER_238_1328 ();
 b15zdnd00an1n01x5 FILLER_238_1330 ();
 b15zdnd11an1n64x5 FILLER_238_1347 ();
 b15zdnd11an1n04x5 FILLER_238_1411 ();
 b15zdnd00an1n02x5 FILLER_238_1415 ();
 b15zdnd11an1n16x5 FILLER_238_1425 ();
 b15zdnd11an1n08x5 FILLER_238_1441 ();
 b15zdnd11an1n04x5 FILLER_238_1449 ();
 b15zdnd00an1n01x5 FILLER_238_1453 ();
 b15zdnd11an1n64x5 FILLER_238_1461 ();
 b15zdnd11an1n64x5 FILLER_238_1525 ();
 b15zdnd11an1n16x5 FILLER_238_1589 ();
 b15zdnd11an1n04x5 FILLER_238_1605 ();
 b15zdnd00an1n02x5 FILLER_238_1609 ();
 b15zdnd11an1n08x5 FILLER_238_1618 ();
 b15zdnd00an1n02x5 FILLER_238_1626 ();
 b15zdnd11an1n16x5 FILLER_238_1635 ();
 b15zdnd00an1n02x5 FILLER_238_1651 ();
 b15zdnd11an1n08x5 FILLER_238_1665 ();
 b15zdnd00an1n02x5 FILLER_238_1673 ();
 b15zdnd00an1n01x5 FILLER_238_1675 ();
 b15zdnd11an1n04x5 FILLER_238_1681 ();
 b15zdnd11an1n08x5 FILLER_238_1692 ();
 b15zdnd11an1n04x5 FILLER_238_1700 ();
 b15zdnd00an1n02x5 FILLER_238_1704 ();
 b15zdnd00an1n01x5 FILLER_238_1706 ();
 b15zdnd11an1n04x5 FILLER_238_1715 ();
 b15zdnd11an1n32x5 FILLER_238_1727 ();
 b15zdnd11an1n08x5 FILLER_238_1759 ();
 b15zdnd00an1n02x5 FILLER_238_1767 ();
 b15zdnd11an1n16x5 FILLER_238_1781 ();
 b15zdnd11an1n08x5 FILLER_238_1797 ();
 b15zdnd11an1n04x5 FILLER_238_1805 ();
 b15zdnd11an1n64x5 FILLER_238_1814 ();
 b15zdnd11an1n08x5 FILLER_238_1878 ();
 b15zdnd11an1n32x5 FILLER_238_1902 ();
 b15zdnd11an1n04x5 FILLER_238_1934 ();
 b15zdnd00an1n01x5 FILLER_238_1938 ();
 b15zdnd11an1n08x5 FILLER_238_1955 ();
 b15zdnd11an1n04x5 FILLER_238_1963 ();
 b15zdnd11an1n08x5 FILLER_238_1976 ();
 b15zdnd11an1n04x5 FILLER_238_1984 ();
 b15zdnd00an1n02x5 FILLER_238_1988 ();
 b15zdnd11an1n08x5 FILLER_238_1996 ();
 b15zdnd11an1n04x5 FILLER_238_2004 ();
 b15zdnd00an1n02x5 FILLER_238_2008 ();
 b15zdnd11an1n16x5 FILLER_238_2017 ();
 b15zdnd11an1n08x5 FILLER_238_2033 ();
 b15zdnd11an1n04x5 FILLER_238_2041 ();
 b15zdnd00an1n02x5 FILLER_238_2045 ();
 b15zdnd11an1n16x5 FILLER_238_2053 ();
 b15zdnd11an1n08x5 FILLER_238_2069 ();
 b15zdnd11an1n16x5 FILLER_238_2084 ();
 b15zdnd11an1n16x5 FILLER_238_2112 ();
 b15zdnd11an1n08x5 FILLER_238_2128 ();
 b15zdnd11an1n04x5 FILLER_238_2136 ();
 b15zdnd00an1n02x5 FILLER_238_2140 ();
 b15zdnd11an1n08x5 FILLER_238_2146 ();
 b15zdnd11an1n08x5 FILLER_238_2162 ();
 b15zdnd11an1n64x5 FILLER_238_2182 ();
 b15zdnd11an1n16x5 FILLER_238_2246 ();
 b15zdnd11an1n08x5 FILLER_238_2262 ();
 b15zdnd11an1n04x5 FILLER_238_2270 ();
 b15zdnd00an1n02x5 FILLER_238_2274 ();
 b15zdnd11an1n32x5 FILLER_239_0 ();
 b15zdnd11an1n16x5 FILLER_239_32 ();
 b15zdnd00an1n02x5 FILLER_239_48 ();
 b15zdnd00an1n01x5 FILLER_239_50 ();
 b15zdnd11an1n32x5 FILLER_239_61 ();
 b15zdnd11an1n16x5 FILLER_239_93 ();
 b15zdnd00an1n02x5 FILLER_239_109 ();
 b15zdnd00an1n01x5 FILLER_239_111 ();
 b15zdnd11an1n64x5 FILLER_239_126 ();
 b15zdnd11an1n16x5 FILLER_239_190 ();
 b15zdnd11an1n16x5 FILLER_239_212 ();
 b15zdnd11an1n04x5 FILLER_239_248 ();
 b15zdnd11an1n16x5 FILLER_239_257 ();
 b15zdnd11an1n16x5 FILLER_239_278 ();
 b15zdnd11an1n08x5 FILLER_239_294 ();
 b15zdnd11an1n04x5 FILLER_239_302 ();
 b15zdnd00an1n02x5 FILLER_239_306 ();
 b15zdnd11an1n04x5 FILLER_239_314 ();
 b15zdnd11an1n04x5 FILLER_239_328 ();
 b15zdnd11an1n16x5 FILLER_239_337 ();
 b15zdnd11an1n08x5 FILLER_239_353 ();
 b15zdnd11an1n32x5 FILLER_239_371 ();
 b15zdnd11an1n16x5 FILLER_239_403 ();
 b15zdnd11an1n04x5 FILLER_239_419 ();
 b15zdnd00an1n02x5 FILLER_239_423 ();
 b15zdnd11an1n04x5 FILLER_239_446 ();
 b15zdnd11an1n08x5 FILLER_239_454 ();
 b15zdnd00an1n01x5 FILLER_239_462 ();
 b15zdnd11an1n64x5 FILLER_239_468 ();
 b15zdnd11an1n32x5 FILLER_239_532 ();
 b15zdnd11an1n16x5 FILLER_239_564 ();
 b15zdnd11an1n08x5 FILLER_239_580 ();
 b15zdnd00an1n02x5 FILLER_239_588 ();
 b15zdnd00an1n01x5 FILLER_239_590 ();
 b15zdnd11an1n08x5 FILLER_239_603 ();
 b15zdnd11an1n64x5 FILLER_239_619 ();
 b15zdnd11an1n32x5 FILLER_239_683 ();
 b15zdnd11an1n16x5 FILLER_239_715 ();
 b15zdnd11an1n04x5 FILLER_239_731 ();
 b15zdnd00an1n02x5 FILLER_239_735 ();
 b15zdnd11an1n32x5 FILLER_239_744 ();
 b15zdnd11an1n16x5 FILLER_239_776 ();
 b15zdnd00an1n01x5 FILLER_239_792 ();
 b15zdnd11an1n04x5 FILLER_239_814 ();
 b15zdnd11an1n08x5 FILLER_239_844 ();
 b15zdnd11an1n04x5 FILLER_239_852 ();
 b15zdnd00an1n01x5 FILLER_239_856 ();
 b15zdnd11an1n16x5 FILLER_239_883 ();
 b15zdnd11an1n08x5 FILLER_239_899 ();
 b15zdnd11an1n04x5 FILLER_239_907 ();
 b15zdnd11an1n32x5 FILLER_239_920 ();
 b15zdnd11an1n16x5 FILLER_239_952 ();
 b15zdnd11an1n08x5 FILLER_239_968 ();
 b15zdnd00an1n02x5 FILLER_239_976 ();
 b15zdnd00an1n01x5 FILLER_239_978 ();
 b15zdnd11an1n04x5 FILLER_239_997 ();
 b15zdnd11an1n64x5 FILLER_239_1010 ();
 b15zdnd11an1n08x5 FILLER_239_1074 ();
 b15zdnd11an1n04x5 FILLER_239_1082 ();
 b15zdnd00an1n02x5 FILLER_239_1086 ();
 b15zdnd11an1n04x5 FILLER_239_1106 ();
 b15zdnd11an1n16x5 FILLER_239_1116 ();
 b15zdnd11an1n08x5 FILLER_239_1132 ();
 b15zdnd11an1n04x5 FILLER_239_1140 ();
 b15zdnd11an1n04x5 FILLER_239_1150 ();
 b15zdnd00an1n02x5 FILLER_239_1154 ();
 b15zdnd11an1n64x5 FILLER_239_1169 ();
 b15zdnd11an1n08x5 FILLER_239_1233 ();
 b15zdnd00an1n02x5 FILLER_239_1241 ();
 b15zdnd00an1n01x5 FILLER_239_1243 ();
 b15zdnd11an1n32x5 FILLER_239_1251 ();
 b15zdnd11an1n08x5 FILLER_239_1283 ();
 b15zdnd00an1n01x5 FILLER_239_1291 ();
 b15zdnd11an1n64x5 FILLER_239_1323 ();
 b15zdnd11an1n64x5 FILLER_239_1387 ();
 b15zdnd11an1n64x5 FILLER_239_1451 ();
 b15zdnd11an1n64x5 FILLER_239_1515 ();
 b15zdnd11an1n16x5 FILLER_239_1579 ();
 b15zdnd11an1n08x5 FILLER_239_1595 ();
 b15zdnd00an1n02x5 FILLER_239_1603 ();
 b15zdnd11an1n04x5 FILLER_239_1615 ();
 b15zdnd11an1n16x5 FILLER_239_1629 ();
 b15zdnd11an1n04x5 FILLER_239_1645 ();
 b15zdnd11an1n16x5 FILLER_239_1654 ();
 b15zdnd11an1n08x5 FILLER_239_1670 ();
 b15zdnd11an1n04x5 FILLER_239_1678 ();
 b15zdnd00an1n02x5 FILLER_239_1682 ();
 b15zdnd00an1n01x5 FILLER_239_1684 ();
 b15zdnd11an1n04x5 FILLER_239_1697 ();
 b15zdnd00an1n02x5 FILLER_239_1701 ();
 b15zdnd11an1n04x5 FILLER_239_1712 ();
 b15zdnd11an1n04x5 FILLER_239_1721 ();
 b15zdnd00an1n02x5 FILLER_239_1725 ();
 b15zdnd00an1n01x5 FILLER_239_1727 ();
 b15zdnd11an1n16x5 FILLER_239_1736 ();
 b15zdnd11an1n04x5 FILLER_239_1752 ();
 b15zdnd00an1n02x5 FILLER_239_1756 ();
 b15zdnd00an1n01x5 FILLER_239_1758 ();
 b15zdnd11an1n32x5 FILLER_239_1775 ();
 b15zdnd11an1n16x5 FILLER_239_1807 ();
 b15zdnd11an1n08x5 FILLER_239_1823 ();
 b15zdnd00an1n02x5 FILLER_239_1831 ();
 b15zdnd11an1n04x5 FILLER_239_1859 ();
 b15zdnd11an1n04x5 FILLER_239_1894 ();
 b15zdnd11an1n08x5 FILLER_239_1902 ();
 b15zdnd00an1n01x5 FILLER_239_1910 ();
 b15zdnd11an1n32x5 FILLER_239_1928 ();
 b15zdnd11an1n16x5 FILLER_239_1991 ();
 b15zdnd00an1n02x5 FILLER_239_2007 ();
 b15zdnd00an1n01x5 FILLER_239_2009 ();
 b15zdnd11an1n32x5 FILLER_239_2017 ();
 b15zdnd00an1n02x5 FILLER_239_2049 ();
 b15zdnd11an1n08x5 FILLER_239_2057 ();
 b15zdnd11an1n08x5 FILLER_239_2074 ();
 b15zdnd00an1n02x5 FILLER_239_2082 ();
 b15zdnd11an1n04x5 FILLER_239_2090 ();
 b15zdnd11an1n04x5 FILLER_239_2115 ();
 b15zdnd00an1n02x5 FILLER_239_2119 ();
 b15zdnd11an1n32x5 FILLER_239_2133 ();
 b15zdnd11an1n08x5 FILLER_239_2165 ();
 b15zdnd00an1n02x5 FILLER_239_2173 ();
 b15zdnd11an1n04x5 FILLER_239_2180 ();
 b15zdnd11an1n16x5 FILLER_239_2189 ();
 b15zdnd11an1n32x5 FILLER_239_2221 ();
 b15zdnd11an1n16x5 FILLER_239_2253 ();
 b15zdnd11an1n08x5 FILLER_239_2269 ();
 b15zdnd11an1n04x5 FILLER_239_2277 ();
 b15zdnd00an1n02x5 FILLER_239_2281 ();
 b15zdnd00an1n01x5 FILLER_239_2283 ();
 b15zdnd11an1n32x5 FILLER_240_8 ();
 b15zdnd11an1n08x5 FILLER_240_40 ();
 b15zdnd00an1n02x5 FILLER_240_48 ();
 b15zdnd00an1n01x5 FILLER_240_50 ();
 b15zdnd11an1n04x5 FILLER_240_56 ();
 b15zdnd00an1n02x5 FILLER_240_60 ();
 b15zdnd11an1n32x5 FILLER_240_78 ();
 b15zdnd00an1n01x5 FILLER_240_110 ();
 b15zdnd11an1n04x5 FILLER_240_120 ();
 b15zdnd11an1n16x5 FILLER_240_141 ();
 b15zdnd11an1n08x5 FILLER_240_157 ();
 b15zdnd11an1n04x5 FILLER_240_165 ();
 b15zdnd11an1n04x5 FILLER_240_195 ();
 b15zdnd00an1n02x5 FILLER_240_199 ();
 b15zdnd00an1n01x5 FILLER_240_201 ();
 b15zdnd11an1n16x5 FILLER_240_208 ();
 b15zdnd11an1n08x5 FILLER_240_239 ();
 b15zdnd11an1n04x5 FILLER_240_247 ();
 b15zdnd00an1n02x5 FILLER_240_251 ();
 b15zdnd00an1n01x5 FILLER_240_253 ();
 b15zdnd11an1n32x5 FILLER_240_261 ();
 b15zdnd11an1n16x5 FILLER_240_293 ();
 b15zdnd00an1n02x5 FILLER_240_309 ();
 b15zdnd11an1n08x5 FILLER_240_329 ();
 b15zdnd11an1n04x5 FILLER_240_347 ();
 b15zdnd11an1n32x5 FILLER_240_363 ();
 b15zdnd11an1n16x5 FILLER_240_395 ();
 b15zdnd11an1n08x5 FILLER_240_411 ();
 b15zdnd11an1n04x5 FILLER_240_419 ();
 b15zdnd00an1n02x5 FILLER_240_423 ();
 b15zdnd11an1n04x5 FILLER_240_433 ();
 b15zdnd11an1n04x5 FILLER_240_455 ();
 b15zdnd11an1n08x5 FILLER_240_468 ();
 b15zdnd00an1n01x5 FILLER_240_476 ();
 b15zdnd11an1n04x5 FILLER_240_483 ();
 b15zdnd11an1n08x5 FILLER_240_499 ();
 b15zdnd11an1n04x5 FILLER_240_507 ();
 b15zdnd00an1n02x5 FILLER_240_511 ();
 b15zdnd11an1n64x5 FILLER_240_528 ();
 b15zdnd11an1n04x5 FILLER_240_592 ();
 b15zdnd00an1n02x5 FILLER_240_596 ();
 b15zdnd00an1n01x5 FILLER_240_598 ();
 b15zdnd11an1n04x5 FILLER_240_604 ();
 b15zdnd11an1n32x5 FILLER_240_614 ();
 b15zdnd11an1n04x5 FILLER_240_646 ();
 b15zdnd00an1n02x5 FILLER_240_650 ();
 b15zdnd00an1n01x5 FILLER_240_652 ();
 b15zdnd11an1n08x5 FILLER_240_663 ();
 b15zdnd00an1n02x5 FILLER_240_671 ();
 b15zdnd00an1n01x5 FILLER_240_673 ();
 b15zdnd11an1n16x5 FILLER_240_679 ();
 b15zdnd11an1n04x5 FILLER_240_695 ();
 b15zdnd00an1n02x5 FILLER_240_699 ();
 b15zdnd00an1n01x5 FILLER_240_701 ();
 b15zdnd00an1n02x5 FILLER_240_716 ();
 b15zdnd11an1n08x5 FILLER_240_726 ();
 b15zdnd11an1n32x5 FILLER_240_744 ();
 b15zdnd11an1n16x5 FILLER_240_776 ();
 b15zdnd11an1n08x5 FILLER_240_792 ();
 b15zdnd11an1n04x5 FILLER_240_800 ();
 b15zdnd00an1n01x5 FILLER_240_804 ();
 b15zdnd11an1n32x5 FILLER_240_831 ();
 b15zdnd11an1n08x5 FILLER_240_863 ();
 b15zdnd11an1n04x5 FILLER_240_871 ();
 b15zdnd00an1n01x5 FILLER_240_875 ();
 b15zdnd11an1n32x5 FILLER_240_896 ();
 b15zdnd11an1n16x5 FILLER_240_928 ();
 b15zdnd11an1n08x5 FILLER_240_944 ();
 b15zdnd00an1n02x5 FILLER_240_952 ();
 b15zdnd00an1n01x5 FILLER_240_954 ();
 b15zdnd11an1n04x5 FILLER_240_971 ();
 b15zdnd00an1n01x5 FILLER_240_975 ();
 b15zdnd11an1n32x5 FILLER_240_982 ();
 b15zdnd11an1n08x5 FILLER_240_1014 ();
 b15zdnd00an1n02x5 FILLER_240_1022 ();
 b15zdnd11an1n04x5 FILLER_240_1030 ();
 b15zdnd00an1n02x5 FILLER_240_1034 ();
 b15zdnd00an1n01x5 FILLER_240_1036 ();
 b15zdnd11an1n04x5 FILLER_240_1042 ();
 b15zdnd11an1n08x5 FILLER_240_1051 ();
 b15zdnd00an1n01x5 FILLER_240_1059 ();
 b15zdnd11an1n04x5 FILLER_240_1076 ();
 b15zdnd00an1n01x5 FILLER_240_1080 ();
 b15zdnd11an1n08x5 FILLER_240_1086 ();
 b15zdnd00an1n02x5 FILLER_240_1094 ();
 b15zdnd00an1n01x5 FILLER_240_1096 ();
 b15zdnd11an1n16x5 FILLER_240_1104 ();
 b15zdnd00an1n02x5 FILLER_240_1120 ();
 b15zdnd11an1n04x5 FILLER_240_1140 ();
 b15zdnd00an1n02x5 FILLER_240_1144 ();
 b15zdnd00an1n01x5 FILLER_240_1146 ();
 b15zdnd11an1n04x5 FILLER_240_1159 ();
 b15zdnd00an1n01x5 FILLER_240_1163 ();
 b15zdnd11an1n16x5 FILLER_240_1170 ();
 b15zdnd11an1n08x5 FILLER_240_1186 ();
 b15zdnd11an1n04x5 FILLER_240_1194 ();
 b15zdnd00an1n02x5 FILLER_240_1198 ();
 b15zdnd00an1n01x5 FILLER_240_1200 ();
 b15zdnd11an1n64x5 FILLER_240_1206 ();
 b15zdnd11an1n32x5 FILLER_240_1270 ();
 b15zdnd11an1n04x5 FILLER_240_1302 ();
 b15zdnd00an1n01x5 FILLER_240_1306 ();
 b15zdnd11an1n16x5 FILLER_240_1330 ();
 b15zdnd11an1n08x5 FILLER_240_1346 ();
 b15zdnd00an1n02x5 FILLER_240_1354 ();
 b15zdnd00an1n01x5 FILLER_240_1356 ();
 b15zdnd11an1n64x5 FILLER_240_1381 ();
 b15zdnd11an1n32x5 FILLER_240_1445 ();
 b15zdnd11an1n08x5 FILLER_240_1477 ();
 b15zdnd11an1n04x5 FILLER_240_1485 ();
 b15zdnd00an1n01x5 FILLER_240_1489 ();
 b15zdnd11an1n64x5 FILLER_240_1500 ();
 b15zdnd11an1n16x5 FILLER_240_1564 ();
 b15zdnd00an1n02x5 FILLER_240_1580 ();
 b15zdnd00an1n01x5 FILLER_240_1582 ();
 b15zdnd11an1n32x5 FILLER_240_1587 ();
 b15zdnd11an1n16x5 FILLER_240_1619 ();
 b15zdnd11an1n08x5 FILLER_240_1635 ();
 b15zdnd00an1n02x5 FILLER_240_1643 ();
 b15zdnd00an1n01x5 FILLER_240_1645 ();
 b15zdnd11an1n16x5 FILLER_240_1651 ();
 b15zdnd11an1n08x5 FILLER_240_1667 ();
 b15zdnd11an1n04x5 FILLER_240_1675 ();
 b15zdnd00an1n02x5 FILLER_240_1679 ();
 b15zdnd00an1n01x5 FILLER_240_1681 ();
 b15zdnd11an1n64x5 FILLER_240_1689 ();
 b15zdnd11an1n16x5 FILLER_240_1753 ();
 b15zdnd11an1n04x5 FILLER_240_1769 ();
 b15zdnd11an1n64x5 FILLER_240_1786 ();
 b15zdnd11an1n32x5 FILLER_240_1850 ();
 b15zdnd11an1n08x5 FILLER_240_1882 ();
 b15zdnd11an1n04x5 FILLER_240_1890 ();
 b15zdnd00an1n02x5 FILLER_240_1894 ();
 b15zdnd00an1n01x5 FILLER_240_1896 ();
 b15zdnd11an1n16x5 FILLER_240_1904 ();
 b15zdnd00an1n02x5 FILLER_240_1920 ();
 b15zdnd11an1n08x5 FILLER_240_1936 ();
 b15zdnd00an1n01x5 FILLER_240_1944 ();
 b15zdnd11an1n04x5 FILLER_240_1955 ();
 b15zdnd11an1n16x5 FILLER_240_1971 ();
 b15zdnd00an1n01x5 FILLER_240_1987 ();
 b15zdnd11an1n64x5 FILLER_240_2020 ();
 b15zdnd11an1n16x5 FILLER_240_2084 ();
 b15zdnd00an1n02x5 FILLER_240_2100 ();
 b15zdnd00an1n01x5 FILLER_240_2102 ();
 b15zdnd11an1n08x5 FILLER_240_2115 ();
 b15zdnd11an1n04x5 FILLER_240_2123 ();
 b15zdnd11an1n08x5 FILLER_240_2143 ();
 b15zdnd00an1n02x5 FILLER_240_2151 ();
 b15zdnd00an1n01x5 FILLER_240_2153 ();
 b15zdnd11an1n16x5 FILLER_240_2162 ();
 b15zdnd11an1n04x5 FILLER_240_2178 ();
 b15zdnd11an1n16x5 FILLER_240_2188 ();
 b15zdnd11an1n04x5 FILLER_240_2220 ();
 b15zdnd00an1n01x5 FILLER_240_2224 ();
 b15zdnd11an1n08x5 FILLER_240_2241 ();
 b15zdnd11an1n04x5 FILLER_240_2249 ();
 b15zdnd00an1n01x5 FILLER_240_2253 ();
 b15zdnd00an1n02x5 FILLER_240_2274 ();
 b15zdnd11an1n32x5 FILLER_241_0 ();
 b15zdnd11an1n04x5 FILLER_241_32 ();
 b15zdnd00an1n01x5 FILLER_241_36 ();
 b15zdnd11an1n64x5 FILLER_241_53 ();
 b15zdnd11an1n64x5 FILLER_241_117 ();
 b15zdnd11an1n32x5 FILLER_241_181 ();
 b15zdnd11an1n08x5 FILLER_241_213 ();
 b15zdnd11an1n04x5 FILLER_241_221 ();
 b15zdnd00an1n02x5 FILLER_241_225 ();
 b15zdnd11an1n16x5 FILLER_241_233 ();
 b15zdnd11an1n04x5 FILLER_241_249 ();
 b15zdnd11an1n16x5 FILLER_241_258 ();
 b15zdnd11an1n04x5 FILLER_241_274 ();
 b15zdnd00an1n02x5 FILLER_241_278 ();
 b15zdnd11an1n04x5 FILLER_241_284 ();
 b15zdnd11an1n08x5 FILLER_241_299 ();
 b15zdnd11an1n04x5 FILLER_241_307 ();
 b15zdnd11an1n64x5 FILLER_241_327 ();
 b15zdnd11an1n64x5 FILLER_241_391 ();
 b15zdnd11an1n16x5 FILLER_241_455 ();
 b15zdnd11an1n08x5 FILLER_241_475 ();
 b15zdnd00an1n01x5 FILLER_241_483 ();
 b15zdnd11an1n04x5 FILLER_241_490 ();
 b15zdnd00an1n02x5 FILLER_241_494 ();
 b15zdnd00an1n01x5 FILLER_241_496 ();
 b15zdnd11an1n04x5 FILLER_241_503 ();
 b15zdnd00an1n01x5 FILLER_241_507 ();
 b15zdnd11an1n04x5 FILLER_241_514 ();
 b15zdnd00an1n01x5 FILLER_241_518 ();
 b15zdnd11an1n04x5 FILLER_241_524 ();
 b15zdnd11an1n16x5 FILLER_241_534 ();
 b15zdnd11an1n08x5 FILLER_241_550 ();
 b15zdnd00an1n01x5 FILLER_241_558 ();
 b15zdnd11an1n04x5 FILLER_241_572 ();
 b15zdnd11an1n16x5 FILLER_241_581 ();
 b15zdnd11an1n04x5 FILLER_241_597 ();
 b15zdnd11an1n16x5 FILLER_241_613 ();
 b15zdnd00an1n02x5 FILLER_241_629 ();
 b15zdnd00an1n01x5 FILLER_241_631 ();
 b15zdnd11an1n16x5 FILLER_241_648 ();
 b15zdnd11an1n08x5 FILLER_241_664 ();
 b15zdnd11an1n04x5 FILLER_241_672 ();
 b15zdnd00an1n02x5 FILLER_241_676 ();
 b15zdnd11an1n04x5 FILLER_241_684 ();
 b15zdnd00an1n02x5 FILLER_241_688 ();
 b15zdnd00an1n01x5 FILLER_241_690 ();
 b15zdnd11an1n04x5 FILLER_241_696 ();
 b15zdnd11an1n16x5 FILLER_241_719 ();
 b15zdnd11an1n04x5 FILLER_241_743 ();
 b15zdnd00an1n02x5 FILLER_241_747 ();
 b15zdnd11an1n16x5 FILLER_241_753 ();
 b15zdnd11an1n08x5 FILLER_241_769 ();
 b15zdnd00an1n02x5 FILLER_241_777 ();
 b15zdnd11an1n16x5 FILLER_241_787 ();
 b15zdnd11an1n08x5 FILLER_241_803 ();
 b15zdnd00an1n02x5 FILLER_241_811 ();
 b15zdnd00an1n01x5 FILLER_241_813 ();
 b15zdnd11an1n04x5 FILLER_241_830 ();
 b15zdnd11an1n08x5 FILLER_241_860 ();
 b15zdnd11an1n04x5 FILLER_241_868 ();
 b15zdnd00an1n02x5 FILLER_241_872 ();
 b15zdnd11an1n08x5 FILLER_241_879 ();
 b15zdnd11an1n64x5 FILLER_241_891 ();
 b15zdnd11an1n16x5 FILLER_241_955 ();
 b15zdnd11an1n08x5 FILLER_241_971 ();
 b15zdnd11an1n04x5 FILLER_241_979 ();
 b15zdnd11an1n08x5 FILLER_241_989 ();
 b15zdnd00an1n02x5 FILLER_241_997 ();
 b15zdnd00an1n01x5 FILLER_241_999 ();
 b15zdnd11an1n08x5 FILLER_241_1012 ();
 b15zdnd00an1n01x5 FILLER_241_1020 ();
 b15zdnd11an1n32x5 FILLER_241_1033 ();
 b15zdnd00an1n01x5 FILLER_241_1065 ();
 b15zdnd11an1n04x5 FILLER_241_1077 ();
 b15zdnd00an1n02x5 FILLER_241_1081 ();
 b15zdnd11an1n04x5 FILLER_241_1097 ();
 b15zdnd00an1n02x5 FILLER_241_1101 ();
 b15zdnd11an1n16x5 FILLER_241_1109 ();
 b15zdnd11an1n08x5 FILLER_241_1129 ();
 b15zdnd11an1n04x5 FILLER_241_1137 ();
 b15zdnd00an1n02x5 FILLER_241_1141 ();
 b15zdnd11an1n08x5 FILLER_241_1149 ();
 b15zdnd11an1n04x5 FILLER_241_1157 ();
 b15zdnd11an1n08x5 FILLER_241_1187 ();
 b15zdnd11an1n04x5 FILLER_241_1195 ();
 b15zdnd00an1n02x5 FILLER_241_1199 ();
 b15zdnd00an1n01x5 FILLER_241_1201 ();
 b15zdnd11an1n16x5 FILLER_241_1208 ();
 b15zdnd11an1n08x5 FILLER_241_1224 ();
 b15zdnd00an1n01x5 FILLER_241_1232 ();
 b15zdnd11an1n04x5 FILLER_241_1242 ();
 b15zdnd11an1n16x5 FILLER_241_1250 ();
 b15zdnd11an1n08x5 FILLER_241_1266 ();
 b15zdnd00an1n01x5 FILLER_241_1274 ();
 b15zdnd11an1n16x5 FILLER_241_1280 ();
 b15zdnd00an1n02x5 FILLER_241_1296 ();
 b15zdnd11an1n32x5 FILLER_241_1315 ();
 b15zdnd00an1n02x5 FILLER_241_1347 ();
 b15zdnd00an1n01x5 FILLER_241_1349 ();
 b15zdnd11an1n04x5 FILLER_241_1382 ();
 b15zdnd11an1n04x5 FILLER_241_1417 ();
 b15zdnd11an1n64x5 FILLER_241_1452 ();
 b15zdnd11an1n08x5 FILLER_241_1516 ();
 b15zdnd00an1n02x5 FILLER_241_1524 ();
 b15zdnd00an1n01x5 FILLER_241_1526 ();
 b15zdnd11an1n16x5 FILLER_241_1536 ();
 b15zdnd11an1n04x5 FILLER_241_1552 ();
 b15zdnd00an1n01x5 FILLER_241_1556 ();
 b15zdnd11an1n16x5 FILLER_241_1565 ();
 b15zdnd11an1n08x5 FILLER_241_1581 ();
 b15zdnd11an1n04x5 FILLER_241_1589 ();
 b15zdnd00an1n02x5 FILLER_241_1593 ();
 b15zdnd00an1n01x5 FILLER_241_1595 ();
 b15zdnd11an1n04x5 FILLER_241_1602 ();
 b15zdnd00an1n01x5 FILLER_241_1606 ();
 b15zdnd11an1n64x5 FILLER_241_1613 ();
 b15zdnd11an1n64x5 FILLER_241_1677 ();
 b15zdnd11an1n64x5 FILLER_241_1741 ();
 b15zdnd11an1n64x5 FILLER_241_1805 ();
 b15zdnd11an1n16x5 FILLER_241_1869 ();
 b15zdnd00an1n01x5 FILLER_241_1885 ();
 b15zdnd11an1n04x5 FILLER_241_1891 ();
 b15zdnd11an1n04x5 FILLER_241_1910 ();
 b15zdnd11an1n04x5 FILLER_241_1924 ();
 b15zdnd00an1n02x5 FILLER_241_1928 ();
 b15zdnd11an1n64x5 FILLER_241_1940 ();
 b15zdnd11an1n32x5 FILLER_241_2004 ();
 b15zdnd11an1n08x5 FILLER_241_2036 ();
 b15zdnd00an1n01x5 FILLER_241_2044 ();
 b15zdnd11an1n64x5 FILLER_241_2052 ();
 b15zdnd11an1n64x5 FILLER_241_2116 ();
 b15zdnd11an1n04x5 FILLER_241_2180 ();
 b15zdnd00an1n01x5 FILLER_241_2184 ();
 b15zdnd11an1n32x5 FILLER_241_2190 ();
 b15zdnd11an1n08x5 FILLER_241_2222 ();
 b15zdnd11an1n32x5 FILLER_241_2246 ();
 b15zdnd11an1n04x5 FILLER_241_2278 ();
 b15zdnd00an1n02x5 FILLER_241_2282 ();
 b15zdnd11an1n16x5 FILLER_242_8 ();
 b15zdnd11an1n08x5 FILLER_242_24 ();
 b15zdnd11an1n16x5 FILLER_242_40 ();
 b15zdnd11an1n08x5 FILLER_242_56 ();
 b15zdnd11an1n04x5 FILLER_242_64 ();
 b15zdnd00an1n02x5 FILLER_242_68 ();
 b15zdnd00an1n01x5 FILLER_242_70 ();
 b15zdnd11an1n04x5 FILLER_242_75 ();
 b15zdnd11an1n64x5 FILLER_242_86 ();
 b15zdnd11an1n04x5 FILLER_242_150 ();
 b15zdnd00an1n01x5 FILLER_242_154 ();
 b15zdnd11an1n04x5 FILLER_242_169 ();
 b15zdnd11an1n64x5 FILLER_242_177 ();
 b15zdnd11an1n64x5 FILLER_242_241 ();
 b15zdnd11an1n16x5 FILLER_242_305 ();
 b15zdnd00an1n02x5 FILLER_242_321 ();
 b15zdnd11an1n64x5 FILLER_242_344 ();
 b15zdnd11an1n32x5 FILLER_242_408 ();
 b15zdnd11an1n08x5 FILLER_242_440 ();
 b15zdnd11an1n04x5 FILLER_242_448 ();
 b15zdnd00an1n02x5 FILLER_242_452 ();
 b15zdnd11an1n16x5 FILLER_242_459 ();
 b15zdnd11an1n08x5 FILLER_242_475 ();
 b15zdnd00an1n02x5 FILLER_242_483 ();
 b15zdnd00an1n01x5 FILLER_242_485 ();
 b15zdnd11an1n32x5 FILLER_242_492 ();
 b15zdnd11an1n08x5 FILLER_242_524 ();
 b15zdnd11an1n04x5 FILLER_242_532 ();
 b15zdnd00an1n02x5 FILLER_242_536 ();
 b15zdnd00an1n01x5 FILLER_242_538 ();
 b15zdnd11an1n32x5 FILLER_242_543 ();
 b15zdnd11an1n04x5 FILLER_242_575 ();
 b15zdnd00an1n01x5 FILLER_242_579 ();
 b15zdnd11an1n16x5 FILLER_242_584 ();
 b15zdnd11an1n04x5 FILLER_242_600 ();
 b15zdnd11an1n08x5 FILLER_242_614 ();
 b15zdnd00an1n01x5 FILLER_242_622 ();
 b15zdnd11an1n08x5 FILLER_242_641 ();
 b15zdnd00an1n02x5 FILLER_242_649 ();
 b15zdnd00an1n01x5 FILLER_242_651 ();
 b15zdnd11an1n16x5 FILLER_242_668 ();
 b15zdnd11an1n16x5 FILLER_242_691 ();
 b15zdnd11an1n08x5 FILLER_242_707 ();
 b15zdnd00an1n02x5 FILLER_242_715 ();
 b15zdnd00an1n01x5 FILLER_242_717 ();
 b15zdnd11an1n08x5 FILLER_242_726 ();
 b15zdnd11an1n04x5 FILLER_242_734 ();
 b15zdnd00an1n02x5 FILLER_242_738 ();
 b15zdnd00an1n01x5 FILLER_242_740 ();
 b15zdnd11an1n04x5 FILLER_242_751 ();
 b15zdnd11an1n04x5 FILLER_242_774 ();
 b15zdnd11an1n04x5 FILLER_242_785 ();
 b15zdnd00an1n02x5 FILLER_242_789 ();
 b15zdnd00an1n01x5 FILLER_242_791 ();
 b15zdnd11an1n16x5 FILLER_242_808 ();
 b15zdnd11an1n64x5 FILLER_242_850 ();
 b15zdnd11an1n32x5 FILLER_242_914 ();
 b15zdnd11an1n16x5 FILLER_242_946 ();
 b15zdnd11an1n08x5 FILLER_242_962 ();
 b15zdnd00an1n01x5 FILLER_242_970 ();
 b15zdnd11an1n04x5 FILLER_242_989 ();
 b15zdnd11an1n16x5 FILLER_242_1009 ();
 b15zdnd11an1n08x5 FILLER_242_1025 ();
 b15zdnd11an1n04x5 FILLER_242_1033 ();
 b15zdnd00an1n02x5 FILLER_242_1037 ();
 b15zdnd11an1n04x5 FILLER_242_1057 ();
 b15zdnd11an1n16x5 FILLER_242_1079 ();
 b15zdnd11an1n08x5 FILLER_242_1095 ();
 b15zdnd11an1n04x5 FILLER_242_1103 ();
 b15zdnd00an1n01x5 FILLER_242_1107 ();
 b15zdnd11an1n08x5 FILLER_242_1115 ();
 b15zdnd00an1n02x5 FILLER_242_1123 ();
 b15zdnd00an1n01x5 FILLER_242_1125 ();
 b15zdnd11an1n32x5 FILLER_242_1133 ();
 b15zdnd11an1n04x5 FILLER_242_1165 ();
 b15zdnd00an1n02x5 FILLER_242_1169 ();
 b15zdnd11an1n16x5 FILLER_242_1175 ();
 b15zdnd11an1n04x5 FILLER_242_1191 ();
 b15zdnd11an1n04x5 FILLER_242_1202 ();
 b15zdnd00an1n02x5 FILLER_242_1206 ();
 b15zdnd11an1n04x5 FILLER_242_1213 ();
 b15zdnd00an1n02x5 FILLER_242_1217 ();
 b15zdnd11an1n16x5 FILLER_242_1229 ();
 b15zdnd11an1n04x5 FILLER_242_1245 ();
 b15zdnd00an1n02x5 FILLER_242_1249 ();
 b15zdnd11an1n04x5 FILLER_242_1275 ();
 b15zdnd11an1n16x5 FILLER_242_1293 ();
 b15zdnd11an1n08x5 FILLER_242_1309 ();
 b15zdnd11an1n04x5 FILLER_242_1317 ();
 b15zdnd00an1n02x5 FILLER_242_1321 ();
 b15zdnd00an1n01x5 FILLER_242_1323 ();
 b15zdnd11an1n16x5 FILLER_242_1329 ();
 b15zdnd11an1n04x5 FILLER_242_1345 ();
 b15zdnd00an1n02x5 FILLER_242_1349 ();
 b15zdnd00an1n01x5 FILLER_242_1351 ();
 b15zdnd11an1n64x5 FILLER_242_1383 ();
 b15zdnd11an1n16x5 FILLER_242_1447 ();
 b15zdnd11an1n08x5 FILLER_242_1463 ();
 b15zdnd00an1n02x5 FILLER_242_1471 ();
 b15zdnd00an1n01x5 FILLER_242_1473 ();
 b15zdnd11an1n04x5 FILLER_242_1500 ();
 b15zdnd11an1n16x5 FILLER_242_1514 ();
 b15zdnd11an1n08x5 FILLER_242_1530 ();
 b15zdnd11an1n04x5 FILLER_242_1544 ();
 b15zdnd11an1n04x5 FILLER_242_1574 ();
 b15zdnd11an1n08x5 FILLER_242_1582 ();
 b15zdnd00an1n01x5 FILLER_242_1590 ();
 b15zdnd11an1n08x5 FILLER_242_1600 ();
 b15zdnd11an1n64x5 FILLER_242_1624 ();
 b15zdnd11an1n32x5 FILLER_242_1688 ();
 b15zdnd00an1n01x5 FILLER_242_1720 ();
 b15zdnd11an1n16x5 FILLER_242_1729 ();
 b15zdnd11an1n08x5 FILLER_242_1745 ();
 b15zdnd00an1n01x5 FILLER_242_1753 ();
 b15zdnd11an1n04x5 FILLER_242_1770 ();
 b15zdnd11an1n16x5 FILLER_242_1779 ();
 b15zdnd11an1n08x5 FILLER_242_1795 ();
 b15zdnd00an1n02x5 FILLER_242_1803 ();
 b15zdnd11an1n04x5 FILLER_242_1810 ();
 b15zdnd11an1n16x5 FILLER_242_1823 ();
 b15zdnd00an1n01x5 FILLER_242_1839 ();
 b15zdnd11an1n16x5 FILLER_242_1860 ();
 b15zdnd11an1n16x5 FILLER_242_1902 ();
 b15zdnd11an1n08x5 FILLER_242_1918 ();
 b15zdnd11an1n04x5 FILLER_242_1926 ();
 b15zdnd00an1n01x5 FILLER_242_1930 ();
 b15zdnd11an1n32x5 FILLER_242_1943 ();
 b15zdnd11an1n16x5 FILLER_242_1975 ();
 b15zdnd11an1n08x5 FILLER_242_1991 ();
 b15zdnd11an1n04x5 FILLER_242_1999 ();
 b15zdnd00an1n01x5 FILLER_242_2003 ();
 b15zdnd11an1n04x5 FILLER_242_2009 ();
 b15zdnd00an1n01x5 FILLER_242_2013 ();
 b15zdnd11an1n32x5 FILLER_242_2022 ();
 b15zdnd11an1n32x5 FILLER_242_2060 ();
 b15zdnd11an1n16x5 FILLER_242_2092 ();
 b15zdnd11an1n08x5 FILLER_242_2108 ();
 b15zdnd11an1n16x5 FILLER_242_2122 ();
 b15zdnd11an1n04x5 FILLER_242_2138 ();
 b15zdnd11an1n04x5 FILLER_242_2150 ();
 b15zdnd11an1n64x5 FILLER_242_2162 ();
 b15zdnd11an1n32x5 FILLER_242_2226 ();
 b15zdnd11an1n16x5 FILLER_242_2258 ();
 b15zdnd00an1n02x5 FILLER_242_2274 ();
 b15zdnd11an1n64x5 FILLER_243_0 ();
 b15zdnd11an1n16x5 FILLER_243_64 ();
 b15zdnd00an1n01x5 FILLER_243_80 ();
 b15zdnd11an1n08x5 FILLER_243_95 ();
 b15zdnd11an1n04x5 FILLER_243_103 ();
 b15zdnd00an1n01x5 FILLER_243_107 ();
 b15zdnd11an1n16x5 FILLER_243_120 ();
 b15zdnd00an1n02x5 FILLER_243_136 ();
 b15zdnd00an1n01x5 FILLER_243_138 ();
 b15zdnd11an1n08x5 FILLER_243_144 ();
 b15zdnd11an1n04x5 FILLER_243_161 ();
 b15zdnd00an1n02x5 FILLER_243_165 ();
 b15zdnd11an1n16x5 FILLER_243_183 ();
 b15zdnd11an1n08x5 FILLER_243_199 ();
 b15zdnd11an1n04x5 FILLER_243_207 ();
 b15zdnd00an1n02x5 FILLER_243_211 ();
 b15zdnd00an1n01x5 FILLER_243_213 ();
 b15zdnd11an1n32x5 FILLER_243_225 ();
 b15zdnd11an1n16x5 FILLER_243_257 ();
 b15zdnd11an1n08x5 FILLER_243_273 ();
 b15zdnd11an1n04x5 FILLER_243_281 ();
 b15zdnd00an1n02x5 FILLER_243_285 ();
 b15zdnd11an1n16x5 FILLER_243_292 ();
 b15zdnd11an1n04x5 FILLER_243_308 ();
 b15zdnd00an1n02x5 FILLER_243_312 ();
 b15zdnd00an1n01x5 FILLER_243_314 ();
 b15zdnd11an1n64x5 FILLER_243_331 ();
 b15zdnd11an1n64x5 FILLER_243_395 ();
 b15zdnd11an1n64x5 FILLER_243_459 ();
 b15zdnd11an1n08x5 FILLER_243_523 ();
 b15zdnd11an1n04x5 FILLER_243_531 ();
 b15zdnd00an1n02x5 FILLER_243_535 ();
 b15zdnd00an1n01x5 FILLER_243_537 ();
 b15zdnd11an1n64x5 FILLER_243_550 ();
 b15zdnd11an1n32x5 FILLER_243_614 ();
 b15zdnd11an1n08x5 FILLER_243_646 ();
 b15zdnd11an1n04x5 FILLER_243_654 ();
 b15zdnd00an1n02x5 FILLER_243_658 ();
 b15zdnd11an1n64x5 FILLER_243_670 ();
 b15zdnd11an1n16x5 FILLER_243_734 ();
 b15zdnd11an1n08x5 FILLER_243_750 ();
 b15zdnd00an1n02x5 FILLER_243_758 ();
 b15zdnd00an1n01x5 FILLER_243_760 ();
 b15zdnd11an1n08x5 FILLER_243_771 ();
 b15zdnd11an1n16x5 FILLER_243_784 ();
 b15zdnd11an1n04x5 FILLER_243_800 ();
 b15zdnd00an1n02x5 FILLER_243_804 ();
 b15zdnd00an1n01x5 FILLER_243_806 ();
 b15zdnd11an1n08x5 FILLER_243_817 ();
 b15zdnd11an1n04x5 FILLER_243_825 ();
 b15zdnd00an1n02x5 FILLER_243_829 ();
 b15zdnd11an1n64x5 FILLER_243_857 ();
 b15zdnd11an1n64x5 FILLER_243_921 ();
 b15zdnd11an1n64x5 FILLER_243_985 ();
 b15zdnd11an1n64x5 FILLER_243_1049 ();
 b15zdnd11an1n32x5 FILLER_243_1113 ();
 b15zdnd11an1n16x5 FILLER_243_1145 ();
 b15zdnd11an1n04x5 FILLER_243_1161 ();
 b15zdnd11an1n32x5 FILLER_243_1180 ();
 b15zdnd11an1n04x5 FILLER_243_1212 ();
 b15zdnd00an1n02x5 FILLER_243_1216 ();
 b15zdnd00an1n01x5 FILLER_243_1218 ();
 b15zdnd11an1n64x5 FILLER_243_1229 ();
 b15zdnd11an1n16x5 FILLER_243_1293 ();
 b15zdnd00an1n01x5 FILLER_243_1309 ();
 b15zdnd11an1n04x5 FILLER_243_1319 ();
 b15zdnd11an1n16x5 FILLER_243_1330 ();
 b15zdnd11an1n04x5 FILLER_243_1346 ();
 b15zdnd11an1n64x5 FILLER_243_1382 ();
 b15zdnd11an1n16x5 FILLER_243_1446 ();
 b15zdnd11an1n08x5 FILLER_243_1462 ();
 b15zdnd11an1n04x5 FILLER_243_1470 ();
 b15zdnd00an1n02x5 FILLER_243_1474 ();
 b15zdnd11an1n04x5 FILLER_243_1502 ();
 b15zdnd11an1n16x5 FILLER_243_1513 ();
 b15zdnd00an1n02x5 FILLER_243_1529 ();
 b15zdnd00an1n01x5 FILLER_243_1531 ();
 b15zdnd11an1n32x5 FILLER_243_1537 ();
 b15zdnd00an1n01x5 FILLER_243_1569 ();
 b15zdnd11an1n32x5 FILLER_243_1582 ();
 b15zdnd11an1n16x5 FILLER_243_1614 ();
 b15zdnd11an1n08x5 FILLER_243_1630 ();
 b15zdnd00an1n02x5 FILLER_243_1638 ();
 b15zdnd00an1n01x5 FILLER_243_1640 ();
 b15zdnd11an1n32x5 FILLER_243_1650 ();
 b15zdnd00an1n02x5 FILLER_243_1682 ();
 b15zdnd11an1n16x5 FILLER_243_1698 ();
 b15zdnd11an1n04x5 FILLER_243_1719 ();
 b15zdnd11an1n04x5 FILLER_243_1737 ();
 b15zdnd11an1n04x5 FILLER_243_1746 ();
 b15zdnd11an1n04x5 FILLER_243_1776 ();
 b15zdnd11an1n04x5 FILLER_243_1785 ();
 b15zdnd11an1n64x5 FILLER_243_1794 ();
 b15zdnd11an1n64x5 FILLER_243_1858 ();
 b15zdnd11an1n64x5 FILLER_243_1922 ();
 b15zdnd11an1n16x5 FILLER_243_1986 ();
 b15zdnd00an1n01x5 FILLER_243_2002 ();
 b15zdnd11an1n32x5 FILLER_243_2010 ();
 b15zdnd11an1n04x5 FILLER_243_2042 ();
 b15zdnd00an1n02x5 FILLER_243_2046 ();
 b15zdnd00an1n01x5 FILLER_243_2048 ();
 b15zdnd11an1n04x5 FILLER_243_2061 ();
 b15zdnd11an1n32x5 FILLER_243_2073 ();
 b15zdnd11an1n08x5 FILLER_243_2105 ();
 b15zdnd11an1n04x5 FILLER_243_2113 ();
 b15zdnd00an1n02x5 FILLER_243_2117 ();
 b15zdnd00an1n01x5 FILLER_243_2119 ();
 b15zdnd11an1n16x5 FILLER_243_2124 ();
 b15zdnd11an1n08x5 FILLER_243_2140 ();
 b15zdnd00an1n01x5 FILLER_243_2148 ();
 b15zdnd11an1n04x5 FILLER_243_2170 ();
 b15zdnd11an1n04x5 FILLER_243_2188 ();
 b15zdnd00an1n02x5 FILLER_243_2192 ();
 b15zdnd00an1n01x5 FILLER_243_2194 ();
 b15zdnd11an1n04x5 FILLER_243_2201 ();
 b15zdnd11an1n64x5 FILLER_243_2211 ();
 b15zdnd11an1n08x5 FILLER_243_2275 ();
 b15zdnd00an1n01x5 FILLER_243_2283 ();
 b15zdnd11an1n16x5 FILLER_244_8 ();
 b15zdnd00an1n02x5 FILLER_244_24 ();
 b15zdnd11an1n32x5 FILLER_244_30 ();
 b15zdnd11an1n16x5 FILLER_244_62 ();
 b15zdnd11an1n08x5 FILLER_244_78 ();
 b15zdnd11an1n04x5 FILLER_244_96 ();
 b15zdnd00an1n02x5 FILLER_244_100 ();
 b15zdnd11an1n04x5 FILLER_244_116 ();
 b15zdnd11an1n08x5 FILLER_244_127 ();
 b15zdnd11an1n04x5 FILLER_244_147 ();
 b15zdnd11an1n16x5 FILLER_244_159 ();
 b15zdnd00an1n02x5 FILLER_244_175 ();
 b15zdnd00an1n01x5 FILLER_244_177 ();
 b15zdnd11an1n16x5 FILLER_244_187 ();
 b15zdnd11an1n08x5 FILLER_244_203 ();
 b15zdnd11an1n04x5 FILLER_244_211 ();
 b15zdnd11an1n16x5 FILLER_244_221 ();
 b15zdnd11an1n08x5 FILLER_244_237 ();
 b15zdnd11an1n04x5 FILLER_244_245 ();
 b15zdnd00an1n02x5 FILLER_244_249 ();
 b15zdnd11an1n04x5 FILLER_244_257 ();
 b15zdnd11an1n16x5 FILLER_244_273 ();
 b15zdnd11an1n08x5 FILLER_244_289 ();
 b15zdnd11an1n04x5 FILLER_244_297 ();
 b15zdnd11an1n64x5 FILLER_244_309 ();
 b15zdnd11an1n64x5 FILLER_244_373 ();
 b15zdnd11an1n64x5 FILLER_244_437 ();
 b15zdnd11an1n16x5 FILLER_244_501 ();
 b15zdnd11an1n04x5 FILLER_244_517 ();
 b15zdnd00an1n02x5 FILLER_244_521 ();
 b15zdnd11an1n64x5 FILLER_244_534 ();
 b15zdnd11an1n64x5 FILLER_244_598 ();
 b15zdnd11an1n32x5 FILLER_244_662 ();
 b15zdnd11an1n16x5 FILLER_244_694 ();
 b15zdnd11an1n08x5 FILLER_244_710 ();
 b15zdnd11an1n16x5 FILLER_244_726 ();
 b15zdnd11an1n04x5 FILLER_244_742 ();
 b15zdnd00an1n02x5 FILLER_244_746 ();
 b15zdnd00an1n01x5 FILLER_244_748 ();
 b15zdnd11an1n04x5 FILLER_244_769 ();
 b15zdnd00an1n02x5 FILLER_244_773 ();
 b15zdnd00an1n01x5 FILLER_244_775 ();
 b15zdnd11an1n64x5 FILLER_244_786 ();
 b15zdnd11an1n32x5 FILLER_244_850 ();
 b15zdnd11an1n16x5 FILLER_244_882 ();
 b15zdnd11an1n08x5 FILLER_244_898 ();
 b15zdnd00an1n02x5 FILLER_244_906 ();
 b15zdnd00an1n01x5 FILLER_244_908 ();
 b15zdnd11an1n64x5 FILLER_244_920 ();
 b15zdnd11an1n08x5 FILLER_244_984 ();
 b15zdnd00an1n01x5 FILLER_244_992 ();
 b15zdnd11an1n64x5 FILLER_244_1025 ();
 b15zdnd11an1n64x5 FILLER_244_1089 ();
 b15zdnd11an1n32x5 FILLER_244_1153 ();
 b15zdnd11an1n08x5 FILLER_244_1185 ();
 b15zdnd11an1n16x5 FILLER_244_1197 ();
 b15zdnd11an1n08x5 FILLER_244_1213 ();
 b15zdnd00an1n01x5 FILLER_244_1221 ();
 b15zdnd11an1n64x5 FILLER_244_1236 ();
 b15zdnd00an1n02x5 FILLER_244_1300 ();
 b15zdnd11an1n04x5 FILLER_244_1323 ();
 b15zdnd11an1n32x5 FILLER_244_1332 ();
 b15zdnd11an1n16x5 FILLER_244_1364 ();
 b15zdnd11an1n08x5 FILLER_244_1380 ();
 b15zdnd11an1n04x5 FILLER_244_1388 ();
 b15zdnd00an1n01x5 FILLER_244_1392 ();
 b15zdnd11an1n64x5 FILLER_244_1408 ();
 b15zdnd11an1n04x5 FILLER_244_1472 ();
 b15zdnd00an1n02x5 FILLER_244_1476 ();
 b15zdnd11an1n04x5 FILLER_244_1496 ();
 b15zdnd00an1n02x5 FILLER_244_1500 ();
 b15zdnd11an1n04x5 FILLER_244_1508 ();
 b15zdnd11an1n16x5 FILLER_244_1520 ();
 b15zdnd11an1n04x5 FILLER_244_1536 ();
 b15zdnd00an1n02x5 FILLER_244_1540 ();
 b15zdnd00an1n01x5 FILLER_244_1542 ();
 b15zdnd11an1n08x5 FILLER_244_1552 ();
 b15zdnd00an1n02x5 FILLER_244_1560 ();
 b15zdnd00an1n01x5 FILLER_244_1562 ();
 b15zdnd11an1n08x5 FILLER_244_1572 ();
 b15zdnd00an1n02x5 FILLER_244_1580 ();
 b15zdnd00an1n01x5 FILLER_244_1582 ();
 b15zdnd11an1n04x5 FILLER_244_1597 ();
 b15zdnd11an1n16x5 FILLER_244_1606 ();
 b15zdnd11an1n08x5 FILLER_244_1622 ();
 b15zdnd11an1n04x5 FILLER_244_1630 ();
 b15zdnd00an1n02x5 FILLER_244_1634 ();
 b15zdnd11an1n32x5 FILLER_244_1650 ();
 b15zdnd11an1n08x5 FILLER_244_1682 ();
 b15zdnd11an1n04x5 FILLER_244_1690 ();
 b15zdnd11an1n04x5 FILLER_244_1716 ();
 b15zdnd11an1n64x5 FILLER_244_1726 ();
 b15zdnd11an1n64x5 FILLER_244_1790 ();
 b15zdnd11an1n64x5 FILLER_244_1854 ();
 b15zdnd11an1n04x5 FILLER_244_1918 ();
 b15zdnd00an1n02x5 FILLER_244_1922 ();
 b15zdnd11an1n32x5 FILLER_244_1943 ();
 b15zdnd11an1n16x5 FILLER_244_1975 ();
 b15zdnd00an1n02x5 FILLER_244_1991 ();
 b15zdnd11an1n04x5 FILLER_244_1999 ();
 b15zdnd11an1n08x5 FILLER_244_2015 ();
 b15zdnd00an1n01x5 FILLER_244_2023 ();
 b15zdnd11an1n04x5 FILLER_244_2046 ();
 b15zdnd00an1n01x5 FILLER_244_2050 ();
 b15zdnd11an1n16x5 FILLER_244_2063 ();
 b15zdnd11an1n08x5 FILLER_244_2079 ();
 b15zdnd11an1n04x5 FILLER_244_2087 ();
 b15zdnd11an1n16x5 FILLER_244_2103 ();
 b15zdnd11an1n08x5 FILLER_244_2119 ();
 b15zdnd00an1n01x5 FILLER_244_2127 ();
 b15zdnd11an1n16x5 FILLER_244_2137 ();
 b15zdnd00an1n01x5 FILLER_244_2153 ();
 b15zdnd11an1n32x5 FILLER_244_2162 ();
 b15zdnd11an1n04x5 FILLER_244_2194 ();
 b15zdnd00an1n01x5 FILLER_244_2198 ();
 b15zdnd11an1n64x5 FILLER_244_2203 ();
 b15zdnd11an1n08x5 FILLER_244_2267 ();
 b15zdnd00an1n01x5 FILLER_244_2275 ();
 b15zdnd11an1n32x5 FILLER_245_0 ();
 b15zdnd11an1n04x5 FILLER_245_32 ();
 b15zdnd00an1n01x5 FILLER_245_36 ();
 b15zdnd11an1n04x5 FILLER_245_41 ();
 b15zdnd11an1n16x5 FILLER_245_57 ();
 b15zdnd11an1n64x5 FILLER_245_86 ();
 b15zdnd11an1n16x5 FILLER_245_150 ();
 b15zdnd11an1n08x5 FILLER_245_166 ();
 b15zdnd11an1n04x5 FILLER_245_174 ();
 b15zdnd00an1n02x5 FILLER_245_178 ();
 b15zdnd11an1n32x5 FILLER_245_196 ();
 b15zdnd11an1n16x5 FILLER_245_228 ();
 b15zdnd11an1n08x5 FILLER_245_244 ();
 b15zdnd11an1n04x5 FILLER_245_252 ();
 b15zdnd00an1n02x5 FILLER_245_256 ();
 b15zdnd11an1n16x5 FILLER_245_263 ();
 b15zdnd11an1n08x5 FILLER_245_279 ();
 b15zdnd00an1n02x5 FILLER_245_287 ();
 b15zdnd00an1n01x5 FILLER_245_289 ();
 b15zdnd11an1n16x5 FILLER_245_304 ();
 b15zdnd11an1n16x5 FILLER_245_333 ();
 b15zdnd11an1n04x5 FILLER_245_349 ();
 b15zdnd00an1n01x5 FILLER_245_353 ();
 b15zdnd11an1n64x5 FILLER_245_364 ();
 b15zdnd11an1n08x5 FILLER_245_428 ();
 b15zdnd11an1n32x5 FILLER_245_444 ();
 b15zdnd11an1n16x5 FILLER_245_476 ();
 b15zdnd11an1n08x5 FILLER_245_492 ();
 b15zdnd11an1n08x5 FILLER_245_505 ();
 b15zdnd00an1n02x5 FILLER_245_513 ();
 b15zdnd11an1n32x5 FILLER_245_531 ();
 b15zdnd11an1n08x5 FILLER_245_563 ();
 b15zdnd11an1n04x5 FILLER_245_571 ();
 b15zdnd11an1n08x5 FILLER_245_595 ();
 b15zdnd00an1n02x5 FILLER_245_603 ();
 b15zdnd00an1n01x5 FILLER_245_605 ();
 b15zdnd11an1n32x5 FILLER_245_612 ();
 b15zdnd11an1n16x5 FILLER_245_644 ();
 b15zdnd00an1n01x5 FILLER_245_660 ();
 b15zdnd11an1n04x5 FILLER_245_682 ();
 b15zdnd11an1n04x5 FILLER_245_692 ();
 b15zdnd00an1n02x5 FILLER_245_696 ();
 b15zdnd11an1n64x5 FILLER_245_703 ();
 b15zdnd11an1n32x5 FILLER_245_767 ();
 b15zdnd11an1n08x5 FILLER_245_799 ();
 b15zdnd11an1n04x5 FILLER_245_807 ();
 b15zdnd00an1n02x5 FILLER_245_811 ();
 b15zdnd11an1n04x5 FILLER_245_829 ();
 b15zdnd11an1n04x5 FILLER_245_853 ();
 b15zdnd00an1n02x5 FILLER_245_857 ();
 b15zdnd11an1n64x5 FILLER_245_863 ();
 b15zdnd11an1n32x5 FILLER_245_927 ();
 b15zdnd11an1n16x5 FILLER_245_959 ();
 b15zdnd11an1n04x5 FILLER_245_975 ();
 b15zdnd00an1n02x5 FILLER_245_979 ();
 b15zdnd00an1n01x5 FILLER_245_981 ();
 b15zdnd11an1n16x5 FILLER_245_1002 ();
 b15zdnd11an1n08x5 FILLER_245_1018 ();
 b15zdnd11an1n04x5 FILLER_245_1026 ();
 b15zdnd00an1n02x5 FILLER_245_1030 ();
 b15zdnd11an1n04x5 FILLER_245_1045 ();
 b15zdnd11an1n64x5 FILLER_245_1054 ();
 b15zdnd11an1n08x5 FILLER_245_1118 ();
 b15zdnd11an1n04x5 FILLER_245_1126 ();
 b15zdnd11an1n32x5 FILLER_245_1135 ();
 b15zdnd11an1n08x5 FILLER_245_1172 ();
 b15zdnd11an1n04x5 FILLER_245_1180 ();
 b15zdnd11an1n16x5 FILLER_245_1199 ();
 b15zdnd11an1n08x5 FILLER_245_1215 ();
 b15zdnd11an1n04x5 FILLER_245_1223 ();
 b15zdnd00an1n02x5 FILLER_245_1227 ();
 b15zdnd00an1n01x5 FILLER_245_1229 ();
 b15zdnd11an1n16x5 FILLER_245_1237 ();
 b15zdnd11an1n04x5 FILLER_245_1253 ();
 b15zdnd11an1n08x5 FILLER_245_1269 ();
 b15zdnd11an1n16x5 FILLER_245_1285 ();
 b15zdnd11an1n08x5 FILLER_245_1301 ();
 b15zdnd00an1n02x5 FILLER_245_1309 ();
 b15zdnd00an1n01x5 FILLER_245_1311 ();
 b15zdnd11an1n08x5 FILLER_245_1328 ();
 b15zdnd11an1n04x5 FILLER_245_1336 ();
 b15zdnd00an1n01x5 FILLER_245_1340 ();
 b15zdnd11an1n04x5 FILLER_245_1367 ();
 b15zdnd11an1n04x5 FILLER_245_1389 ();
 b15zdnd11an1n08x5 FILLER_245_1419 ();
 b15zdnd11an1n04x5 FILLER_245_1427 ();
 b15zdnd11an1n16x5 FILLER_245_1449 ();
 b15zdnd11an1n08x5 FILLER_245_1465 ();
 b15zdnd00an1n02x5 FILLER_245_1473 ();
 b15zdnd00an1n01x5 FILLER_245_1475 ();
 b15zdnd11an1n32x5 FILLER_245_1492 ();
 b15zdnd11an1n08x5 FILLER_245_1524 ();
 b15zdnd00an1n01x5 FILLER_245_1532 ();
 b15zdnd11an1n64x5 FILLER_245_1545 ();
 b15zdnd11an1n16x5 FILLER_245_1609 ();
 b15zdnd11an1n04x5 FILLER_245_1625 ();
 b15zdnd00an1n01x5 FILLER_245_1629 ();
 b15zdnd11an1n04x5 FILLER_245_1639 ();
 b15zdnd00an1n01x5 FILLER_245_1643 ();
 b15zdnd11an1n16x5 FILLER_245_1650 ();
 b15zdnd00an1n01x5 FILLER_245_1666 ();
 b15zdnd11an1n04x5 FILLER_245_1671 ();
 b15zdnd11an1n32x5 FILLER_245_1682 ();
 b15zdnd11an1n64x5 FILLER_245_1719 ();
 b15zdnd11an1n64x5 FILLER_245_1783 ();
 b15zdnd11an1n64x5 FILLER_245_1847 ();
 b15zdnd11an1n16x5 FILLER_245_1911 ();
 b15zdnd11an1n04x5 FILLER_245_1931 ();
 b15zdnd00an1n01x5 FILLER_245_1935 ();
 b15zdnd11an1n16x5 FILLER_245_1946 ();
 b15zdnd11an1n04x5 FILLER_245_1967 ();
 b15zdnd11an1n08x5 FILLER_245_1978 ();
 b15zdnd11an1n04x5 FILLER_245_1986 ();
 b15zdnd00an1n02x5 FILLER_245_1990 ();
 b15zdnd00an1n01x5 FILLER_245_1992 ();
 b15zdnd11an1n16x5 FILLER_245_2008 ();
 b15zdnd11an1n08x5 FILLER_245_2024 ();
 b15zdnd11an1n04x5 FILLER_245_2042 ();
 b15zdnd00an1n02x5 FILLER_245_2046 ();
 b15zdnd11an1n32x5 FILLER_245_2053 ();
 b15zdnd11an1n08x5 FILLER_245_2085 ();
 b15zdnd11an1n04x5 FILLER_245_2093 ();
 b15zdnd00an1n02x5 FILLER_245_2097 ();
 b15zdnd00an1n01x5 FILLER_245_2099 ();
 b15zdnd11an1n08x5 FILLER_245_2106 ();
 b15zdnd00an1n02x5 FILLER_245_2114 ();
 b15zdnd00an1n01x5 FILLER_245_2116 ();
 b15zdnd11an1n16x5 FILLER_245_2124 ();
 b15zdnd11an1n16x5 FILLER_245_2148 ();
 b15zdnd11an1n04x5 FILLER_245_2164 ();
 b15zdnd00an1n02x5 FILLER_245_2168 ();
 b15zdnd00an1n01x5 FILLER_245_2170 ();
 b15zdnd11an1n04x5 FILLER_245_2181 ();
 b15zdnd11an1n04x5 FILLER_245_2189 ();
 b15zdnd11an1n16x5 FILLER_245_2198 ();
 b15zdnd11an1n08x5 FILLER_245_2214 ();
 b15zdnd00an1n02x5 FILLER_245_2222 ();
 b15zdnd11an1n32x5 FILLER_245_2234 ();
 b15zdnd11an1n16x5 FILLER_245_2266 ();
 b15zdnd00an1n02x5 FILLER_245_2282 ();
 b15zdnd11an1n16x5 FILLER_246_8 ();
 b15zdnd11an1n08x5 FILLER_246_24 ();
 b15zdnd11an1n04x5 FILLER_246_32 ();
 b15zdnd00an1n01x5 FILLER_246_36 ();
 b15zdnd11an1n08x5 FILLER_246_68 ();
 b15zdnd11an1n04x5 FILLER_246_76 ();
 b15zdnd00an1n02x5 FILLER_246_80 ();
 b15zdnd11an1n32x5 FILLER_246_98 ();
 b15zdnd11an1n16x5 FILLER_246_130 ();
 b15zdnd11an1n08x5 FILLER_246_152 ();
 b15zdnd11an1n32x5 FILLER_246_179 ();
 b15zdnd11an1n16x5 FILLER_246_211 ();
 b15zdnd00an1n01x5 FILLER_246_227 ();
 b15zdnd11an1n64x5 FILLER_246_238 ();
 b15zdnd11an1n16x5 FILLER_246_302 ();
 b15zdnd11an1n08x5 FILLER_246_318 ();
 b15zdnd11an1n04x5 FILLER_246_326 ();
 b15zdnd00an1n02x5 FILLER_246_330 ();
 b15zdnd11an1n64x5 FILLER_246_337 ();
 b15zdnd11an1n16x5 FILLER_246_401 ();
 b15zdnd11an1n08x5 FILLER_246_417 ();
 b15zdnd11an1n04x5 FILLER_246_425 ();
 b15zdnd00an1n01x5 FILLER_246_429 ();
 b15zdnd11an1n08x5 FILLER_246_440 ();
 b15zdnd11an1n16x5 FILLER_246_453 ();
 b15zdnd11an1n04x5 FILLER_246_469 ();
 b15zdnd11an1n64x5 FILLER_246_485 ();
 b15zdnd11an1n16x5 FILLER_246_549 ();
 b15zdnd11an1n04x5 FILLER_246_565 ();
 b15zdnd00an1n02x5 FILLER_246_569 ();
 b15zdnd11an1n08x5 FILLER_246_575 ();
 b15zdnd00an1n01x5 FILLER_246_583 ();
 b15zdnd11an1n08x5 FILLER_246_598 ();
 b15zdnd00an1n01x5 FILLER_246_606 ();
 b15zdnd11an1n16x5 FILLER_246_617 ();
 b15zdnd00an1n01x5 FILLER_246_633 ();
 b15zdnd11an1n08x5 FILLER_246_646 ();
 b15zdnd00an1n01x5 FILLER_246_654 ();
 b15zdnd11an1n32x5 FILLER_246_668 ();
 b15zdnd00an1n02x5 FILLER_246_700 ();
 b15zdnd11an1n04x5 FILLER_246_712 ();
 b15zdnd00an1n02x5 FILLER_246_716 ();
 b15zdnd00an1n02x5 FILLER_246_726 ();
 b15zdnd11an1n08x5 FILLER_246_754 ();
 b15zdnd11an1n04x5 FILLER_246_762 ();
 b15zdnd11an1n64x5 FILLER_246_778 ();
 b15zdnd11an1n16x5 FILLER_246_842 ();
 b15zdnd11an1n04x5 FILLER_246_858 ();
 b15zdnd00an1n01x5 FILLER_246_862 ();
 b15zdnd11an1n32x5 FILLER_246_868 ();
 b15zdnd11an1n04x5 FILLER_246_900 ();
 b15zdnd00an1n01x5 FILLER_246_904 ();
 b15zdnd11an1n04x5 FILLER_246_910 ();
 b15zdnd11an1n32x5 FILLER_246_917 ();
 b15zdnd11an1n08x5 FILLER_246_949 ();
 b15zdnd11an1n04x5 FILLER_246_957 ();
 b15zdnd00an1n02x5 FILLER_246_961 ();
 b15zdnd00an1n01x5 FILLER_246_963 ();
 b15zdnd11an1n04x5 FILLER_246_971 ();
 b15zdnd11an1n16x5 FILLER_246_984 ();
 b15zdnd11an1n16x5 FILLER_246_1004 ();
 b15zdnd11an1n08x5 FILLER_246_1020 ();
 b15zdnd11an1n04x5 FILLER_246_1028 ();
 b15zdnd00an1n02x5 FILLER_246_1032 ();
 b15zdnd11an1n08x5 FILLER_246_1039 ();
 b15zdnd00an1n01x5 FILLER_246_1047 ();
 b15zdnd11an1n04x5 FILLER_246_1055 ();
 b15zdnd00an1n02x5 FILLER_246_1059 ();
 b15zdnd00an1n01x5 FILLER_246_1061 ();
 b15zdnd11an1n04x5 FILLER_246_1072 ();
 b15zdnd11an1n04x5 FILLER_246_1080 ();
 b15zdnd00an1n02x5 FILLER_246_1084 ();
 b15zdnd00an1n01x5 FILLER_246_1086 ();
 b15zdnd11an1n08x5 FILLER_246_1100 ();
 b15zdnd11an1n04x5 FILLER_246_1108 ();
 b15zdnd00an1n02x5 FILLER_246_1112 ();
 b15zdnd11an1n08x5 FILLER_246_1118 ();
 b15zdnd00an1n02x5 FILLER_246_1126 ();
 b15zdnd11an1n16x5 FILLER_246_1133 ();
 b15zdnd11an1n08x5 FILLER_246_1149 ();
 b15zdnd11an1n04x5 FILLER_246_1157 ();
 b15zdnd00an1n01x5 FILLER_246_1161 ();
 b15zdnd11an1n16x5 FILLER_246_1169 ();
 b15zdnd11an1n16x5 FILLER_246_1192 ();
 b15zdnd11an1n08x5 FILLER_246_1208 ();
 b15zdnd11an1n16x5 FILLER_246_1225 ();
 b15zdnd11an1n08x5 FILLER_246_1241 ();
 b15zdnd11an1n04x5 FILLER_246_1249 ();
 b15zdnd00an1n02x5 FILLER_246_1253 ();
 b15zdnd00an1n01x5 FILLER_246_1255 ();
 b15zdnd11an1n08x5 FILLER_246_1270 ();
 b15zdnd11an1n04x5 FILLER_246_1278 ();
 b15zdnd00an1n01x5 FILLER_246_1282 ();
 b15zdnd11an1n32x5 FILLER_246_1291 ();
 b15zdnd11an1n08x5 FILLER_246_1323 ();
 b15zdnd11an1n04x5 FILLER_246_1331 ();
 b15zdnd00an1n02x5 FILLER_246_1335 ();
 b15zdnd00an1n01x5 FILLER_246_1337 ();
 b15zdnd11an1n04x5 FILLER_246_1370 ();
 b15zdnd11an1n04x5 FILLER_246_1384 ();
 b15zdnd11an1n04x5 FILLER_246_1414 ();
 b15zdnd11an1n04x5 FILLER_246_1444 ();
 b15zdnd00an1n02x5 FILLER_246_1448 ();
 b15zdnd00an1n01x5 FILLER_246_1450 ();
 b15zdnd11an1n32x5 FILLER_246_1477 ();
 b15zdnd11an1n16x5 FILLER_246_1509 ();
 b15zdnd11an1n04x5 FILLER_246_1525 ();
 b15zdnd11an1n32x5 FILLER_246_1547 ();
 b15zdnd11an1n08x5 FILLER_246_1579 ();
 b15zdnd11an1n04x5 FILLER_246_1587 ();
 b15zdnd11an1n04x5 FILLER_246_1596 ();
 b15zdnd11an1n16x5 FILLER_246_1613 ();
 b15zdnd11an1n08x5 FILLER_246_1629 ();
 b15zdnd11an1n16x5 FILLER_246_1642 ();
 b15zdnd11an1n08x5 FILLER_246_1658 ();
 b15zdnd11an1n04x5 FILLER_246_1666 ();
 b15zdnd00an1n02x5 FILLER_246_1670 ();
 b15zdnd11an1n32x5 FILLER_246_1684 ();
 b15zdnd11an1n16x5 FILLER_246_1716 ();
 b15zdnd11an1n04x5 FILLER_246_1732 ();
 b15zdnd00an1n01x5 FILLER_246_1736 ();
 b15zdnd11an1n04x5 FILLER_246_1742 ();
 b15zdnd11an1n16x5 FILLER_246_1758 ();
 b15zdnd11an1n08x5 FILLER_246_1774 ();
 b15zdnd00an1n02x5 FILLER_246_1782 ();
 b15zdnd11an1n08x5 FILLER_246_1790 ();
 b15zdnd11an1n32x5 FILLER_246_1830 ();
 b15zdnd11an1n16x5 FILLER_246_1862 ();
 b15zdnd11an1n08x5 FILLER_246_1878 ();
 b15zdnd00an1n01x5 FILLER_246_1886 ();
 b15zdnd11an1n08x5 FILLER_246_1901 ();
 b15zdnd11an1n04x5 FILLER_246_1909 ();
 b15zdnd00an1n02x5 FILLER_246_1913 ();
 b15zdnd11an1n04x5 FILLER_246_1921 ();
 b15zdnd11an1n32x5 FILLER_246_1932 ();
 b15zdnd11an1n16x5 FILLER_246_1964 ();
 b15zdnd11an1n04x5 FILLER_246_1980 ();
 b15zdnd00an1n01x5 FILLER_246_1984 ();
 b15zdnd11an1n32x5 FILLER_246_2001 ();
 b15zdnd11an1n16x5 FILLER_246_2033 ();
 b15zdnd11an1n08x5 FILLER_246_2049 ();
 b15zdnd00an1n02x5 FILLER_246_2057 ();
 b15zdnd00an1n01x5 FILLER_246_2059 ();
 b15zdnd11an1n08x5 FILLER_246_2069 ();
 b15zdnd11an1n32x5 FILLER_246_2083 ();
 b15zdnd11an1n08x5 FILLER_246_2115 ();
 b15zdnd00an1n02x5 FILLER_246_2123 ();
 b15zdnd11an1n08x5 FILLER_246_2141 ();
 b15zdnd11an1n04x5 FILLER_246_2149 ();
 b15zdnd00an1n01x5 FILLER_246_2153 ();
 b15zdnd11an1n08x5 FILLER_246_2162 ();
 b15zdnd11an1n04x5 FILLER_246_2170 ();
 b15zdnd00an1n02x5 FILLER_246_2174 ();
 b15zdnd11an1n32x5 FILLER_246_2191 ();
 b15zdnd11an1n32x5 FILLER_246_2233 ();
 b15zdnd11an1n08x5 FILLER_246_2265 ();
 b15zdnd00an1n02x5 FILLER_246_2273 ();
 b15zdnd00an1n01x5 FILLER_246_2275 ();
 b15zdnd11an1n64x5 FILLER_247_0 ();
 b15zdnd11an1n32x5 FILLER_247_64 ();
 b15zdnd11an1n08x5 FILLER_247_96 ();
 b15zdnd11an1n04x5 FILLER_247_104 ();
 b15zdnd00an1n02x5 FILLER_247_108 ();
 b15zdnd11an1n16x5 FILLER_247_116 ();
 b15zdnd11an1n64x5 FILLER_247_138 ();
 b15zdnd11an1n32x5 FILLER_247_202 ();
 b15zdnd11an1n16x5 FILLER_247_234 ();
 b15zdnd11an1n04x5 FILLER_247_250 ();
 b15zdnd11an1n32x5 FILLER_247_261 ();
 b15zdnd11an1n16x5 FILLER_247_300 ();
 b15zdnd11an1n16x5 FILLER_247_321 ();
 b15zdnd11an1n04x5 FILLER_247_337 ();
 b15zdnd00an1n02x5 FILLER_247_341 ();
 b15zdnd00an1n01x5 FILLER_247_343 ();
 b15zdnd11an1n04x5 FILLER_247_353 ();
 b15zdnd11an1n32x5 FILLER_247_370 ();
 b15zdnd11an1n16x5 FILLER_247_402 ();
 b15zdnd11an1n08x5 FILLER_247_418 ();
 b15zdnd11an1n04x5 FILLER_247_426 ();
 b15zdnd00an1n02x5 FILLER_247_430 ();
 b15zdnd11an1n08x5 FILLER_247_448 ();
 b15zdnd11an1n04x5 FILLER_247_456 ();
 b15zdnd11an1n04x5 FILLER_247_470 ();
 b15zdnd00an1n01x5 FILLER_247_474 ();
 b15zdnd11an1n16x5 FILLER_247_486 ();
 b15zdnd11an1n04x5 FILLER_247_502 ();
 b15zdnd00an1n02x5 FILLER_247_506 ();
 b15zdnd00an1n01x5 FILLER_247_508 ();
 b15zdnd11an1n04x5 FILLER_247_518 ();
 b15zdnd00an1n02x5 FILLER_247_522 ();
 b15zdnd11an1n04x5 FILLER_247_529 ();
 b15zdnd11an1n16x5 FILLER_247_538 ();
 b15zdnd11an1n08x5 FILLER_247_559 ();
 b15zdnd11an1n04x5 FILLER_247_567 ();
 b15zdnd11an1n08x5 FILLER_247_597 ();
 b15zdnd00an1n02x5 FILLER_247_605 ();
 b15zdnd11an1n16x5 FILLER_247_612 ();
 b15zdnd11an1n08x5 FILLER_247_628 ();
 b15zdnd11an1n04x5 FILLER_247_636 ();
 b15zdnd11an1n08x5 FILLER_247_644 ();
 b15zdnd11an1n04x5 FILLER_247_652 ();
 b15zdnd00an1n01x5 FILLER_247_656 ();
 b15zdnd11an1n32x5 FILLER_247_662 ();
 b15zdnd11an1n16x5 FILLER_247_694 ();
 b15zdnd11an1n04x5 FILLER_247_720 ();
 b15zdnd11an1n08x5 FILLER_247_738 ();
 b15zdnd00an1n01x5 FILLER_247_746 ();
 b15zdnd11an1n04x5 FILLER_247_764 ();
 b15zdnd11an1n64x5 FILLER_247_784 ();
 b15zdnd11an1n16x5 FILLER_247_848 ();
 b15zdnd11an1n16x5 FILLER_247_884 ();
 b15zdnd11an1n32x5 FILLER_247_920 ();
 b15zdnd00an1n02x5 FILLER_247_952 ();
 b15zdnd00an1n01x5 FILLER_247_954 ();
 b15zdnd11an1n04x5 FILLER_247_971 ();
 b15zdnd00an1n02x5 FILLER_247_975 ();
 b15zdnd00an1n01x5 FILLER_247_977 ();
 b15zdnd11an1n08x5 FILLER_247_988 ();
 b15zdnd00an1n01x5 FILLER_247_996 ();
 b15zdnd11an1n32x5 FILLER_247_1021 ();
 b15zdnd11an1n08x5 FILLER_247_1053 ();
 b15zdnd00an1n02x5 FILLER_247_1061 ();
 b15zdnd11an1n04x5 FILLER_247_1074 ();
 b15zdnd11an1n08x5 FILLER_247_1098 ();
 b15zdnd11an1n04x5 FILLER_247_1106 ();
 b15zdnd00an1n02x5 FILLER_247_1110 ();
 b15zdnd11an1n08x5 FILLER_247_1118 ();
 b15zdnd00an1n02x5 FILLER_247_1126 ();
 b15zdnd11an1n04x5 FILLER_247_1140 ();
 b15zdnd11an1n64x5 FILLER_247_1151 ();
 b15zdnd11an1n16x5 FILLER_247_1215 ();
 b15zdnd00an1n02x5 FILLER_247_1231 ();
 b15zdnd00an1n01x5 FILLER_247_1233 ();
 b15zdnd11an1n08x5 FILLER_247_1254 ();
 b15zdnd00an1n02x5 FILLER_247_1262 ();
 b15zdnd11an1n08x5 FILLER_247_1271 ();
 b15zdnd11an1n04x5 FILLER_247_1279 ();
 b15zdnd11an1n64x5 FILLER_247_1290 ();
 b15zdnd11an1n16x5 FILLER_247_1354 ();
 b15zdnd11an1n04x5 FILLER_247_1370 ();
 b15zdnd00an1n01x5 FILLER_247_1374 ();
 b15zdnd11an1n64x5 FILLER_247_1401 ();
 b15zdnd11an1n64x5 FILLER_247_1465 ();
 b15zdnd11an1n16x5 FILLER_247_1529 ();
 b15zdnd11an1n08x5 FILLER_247_1545 ();
 b15zdnd11an1n04x5 FILLER_247_1553 ();
 b15zdnd11an1n16x5 FILLER_247_1572 ();
 b15zdnd11an1n04x5 FILLER_247_1588 ();
 b15zdnd00an1n01x5 FILLER_247_1592 ();
 b15zdnd11an1n64x5 FILLER_247_1611 ();
 b15zdnd11an1n16x5 FILLER_247_1675 ();
 b15zdnd00an1n02x5 FILLER_247_1691 ();
 b15zdnd11an1n04x5 FILLER_247_1699 ();
 b15zdnd11an1n16x5 FILLER_247_1715 ();
 b15zdnd00an1n02x5 FILLER_247_1731 ();
 b15zdnd11an1n16x5 FILLER_247_1739 ();
 b15zdnd11an1n04x5 FILLER_247_1755 ();
 b15zdnd11an1n04x5 FILLER_247_1765 ();
 b15zdnd11an1n08x5 FILLER_247_1785 ();
 b15zdnd11an1n04x5 FILLER_247_1793 ();
 b15zdnd00an1n02x5 FILLER_247_1797 ();
 b15zdnd11an1n64x5 FILLER_247_1815 ();
 b15zdnd11an1n04x5 FILLER_247_1879 ();
 b15zdnd00an1n02x5 FILLER_247_1883 ();
 b15zdnd11an1n04x5 FILLER_247_1903 ();
 b15zdnd11an1n08x5 FILLER_247_1913 ();
 b15zdnd11an1n04x5 FILLER_247_1937 ();
 b15zdnd11an1n32x5 FILLER_247_1946 ();
 b15zdnd11an1n16x5 FILLER_247_1978 ();
 b15zdnd11an1n08x5 FILLER_247_1994 ();
 b15zdnd11an1n04x5 FILLER_247_2002 ();
 b15zdnd00an1n02x5 FILLER_247_2006 ();
 b15zdnd00an1n01x5 FILLER_247_2008 ();
 b15zdnd11an1n16x5 FILLER_247_2018 ();
 b15zdnd11an1n08x5 FILLER_247_2034 ();
 b15zdnd11an1n04x5 FILLER_247_2042 ();
 b15zdnd00an1n02x5 FILLER_247_2046 ();
 b15zdnd11an1n32x5 FILLER_247_2055 ();
 b15zdnd11an1n16x5 FILLER_247_2087 ();
 b15zdnd11an1n08x5 FILLER_247_2103 ();
 b15zdnd11an1n04x5 FILLER_247_2111 ();
 b15zdnd11an1n64x5 FILLER_247_2128 ();
 b15zdnd11an1n64x5 FILLER_247_2192 ();
 b15zdnd11an1n16x5 FILLER_247_2256 ();
 b15zdnd11an1n08x5 FILLER_247_2272 ();
 b15zdnd11an1n04x5 FILLER_247_2280 ();
 b15zdnd11an1n64x5 FILLER_248_8 ();
 b15zdnd11an1n16x5 FILLER_248_72 ();
 b15zdnd11an1n08x5 FILLER_248_88 ();
 b15zdnd11an1n04x5 FILLER_248_96 ();
 b15zdnd00an1n02x5 FILLER_248_100 ();
 b15zdnd00an1n01x5 FILLER_248_102 ();
 b15zdnd11an1n04x5 FILLER_248_125 ();
 b15zdnd11an1n16x5 FILLER_248_139 ();
 b15zdnd11an1n04x5 FILLER_248_155 ();
 b15zdnd11an1n16x5 FILLER_248_164 ();
 b15zdnd11an1n16x5 FILLER_248_199 ();
 b15zdnd11an1n32x5 FILLER_248_230 ();
 b15zdnd11an1n08x5 FILLER_248_262 ();
 b15zdnd00an1n02x5 FILLER_248_270 ();
 b15zdnd11an1n16x5 FILLER_248_276 ();
 b15zdnd11an1n04x5 FILLER_248_292 ();
 b15zdnd11an1n08x5 FILLER_248_306 ();
 b15zdnd00an1n01x5 FILLER_248_314 ();
 b15zdnd11an1n64x5 FILLER_248_321 ();
 b15zdnd11an1n32x5 FILLER_248_385 ();
 b15zdnd11an1n08x5 FILLER_248_417 ();
 b15zdnd11an1n04x5 FILLER_248_425 ();
 b15zdnd11an1n04x5 FILLER_248_449 ();
 b15zdnd11an1n16x5 FILLER_248_457 ();
 b15zdnd11an1n08x5 FILLER_248_473 ();
 b15zdnd11an1n04x5 FILLER_248_481 ();
 b15zdnd00an1n01x5 FILLER_248_485 ();
 b15zdnd11an1n16x5 FILLER_248_498 ();
 b15zdnd11an1n04x5 FILLER_248_519 ();
 b15zdnd00an1n02x5 FILLER_248_523 ();
 b15zdnd11an1n08x5 FILLER_248_530 ();
 b15zdnd11an1n64x5 FILLER_248_549 ();
 b15zdnd11an1n64x5 FILLER_248_613 ();
 b15zdnd11an1n32x5 FILLER_248_677 ();
 b15zdnd11an1n08x5 FILLER_248_709 ();
 b15zdnd00an1n01x5 FILLER_248_717 ();
 b15zdnd11an1n04x5 FILLER_248_726 ();
 b15zdnd11an1n16x5 FILLER_248_739 ();
 b15zdnd11an1n04x5 FILLER_248_755 ();
 b15zdnd00an1n02x5 FILLER_248_759 ();
 b15zdnd00an1n01x5 FILLER_248_761 ();
 b15zdnd11an1n04x5 FILLER_248_769 ();
 b15zdnd11an1n04x5 FILLER_248_799 ();
 b15zdnd00an1n01x5 FILLER_248_803 ();
 b15zdnd11an1n32x5 FILLER_248_822 ();
 b15zdnd11an1n16x5 FILLER_248_854 ();
 b15zdnd00an1n02x5 FILLER_248_870 ();
 b15zdnd00an1n01x5 FILLER_248_872 ();
 b15zdnd11an1n32x5 FILLER_248_876 ();
 b15zdnd00an1n01x5 FILLER_248_908 ();
 b15zdnd11an1n64x5 FILLER_248_913 ();
 b15zdnd00an1n02x5 FILLER_248_977 ();
 b15zdnd11an1n64x5 FILLER_248_985 ();
 b15zdnd11an1n64x5 FILLER_248_1049 ();
 b15zdnd11an1n16x5 FILLER_248_1113 ();
 b15zdnd00an1n02x5 FILLER_248_1129 ();
 b15zdnd11an1n04x5 FILLER_248_1144 ();
 b15zdnd11an1n04x5 FILLER_248_1158 ();
 b15zdnd00an1n01x5 FILLER_248_1162 ();
 b15zdnd11an1n64x5 FILLER_248_1169 ();
 b15zdnd11an1n64x5 FILLER_248_1233 ();
 b15zdnd00an1n02x5 FILLER_248_1297 ();
 b15zdnd11an1n32x5 FILLER_248_1305 ();
 b15zdnd11an1n08x5 FILLER_248_1337 ();
 b15zdnd11an1n08x5 FILLER_248_1349 ();
 b15zdnd11an1n04x5 FILLER_248_1357 ();
 b15zdnd00an1n02x5 FILLER_248_1361 ();
 b15zdnd00an1n01x5 FILLER_248_1363 ();
 b15zdnd11an1n04x5 FILLER_248_1390 ();
 b15zdnd11an1n32x5 FILLER_248_1420 ();
 b15zdnd11an1n04x5 FILLER_248_1452 ();
 b15zdnd00an1n02x5 FILLER_248_1456 ();
 b15zdnd11an1n04x5 FILLER_248_1463 ();
 b15zdnd00an1n01x5 FILLER_248_1467 ();
 b15zdnd11an1n04x5 FILLER_248_1473 ();
 b15zdnd11an1n08x5 FILLER_248_1481 ();
 b15zdnd11an1n04x5 FILLER_248_1489 ();
 b15zdnd11an1n16x5 FILLER_248_1505 ();
 b15zdnd00an1n02x5 FILLER_248_1521 ();
 b15zdnd11an1n16x5 FILLER_248_1539 ();
 b15zdnd11an1n04x5 FILLER_248_1555 ();
 b15zdnd00an1n01x5 FILLER_248_1559 ();
 b15zdnd11an1n04x5 FILLER_248_1572 ();
 b15zdnd00an1n02x5 FILLER_248_1576 ();
 b15zdnd00an1n01x5 FILLER_248_1578 ();
 b15zdnd11an1n64x5 FILLER_248_1589 ();
 b15zdnd11an1n64x5 FILLER_248_1653 ();
 b15zdnd11an1n16x5 FILLER_248_1717 ();
 b15zdnd11an1n04x5 FILLER_248_1733 ();
 b15zdnd00an1n02x5 FILLER_248_1737 ();
 b15zdnd11an1n16x5 FILLER_248_1744 ();
 b15zdnd00an1n02x5 FILLER_248_1760 ();
 b15zdnd11an1n16x5 FILLER_248_1778 ();
 b15zdnd11an1n08x5 FILLER_248_1794 ();
 b15zdnd00an1n01x5 FILLER_248_1802 ();
 b15zdnd11an1n64x5 FILLER_248_1819 ();
 b15zdnd11an1n64x5 FILLER_248_1893 ();
 b15zdnd11an1n32x5 FILLER_248_1957 ();
 b15zdnd11an1n16x5 FILLER_248_1989 ();
 b15zdnd11an1n04x5 FILLER_248_2005 ();
 b15zdnd00an1n01x5 FILLER_248_2009 ();
 b15zdnd11an1n64x5 FILLER_248_2016 ();
 b15zdnd11an1n64x5 FILLER_248_2080 ();
 b15zdnd11an1n08x5 FILLER_248_2144 ();
 b15zdnd00an1n02x5 FILLER_248_2152 ();
 b15zdnd11an1n32x5 FILLER_248_2162 ();
 b15zdnd11an1n16x5 FILLER_248_2194 ();
 b15zdnd11an1n08x5 FILLER_248_2210 ();
 b15zdnd00an1n02x5 FILLER_248_2218 ();
 b15zdnd11an1n16x5 FILLER_248_2230 ();
 b15zdnd11an1n08x5 FILLER_248_2246 ();
 b15zdnd00an1n02x5 FILLER_248_2274 ();
 b15zdnd11an1n32x5 FILLER_249_0 ();
 b15zdnd11an1n16x5 FILLER_249_32 ();
 b15zdnd00an1n01x5 FILLER_249_48 ();
 b15zdnd11an1n32x5 FILLER_249_55 ();
 b15zdnd11an1n16x5 FILLER_249_87 ();
 b15zdnd11an1n04x5 FILLER_249_103 ();
 b15zdnd00an1n02x5 FILLER_249_107 ();
 b15zdnd11an1n16x5 FILLER_249_118 ();
 b15zdnd11an1n08x5 FILLER_249_134 ();
 b15zdnd11an1n08x5 FILLER_249_151 ();
 b15zdnd11an1n04x5 FILLER_249_159 ();
 b15zdnd11an1n04x5 FILLER_249_178 ();
 b15zdnd11an1n04x5 FILLER_249_188 ();
 b15zdnd00an1n01x5 FILLER_249_192 ();
 b15zdnd11an1n08x5 FILLER_249_219 ();
 b15zdnd11an1n04x5 FILLER_249_227 ();
 b15zdnd11an1n32x5 FILLER_249_238 ();
 b15zdnd00an1n01x5 FILLER_249_270 ();
 b15zdnd11an1n08x5 FILLER_249_278 ();
 b15zdnd11an1n04x5 FILLER_249_286 ();
 b15zdnd11an1n64x5 FILLER_249_296 ();
 b15zdnd11an1n64x5 FILLER_249_360 ();
 b15zdnd11an1n32x5 FILLER_249_424 ();
 b15zdnd00an1n02x5 FILLER_249_456 ();
 b15zdnd11an1n64x5 FILLER_249_469 ();
 b15zdnd11an1n04x5 FILLER_249_533 ();
 b15zdnd00an1n02x5 FILLER_249_537 ();
 b15zdnd00an1n01x5 FILLER_249_539 ();
 b15zdnd11an1n32x5 FILLER_249_559 ();
 b15zdnd11an1n16x5 FILLER_249_591 ();
 b15zdnd11an1n08x5 FILLER_249_607 ();
 b15zdnd11an1n04x5 FILLER_249_615 ();
 b15zdnd00an1n01x5 FILLER_249_619 ();
 b15zdnd11an1n16x5 FILLER_249_638 ();
 b15zdnd11an1n08x5 FILLER_249_654 ();
 b15zdnd00an1n01x5 FILLER_249_662 ();
 b15zdnd11an1n04x5 FILLER_249_667 ();
 b15zdnd11an1n64x5 FILLER_249_675 ();
 b15zdnd11an1n32x5 FILLER_249_739 ();
 b15zdnd11an1n08x5 FILLER_249_771 ();
 b15zdnd00an1n01x5 FILLER_249_779 ();
 b15zdnd11an1n16x5 FILLER_249_793 ();
 b15zdnd11an1n04x5 FILLER_249_809 ();
 b15zdnd00an1n01x5 FILLER_249_813 ();
 b15zdnd11an1n64x5 FILLER_249_821 ();
 b15zdnd11an1n64x5 FILLER_249_885 ();
 b15zdnd11an1n64x5 FILLER_249_949 ();
 b15zdnd11an1n32x5 FILLER_249_1013 ();
 b15zdnd11an1n08x5 FILLER_249_1045 ();
 b15zdnd00an1n02x5 FILLER_249_1053 ();
 b15zdnd11an1n64x5 FILLER_249_1071 ();
 b15zdnd11an1n64x5 FILLER_249_1135 ();
 b15zdnd11an1n64x5 FILLER_249_1199 ();
 b15zdnd11an1n32x5 FILLER_249_1263 ();
 b15zdnd11an1n08x5 FILLER_249_1295 ();
 b15zdnd00an1n02x5 FILLER_249_1303 ();
 b15zdnd00an1n01x5 FILLER_249_1305 ();
 b15zdnd11an1n16x5 FILLER_249_1314 ();
 b15zdnd11an1n04x5 FILLER_249_1330 ();
 b15zdnd00an1n01x5 FILLER_249_1334 ();
 b15zdnd11an1n32x5 FILLER_249_1342 ();
 b15zdnd11an1n08x5 FILLER_249_1374 ();
 b15zdnd00an1n02x5 FILLER_249_1382 ();
 b15zdnd11an1n32x5 FILLER_249_1410 ();
 b15zdnd11an1n16x5 FILLER_249_1442 ();
 b15zdnd00an1n02x5 FILLER_249_1458 ();
 b15zdnd11an1n04x5 FILLER_249_1472 ();
 b15zdnd11an1n04x5 FILLER_249_1489 ();
 b15zdnd11an1n32x5 FILLER_249_1507 ();
 b15zdnd11an1n16x5 FILLER_249_1539 ();
 b15zdnd11an1n08x5 FILLER_249_1555 ();
 b15zdnd11an1n04x5 FILLER_249_1563 ();
 b15zdnd11an1n32x5 FILLER_249_1587 ();
 b15zdnd00an1n01x5 FILLER_249_1619 ();
 b15zdnd11an1n16x5 FILLER_249_1626 ();
 b15zdnd11an1n08x5 FILLER_249_1642 ();
 b15zdnd00an1n02x5 FILLER_249_1650 ();
 b15zdnd11an1n16x5 FILLER_249_1663 ();
 b15zdnd00an1n01x5 FILLER_249_1679 ();
 b15zdnd11an1n04x5 FILLER_249_1685 ();
 b15zdnd11an1n32x5 FILLER_249_1703 ();
 b15zdnd11an1n16x5 FILLER_249_1735 ();
 b15zdnd11an1n08x5 FILLER_249_1751 ();
 b15zdnd11an1n04x5 FILLER_249_1759 ();
 b15zdnd00an1n02x5 FILLER_249_1763 ();
 b15zdnd11an1n64x5 FILLER_249_1778 ();
 b15zdnd11an1n64x5 FILLER_249_1842 ();
 b15zdnd11an1n64x5 FILLER_249_1906 ();
 b15zdnd11an1n32x5 FILLER_249_1970 ();
 b15zdnd11an1n08x5 FILLER_249_2002 ();
 b15zdnd00an1n02x5 FILLER_249_2010 ();
 b15zdnd11an1n32x5 FILLER_249_2016 ();
 b15zdnd11an1n08x5 FILLER_249_2048 ();
 b15zdnd00an1n02x5 FILLER_249_2056 ();
 b15zdnd11an1n08x5 FILLER_249_2068 ();
 b15zdnd00an1n02x5 FILLER_249_2076 ();
 b15zdnd00an1n01x5 FILLER_249_2078 ();
 b15zdnd11an1n08x5 FILLER_249_2085 ();
 b15zdnd11an1n04x5 FILLER_249_2093 ();
 b15zdnd00an1n02x5 FILLER_249_2097 ();
 b15zdnd11an1n08x5 FILLER_249_2114 ();
 b15zdnd11an1n04x5 FILLER_249_2122 ();
 b15zdnd00an1n02x5 FILLER_249_2126 ();
 b15zdnd11an1n08x5 FILLER_249_2134 ();
 b15zdnd11an1n32x5 FILLER_249_2148 ();
 b15zdnd11an1n08x5 FILLER_249_2180 ();
 b15zdnd00an1n02x5 FILLER_249_2188 ();
 b15zdnd00an1n01x5 FILLER_249_2190 ();
 b15zdnd11an1n04x5 FILLER_249_2198 ();
 b15zdnd11an1n04x5 FILLER_249_2208 ();
 b15zdnd11an1n64x5 FILLER_249_2218 ();
 b15zdnd00an1n02x5 FILLER_249_2282 ();
 b15zdnd11an1n32x5 FILLER_250_8 ();
 b15zdnd11an1n08x5 FILLER_250_40 ();
 b15zdnd11an1n04x5 FILLER_250_48 ();
 b15zdnd00an1n02x5 FILLER_250_52 ();
 b15zdnd11an1n16x5 FILLER_250_66 ();
 b15zdnd11an1n64x5 FILLER_250_87 ();
 b15zdnd11an1n32x5 FILLER_250_151 ();
 b15zdnd00an1n02x5 FILLER_250_183 ();
 b15zdnd00an1n01x5 FILLER_250_185 ();
 b15zdnd11an1n32x5 FILLER_250_191 ();
 b15zdnd00an1n02x5 FILLER_250_223 ();
 b15zdnd11an1n64x5 FILLER_250_239 ();
 b15zdnd11an1n32x5 FILLER_250_303 ();
 b15zdnd11an1n08x5 FILLER_250_335 ();
 b15zdnd11an1n04x5 FILLER_250_343 ();
 b15zdnd00an1n02x5 FILLER_250_347 ();
 b15zdnd00an1n01x5 FILLER_250_349 ();
 b15zdnd11an1n04x5 FILLER_250_358 ();
 b15zdnd11an1n64x5 FILLER_250_368 ();
 b15zdnd11an1n64x5 FILLER_250_432 ();
 b15zdnd11an1n64x5 FILLER_250_496 ();
 b15zdnd11an1n08x5 FILLER_250_560 ();
 b15zdnd11an1n04x5 FILLER_250_568 ();
 b15zdnd00an1n02x5 FILLER_250_572 ();
 b15zdnd11an1n32x5 FILLER_250_583 ();
 b15zdnd11an1n08x5 FILLER_250_615 ();
 b15zdnd00an1n01x5 FILLER_250_623 ();
 b15zdnd11an1n32x5 FILLER_250_628 ();
 b15zdnd11an1n08x5 FILLER_250_660 ();
 b15zdnd00an1n02x5 FILLER_250_668 ();
 b15zdnd11an1n04x5 FILLER_250_679 ();
 b15zdnd11an1n04x5 FILLER_250_697 ();
 b15zdnd11an1n08x5 FILLER_250_710 ();
 b15zdnd11an1n64x5 FILLER_250_726 ();
 b15zdnd11an1n16x5 FILLER_250_790 ();
 b15zdnd11an1n04x5 FILLER_250_806 ();
 b15zdnd00an1n02x5 FILLER_250_810 ();
 b15zdnd11an1n08x5 FILLER_250_822 ();
 b15zdnd11an1n04x5 FILLER_250_830 ();
 b15zdnd00an1n02x5 FILLER_250_834 ();
 b15zdnd00an1n01x5 FILLER_250_836 ();
 b15zdnd11an1n64x5 FILLER_250_863 ();
 b15zdnd11an1n32x5 FILLER_250_927 ();
 b15zdnd11an1n16x5 FILLER_250_959 ();
 b15zdnd11an1n04x5 FILLER_250_975 ();
 b15zdnd00an1n02x5 FILLER_250_979 ();
 b15zdnd11an1n04x5 FILLER_250_994 ();
 b15zdnd11an1n32x5 FILLER_250_1011 ();
 b15zdnd11an1n16x5 FILLER_250_1043 ();
 b15zdnd00an1n01x5 FILLER_250_1059 ();
 b15zdnd11an1n16x5 FILLER_250_1070 ();
 b15zdnd11an1n08x5 FILLER_250_1086 ();
 b15zdnd11an1n04x5 FILLER_250_1094 ();
 b15zdnd00an1n01x5 FILLER_250_1098 ();
 b15zdnd11an1n64x5 FILLER_250_1112 ();
 b15zdnd11an1n08x5 FILLER_250_1176 ();
 b15zdnd11an1n04x5 FILLER_250_1184 ();
 b15zdnd11an1n32x5 FILLER_250_1192 ();
 b15zdnd11an1n04x5 FILLER_250_1224 ();
 b15zdnd11an1n16x5 FILLER_250_1235 ();
 b15zdnd11an1n08x5 FILLER_250_1251 ();
 b15zdnd00an1n01x5 FILLER_250_1259 ();
 b15zdnd11an1n08x5 FILLER_250_1268 ();
 b15zdnd11an1n04x5 FILLER_250_1276 ();
 b15zdnd00an1n01x5 FILLER_250_1280 ();
 b15zdnd11an1n16x5 FILLER_250_1287 ();
 b15zdnd11an1n04x5 FILLER_250_1303 ();
 b15zdnd11an1n16x5 FILLER_250_1319 ();
 b15zdnd11an1n04x5 FILLER_250_1335 ();
 b15zdnd11an1n04x5 FILLER_250_1343 ();
 b15zdnd11an1n16x5 FILLER_250_1353 ();
 b15zdnd00an1n02x5 FILLER_250_1369 ();
 b15zdnd11an1n04x5 FILLER_250_1376 ();
 b15zdnd11an1n64x5 FILLER_250_1384 ();
 b15zdnd11an1n64x5 FILLER_250_1448 ();
 b15zdnd11an1n08x5 FILLER_250_1512 ();
 b15zdnd11an1n04x5 FILLER_250_1520 ();
 b15zdnd00an1n02x5 FILLER_250_1524 ();
 b15zdnd11an1n32x5 FILLER_250_1543 ();
 b15zdnd00an1n01x5 FILLER_250_1575 ();
 b15zdnd11an1n32x5 FILLER_250_1580 ();
 b15zdnd11an1n04x5 FILLER_250_1612 ();
 b15zdnd11an1n32x5 FILLER_250_1621 ();
 b15zdnd11an1n08x5 FILLER_250_1667 ();
 b15zdnd11an1n04x5 FILLER_250_1675 ();
 b15zdnd00an1n02x5 FILLER_250_1679 ();
 b15zdnd11an1n04x5 FILLER_250_1686 ();
 b15zdnd11an1n16x5 FILLER_250_1711 ();
 b15zdnd11an1n08x5 FILLER_250_1727 ();
 b15zdnd00an1n02x5 FILLER_250_1735 ();
 b15zdnd11an1n64x5 FILLER_250_1746 ();
 b15zdnd11an1n32x5 FILLER_250_1826 ();
 b15zdnd11an1n16x5 FILLER_250_1858 ();
 b15zdnd11an1n04x5 FILLER_250_1874 ();
 b15zdnd00an1n02x5 FILLER_250_1878 ();
 b15zdnd11an1n04x5 FILLER_250_1889 ();
 b15zdnd11an1n64x5 FILLER_250_1897 ();
 b15zdnd11an1n16x5 FILLER_250_1961 ();
 b15zdnd11an1n04x5 FILLER_250_1990 ();
 b15zdnd11an1n08x5 FILLER_250_2003 ();
 b15zdnd00an1n01x5 FILLER_250_2011 ();
 b15zdnd11an1n32x5 FILLER_250_2025 ();
 b15zdnd11an1n08x5 FILLER_250_2057 ();
 b15zdnd11an1n08x5 FILLER_250_2086 ();
 b15zdnd00an1n02x5 FILLER_250_2094 ();
 b15zdnd00an1n01x5 FILLER_250_2096 ();
 b15zdnd11an1n16x5 FILLER_250_2103 ();
 b15zdnd11an1n08x5 FILLER_250_2119 ();
 b15zdnd00an1n01x5 FILLER_250_2127 ();
 b15zdnd11an1n08x5 FILLER_250_2140 ();
 b15zdnd11an1n04x5 FILLER_250_2148 ();
 b15zdnd00an1n02x5 FILLER_250_2152 ();
 b15zdnd11an1n16x5 FILLER_250_2162 ();
 b15zdnd11an1n08x5 FILLER_250_2178 ();
 b15zdnd00an1n02x5 FILLER_250_2186 ();
 b15zdnd00an1n01x5 FILLER_250_2188 ();
 b15zdnd11an1n04x5 FILLER_250_2199 ();
 b15zdnd00an1n01x5 FILLER_250_2203 ();
 b15zdnd11an1n04x5 FILLER_250_2210 ();
 b15zdnd11an1n32x5 FILLER_250_2222 ();
 b15zdnd11an1n16x5 FILLER_250_2254 ();
 b15zdnd11an1n04x5 FILLER_250_2270 ();
 b15zdnd00an1n02x5 FILLER_250_2274 ();
 b15zdnd11an1n32x5 FILLER_251_0 ();
 b15zdnd11an1n04x5 FILLER_251_32 ();
 b15zdnd00an1n02x5 FILLER_251_36 ();
 b15zdnd11an1n04x5 FILLER_251_42 ();
 b15zdnd11an1n04x5 FILLER_251_53 ();
 b15zdnd11an1n08x5 FILLER_251_63 ();
 b15zdnd00an1n02x5 FILLER_251_71 ();
 b15zdnd11an1n64x5 FILLER_251_82 ();
 b15zdnd11an1n08x5 FILLER_251_146 ();
 b15zdnd11an1n04x5 FILLER_251_154 ();
 b15zdnd00an1n02x5 FILLER_251_158 ();
 b15zdnd00an1n01x5 FILLER_251_160 ();
 b15zdnd11an1n64x5 FILLER_251_177 ();
 b15zdnd11an1n32x5 FILLER_251_241 ();
 b15zdnd11an1n64x5 FILLER_251_279 ();
 b15zdnd11an1n64x5 FILLER_251_343 ();
 b15zdnd11an1n08x5 FILLER_251_407 ();
 b15zdnd11an1n04x5 FILLER_251_415 ();
 b15zdnd00an1n02x5 FILLER_251_419 ();
 b15zdnd11an1n04x5 FILLER_251_424 ();
 b15zdnd11an1n32x5 FILLER_251_433 ();
 b15zdnd11an1n16x5 FILLER_251_465 ();
 b15zdnd11an1n04x5 FILLER_251_481 ();
 b15zdnd00an1n02x5 FILLER_251_485 ();
 b15zdnd11an1n16x5 FILLER_251_491 ();
 b15zdnd11an1n04x5 FILLER_251_507 ();
 b15zdnd00an1n01x5 FILLER_251_511 ();
 b15zdnd11an1n04x5 FILLER_251_522 ();
 b15zdnd11an1n16x5 FILLER_251_541 ();
 b15zdnd11an1n04x5 FILLER_251_557 ();
 b15zdnd11an1n32x5 FILLER_251_567 ();
 b15zdnd11an1n16x5 FILLER_251_599 ();
 b15zdnd11an1n08x5 FILLER_251_615 ();
 b15zdnd00an1n01x5 FILLER_251_623 ();
 b15zdnd11an1n64x5 FILLER_251_630 ();
 b15zdnd11an1n08x5 FILLER_251_694 ();
 b15zdnd11an1n08x5 FILLER_251_718 ();
 b15zdnd00an1n02x5 FILLER_251_726 ();
 b15zdnd11an1n04x5 FILLER_251_740 ();
 b15zdnd00an1n02x5 FILLER_251_744 ();
 b15zdnd00an1n01x5 FILLER_251_746 ();
 b15zdnd11an1n16x5 FILLER_251_753 ();
 b15zdnd11an1n04x5 FILLER_251_782 ();
 b15zdnd00an1n01x5 FILLER_251_786 ();
 b15zdnd11an1n08x5 FILLER_251_799 ();
 b15zdnd00an1n01x5 FILLER_251_807 ();
 b15zdnd11an1n32x5 FILLER_251_815 ();
 b15zdnd11an1n08x5 FILLER_251_847 ();
 b15zdnd11an1n04x5 FILLER_251_855 ();
 b15zdnd11an1n64x5 FILLER_251_868 ();
 b15zdnd11an1n16x5 FILLER_251_932 ();
 b15zdnd11an1n64x5 FILLER_251_979 ();
 b15zdnd11an1n16x5 FILLER_251_1043 ();
 b15zdnd11an1n08x5 FILLER_251_1059 ();
 b15zdnd11an1n04x5 FILLER_251_1067 ();
 b15zdnd00an1n02x5 FILLER_251_1071 ();
 b15zdnd11an1n32x5 FILLER_251_1083 ();
 b15zdnd11an1n08x5 FILLER_251_1115 ();
 b15zdnd00an1n01x5 FILLER_251_1123 ();
 b15zdnd11an1n64x5 FILLER_251_1128 ();
 b15zdnd11an1n32x5 FILLER_251_1192 ();
 b15zdnd00an1n02x5 FILLER_251_1224 ();
 b15zdnd00an1n01x5 FILLER_251_1226 ();
 b15zdnd11an1n16x5 FILLER_251_1232 ();
 b15zdnd11an1n04x5 FILLER_251_1248 ();
 b15zdnd11an1n32x5 FILLER_251_1262 ();
 b15zdnd11an1n04x5 FILLER_251_1294 ();
 b15zdnd00an1n01x5 FILLER_251_1298 ();
 b15zdnd11an1n32x5 FILLER_251_1313 ();
 b15zdnd00an1n01x5 FILLER_251_1345 ();
 b15zdnd11an1n16x5 FILLER_251_1354 ();
 b15zdnd11an1n04x5 FILLER_251_1370 ();
 b15zdnd11an1n04x5 FILLER_251_1379 ();
 b15zdnd11an1n32x5 FILLER_251_1390 ();
 b15zdnd11an1n08x5 FILLER_251_1422 ();
 b15zdnd11an1n04x5 FILLER_251_1430 ();
 b15zdnd00an1n02x5 FILLER_251_1434 ();
 b15zdnd00an1n01x5 FILLER_251_1436 ();
 b15zdnd11an1n32x5 FILLER_251_1455 ();
 b15zdnd11an1n04x5 FILLER_251_1487 ();
 b15zdnd00an1n01x5 FILLER_251_1491 ();
 b15zdnd11an1n16x5 FILLER_251_1503 ();
 b15zdnd11an1n04x5 FILLER_251_1519 ();
 b15zdnd00an1n02x5 FILLER_251_1523 ();
 b15zdnd00an1n01x5 FILLER_251_1525 ();
 b15zdnd11an1n04x5 FILLER_251_1531 ();
 b15zdnd00an1n02x5 FILLER_251_1535 ();
 b15zdnd00an1n01x5 FILLER_251_1537 ();
 b15zdnd11an1n04x5 FILLER_251_1543 ();
 b15zdnd11an1n32x5 FILLER_251_1553 ();
 b15zdnd11an1n16x5 FILLER_251_1585 ();
 b15zdnd11an1n08x5 FILLER_251_1601 ();
 b15zdnd00an1n02x5 FILLER_251_1609 ();
 b15zdnd11an1n04x5 FILLER_251_1616 ();
 b15zdnd00an1n01x5 FILLER_251_1620 ();
 b15zdnd11an1n16x5 FILLER_251_1634 ();
 b15zdnd11an1n04x5 FILLER_251_1650 ();
 b15zdnd11an1n16x5 FILLER_251_1659 ();
 b15zdnd11an1n04x5 FILLER_251_1675 ();
 b15zdnd00an1n01x5 FILLER_251_1679 ();
 b15zdnd11an1n04x5 FILLER_251_1686 ();
 b15zdnd11an1n32x5 FILLER_251_1699 ();
 b15zdnd11an1n16x5 FILLER_251_1731 ();
 b15zdnd11an1n16x5 FILLER_251_1759 ();
 b15zdnd11an1n04x5 FILLER_251_1775 ();
 b15zdnd00an1n01x5 FILLER_251_1779 ();
 b15zdnd11an1n04x5 FILLER_251_1800 ();
 b15zdnd11an1n64x5 FILLER_251_1811 ();
 b15zdnd11an1n08x5 FILLER_251_1875 ();
 b15zdnd11an1n04x5 FILLER_251_1883 ();
 b15zdnd00an1n02x5 FILLER_251_1887 ();
 b15zdnd11an1n16x5 FILLER_251_1898 ();
 b15zdnd11an1n04x5 FILLER_251_1914 ();
 b15zdnd00an1n02x5 FILLER_251_1918 ();
 b15zdnd00an1n01x5 FILLER_251_1920 ();
 b15zdnd11an1n08x5 FILLER_251_1934 ();
 b15zdnd00an1n02x5 FILLER_251_1942 ();
 b15zdnd00an1n01x5 FILLER_251_1944 ();
 b15zdnd11an1n16x5 FILLER_251_1951 ();
 b15zdnd11an1n08x5 FILLER_251_1967 ();
 b15zdnd00an1n02x5 FILLER_251_1975 ();
 b15zdnd00an1n01x5 FILLER_251_1977 ();
 b15zdnd11an1n04x5 FILLER_251_1985 ();
 b15zdnd00an1n02x5 FILLER_251_1989 ();
 b15zdnd11an1n32x5 FILLER_251_2001 ();
 b15zdnd11an1n16x5 FILLER_251_2033 ();
 b15zdnd11an1n08x5 FILLER_251_2049 ();
 b15zdnd00an1n02x5 FILLER_251_2057 ();
 b15zdnd00an1n01x5 FILLER_251_2059 ();
 b15zdnd11an1n32x5 FILLER_251_2072 ();
 b15zdnd11an1n16x5 FILLER_251_2104 ();
 b15zdnd11an1n08x5 FILLER_251_2120 ();
 b15zdnd11an1n04x5 FILLER_251_2128 ();
 b15zdnd00an1n01x5 FILLER_251_2132 ();
 b15zdnd11an1n04x5 FILLER_251_2143 ();
 b15zdnd11an1n16x5 FILLER_251_2153 ();
 b15zdnd11an1n08x5 FILLER_251_2169 ();
 b15zdnd00an1n02x5 FILLER_251_2177 ();
 b15zdnd00an1n01x5 FILLER_251_2179 ();
 b15zdnd11an1n64x5 FILLER_251_2184 ();
 b15zdnd11an1n32x5 FILLER_251_2248 ();
 b15zdnd11an1n04x5 FILLER_251_2280 ();
 b15zdnd11an1n64x5 FILLER_252_8 ();
 b15zdnd11an1n64x5 FILLER_252_72 ();
 b15zdnd11an1n16x5 FILLER_252_136 ();
 b15zdnd11an1n04x5 FILLER_252_152 ();
 b15zdnd00an1n01x5 FILLER_252_156 ();
 b15zdnd11an1n16x5 FILLER_252_167 ();
 b15zdnd11an1n08x5 FILLER_252_183 ();
 b15zdnd11an1n04x5 FILLER_252_191 ();
 b15zdnd11an1n04x5 FILLER_252_201 ();
 b15zdnd11an1n16x5 FILLER_252_211 ();
 b15zdnd11an1n08x5 FILLER_252_227 ();
 b15zdnd00an1n01x5 FILLER_252_235 ();
 b15zdnd11an1n08x5 FILLER_252_243 ();
 b15zdnd00an1n02x5 FILLER_252_251 ();
 b15zdnd11an1n32x5 FILLER_252_259 ();
 b15zdnd11an1n16x5 FILLER_252_291 ();
 b15zdnd11an1n04x5 FILLER_252_307 ();
 b15zdnd00an1n01x5 FILLER_252_311 ();
 b15zdnd11an1n04x5 FILLER_252_318 ();
 b15zdnd11an1n64x5 FILLER_252_326 ();
 b15zdnd11an1n32x5 FILLER_252_390 ();
 b15zdnd00an1n02x5 FILLER_252_422 ();
 b15zdnd11an1n16x5 FILLER_252_433 ();
 b15zdnd00an1n02x5 FILLER_252_449 ();
 b15zdnd00an1n01x5 FILLER_252_451 ();
 b15zdnd11an1n16x5 FILLER_252_458 ();
 b15zdnd11an1n08x5 FILLER_252_474 ();
 b15zdnd11an1n04x5 FILLER_252_482 ();
 b15zdnd00an1n02x5 FILLER_252_486 ();
 b15zdnd11an1n08x5 FILLER_252_494 ();
 b15zdnd11an1n04x5 FILLER_252_502 ();
 b15zdnd00an1n01x5 FILLER_252_506 ();
 b15zdnd11an1n64x5 FILLER_252_517 ();
 b15zdnd11an1n04x5 FILLER_252_581 ();
 b15zdnd11an1n04x5 FILLER_252_591 ();
 b15zdnd11an1n04x5 FILLER_252_600 ();
 b15zdnd11an1n16x5 FILLER_252_610 ();
 b15zdnd11an1n08x5 FILLER_252_626 ();
 b15zdnd11an1n04x5 FILLER_252_634 ();
 b15zdnd00an1n02x5 FILLER_252_638 ();
 b15zdnd11an1n04x5 FILLER_252_646 ();
 b15zdnd11an1n08x5 FILLER_252_666 ();
 b15zdnd00an1n01x5 FILLER_252_674 ();
 b15zdnd11an1n04x5 FILLER_252_682 ();
 b15zdnd00an1n02x5 FILLER_252_686 ();
 b15zdnd00an1n01x5 FILLER_252_688 ();
 b15zdnd11an1n16x5 FILLER_252_699 ();
 b15zdnd00an1n02x5 FILLER_252_715 ();
 b15zdnd00an1n01x5 FILLER_252_717 ();
 b15zdnd11an1n16x5 FILLER_252_726 ();
 b15zdnd00an1n02x5 FILLER_252_742 ();
 b15zdnd11an1n04x5 FILLER_252_748 ();
 b15zdnd11an1n16x5 FILLER_252_764 ();
 b15zdnd00an1n02x5 FILLER_252_780 ();
 b15zdnd11an1n32x5 FILLER_252_787 ();
 b15zdnd11an1n16x5 FILLER_252_819 ();
 b15zdnd11an1n08x5 FILLER_252_835 ();
 b15zdnd11an1n04x5 FILLER_252_843 ();
 b15zdnd00an1n02x5 FILLER_252_847 ();
 b15zdnd11an1n64x5 FILLER_252_869 ();
 b15zdnd11an1n16x5 FILLER_252_933 ();
 b15zdnd11an1n08x5 FILLER_252_949 ();
 b15zdnd00an1n02x5 FILLER_252_957 ();
 b15zdnd11an1n16x5 FILLER_252_964 ();
 b15zdnd11an1n04x5 FILLER_252_980 ();
 b15zdnd00an1n01x5 FILLER_252_984 ();
 b15zdnd11an1n04x5 FILLER_252_996 ();
 b15zdnd11an1n08x5 FILLER_252_1007 ();
 b15zdnd11an1n04x5 FILLER_252_1032 ();
 b15zdnd11an1n16x5 FILLER_252_1048 ();
 b15zdnd11an1n04x5 FILLER_252_1064 ();
 b15zdnd00an1n02x5 FILLER_252_1068 ();
 b15zdnd11an1n64x5 FILLER_252_1081 ();
 b15zdnd11an1n08x5 FILLER_252_1154 ();
 b15zdnd00an1n01x5 FILLER_252_1162 ();
 b15zdnd11an1n16x5 FILLER_252_1170 ();
 b15zdnd11an1n04x5 FILLER_252_1190 ();
 b15zdnd00an1n01x5 FILLER_252_1194 ();
 b15zdnd11an1n32x5 FILLER_252_1202 ();
 b15zdnd11an1n16x5 FILLER_252_1234 ();
 b15zdnd11an1n04x5 FILLER_252_1250 ();
 b15zdnd00an1n01x5 FILLER_252_1254 ();
 b15zdnd11an1n16x5 FILLER_252_1268 ();
 b15zdnd11an1n04x5 FILLER_252_1284 ();
 b15zdnd00an1n02x5 FILLER_252_1288 ();
 b15zdnd11an1n64x5 FILLER_252_1308 ();
 b15zdnd11an1n64x5 FILLER_252_1372 ();
 b15zdnd11an1n64x5 FILLER_252_1436 ();
 b15zdnd11an1n32x5 FILLER_252_1500 ();
 b15zdnd11an1n08x5 FILLER_252_1532 ();
 b15zdnd00an1n01x5 FILLER_252_1540 ();
 b15zdnd11an1n04x5 FILLER_252_1553 ();
 b15zdnd00an1n01x5 FILLER_252_1557 ();
 b15zdnd11an1n32x5 FILLER_252_1563 ();
 b15zdnd11an1n16x5 FILLER_252_1595 ();
 b15zdnd11an1n08x5 FILLER_252_1611 ();
 b15zdnd11an1n04x5 FILLER_252_1619 ();
 b15zdnd11an1n32x5 FILLER_252_1628 ();
 b15zdnd11an1n16x5 FILLER_252_1660 ();
 b15zdnd11an1n08x5 FILLER_252_1676 ();
 b15zdnd11an1n04x5 FILLER_252_1684 ();
 b15zdnd00an1n02x5 FILLER_252_1688 ();
 b15zdnd00an1n01x5 FILLER_252_1690 ();
 b15zdnd11an1n04x5 FILLER_252_1702 ();
 b15zdnd11an1n16x5 FILLER_252_1711 ();
 b15zdnd11an1n08x5 FILLER_252_1727 ();
 b15zdnd11an1n08x5 FILLER_252_1747 ();
 b15zdnd11an1n04x5 FILLER_252_1761 ();
 b15zdnd11an1n04x5 FILLER_252_1779 ();
 b15zdnd00an1n01x5 FILLER_252_1783 ();
 b15zdnd11an1n04x5 FILLER_252_1795 ();
 b15zdnd00an1n01x5 FILLER_252_1799 ();
 b15zdnd11an1n16x5 FILLER_252_1806 ();
 b15zdnd00an1n02x5 FILLER_252_1822 ();
 b15zdnd00an1n01x5 FILLER_252_1824 ();
 b15zdnd11an1n32x5 FILLER_252_1841 ();
 b15zdnd11an1n08x5 FILLER_252_1873 ();
 b15zdnd11an1n04x5 FILLER_252_1881 ();
 b15zdnd00an1n02x5 FILLER_252_1885 ();
 b15zdnd00an1n01x5 FILLER_252_1887 ();
 b15zdnd11an1n16x5 FILLER_252_1903 ();
 b15zdnd00an1n02x5 FILLER_252_1919 ();
 b15zdnd00an1n01x5 FILLER_252_1921 ();
 b15zdnd11an1n16x5 FILLER_252_1927 ();
 b15zdnd11an1n04x5 FILLER_252_1943 ();
 b15zdnd00an1n01x5 FILLER_252_1947 ();
 b15zdnd11an1n32x5 FILLER_252_1954 ();
 b15zdnd11an1n08x5 FILLER_252_1986 ();
 b15zdnd11an1n32x5 FILLER_252_2000 ();
 b15zdnd11an1n08x5 FILLER_252_2051 ();
 b15zdnd00an1n02x5 FILLER_252_2059 ();
 b15zdnd11an1n32x5 FILLER_252_2067 ();
 b15zdnd11an1n04x5 FILLER_252_2099 ();
 b15zdnd00an1n02x5 FILLER_252_2103 ();
 b15zdnd00an1n01x5 FILLER_252_2105 ();
 b15zdnd11an1n16x5 FILLER_252_2120 ();
 b15zdnd11an1n08x5 FILLER_252_2136 ();
 b15zdnd00an1n02x5 FILLER_252_2144 ();
 b15zdnd00an1n02x5 FILLER_252_2152 ();
 b15zdnd11an1n16x5 FILLER_252_2162 ();
 b15zdnd11an1n08x5 FILLER_252_2178 ();
 b15zdnd00an1n02x5 FILLER_252_2186 ();
 b15zdnd00an1n01x5 FILLER_252_2188 ();
 b15zdnd11an1n16x5 FILLER_252_2213 ();
 b15zdnd11an1n08x5 FILLER_252_2229 ();
 b15zdnd11an1n16x5 FILLER_252_2245 ();
 b15zdnd11an1n08x5 FILLER_252_2261 ();
 b15zdnd11an1n04x5 FILLER_252_2269 ();
 b15zdnd00an1n02x5 FILLER_252_2273 ();
 b15zdnd00an1n01x5 FILLER_252_2275 ();
 b15zdnd11an1n64x5 FILLER_253_0 ();
 b15zdnd11an1n32x5 FILLER_253_64 ();
 b15zdnd00an1n02x5 FILLER_253_96 ();
 b15zdnd00an1n01x5 FILLER_253_98 ();
 b15zdnd11an1n04x5 FILLER_253_112 ();
 b15zdnd11an1n32x5 FILLER_253_147 ();
 b15zdnd11an1n08x5 FILLER_253_179 ();
 b15zdnd00an1n01x5 FILLER_253_187 ();
 b15zdnd11an1n08x5 FILLER_253_198 ();
 b15zdnd11an1n04x5 FILLER_253_206 ();
 b15zdnd00an1n02x5 FILLER_253_210 ();
 b15zdnd00an1n01x5 FILLER_253_212 ();
 b15zdnd11an1n64x5 FILLER_253_217 ();
 b15zdnd00an1n02x5 FILLER_253_281 ();
 b15zdnd11an1n16x5 FILLER_253_289 ();
 b15zdnd11an1n08x5 FILLER_253_305 ();
 b15zdnd00an1n02x5 FILLER_253_313 ();
 b15zdnd00an1n01x5 FILLER_253_315 ();
 b15zdnd11an1n04x5 FILLER_253_322 ();
 b15zdnd00an1n01x5 FILLER_253_326 ();
 b15zdnd11an1n08x5 FILLER_253_332 ();
 b15zdnd11an1n04x5 FILLER_253_340 ();
 b15zdnd11an1n64x5 FILLER_253_352 ();
 b15zdnd11an1n32x5 FILLER_253_416 ();
 b15zdnd00an1n02x5 FILLER_253_448 ();
 b15zdnd11an1n04x5 FILLER_253_454 ();
 b15zdnd11an1n08x5 FILLER_253_465 ();
 b15zdnd11an1n04x5 FILLER_253_473 ();
 b15zdnd00an1n02x5 FILLER_253_477 ();
 b15zdnd11an1n64x5 FILLER_253_484 ();
 b15zdnd11an1n32x5 FILLER_253_548 ();
 b15zdnd11an1n08x5 FILLER_253_580 ();
 b15zdnd11an1n04x5 FILLER_253_588 ();
 b15zdnd00an1n02x5 FILLER_253_592 ();
 b15zdnd00an1n01x5 FILLER_253_594 ();
 b15zdnd11an1n04x5 FILLER_253_602 ();
 b15zdnd11an1n32x5 FILLER_253_613 ();
 b15zdnd11an1n08x5 FILLER_253_645 ();
 b15zdnd11an1n04x5 FILLER_253_653 ();
 b15zdnd00an1n02x5 FILLER_253_657 ();
 b15zdnd00an1n01x5 FILLER_253_659 ();
 b15zdnd11an1n64x5 FILLER_253_670 ();
 b15zdnd11an1n04x5 FILLER_253_734 ();
 b15zdnd00an1n01x5 FILLER_253_738 ();
 b15zdnd11an1n08x5 FILLER_253_758 ();
 b15zdnd11an1n04x5 FILLER_253_766 ();
 b15zdnd00an1n02x5 FILLER_253_770 ();
 b15zdnd11an1n04x5 FILLER_253_777 ();
 b15zdnd11an1n16x5 FILLER_253_793 ();
 b15zdnd11an1n04x5 FILLER_253_809 ();
 b15zdnd11an1n64x5 FILLER_253_833 ();
 b15zdnd11an1n64x5 FILLER_253_897 ();
 b15zdnd11an1n32x5 FILLER_253_961 ();
 b15zdnd11an1n04x5 FILLER_253_993 ();
 b15zdnd00an1n02x5 FILLER_253_997 ();
 b15zdnd00an1n01x5 FILLER_253_999 ();
 b15zdnd11an1n08x5 FILLER_253_1006 ();
 b15zdnd11an1n32x5 FILLER_253_1030 ();
 b15zdnd11an1n04x5 FILLER_253_1062 ();
 b15zdnd00an1n02x5 FILLER_253_1066 ();
 b15zdnd00an1n01x5 FILLER_253_1068 ();
 b15zdnd11an1n16x5 FILLER_253_1073 ();
 b15zdnd11an1n04x5 FILLER_253_1089 ();
 b15zdnd00an1n02x5 FILLER_253_1093 ();
 b15zdnd00an1n01x5 FILLER_253_1095 ();
 b15zdnd11an1n04x5 FILLER_253_1102 ();
 b15zdnd11an1n08x5 FILLER_253_1115 ();
 b15zdnd00an1n02x5 FILLER_253_1123 ();
 b15zdnd11an1n32x5 FILLER_253_1131 ();
 b15zdnd11an1n16x5 FILLER_253_1169 ();
 b15zdnd11an1n08x5 FILLER_253_1185 ();
 b15zdnd00an1n02x5 FILLER_253_1193 ();
 b15zdnd11an1n04x5 FILLER_253_1210 ();
 b15zdnd00an1n02x5 FILLER_253_1214 ();
 b15zdnd00an1n01x5 FILLER_253_1216 ();
 b15zdnd11an1n16x5 FILLER_253_1227 ();
 b15zdnd11an1n04x5 FILLER_253_1243 ();
 b15zdnd00an1n02x5 FILLER_253_1247 ();
 b15zdnd11an1n04x5 FILLER_253_1263 ();
 b15zdnd00an1n02x5 FILLER_253_1267 ();
 b15zdnd00an1n01x5 FILLER_253_1269 ();
 b15zdnd11an1n64x5 FILLER_253_1280 ();
 b15zdnd11an1n64x5 FILLER_253_1344 ();
 b15zdnd11an1n32x5 FILLER_253_1408 ();
 b15zdnd11an1n04x5 FILLER_253_1440 ();
 b15zdnd11an1n16x5 FILLER_253_1457 ();
 b15zdnd11an1n08x5 FILLER_253_1473 ();
 b15zdnd11an1n04x5 FILLER_253_1481 ();
 b15zdnd00an1n02x5 FILLER_253_1485 ();
 b15zdnd00an1n01x5 FILLER_253_1487 ();
 b15zdnd11an1n04x5 FILLER_253_1513 ();
 b15zdnd11an1n64x5 FILLER_253_1543 ();
 b15zdnd11an1n64x5 FILLER_253_1607 ();
 b15zdnd11an1n64x5 FILLER_253_1671 ();
 b15zdnd00an1n02x5 FILLER_253_1735 ();
 b15zdnd11an1n08x5 FILLER_253_1744 ();
 b15zdnd00an1n02x5 FILLER_253_1752 ();
 b15zdnd11an1n64x5 FILLER_253_1758 ();
 b15zdnd11an1n64x5 FILLER_253_1822 ();
 b15zdnd11an1n04x5 FILLER_253_1886 ();
 b15zdnd00an1n02x5 FILLER_253_1890 ();
 b15zdnd00an1n01x5 FILLER_253_1892 ();
 b15zdnd11an1n32x5 FILLER_253_1900 ();
 b15zdnd00an1n02x5 FILLER_253_1932 ();
 b15zdnd11an1n64x5 FILLER_253_1942 ();
 b15zdnd11an1n04x5 FILLER_253_2006 ();
 b15zdnd00an1n02x5 FILLER_253_2010 ();
 b15zdnd11an1n64x5 FILLER_253_2018 ();
 b15zdnd11an1n64x5 FILLER_253_2082 ();
 b15zdnd11an1n32x5 FILLER_253_2146 ();
 b15zdnd11an1n16x5 FILLER_253_2178 ();
 b15zdnd00an1n02x5 FILLER_253_2194 ();
 b15zdnd00an1n01x5 FILLER_253_2196 ();
 b15zdnd11an1n16x5 FILLER_253_2205 ();
 b15zdnd00an1n01x5 FILLER_253_2221 ();
 b15zdnd11an1n04x5 FILLER_253_2231 ();
 b15zdnd11an1n04x5 FILLER_253_2251 ();
 b15zdnd11an1n16x5 FILLER_253_2259 ();
 b15zdnd11an1n08x5 FILLER_253_2275 ();
 b15zdnd00an1n01x5 FILLER_253_2283 ();
 b15zdnd11an1n64x5 FILLER_254_8 ();
 b15zdnd11an1n08x5 FILLER_254_72 ();
 b15zdnd00an1n02x5 FILLER_254_80 ();
 b15zdnd11an1n04x5 FILLER_254_89 ();
 b15zdnd11an1n32x5 FILLER_254_102 ();
 b15zdnd11an1n16x5 FILLER_254_134 ();
 b15zdnd11an1n08x5 FILLER_254_150 ();
 b15zdnd00an1n01x5 FILLER_254_158 ();
 b15zdnd11an1n16x5 FILLER_254_163 ();
 b15zdnd00an1n02x5 FILLER_254_179 ();
 b15zdnd11an1n16x5 FILLER_254_193 ();
 b15zdnd11an1n04x5 FILLER_254_209 ();
 b15zdnd00an1n02x5 FILLER_254_213 ();
 b15zdnd11an1n08x5 FILLER_254_221 ();
 b15zdnd11an1n04x5 FILLER_254_229 ();
 b15zdnd00an1n01x5 FILLER_254_233 ();
 b15zdnd11an1n08x5 FILLER_254_241 ();
 b15zdnd11an1n04x5 FILLER_254_249 ();
 b15zdnd11an1n04x5 FILLER_254_279 ();
 b15zdnd11an1n16x5 FILLER_254_288 ();
 b15zdnd11an1n08x5 FILLER_254_304 ();
 b15zdnd11an1n04x5 FILLER_254_312 ();
 b15zdnd00an1n01x5 FILLER_254_316 ();
 b15zdnd11an1n08x5 FILLER_254_323 ();
 b15zdnd11an1n04x5 FILLER_254_331 ();
 b15zdnd00an1n02x5 FILLER_254_335 ();
 b15zdnd11an1n08x5 FILLER_254_345 ();
 b15zdnd11an1n04x5 FILLER_254_353 ();
 b15zdnd00an1n02x5 FILLER_254_357 ();
 b15zdnd11an1n32x5 FILLER_254_368 ();
 b15zdnd11an1n16x5 FILLER_254_400 ();
 b15zdnd00an1n02x5 FILLER_254_416 ();
 b15zdnd00an1n01x5 FILLER_254_418 ();
 b15zdnd11an1n08x5 FILLER_254_435 ();
 b15zdnd11an1n04x5 FILLER_254_443 ();
 b15zdnd00an1n01x5 FILLER_254_447 ();
 b15zdnd11an1n16x5 FILLER_254_464 ();
 b15zdnd11an1n08x5 FILLER_254_480 ();
 b15zdnd00an1n02x5 FILLER_254_488 ();
 b15zdnd00an1n01x5 FILLER_254_490 ();
 b15zdnd11an1n16x5 FILLER_254_497 ();
 b15zdnd11an1n08x5 FILLER_254_513 ();
 b15zdnd00an1n02x5 FILLER_254_521 ();
 b15zdnd11an1n04x5 FILLER_254_529 ();
 b15zdnd00an1n01x5 FILLER_254_533 ();
 b15zdnd11an1n04x5 FILLER_254_548 ();
 b15zdnd11an1n08x5 FILLER_254_560 ();
 b15zdnd11an1n32x5 FILLER_254_583 ();
 b15zdnd11an1n08x5 FILLER_254_615 ();
 b15zdnd11an1n04x5 FILLER_254_623 ();
 b15zdnd11an1n16x5 FILLER_254_639 ();
 b15zdnd11an1n08x5 FILLER_254_655 ();
 b15zdnd00an1n02x5 FILLER_254_663 ();
 b15zdnd11an1n32x5 FILLER_254_681 ();
 b15zdnd11an1n04x5 FILLER_254_713 ();
 b15zdnd00an1n01x5 FILLER_254_717 ();
 b15zdnd11an1n08x5 FILLER_254_726 ();
 b15zdnd00an1n02x5 FILLER_254_734 ();
 b15zdnd00an1n01x5 FILLER_254_736 ();
 b15zdnd11an1n16x5 FILLER_254_741 ();
 b15zdnd11an1n08x5 FILLER_254_757 ();
 b15zdnd00an1n02x5 FILLER_254_765 ();
 b15zdnd11an1n16x5 FILLER_254_771 ();
 b15zdnd11an1n04x5 FILLER_254_787 ();
 b15zdnd00an1n01x5 FILLER_254_791 ();
 b15zdnd11an1n64x5 FILLER_254_799 ();
 b15zdnd11an1n08x5 FILLER_254_863 ();
 b15zdnd11an1n16x5 FILLER_254_880 ();
 b15zdnd00an1n02x5 FILLER_254_896 ();
 b15zdnd00an1n01x5 FILLER_254_898 ();
 b15zdnd11an1n04x5 FILLER_254_930 ();
 b15zdnd11an1n32x5 FILLER_254_949 ();
 b15zdnd11an1n08x5 FILLER_254_981 ();
 b15zdnd11an1n32x5 FILLER_254_1001 ();
 b15zdnd00an1n02x5 FILLER_254_1033 ();
 b15zdnd00an1n01x5 FILLER_254_1035 ();
 b15zdnd11an1n16x5 FILLER_254_1042 ();
 b15zdnd11an1n04x5 FILLER_254_1064 ();
 b15zdnd00an1n02x5 FILLER_254_1068 ();
 b15zdnd11an1n04x5 FILLER_254_1076 ();
 b15zdnd00an1n02x5 FILLER_254_1080 ();
 b15zdnd00an1n01x5 FILLER_254_1082 ();
 b15zdnd11an1n04x5 FILLER_254_1087 ();
 b15zdnd11an1n32x5 FILLER_254_1103 ();
 b15zdnd11an1n16x5 FILLER_254_1135 ();
 b15zdnd11an1n08x5 FILLER_254_1151 ();
 b15zdnd11an1n16x5 FILLER_254_1172 ();
 b15zdnd11an1n08x5 FILLER_254_1188 ();
 b15zdnd00an1n02x5 FILLER_254_1196 ();
 b15zdnd11an1n08x5 FILLER_254_1208 ();
 b15zdnd11an1n04x5 FILLER_254_1216 ();
 b15zdnd11an1n04x5 FILLER_254_1225 ();
 b15zdnd11an1n32x5 FILLER_254_1234 ();
 b15zdnd11an1n16x5 FILLER_254_1291 ();
 b15zdnd11an1n08x5 FILLER_254_1307 ();
 b15zdnd11an1n64x5 FILLER_254_1320 ();
 b15zdnd11an1n32x5 FILLER_254_1384 ();
 b15zdnd11an1n16x5 FILLER_254_1416 ();
 b15zdnd11an1n04x5 FILLER_254_1432 ();
 b15zdnd00an1n02x5 FILLER_254_1436 ();
 b15zdnd11an1n04x5 FILLER_254_1446 ();
 b15zdnd11an1n04x5 FILLER_254_1462 ();
 b15zdnd11an1n04x5 FILLER_254_1472 ();
 b15zdnd11an1n32x5 FILLER_254_1492 ();
 b15zdnd00an1n01x5 FILLER_254_1524 ();
 b15zdnd11an1n32x5 FILLER_254_1534 ();
 b15zdnd11an1n08x5 FILLER_254_1566 ();
 b15zdnd00an1n02x5 FILLER_254_1574 ();
 b15zdnd00an1n01x5 FILLER_254_1576 ();
 b15zdnd11an1n16x5 FILLER_254_1583 ();
 b15zdnd11an1n08x5 FILLER_254_1599 ();
 b15zdnd00an1n02x5 FILLER_254_1607 ();
 b15zdnd11an1n32x5 FILLER_254_1621 ();
 b15zdnd11an1n04x5 FILLER_254_1653 ();
 b15zdnd00an1n02x5 FILLER_254_1657 ();
 b15zdnd11an1n32x5 FILLER_254_1669 ();
 b15zdnd11an1n16x5 FILLER_254_1701 ();
 b15zdnd00an1n01x5 FILLER_254_1717 ();
 b15zdnd11an1n32x5 FILLER_254_1723 ();
 b15zdnd11an1n16x5 FILLER_254_1755 ();
 b15zdnd11an1n08x5 FILLER_254_1771 ();
 b15zdnd11an1n04x5 FILLER_254_1779 ();
 b15zdnd00an1n01x5 FILLER_254_1783 ();
 b15zdnd11an1n64x5 FILLER_254_1804 ();
 b15zdnd11an1n16x5 FILLER_254_1868 ();
 b15zdnd11an1n04x5 FILLER_254_1884 ();
 b15zdnd11an1n32x5 FILLER_254_1904 ();
 b15zdnd11an1n08x5 FILLER_254_1936 ();
 b15zdnd11an1n32x5 FILLER_254_1955 ();
 b15zdnd11an1n08x5 FILLER_254_1987 ();
 b15zdnd11an1n04x5 FILLER_254_1995 ();
 b15zdnd00an1n02x5 FILLER_254_1999 ();
 b15zdnd00an1n01x5 FILLER_254_2001 ();
 b15zdnd11an1n04x5 FILLER_254_2008 ();
 b15zdnd11an1n32x5 FILLER_254_2022 ();
 b15zdnd11an1n08x5 FILLER_254_2054 ();
 b15zdnd00an1n02x5 FILLER_254_2062 ();
 b15zdnd00an1n01x5 FILLER_254_2064 ();
 b15zdnd11an1n16x5 FILLER_254_2076 ();
 b15zdnd11an1n08x5 FILLER_254_2092 ();
 b15zdnd11an1n04x5 FILLER_254_2100 ();
 b15zdnd11an1n08x5 FILLER_254_2109 ();
 b15zdnd11an1n04x5 FILLER_254_2117 ();
 b15zdnd11an1n08x5 FILLER_254_2133 ();
 b15zdnd11an1n04x5 FILLER_254_2141 ();
 b15zdnd00an1n01x5 FILLER_254_2145 ();
 b15zdnd11an1n04x5 FILLER_254_2150 ();
 b15zdnd11an1n16x5 FILLER_254_2162 ();
 b15zdnd11an1n08x5 FILLER_254_2178 ();
 b15zdnd11an1n04x5 FILLER_254_2186 ();
 b15zdnd00an1n01x5 FILLER_254_2190 ();
 b15zdnd11an1n04x5 FILLER_254_2196 ();
 b15zdnd11an1n16x5 FILLER_254_2213 ();
 b15zdnd11an1n04x5 FILLER_254_2229 ();
 b15zdnd11an1n08x5 FILLER_254_2239 ();
 b15zdnd00an1n01x5 FILLER_254_2247 ();
 b15zdnd11an1n16x5 FILLER_254_2253 ();
 b15zdnd11an1n04x5 FILLER_254_2269 ();
 b15zdnd00an1n02x5 FILLER_254_2273 ();
 b15zdnd00an1n01x5 FILLER_254_2275 ();
 b15zdnd11an1n32x5 FILLER_255_0 ();
 b15zdnd11an1n04x5 FILLER_255_32 ();
 b15zdnd00an1n02x5 FILLER_255_36 ();
 b15zdnd11an1n04x5 FILLER_255_44 ();
 b15zdnd11an1n16x5 FILLER_255_53 ();
 b15zdnd00an1n01x5 FILLER_255_69 ();
 b15zdnd11an1n16x5 FILLER_255_85 ();
 b15zdnd11an1n08x5 FILLER_255_101 ();
 b15zdnd11an1n04x5 FILLER_255_109 ();
 b15zdnd00an1n02x5 FILLER_255_113 ();
 b15zdnd00an1n01x5 FILLER_255_115 ();
 b15zdnd11an1n16x5 FILLER_255_126 ();
 b15zdnd11an1n64x5 FILLER_255_157 ();
 b15zdnd11an1n16x5 FILLER_255_221 ();
 b15zdnd11an1n08x5 FILLER_255_237 ();
 b15zdnd11an1n04x5 FILLER_255_245 ();
 b15zdnd00an1n02x5 FILLER_255_249 ();
 b15zdnd00an1n01x5 FILLER_255_251 ();
 b15zdnd11an1n16x5 FILLER_255_258 ();
 b15zdnd11an1n08x5 FILLER_255_274 ();
 b15zdnd11an1n04x5 FILLER_255_282 ();
 b15zdnd00an1n01x5 FILLER_255_286 ();
 b15zdnd11an1n16x5 FILLER_255_295 ();
 b15zdnd00an1n01x5 FILLER_255_311 ();
 b15zdnd11an1n64x5 FILLER_255_326 ();
 b15zdnd11an1n32x5 FILLER_255_390 ();
 b15zdnd00an1n01x5 FILLER_255_422 ();
 b15zdnd11an1n32x5 FILLER_255_429 ();
 b15zdnd11an1n16x5 FILLER_255_461 ();
 b15zdnd11an1n08x5 FILLER_255_477 ();
 b15zdnd11an1n04x5 FILLER_255_485 ();
 b15zdnd00an1n01x5 FILLER_255_489 ();
 b15zdnd11an1n16x5 FILLER_255_522 ();
 b15zdnd11an1n04x5 FILLER_255_538 ();
 b15zdnd00an1n02x5 FILLER_255_542 ();
 b15zdnd00an1n01x5 FILLER_255_544 ();
 b15zdnd11an1n04x5 FILLER_255_558 ();
 b15zdnd00an1n01x5 FILLER_255_562 ();
 b15zdnd11an1n08x5 FILLER_255_580 ();
 b15zdnd11an1n04x5 FILLER_255_588 ();
 b15zdnd00an1n02x5 FILLER_255_592 ();
 b15zdnd11an1n32x5 FILLER_255_600 ();
 b15zdnd11an1n16x5 FILLER_255_632 ();
 b15zdnd11an1n08x5 FILLER_255_648 ();
 b15zdnd11an1n04x5 FILLER_255_656 ();
 b15zdnd00an1n02x5 FILLER_255_660 ();
 b15zdnd11an1n16x5 FILLER_255_666 ();
 b15zdnd00an1n02x5 FILLER_255_682 ();
 b15zdnd00an1n01x5 FILLER_255_684 ();
 b15zdnd11an1n16x5 FILLER_255_705 ();
 b15zdnd11an1n04x5 FILLER_255_721 ();
 b15zdnd00an1n02x5 FILLER_255_725 ();
 b15zdnd11an1n04x5 FILLER_255_732 ();
 b15zdnd11an1n64x5 FILLER_255_748 ();
 b15zdnd11an1n16x5 FILLER_255_812 ();
 b15zdnd11an1n04x5 FILLER_255_828 ();
 b15zdnd00an1n01x5 FILLER_255_832 ();
 b15zdnd11an1n32x5 FILLER_255_843 ();
 b15zdnd11an1n08x5 FILLER_255_875 ();
 b15zdnd11an1n04x5 FILLER_255_883 ();
 b15zdnd00an1n02x5 FILLER_255_887 ();
 b15zdnd00an1n01x5 FILLER_255_889 ();
 b15zdnd11an1n32x5 FILLER_255_915 ();
 b15zdnd11an1n16x5 FILLER_255_947 ();
 b15zdnd11an1n08x5 FILLER_255_963 ();
 b15zdnd11an1n04x5 FILLER_255_971 ();
 b15zdnd00an1n02x5 FILLER_255_975 ();
 b15zdnd00an1n01x5 FILLER_255_977 ();
 b15zdnd11an1n64x5 FILLER_255_988 ();
 b15zdnd11an1n16x5 FILLER_255_1052 ();
 b15zdnd00an1n01x5 FILLER_255_1068 ();
 b15zdnd11an1n64x5 FILLER_255_1074 ();
 b15zdnd00an1n02x5 FILLER_255_1138 ();
 b15zdnd00an1n01x5 FILLER_255_1140 ();
 b15zdnd11an1n08x5 FILLER_255_1147 ();
 b15zdnd11an1n04x5 FILLER_255_1155 ();
 b15zdnd00an1n02x5 FILLER_255_1159 ();
 b15zdnd00an1n01x5 FILLER_255_1161 ();
 b15zdnd11an1n16x5 FILLER_255_1176 ();
 b15zdnd11an1n04x5 FILLER_255_1197 ();
 b15zdnd11an1n16x5 FILLER_255_1206 ();
 b15zdnd11an1n08x5 FILLER_255_1222 ();
 b15zdnd11an1n64x5 FILLER_255_1241 ();
 b15zdnd11an1n04x5 FILLER_255_1305 ();
 b15zdnd00an1n02x5 FILLER_255_1309 ();
 b15zdnd00an1n01x5 FILLER_255_1311 ();
 b15zdnd11an1n04x5 FILLER_255_1317 ();
 b15zdnd11an1n04x5 FILLER_255_1326 ();
 b15zdnd11an1n08x5 FILLER_255_1335 ();
 b15zdnd00an1n01x5 FILLER_255_1343 ();
 b15zdnd11an1n04x5 FILLER_255_1365 ();
 b15zdnd11an1n64x5 FILLER_255_1381 ();
 b15zdnd11an1n32x5 FILLER_255_1445 ();
 b15zdnd11an1n04x5 FILLER_255_1477 ();
 b15zdnd11an1n16x5 FILLER_255_1487 ();
 b15zdnd11an1n04x5 FILLER_255_1503 ();
 b15zdnd00an1n01x5 FILLER_255_1507 ();
 b15zdnd11an1n04x5 FILLER_255_1524 ();
 b15zdnd11an1n32x5 FILLER_255_1534 ();
 b15zdnd11an1n08x5 FILLER_255_1566 ();
 b15zdnd11an1n04x5 FILLER_255_1579 ();
 b15zdnd00an1n01x5 FILLER_255_1583 ();
 b15zdnd11an1n16x5 FILLER_255_1598 ();
 b15zdnd11an1n08x5 FILLER_255_1614 ();
 b15zdnd11an1n04x5 FILLER_255_1622 ();
 b15zdnd00an1n02x5 FILLER_255_1626 ();
 b15zdnd00an1n01x5 FILLER_255_1628 ();
 b15zdnd11an1n08x5 FILLER_255_1643 ();
 b15zdnd11an1n04x5 FILLER_255_1651 ();
 b15zdnd00an1n02x5 FILLER_255_1655 ();
 b15zdnd00an1n01x5 FILLER_255_1657 ();
 b15zdnd11an1n08x5 FILLER_255_1674 ();
 b15zdnd11an1n04x5 FILLER_255_1682 ();
 b15zdnd00an1n02x5 FILLER_255_1686 ();
 b15zdnd11an1n32x5 FILLER_255_1694 ();
 b15zdnd11an1n16x5 FILLER_255_1726 ();
 b15zdnd11an1n08x5 FILLER_255_1742 ();
 b15zdnd00an1n01x5 FILLER_255_1750 ();
 b15zdnd11an1n32x5 FILLER_255_1767 ();
 b15zdnd11an1n16x5 FILLER_255_1799 ();
 b15zdnd11an1n04x5 FILLER_255_1815 ();
 b15zdnd00an1n02x5 FILLER_255_1819 ();
 b15zdnd00an1n01x5 FILLER_255_1821 ();
 b15zdnd11an1n32x5 FILLER_255_1827 ();
 b15zdnd11an1n04x5 FILLER_255_1859 ();
 b15zdnd11an1n32x5 FILLER_255_1889 ();
 b15zdnd11an1n16x5 FILLER_255_1921 ();
 b15zdnd11an1n08x5 FILLER_255_1937 ();
 b15zdnd11an1n16x5 FILLER_255_1951 ();
 b15zdnd11an1n04x5 FILLER_255_1967 ();
 b15zdnd11an1n08x5 FILLER_255_1978 ();
 b15zdnd11an1n04x5 FILLER_255_1986 ();
 b15zdnd00an1n02x5 FILLER_255_1990 ();
 b15zdnd00an1n01x5 FILLER_255_1992 ();
 b15zdnd11an1n08x5 FILLER_255_1999 ();
 b15zdnd11an1n04x5 FILLER_255_2007 ();
 b15zdnd00an1n02x5 FILLER_255_2011 ();
 b15zdnd11an1n16x5 FILLER_255_2029 ();
 b15zdnd11an1n08x5 FILLER_255_2045 ();
 b15zdnd11an1n04x5 FILLER_255_2053 ();
 b15zdnd11an1n16x5 FILLER_255_2072 ();
 b15zdnd11an1n08x5 FILLER_255_2088 ();
 b15zdnd00an1n02x5 FILLER_255_2096 ();
 b15zdnd11an1n64x5 FILLER_255_2103 ();
 b15zdnd11an1n64x5 FILLER_255_2167 ();
 b15zdnd11an1n32x5 FILLER_255_2231 ();
 b15zdnd11an1n16x5 FILLER_255_2263 ();
 b15zdnd11an1n04x5 FILLER_255_2279 ();
 b15zdnd00an1n01x5 FILLER_255_2283 ();
 b15zdnd11an1n16x5 FILLER_256_8 ();
 b15zdnd11an1n08x5 FILLER_256_24 ();
 b15zdnd11an1n04x5 FILLER_256_32 ();
 b15zdnd00an1n01x5 FILLER_256_36 ();
 b15zdnd11an1n04x5 FILLER_256_41 ();
 b15zdnd11an1n04x5 FILLER_256_60 ();
 b15zdnd11an1n32x5 FILLER_256_85 ();
 b15zdnd11an1n16x5 FILLER_256_117 ();
 b15zdnd11an1n08x5 FILLER_256_133 ();
 b15zdnd11an1n08x5 FILLER_256_145 ();
 b15zdnd11an1n04x5 FILLER_256_153 ();
 b15zdnd11an1n16x5 FILLER_256_162 ();
 b15zdnd00an1n02x5 FILLER_256_178 ();
 b15zdnd11an1n16x5 FILLER_256_187 ();
 b15zdnd11an1n04x5 FILLER_256_203 ();
 b15zdnd11an1n32x5 FILLER_256_212 ();
 b15zdnd00an1n02x5 FILLER_256_244 ();
 b15zdnd11an1n16x5 FILLER_256_252 ();
 b15zdnd00an1n01x5 FILLER_256_268 ();
 b15zdnd11an1n32x5 FILLER_256_281 ();
 b15zdnd11an1n16x5 FILLER_256_313 ();
 b15zdnd00an1n02x5 FILLER_256_329 ();
 b15zdnd00an1n01x5 FILLER_256_331 ();
 b15zdnd11an1n64x5 FILLER_256_338 ();
 b15zdnd11an1n64x5 FILLER_256_402 ();
 b15zdnd11an1n16x5 FILLER_256_466 ();
 b15zdnd00an1n02x5 FILLER_256_482 ();
 b15zdnd11an1n08x5 FILLER_256_496 ();
 b15zdnd11an1n04x5 FILLER_256_504 ();
 b15zdnd00an1n01x5 FILLER_256_508 ();
 b15zdnd11an1n32x5 FILLER_256_518 ();
 b15zdnd11an1n04x5 FILLER_256_550 ();
 b15zdnd00an1n02x5 FILLER_256_554 ();
 b15zdnd11an1n32x5 FILLER_256_565 ();
 b15zdnd11an1n08x5 FILLER_256_597 ();
 b15zdnd11an1n04x5 FILLER_256_605 ();
 b15zdnd00an1n02x5 FILLER_256_609 ();
 b15zdnd00an1n01x5 FILLER_256_611 ();
 b15zdnd11an1n04x5 FILLER_256_624 ();
 b15zdnd11an1n16x5 FILLER_256_639 ();
 b15zdnd11an1n08x5 FILLER_256_655 ();
 b15zdnd11an1n08x5 FILLER_256_669 ();
 b15zdnd11an1n04x5 FILLER_256_677 ();
 b15zdnd11an1n08x5 FILLER_256_697 ();
 b15zdnd11an1n04x5 FILLER_256_705 ();
 b15zdnd00an1n02x5 FILLER_256_709 ();
 b15zdnd00an1n01x5 FILLER_256_711 ();
 b15zdnd00an1n02x5 FILLER_256_716 ();
 b15zdnd11an1n64x5 FILLER_256_726 ();
 b15zdnd00an1n02x5 FILLER_256_790 ();
 b15zdnd11an1n04x5 FILLER_256_804 ();
 b15zdnd11an1n16x5 FILLER_256_812 ();
 b15zdnd11an1n08x5 FILLER_256_828 ();
 b15zdnd11an1n04x5 FILLER_256_836 ();
 b15zdnd00an1n02x5 FILLER_256_840 ();
 b15zdnd11an1n64x5 FILLER_256_851 ();
 b15zdnd11an1n64x5 FILLER_256_915 ();
 b15zdnd11an1n16x5 FILLER_256_979 ();
 b15zdnd00an1n02x5 FILLER_256_995 ();
 b15zdnd00an1n01x5 FILLER_256_997 ();
 b15zdnd11an1n16x5 FILLER_256_1010 ();
 b15zdnd11an1n64x5 FILLER_256_1030 ();
 b15zdnd11an1n64x5 FILLER_256_1094 ();
 b15zdnd11an1n64x5 FILLER_256_1158 ();
 b15zdnd11an1n32x5 FILLER_256_1222 ();
 b15zdnd11an1n04x5 FILLER_256_1254 ();
 b15zdnd00an1n02x5 FILLER_256_1258 ();
 b15zdnd11an1n64x5 FILLER_256_1265 ();
 b15zdnd11an1n04x5 FILLER_256_1329 ();
 b15zdnd00an1n02x5 FILLER_256_1333 ();
 b15zdnd00an1n01x5 FILLER_256_1335 ();
 b15zdnd11an1n64x5 FILLER_256_1350 ();
 b15zdnd11an1n08x5 FILLER_256_1414 ();
 b15zdnd11an1n04x5 FILLER_256_1422 ();
 b15zdnd00an1n02x5 FILLER_256_1426 ();
 b15zdnd00an1n01x5 FILLER_256_1428 ();
 b15zdnd11an1n32x5 FILLER_256_1435 ();
 b15zdnd11an1n04x5 FILLER_256_1467 ();
 b15zdnd00an1n02x5 FILLER_256_1471 ();
 b15zdnd11an1n32x5 FILLER_256_1487 ();
 b15zdnd11an1n08x5 FILLER_256_1519 ();
 b15zdnd00an1n02x5 FILLER_256_1527 ();
 b15zdnd11an1n04x5 FILLER_256_1536 ();
 b15zdnd00an1n02x5 FILLER_256_1540 ();
 b15zdnd11an1n32x5 FILLER_256_1552 ();
 b15zdnd11an1n16x5 FILLER_256_1584 ();
 b15zdnd00an1n01x5 FILLER_256_1600 ();
 b15zdnd11an1n16x5 FILLER_256_1610 ();
 b15zdnd11an1n04x5 FILLER_256_1633 ();
 b15zdnd11an1n04x5 FILLER_256_1657 ();
 b15zdnd11an1n04x5 FILLER_256_1672 ();
 b15zdnd11an1n08x5 FILLER_256_1682 ();
 b15zdnd11an1n32x5 FILLER_256_1702 ();
 b15zdnd11an1n04x5 FILLER_256_1734 ();
 b15zdnd00an1n02x5 FILLER_256_1738 ();
 b15zdnd00an1n01x5 FILLER_256_1740 ();
 b15zdnd11an1n04x5 FILLER_256_1747 ();
 b15zdnd11an1n64x5 FILLER_256_1757 ();
 b15zdnd11an1n32x5 FILLER_256_1830 ();
 b15zdnd11an1n08x5 FILLER_256_1862 ();
 b15zdnd11an1n04x5 FILLER_256_1870 ();
 b15zdnd11an1n32x5 FILLER_256_1900 ();
 b15zdnd11an1n16x5 FILLER_256_1932 ();
 b15zdnd00an1n02x5 FILLER_256_1948 ();
 b15zdnd00an1n01x5 FILLER_256_1950 ();
 b15zdnd11an1n16x5 FILLER_256_1955 ();
 b15zdnd11an1n04x5 FILLER_256_1971 ();
 b15zdnd11an1n64x5 FILLER_256_1983 ();
 b15zdnd11an1n32x5 FILLER_256_2047 ();
 b15zdnd11an1n16x5 FILLER_256_2079 ();
 b15zdnd11an1n04x5 FILLER_256_2095 ();
 b15zdnd00an1n02x5 FILLER_256_2099 ();
 b15zdnd11an1n32x5 FILLER_256_2107 ();
 b15zdnd11an1n08x5 FILLER_256_2139 ();
 b15zdnd11an1n04x5 FILLER_256_2147 ();
 b15zdnd00an1n02x5 FILLER_256_2151 ();
 b15zdnd00an1n01x5 FILLER_256_2153 ();
 b15zdnd00an1n02x5 FILLER_256_2162 ();
 b15zdnd00an1n01x5 FILLER_256_2164 ();
 b15zdnd11an1n04x5 FILLER_256_2174 ();
 b15zdnd11an1n04x5 FILLER_256_2189 ();
 b15zdnd11an1n04x5 FILLER_256_2201 ();
 b15zdnd11an1n32x5 FILLER_256_2217 ();
 b15zdnd11an1n16x5 FILLER_256_2249 ();
 b15zdnd11an1n08x5 FILLER_256_2265 ();
 b15zdnd00an1n02x5 FILLER_256_2273 ();
 b15zdnd00an1n01x5 FILLER_256_2275 ();
 b15zdnd11an1n32x5 FILLER_257_0 ();
 b15zdnd00an1n02x5 FILLER_257_32 ();
 b15zdnd00an1n01x5 FILLER_257_34 ();
 b15zdnd11an1n16x5 FILLER_257_40 ();
 b15zdnd11an1n08x5 FILLER_257_56 ();
 b15zdnd00an1n02x5 FILLER_257_64 ();
 b15zdnd00an1n01x5 FILLER_257_66 ();
 b15zdnd11an1n08x5 FILLER_257_80 ();
 b15zdnd00an1n02x5 FILLER_257_88 ();
 b15zdnd11an1n64x5 FILLER_257_96 ();
 b15zdnd11an1n16x5 FILLER_257_160 ();
 b15zdnd11an1n16x5 FILLER_257_185 ();
 b15zdnd00an1n01x5 FILLER_257_201 ();
 b15zdnd11an1n64x5 FILLER_257_209 ();
 b15zdnd11an1n08x5 FILLER_257_273 ();
 b15zdnd11an1n04x5 FILLER_257_281 ();
 b15zdnd00an1n02x5 FILLER_257_285 ();
 b15zdnd11an1n08x5 FILLER_257_303 ();
 b15zdnd11an1n04x5 FILLER_257_311 ();
 b15zdnd00an1n02x5 FILLER_257_315 ();
 b15zdnd11an1n64x5 FILLER_257_326 ();
 b15zdnd11an1n32x5 FILLER_257_390 ();
 b15zdnd11an1n08x5 FILLER_257_422 ();
 b15zdnd00an1n02x5 FILLER_257_430 ();
 b15zdnd00an1n01x5 FILLER_257_432 ();
 b15zdnd11an1n64x5 FILLER_257_439 ();
 b15zdnd11an1n04x5 FILLER_257_503 ();
 b15zdnd11an1n64x5 FILLER_257_512 ();
 b15zdnd11an1n64x5 FILLER_257_576 ();
 b15zdnd00an1n01x5 FILLER_257_640 ();
 b15zdnd11an1n04x5 FILLER_257_646 ();
 b15zdnd00an1n01x5 FILLER_257_650 ();
 b15zdnd11an1n16x5 FILLER_257_659 ();
 b15zdnd11an1n08x5 FILLER_257_675 ();
 b15zdnd00an1n02x5 FILLER_257_683 ();
 b15zdnd00an1n01x5 FILLER_257_685 ();
 b15zdnd11an1n04x5 FILLER_257_706 ();
 b15zdnd11an1n64x5 FILLER_257_717 ();
 b15zdnd11an1n16x5 FILLER_257_781 ();
 b15zdnd11an1n64x5 FILLER_257_804 ();
 b15zdnd11an1n64x5 FILLER_257_868 ();
 b15zdnd11an1n08x5 FILLER_257_932 ();
 b15zdnd11an1n04x5 FILLER_257_940 ();
 b15zdnd00an1n02x5 FILLER_257_944 ();
 b15zdnd11an1n04x5 FILLER_257_951 ();
 b15zdnd11an1n32x5 FILLER_257_960 ();
 b15zdnd11an1n16x5 FILLER_257_1010 ();
 b15zdnd00an1n02x5 FILLER_257_1026 ();
 b15zdnd00an1n01x5 FILLER_257_1028 ();
 b15zdnd11an1n04x5 FILLER_257_1034 ();
 b15zdnd11an1n32x5 FILLER_257_1044 ();
 b15zdnd11an1n16x5 FILLER_257_1076 ();
 b15zdnd11an1n04x5 FILLER_257_1092 ();
 b15zdnd11an1n16x5 FILLER_257_1101 ();
 b15zdnd11an1n08x5 FILLER_257_1117 ();
 b15zdnd11an1n04x5 FILLER_257_1125 ();
 b15zdnd00an1n02x5 FILLER_257_1129 ();
 b15zdnd00an1n01x5 FILLER_257_1131 ();
 b15zdnd11an1n04x5 FILLER_257_1141 ();
 b15zdnd00an1n02x5 FILLER_257_1145 ();
 b15zdnd00an1n01x5 FILLER_257_1147 ();
 b15zdnd11an1n32x5 FILLER_257_1160 ();
 b15zdnd11an1n16x5 FILLER_257_1192 ();
 b15zdnd11an1n08x5 FILLER_257_1208 ();
 b15zdnd11an1n04x5 FILLER_257_1216 ();
 b15zdnd00an1n02x5 FILLER_257_1220 ();
 b15zdnd11an1n64x5 FILLER_257_1226 ();
 b15zdnd11an1n04x5 FILLER_257_1290 ();
 b15zdnd11an1n16x5 FILLER_257_1305 ();
 b15zdnd00an1n02x5 FILLER_257_1321 ();
 b15zdnd00an1n01x5 FILLER_257_1323 ();
 b15zdnd11an1n16x5 FILLER_257_1331 ();
 b15zdnd11an1n08x5 FILLER_257_1347 ();
 b15zdnd11an1n04x5 FILLER_257_1355 ();
 b15zdnd00an1n01x5 FILLER_257_1359 ();
 b15zdnd11an1n64x5 FILLER_257_1366 ();
 b15zdnd00an1n02x5 FILLER_257_1430 ();
 b15zdnd00an1n01x5 FILLER_257_1432 ();
 b15zdnd11an1n32x5 FILLER_257_1443 ();
 b15zdnd11an1n04x5 FILLER_257_1475 ();
 b15zdnd00an1n02x5 FILLER_257_1479 ();
 b15zdnd11an1n16x5 FILLER_257_1485 ();
 b15zdnd11an1n08x5 FILLER_257_1501 ();
 b15zdnd11an1n04x5 FILLER_257_1509 ();
 b15zdnd00an1n02x5 FILLER_257_1513 ();
 b15zdnd00an1n01x5 FILLER_257_1515 ();
 b15zdnd11an1n08x5 FILLER_257_1522 ();
 b15zdnd00an1n01x5 FILLER_257_1530 ();
 b15zdnd11an1n32x5 FILLER_257_1542 ();
 b15zdnd11an1n16x5 FILLER_257_1574 ();
 b15zdnd11an1n04x5 FILLER_257_1590 ();
 b15zdnd00an1n02x5 FILLER_257_1594 ();
 b15zdnd11an1n04x5 FILLER_257_1602 ();
 b15zdnd00an1n02x5 FILLER_257_1606 ();
 b15zdnd11an1n04x5 FILLER_257_1614 ();
 b15zdnd11an1n16x5 FILLER_257_1639 ();
 b15zdnd11an1n08x5 FILLER_257_1655 ();
 b15zdnd11an1n64x5 FILLER_257_1676 ();
 b15zdnd11an1n08x5 FILLER_257_1740 ();
 b15zdnd00an1n01x5 FILLER_257_1748 ();
 b15zdnd11an1n04x5 FILLER_257_1755 ();
 b15zdnd00an1n01x5 FILLER_257_1759 ();
 b15zdnd11an1n04x5 FILLER_257_1778 ();
 b15zdnd11an1n64x5 FILLER_257_1794 ();
 b15zdnd11an1n32x5 FILLER_257_1858 ();
 b15zdnd11an1n16x5 FILLER_257_1890 ();
 b15zdnd11an1n04x5 FILLER_257_1906 ();
 b15zdnd00an1n02x5 FILLER_257_1910 ();
 b15zdnd00an1n01x5 FILLER_257_1912 ();
 b15zdnd11an1n16x5 FILLER_257_1922 ();
 b15zdnd00an1n02x5 FILLER_257_1938 ();
 b15zdnd00an1n01x5 FILLER_257_1940 ();
 b15zdnd11an1n64x5 FILLER_257_1953 ();
 b15zdnd11an1n32x5 FILLER_257_2017 ();
 b15zdnd00an1n02x5 FILLER_257_2049 ();
 b15zdnd11an1n04x5 FILLER_257_2058 ();
 b15zdnd11an1n04x5 FILLER_257_2077 ();
 b15zdnd00an1n01x5 FILLER_257_2081 ();
 b15zdnd11an1n04x5 FILLER_257_2087 ();
 b15zdnd11an1n32x5 FILLER_257_2097 ();
 b15zdnd11an1n08x5 FILLER_257_2129 ();
 b15zdnd00an1n02x5 FILLER_257_2137 ();
 b15zdnd11an1n16x5 FILLER_257_2145 ();
 b15zdnd11an1n04x5 FILLER_257_2161 ();
 b15zdnd00an1n01x5 FILLER_257_2165 ();
 b15zdnd11an1n16x5 FILLER_257_2178 ();
 b15zdnd00an1n01x5 FILLER_257_2194 ();
 b15zdnd11an1n16x5 FILLER_257_2200 ();
 b15zdnd11an1n08x5 FILLER_257_2230 ();
 b15zdnd00an1n02x5 FILLER_257_2238 ();
 b15zdnd11an1n32x5 FILLER_257_2244 ();
 b15zdnd11an1n08x5 FILLER_257_2276 ();
 b15zdnd11an1n64x5 FILLER_258_8 ();
 b15zdnd11an1n32x5 FILLER_258_72 ();
 b15zdnd11an1n04x5 FILLER_258_104 ();
 b15zdnd00an1n02x5 FILLER_258_108 ();
 b15zdnd11an1n16x5 FILLER_258_119 ();
 b15zdnd11an1n04x5 FILLER_258_135 ();
 b15zdnd00an1n02x5 FILLER_258_139 ();
 b15zdnd11an1n32x5 FILLER_258_161 ();
 b15zdnd11an1n16x5 FILLER_258_193 ();
 b15zdnd11an1n08x5 FILLER_258_209 ();
 b15zdnd11an1n04x5 FILLER_258_217 ();
 b15zdnd00an1n02x5 FILLER_258_221 ();
 b15zdnd00an1n01x5 FILLER_258_223 ();
 b15zdnd11an1n04x5 FILLER_258_229 ();
 b15zdnd11an1n04x5 FILLER_258_238 ();
 b15zdnd11an1n08x5 FILLER_258_248 ();
 b15zdnd11an1n04x5 FILLER_258_256 ();
 b15zdnd00an1n02x5 FILLER_258_260 ();
 b15zdnd00an1n01x5 FILLER_258_262 ();
 b15zdnd11an1n04x5 FILLER_258_273 ();
 b15zdnd11an1n16x5 FILLER_258_287 ();
 b15zdnd11an1n04x5 FILLER_258_303 ();
 b15zdnd00an1n02x5 FILLER_258_307 ();
 b15zdnd11an1n32x5 FILLER_258_323 ();
 b15zdnd11an1n04x5 FILLER_258_355 ();
 b15zdnd00an1n01x5 FILLER_258_359 ();
 b15zdnd11an1n32x5 FILLER_258_371 ();
 b15zdnd11an1n08x5 FILLER_258_403 ();
 b15zdnd11an1n04x5 FILLER_258_411 ();
 b15zdnd00an1n01x5 FILLER_258_415 ();
 b15zdnd11an1n04x5 FILLER_258_423 ();
 b15zdnd00an1n02x5 FILLER_258_427 ();
 b15zdnd00an1n01x5 FILLER_258_429 ();
 b15zdnd11an1n04x5 FILLER_258_435 ();
 b15zdnd11an1n32x5 FILLER_258_448 ();
 b15zdnd11an1n08x5 FILLER_258_480 ();
 b15zdnd00an1n01x5 FILLER_258_488 ();
 b15zdnd11an1n64x5 FILLER_258_495 ();
 b15zdnd11an1n64x5 FILLER_258_559 ();
 b15zdnd11an1n32x5 FILLER_258_623 ();
 b15zdnd11an1n16x5 FILLER_258_655 ();
 b15zdnd11an1n08x5 FILLER_258_671 ();
 b15zdnd11an1n04x5 FILLER_258_679 ();
 b15zdnd11an1n16x5 FILLER_258_688 ();
 b15zdnd11an1n08x5 FILLER_258_704 ();
 b15zdnd11an1n04x5 FILLER_258_712 ();
 b15zdnd00an1n02x5 FILLER_258_716 ();
 b15zdnd11an1n08x5 FILLER_258_726 ();
 b15zdnd00an1n01x5 FILLER_258_734 ();
 b15zdnd11an1n04x5 FILLER_258_749 ();
 b15zdnd11an1n16x5 FILLER_258_757 ();
 b15zdnd11an1n04x5 FILLER_258_773 ();
 b15zdnd00an1n02x5 FILLER_258_777 ();
 b15zdnd00an1n01x5 FILLER_258_779 ();
 b15zdnd11an1n04x5 FILLER_258_796 ();
 b15zdnd11an1n64x5 FILLER_258_809 ();
 b15zdnd11an1n16x5 FILLER_258_873 ();
 b15zdnd00an1n02x5 FILLER_258_889 ();
 b15zdnd00an1n01x5 FILLER_258_891 ();
 b15zdnd11an1n32x5 FILLER_258_910 ();
 b15zdnd11an1n16x5 FILLER_258_942 ();
 b15zdnd11an1n04x5 FILLER_258_958 ();
 b15zdnd11an1n08x5 FILLER_258_975 ();
 b15zdnd11an1n04x5 FILLER_258_983 ();
 b15zdnd00an1n01x5 FILLER_258_987 ();
 b15zdnd11an1n04x5 FILLER_258_993 ();
 b15zdnd11an1n08x5 FILLER_258_1003 ();
 b15zdnd00an1n02x5 FILLER_258_1011 ();
 b15zdnd11an1n16x5 FILLER_258_1027 ();
 b15zdnd11an1n08x5 FILLER_258_1043 ();
 b15zdnd00an1n02x5 FILLER_258_1051 ();
 b15zdnd11an1n32x5 FILLER_258_1058 ();
 b15zdnd11an1n04x5 FILLER_258_1090 ();
 b15zdnd11an1n32x5 FILLER_258_1100 ();
 b15zdnd11an1n16x5 FILLER_258_1132 ();
 b15zdnd11an1n04x5 FILLER_258_1148 ();
 b15zdnd00an1n01x5 FILLER_258_1152 ();
 b15zdnd11an1n08x5 FILLER_258_1158 ();
 b15zdnd00an1n01x5 FILLER_258_1166 ();
 b15zdnd11an1n16x5 FILLER_258_1173 ();
 b15zdnd11an1n08x5 FILLER_258_1189 ();
 b15zdnd11an1n04x5 FILLER_258_1197 ();
 b15zdnd00an1n02x5 FILLER_258_1201 ();
 b15zdnd00an1n01x5 FILLER_258_1203 ();
 b15zdnd11an1n04x5 FILLER_258_1210 ();
 b15zdnd00an1n02x5 FILLER_258_1214 ();
 b15zdnd11an1n08x5 FILLER_258_1222 ();
 b15zdnd00an1n02x5 FILLER_258_1230 ();
 b15zdnd00an1n01x5 FILLER_258_1232 ();
 b15zdnd11an1n04x5 FILLER_258_1241 ();
 b15zdnd00an1n02x5 FILLER_258_1245 ();
 b15zdnd00an1n01x5 FILLER_258_1247 ();
 b15zdnd11an1n16x5 FILLER_258_1255 ();
 b15zdnd11an1n08x5 FILLER_258_1271 ();
 b15zdnd00an1n02x5 FILLER_258_1279 ();
 b15zdnd00an1n01x5 FILLER_258_1281 ();
 b15zdnd11an1n08x5 FILLER_258_1286 ();
 b15zdnd11an1n04x5 FILLER_258_1294 ();
 b15zdnd00an1n01x5 FILLER_258_1298 ();
 b15zdnd11an1n32x5 FILLER_258_1312 ();
 b15zdnd11an1n08x5 FILLER_258_1344 ();
 b15zdnd11an1n04x5 FILLER_258_1352 ();
 b15zdnd00an1n02x5 FILLER_258_1356 ();
 b15zdnd11an1n04x5 FILLER_258_1363 ();
 b15zdnd11an1n32x5 FILLER_258_1387 ();
 b15zdnd11an1n08x5 FILLER_258_1419 ();
 b15zdnd00an1n02x5 FILLER_258_1427 ();
 b15zdnd00an1n01x5 FILLER_258_1429 ();
 b15zdnd11an1n64x5 FILLER_258_1444 ();
 b15zdnd00an1n02x5 FILLER_258_1508 ();
 b15zdnd00an1n01x5 FILLER_258_1510 ();
 b15zdnd11an1n04x5 FILLER_258_1528 ();
 b15zdnd11an1n16x5 FILLER_258_1537 ();
 b15zdnd11an1n04x5 FILLER_258_1553 ();
 b15zdnd11an1n64x5 FILLER_258_1569 ();
 b15zdnd11an1n64x5 FILLER_258_1633 ();
 b15zdnd11an1n16x5 FILLER_258_1697 ();
 b15zdnd11an1n04x5 FILLER_258_1713 ();
 b15zdnd00an1n02x5 FILLER_258_1717 ();
 b15zdnd00an1n01x5 FILLER_258_1719 ();
 b15zdnd11an1n64x5 FILLER_258_1725 ();
 b15zdnd11an1n08x5 FILLER_258_1789 ();
 b15zdnd11an1n04x5 FILLER_258_1797 ();
 b15zdnd11an1n04x5 FILLER_258_1807 ();
 b15zdnd00an1n02x5 FILLER_258_1811 ();
 b15zdnd11an1n04x5 FILLER_258_1817 ();
 b15zdnd11an1n32x5 FILLER_258_1834 ();
 b15zdnd11an1n08x5 FILLER_258_1866 ();
 b15zdnd11an1n04x5 FILLER_258_1874 ();
 b15zdnd00an1n02x5 FILLER_258_1878 ();
 b15zdnd00an1n01x5 FILLER_258_1880 ();
 b15zdnd11an1n04x5 FILLER_258_1887 ();
 b15zdnd11an1n16x5 FILLER_258_1895 ();
 b15zdnd11an1n08x5 FILLER_258_1911 ();
 b15zdnd00an1n02x5 FILLER_258_1919 ();
 b15zdnd11an1n08x5 FILLER_258_1947 ();
 b15zdnd11an1n04x5 FILLER_258_1955 ();
 b15zdnd00an1n02x5 FILLER_258_1959 ();
 b15zdnd11an1n32x5 FILLER_258_1970 ();
 b15zdnd11an1n16x5 FILLER_258_2002 ();
 b15zdnd11an1n08x5 FILLER_258_2018 ();
 b15zdnd00an1n02x5 FILLER_258_2026 ();
 b15zdnd00an1n01x5 FILLER_258_2028 ();
 b15zdnd11an1n32x5 FILLER_258_2036 ();
 b15zdnd11an1n08x5 FILLER_258_2068 ();
 b15zdnd11an1n32x5 FILLER_258_2095 ();
 b15zdnd11an1n08x5 FILLER_258_2127 ();
 b15zdnd11an1n04x5 FILLER_258_2135 ();
 b15zdnd00an1n01x5 FILLER_258_2139 ();
 b15zdnd11an1n08x5 FILLER_258_2144 ();
 b15zdnd00an1n02x5 FILLER_258_2152 ();
 b15zdnd11an1n64x5 FILLER_258_2162 ();
 b15zdnd11an1n08x5 FILLER_258_2226 ();
 b15zdnd11an1n04x5 FILLER_258_2234 ();
 b15zdnd00an1n02x5 FILLER_258_2238 ();
 b15zdnd00an1n01x5 FILLER_258_2240 ();
 b15zdnd11an1n16x5 FILLER_258_2245 ();
 b15zdnd11an1n08x5 FILLER_258_2261 ();
 b15zdnd11an1n04x5 FILLER_258_2269 ();
 b15zdnd00an1n02x5 FILLER_258_2273 ();
 b15zdnd00an1n01x5 FILLER_258_2275 ();
 b15zdnd11an1n64x5 FILLER_259_0 ();
 b15zdnd11an1n16x5 FILLER_259_64 ();
 b15zdnd11an1n04x5 FILLER_259_80 ();
 b15zdnd00an1n02x5 FILLER_259_84 ();
 b15zdnd11an1n04x5 FILLER_259_93 ();
 b15zdnd11an1n16x5 FILLER_259_101 ();
 b15zdnd11an1n04x5 FILLER_259_117 ();
 b15zdnd11an1n08x5 FILLER_259_131 ();
 b15zdnd11an1n32x5 FILLER_259_147 ();
 b15zdnd11an1n16x5 FILLER_259_189 ();
 b15zdnd11an1n08x5 FILLER_259_205 ();
 b15zdnd11an1n04x5 FILLER_259_213 ();
 b15zdnd00an1n02x5 FILLER_259_217 ();
 b15zdnd11an1n04x5 FILLER_259_233 ();
 b15zdnd11an1n64x5 FILLER_259_242 ();
 b15zdnd11an1n04x5 FILLER_259_306 ();
 b15zdnd00an1n02x5 FILLER_259_310 ();
 b15zdnd11an1n04x5 FILLER_259_318 ();
 b15zdnd00an1n02x5 FILLER_259_322 ();
 b15zdnd00an1n01x5 FILLER_259_324 ();
 b15zdnd11an1n16x5 FILLER_259_329 ();
 b15zdnd00an1n02x5 FILLER_259_345 ();
 b15zdnd11an1n64x5 FILLER_259_356 ();
 b15zdnd11an1n16x5 FILLER_259_425 ();
 b15zdnd00an1n02x5 FILLER_259_441 ();
 b15zdnd11an1n32x5 FILLER_259_462 ();
 b15zdnd11an1n08x5 FILLER_259_494 ();
 b15zdnd11an1n04x5 FILLER_259_502 ();
 b15zdnd00an1n02x5 FILLER_259_506 ();
 b15zdnd00an1n01x5 FILLER_259_508 ();
 b15zdnd11an1n16x5 FILLER_259_519 ();
 b15zdnd11an1n08x5 FILLER_259_535 ();
 b15zdnd00an1n02x5 FILLER_259_543 ();
 b15zdnd11an1n16x5 FILLER_259_552 ();
 b15zdnd11an1n16x5 FILLER_259_578 ();
 b15zdnd00an1n01x5 FILLER_259_594 ();
 b15zdnd11an1n16x5 FILLER_259_606 ();
 b15zdnd00an1n02x5 FILLER_259_622 ();
 b15zdnd11an1n32x5 FILLER_259_634 ();
 b15zdnd11an1n08x5 FILLER_259_666 ();
 b15zdnd00an1n01x5 FILLER_259_674 ();
 b15zdnd11an1n04x5 FILLER_259_680 ();
 b15zdnd00an1n01x5 FILLER_259_684 ();
 b15zdnd11an1n08x5 FILLER_259_698 ();
 b15zdnd11an1n04x5 FILLER_259_706 ();
 b15zdnd00an1n01x5 FILLER_259_710 ();
 b15zdnd11an1n04x5 FILLER_259_715 ();
 b15zdnd11an1n04x5 FILLER_259_739 ();
 b15zdnd11an1n64x5 FILLER_259_753 ();
 b15zdnd11an1n08x5 FILLER_259_822 ();
 b15zdnd11an1n04x5 FILLER_259_830 ();
 b15zdnd00an1n01x5 FILLER_259_834 ();
 b15zdnd11an1n04x5 FILLER_259_860 ();
 b15zdnd00an1n02x5 FILLER_259_864 ();
 b15zdnd00an1n01x5 FILLER_259_866 ();
 b15zdnd11an1n08x5 FILLER_259_889 ();
 b15zdnd00an1n02x5 FILLER_259_897 ();
 b15zdnd00an1n01x5 FILLER_259_899 ();
 b15zdnd11an1n64x5 FILLER_259_918 ();
 b15zdnd00an1n02x5 FILLER_259_982 ();
 b15zdnd11an1n32x5 FILLER_259_994 ();
 b15zdnd11an1n16x5 FILLER_259_1026 ();
 b15zdnd11an1n08x5 FILLER_259_1042 ();
 b15zdnd00an1n02x5 FILLER_259_1050 ();
 b15zdnd00an1n01x5 FILLER_259_1052 ();
 b15zdnd11an1n16x5 FILLER_259_1062 ();
 b15zdnd11an1n08x5 FILLER_259_1078 ();
 b15zdnd11an1n04x5 FILLER_259_1086 ();
 b15zdnd00an1n01x5 FILLER_259_1090 ();
 b15zdnd11an1n32x5 FILLER_259_1102 ();
 b15zdnd11an1n04x5 FILLER_259_1134 ();
 b15zdnd00an1n02x5 FILLER_259_1138 ();
 b15zdnd11an1n32x5 FILLER_259_1152 ();
 b15zdnd11an1n04x5 FILLER_259_1184 ();
 b15zdnd11an1n08x5 FILLER_259_1194 ();
 b15zdnd11an1n04x5 FILLER_259_1202 ();
 b15zdnd11an1n32x5 FILLER_259_1217 ();
 b15zdnd00an1n01x5 FILLER_259_1249 ();
 b15zdnd11an1n04x5 FILLER_259_1271 ();
 b15zdnd11an1n64x5 FILLER_259_1289 ();
 b15zdnd11an1n64x5 FILLER_259_1353 ();
 b15zdnd11an1n16x5 FILLER_259_1417 ();
 b15zdnd00an1n02x5 FILLER_259_1433 ();
 b15zdnd00an1n01x5 FILLER_259_1435 ();
 b15zdnd11an1n08x5 FILLER_259_1441 ();
 b15zdnd00an1n02x5 FILLER_259_1449 ();
 b15zdnd00an1n01x5 FILLER_259_1451 ();
 b15zdnd11an1n04x5 FILLER_259_1472 ();
 b15zdnd11an1n64x5 FILLER_259_1489 ();
 b15zdnd11an1n32x5 FILLER_259_1553 ();
 b15zdnd11an1n08x5 FILLER_259_1585 ();
 b15zdnd11an1n16x5 FILLER_259_1598 ();
 b15zdnd11an1n04x5 FILLER_259_1614 ();
 b15zdnd00an1n01x5 FILLER_259_1618 ();
 b15zdnd11an1n32x5 FILLER_259_1628 ();
 b15zdnd00an1n02x5 FILLER_259_1660 ();
 b15zdnd00an1n01x5 FILLER_259_1662 ();
 b15zdnd11an1n32x5 FILLER_259_1675 ();
 b15zdnd11an1n08x5 FILLER_259_1707 ();
 b15zdnd11an1n04x5 FILLER_259_1715 ();
 b15zdnd00an1n01x5 FILLER_259_1719 ();
 b15zdnd11an1n64x5 FILLER_259_1725 ();
 b15zdnd11an1n64x5 FILLER_259_1789 ();
 b15zdnd11an1n32x5 FILLER_259_1853 ();
 b15zdnd11an1n04x5 FILLER_259_1885 ();
 b15zdnd00an1n01x5 FILLER_259_1889 ();
 b15zdnd11an1n04x5 FILLER_259_1900 ();
 b15zdnd11an1n04x5 FILLER_259_1911 ();
 b15zdnd11an1n16x5 FILLER_259_1920 ();
 b15zdnd11an1n16x5 FILLER_259_1940 ();
 b15zdnd11an1n08x5 FILLER_259_1956 ();
 b15zdnd00an1n02x5 FILLER_259_1964 ();
 b15zdnd11an1n08x5 FILLER_259_1996 ();
 b15zdnd00an1n02x5 FILLER_259_2004 ();
 b15zdnd11an1n08x5 FILLER_259_2016 ();
 b15zdnd11an1n04x5 FILLER_259_2024 ();
 b15zdnd00an1n02x5 FILLER_259_2028 ();
 b15zdnd00an1n01x5 FILLER_259_2030 ();
 b15zdnd11an1n04x5 FILLER_259_2037 ();
 b15zdnd00an1n02x5 FILLER_259_2041 ();
 b15zdnd11an1n32x5 FILLER_259_2053 ();
 b15zdnd11an1n16x5 FILLER_259_2085 ();
 b15zdnd00an1n02x5 FILLER_259_2101 ();
 b15zdnd00an1n01x5 FILLER_259_2103 ();
 b15zdnd11an1n16x5 FILLER_259_2120 ();
 b15zdnd11an1n08x5 FILLER_259_2136 ();
 b15zdnd11an1n04x5 FILLER_259_2144 ();
 b15zdnd00an1n01x5 FILLER_259_2148 ();
 b15zdnd11an1n32x5 FILLER_259_2163 ();
 b15zdnd11an1n16x5 FILLER_259_2195 ();
 b15zdnd00an1n02x5 FILLER_259_2211 ();
 b15zdnd00an1n01x5 FILLER_259_2213 ();
 b15zdnd11an1n04x5 FILLER_259_2219 ();
 b15zdnd11an1n32x5 FILLER_259_2228 ();
 b15zdnd11an1n16x5 FILLER_259_2260 ();
 b15zdnd11an1n08x5 FILLER_259_2276 ();
 b15zdnd11an1n32x5 FILLER_260_8 ();
 b15zdnd11an1n16x5 FILLER_260_40 ();
 b15zdnd11an1n08x5 FILLER_260_56 ();
 b15zdnd11an1n04x5 FILLER_260_64 ();
 b15zdnd11an1n08x5 FILLER_260_80 ();
 b15zdnd00an1n01x5 FILLER_260_88 ();
 b15zdnd11an1n32x5 FILLER_260_96 ();
 b15zdnd11an1n08x5 FILLER_260_128 ();
 b15zdnd00an1n01x5 FILLER_260_136 ();
 b15zdnd11an1n04x5 FILLER_260_141 ();
 b15zdnd11an1n32x5 FILLER_260_149 ();
 b15zdnd11an1n08x5 FILLER_260_195 ();
 b15zdnd11an1n04x5 FILLER_260_203 ();
 b15zdnd00an1n01x5 FILLER_260_207 ();
 b15zdnd11an1n64x5 FILLER_260_216 ();
 b15zdnd11an1n16x5 FILLER_260_280 ();
 b15zdnd11an1n08x5 FILLER_260_296 ();
 b15zdnd11an1n04x5 FILLER_260_304 ();
 b15zdnd00an1n01x5 FILLER_260_308 ();
 b15zdnd11an1n08x5 FILLER_260_314 ();
 b15zdnd11an1n04x5 FILLER_260_322 ();
 b15zdnd00an1n02x5 FILLER_260_326 ();
 b15zdnd11an1n04x5 FILLER_260_338 ();
 b15zdnd11an1n08x5 FILLER_260_346 ();
 b15zdnd00an1n02x5 FILLER_260_354 ();
 b15zdnd11an1n64x5 FILLER_260_369 ();
 b15zdnd11an1n08x5 FILLER_260_433 ();
 b15zdnd00an1n02x5 FILLER_260_441 ();
 b15zdnd11an1n16x5 FILLER_260_447 ();
 b15zdnd11an1n08x5 FILLER_260_463 ();
 b15zdnd00an1n01x5 FILLER_260_471 ();
 b15zdnd11an1n32x5 FILLER_260_478 ();
 b15zdnd11an1n16x5 FILLER_260_510 ();
 b15zdnd11an1n08x5 FILLER_260_526 ();
 b15zdnd00an1n01x5 FILLER_260_534 ();
 b15zdnd11an1n08x5 FILLER_260_539 ();
 b15zdnd00an1n02x5 FILLER_260_547 ();
 b15zdnd11an1n04x5 FILLER_260_565 ();
 b15zdnd11an1n16x5 FILLER_260_574 ();
 b15zdnd00an1n02x5 FILLER_260_590 ();
 b15zdnd11an1n32x5 FILLER_260_602 ();
 b15zdnd11an1n08x5 FILLER_260_634 ();
 b15zdnd00an1n02x5 FILLER_260_642 ();
 b15zdnd00an1n01x5 FILLER_260_644 ();
 b15zdnd11an1n32x5 FILLER_260_652 ();
 b15zdnd11an1n04x5 FILLER_260_684 ();
 b15zdnd11an1n08x5 FILLER_260_694 ();
 b15zdnd00an1n01x5 FILLER_260_702 ();
 b15zdnd11an1n04x5 FILLER_260_707 ();
 b15zdnd00an1n02x5 FILLER_260_716 ();
 b15zdnd11an1n16x5 FILLER_260_726 ();
 b15zdnd11an1n08x5 FILLER_260_742 ();
 b15zdnd00an1n02x5 FILLER_260_750 ();
 b15zdnd00an1n01x5 FILLER_260_752 ();
 b15zdnd11an1n08x5 FILLER_260_761 ();
 b15zdnd00an1n02x5 FILLER_260_769 ();
 b15zdnd00an1n01x5 FILLER_260_771 ();
 b15zdnd11an1n04x5 FILLER_260_776 ();
 b15zdnd11an1n08x5 FILLER_260_787 ();
 b15zdnd11an1n08x5 FILLER_260_805 ();
 b15zdnd11an1n04x5 FILLER_260_813 ();
 b15zdnd00an1n01x5 FILLER_260_817 ();
 b15zdnd11an1n32x5 FILLER_260_828 ();
 b15zdnd11an1n08x5 FILLER_260_860 ();
 b15zdnd11an1n04x5 FILLER_260_899 ();
 b15zdnd11an1n32x5 FILLER_260_921 ();
 b15zdnd00an1n02x5 FILLER_260_953 ();
 b15zdnd11an1n64x5 FILLER_260_962 ();
 b15zdnd11an1n16x5 FILLER_260_1026 ();
 b15zdnd11an1n08x5 FILLER_260_1042 ();
 b15zdnd11an1n04x5 FILLER_260_1050 ();
 b15zdnd11an1n04x5 FILLER_260_1064 ();
 b15zdnd11an1n64x5 FILLER_260_1073 ();
 b15zdnd11an1n64x5 FILLER_260_1137 ();
 b15zdnd11an1n64x5 FILLER_260_1201 ();
 b15zdnd11an1n32x5 FILLER_260_1265 ();
 b15zdnd00an1n01x5 FILLER_260_1297 ();
 b15zdnd11an1n16x5 FILLER_260_1308 ();
 b15zdnd11an1n04x5 FILLER_260_1324 ();
 b15zdnd11an1n04x5 FILLER_260_1335 ();
 b15zdnd11an1n64x5 FILLER_260_1349 ();
 b15zdnd11an1n64x5 FILLER_260_1413 ();
 b15zdnd11an1n08x5 FILLER_260_1477 ();
 b15zdnd11an1n16x5 FILLER_260_1490 ();
 b15zdnd11an1n08x5 FILLER_260_1506 ();
 b15zdnd11an1n04x5 FILLER_260_1514 ();
 b15zdnd00an1n01x5 FILLER_260_1518 ();
 b15zdnd11an1n32x5 FILLER_260_1539 ();
 b15zdnd11an1n08x5 FILLER_260_1571 ();
 b15zdnd00an1n02x5 FILLER_260_1579 ();
 b15zdnd00an1n01x5 FILLER_260_1581 ();
 b15zdnd11an1n08x5 FILLER_260_1588 ();
 b15zdnd11an1n04x5 FILLER_260_1596 ();
 b15zdnd11an1n64x5 FILLER_260_1606 ();
 b15zdnd11an1n32x5 FILLER_260_1670 ();
 b15zdnd11an1n16x5 FILLER_260_1702 ();
 b15zdnd11an1n04x5 FILLER_260_1718 ();
 b15zdnd00an1n02x5 FILLER_260_1722 ();
 b15zdnd11an1n32x5 FILLER_260_1730 ();
 b15zdnd11an1n16x5 FILLER_260_1762 ();
 b15zdnd00an1n01x5 FILLER_260_1778 ();
 b15zdnd11an1n08x5 FILLER_260_1786 ();
 b15zdnd11an1n04x5 FILLER_260_1794 ();
 b15zdnd00an1n02x5 FILLER_260_1798 ();
 b15zdnd11an1n64x5 FILLER_260_1804 ();
 b15zdnd11an1n16x5 FILLER_260_1868 ();
 b15zdnd00an1n02x5 FILLER_260_1884 ();
 b15zdnd00an1n01x5 FILLER_260_1886 ();
 b15zdnd11an1n32x5 FILLER_260_1891 ();
 b15zdnd11an1n08x5 FILLER_260_1923 ();
 b15zdnd11an1n04x5 FILLER_260_1931 ();
 b15zdnd00an1n01x5 FILLER_260_1935 ();
 b15zdnd11an1n16x5 FILLER_260_1948 ();
 b15zdnd11an1n08x5 FILLER_260_1964 ();
 b15zdnd11an1n04x5 FILLER_260_1972 ();
 b15zdnd00an1n01x5 FILLER_260_1976 ();
 b15zdnd11an1n16x5 FILLER_260_1986 ();
 b15zdnd11an1n08x5 FILLER_260_2002 ();
 b15zdnd11an1n04x5 FILLER_260_2010 ();
 b15zdnd00an1n02x5 FILLER_260_2014 ();
 b15zdnd11an1n64x5 FILLER_260_2028 ();
 b15zdnd11an1n32x5 FILLER_260_2092 ();
 b15zdnd11an1n16x5 FILLER_260_2124 ();
 b15zdnd11an1n08x5 FILLER_260_2140 ();
 b15zdnd11an1n04x5 FILLER_260_2148 ();
 b15zdnd00an1n02x5 FILLER_260_2152 ();
 b15zdnd11an1n08x5 FILLER_260_2162 ();
 b15zdnd11an1n04x5 FILLER_260_2170 ();
 b15zdnd00an1n02x5 FILLER_260_2174 ();
 b15zdnd11an1n04x5 FILLER_260_2182 ();
 b15zdnd11an1n08x5 FILLER_260_2191 ();
 b15zdnd11an1n04x5 FILLER_260_2199 ();
 b15zdnd11an1n04x5 FILLER_260_2215 ();
 b15zdnd11an1n08x5 FILLER_260_2223 ();
 b15zdnd00an1n02x5 FILLER_260_2231 ();
 b15zdnd11an1n04x5 FILLER_260_2241 ();
 b15zdnd11an1n16x5 FILLER_260_2250 ();
 b15zdnd11an1n08x5 FILLER_260_2266 ();
 b15zdnd00an1n02x5 FILLER_260_2274 ();
 b15zdnd11an1n32x5 FILLER_261_0 ();
 b15zdnd11an1n04x5 FILLER_261_32 ();
 b15zdnd00an1n02x5 FILLER_261_36 ();
 b15zdnd11an1n16x5 FILLER_261_50 ();
 b15zdnd11an1n32x5 FILLER_261_75 ();
 b15zdnd11an1n08x5 FILLER_261_107 ();
 b15zdnd00an1n02x5 FILLER_261_115 ();
 b15zdnd00an1n01x5 FILLER_261_117 ();
 b15zdnd11an1n08x5 FILLER_261_131 ();
 b15zdnd00an1n02x5 FILLER_261_139 ();
 b15zdnd11an1n64x5 FILLER_261_157 ();
 b15zdnd11an1n32x5 FILLER_261_221 ();
 b15zdnd11an1n16x5 FILLER_261_253 ();
 b15zdnd11an1n04x5 FILLER_261_269 ();
 b15zdnd00an1n02x5 FILLER_261_273 ();
 b15zdnd00an1n01x5 FILLER_261_275 ();
 b15zdnd11an1n64x5 FILLER_261_281 ();
 b15zdnd11an1n64x5 FILLER_261_345 ();
 b15zdnd11an1n16x5 FILLER_261_409 ();
 b15zdnd11an1n04x5 FILLER_261_425 ();
 b15zdnd00an1n01x5 FILLER_261_429 ();
 b15zdnd11an1n32x5 FILLER_261_445 ();
 b15zdnd11an1n08x5 FILLER_261_477 ();
 b15zdnd11an1n04x5 FILLER_261_485 ();
 b15zdnd00an1n01x5 FILLER_261_489 ();
 b15zdnd11an1n16x5 FILLER_261_494 ();
 b15zdnd11an1n04x5 FILLER_261_510 ();
 b15zdnd00an1n01x5 FILLER_261_514 ();
 b15zdnd11an1n04x5 FILLER_261_525 ();
 b15zdnd11an1n16x5 FILLER_261_542 ();
 b15zdnd11an1n04x5 FILLER_261_558 ();
 b15zdnd00an1n01x5 FILLER_261_562 ();
 b15zdnd11an1n32x5 FILLER_261_567 ();
 b15zdnd11an1n16x5 FILLER_261_599 ();
 b15zdnd00an1n01x5 FILLER_261_615 ();
 b15zdnd11an1n64x5 FILLER_261_625 ();
 b15zdnd11an1n16x5 FILLER_261_689 ();
 b15zdnd11an1n08x5 FILLER_261_705 ();
 b15zdnd00an1n01x5 FILLER_261_713 ();
 b15zdnd11an1n64x5 FILLER_261_729 ();
 b15zdnd11an1n32x5 FILLER_261_793 ();
 b15zdnd11an1n08x5 FILLER_261_825 ();
 b15zdnd11an1n64x5 FILLER_261_859 ();
 b15zdnd11an1n64x5 FILLER_261_923 ();
 b15zdnd11an1n32x5 FILLER_261_987 ();
 b15zdnd11an1n08x5 FILLER_261_1019 ();
 b15zdnd00an1n02x5 FILLER_261_1027 ();
 b15zdnd11an1n04x5 FILLER_261_1038 ();
 b15zdnd00an1n01x5 FILLER_261_1042 ();
 b15zdnd11an1n08x5 FILLER_261_1049 ();
 b15zdnd00an1n01x5 FILLER_261_1057 ();
 b15zdnd11an1n08x5 FILLER_261_1063 ();
 b15zdnd00an1n02x5 FILLER_261_1071 ();
 b15zdnd11an1n08x5 FILLER_261_1079 ();
 b15zdnd11an1n04x5 FILLER_261_1087 ();
 b15zdnd00an1n01x5 FILLER_261_1091 ();
 b15zdnd11an1n04x5 FILLER_261_1096 ();
 b15zdnd00an1n01x5 FILLER_261_1100 ();
 b15zdnd11an1n04x5 FILLER_261_1121 ();
 b15zdnd11an1n32x5 FILLER_261_1131 ();
 b15zdnd11an1n16x5 FILLER_261_1163 ();
 b15zdnd00an1n01x5 FILLER_261_1179 ();
 b15zdnd11an1n16x5 FILLER_261_1187 ();
 b15zdnd11an1n08x5 FILLER_261_1203 ();
 b15zdnd11an1n04x5 FILLER_261_1211 ();
 b15zdnd00an1n01x5 FILLER_261_1215 ();
 b15zdnd11an1n64x5 FILLER_261_1222 ();
 b15zdnd11an1n32x5 FILLER_261_1286 ();
 b15zdnd11an1n16x5 FILLER_261_1318 ();
 b15zdnd11an1n08x5 FILLER_261_1334 ();
 b15zdnd11an1n08x5 FILLER_261_1351 ();
 b15zdnd11an1n04x5 FILLER_261_1366 ();
 b15zdnd11an1n64x5 FILLER_261_1374 ();
 b15zdnd11an1n32x5 FILLER_261_1438 ();
 b15zdnd11an1n08x5 FILLER_261_1470 ();
 b15zdnd00an1n02x5 FILLER_261_1478 ();
 b15zdnd00an1n01x5 FILLER_261_1480 ();
 b15zdnd11an1n32x5 FILLER_261_1492 ();
 b15zdnd11an1n04x5 FILLER_261_1524 ();
 b15zdnd00an1n02x5 FILLER_261_1528 ();
 b15zdnd11an1n16x5 FILLER_261_1536 ();
 b15zdnd11an1n08x5 FILLER_261_1552 ();
 b15zdnd11an1n04x5 FILLER_261_1560 ();
 b15zdnd00an1n01x5 FILLER_261_1564 ();
 b15zdnd11an1n04x5 FILLER_261_1572 ();
 b15zdnd00an1n01x5 FILLER_261_1576 ();
 b15zdnd11an1n32x5 FILLER_261_1590 ();
 b15zdnd11an1n04x5 FILLER_261_1622 ();
 b15zdnd00an1n01x5 FILLER_261_1626 ();
 b15zdnd11an1n16x5 FILLER_261_1637 ();
 b15zdnd11an1n04x5 FILLER_261_1653 ();
 b15zdnd11an1n16x5 FILLER_261_1664 ();
 b15zdnd11an1n04x5 FILLER_261_1680 ();
 b15zdnd11an1n04x5 FILLER_261_1715 ();
 b15zdnd11an1n04x5 FILLER_261_1728 ();
 b15zdnd00an1n02x5 FILLER_261_1732 ();
 b15zdnd11an1n64x5 FILLER_261_1742 ();
 b15zdnd11an1n64x5 FILLER_261_1806 ();
 b15zdnd11an1n64x5 FILLER_261_1870 ();
 b15zdnd00an1n01x5 FILLER_261_1934 ();
 b15zdnd11an1n04x5 FILLER_261_1957 ();
 b15zdnd00an1n02x5 FILLER_261_1961 ();
 b15zdnd00an1n01x5 FILLER_261_1963 ();
 b15zdnd11an1n16x5 FILLER_261_1976 ();
 b15zdnd11an1n08x5 FILLER_261_1992 ();
 b15zdnd11an1n04x5 FILLER_261_2000 ();
 b15zdnd00an1n01x5 FILLER_261_2004 ();
 b15zdnd11an1n32x5 FILLER_261_2012 ();
 b15zdnd11an1n16x5 FILLER_261_2044 ();
 b15zdnd11an1n08x5 FILLER_261_2060 ();
 b15zdnd11an1n04x5 FILLER_261_2068 ();
 b15zdnd00an1n02x5 FILLER_261_2072 ();
 b15zdnd11an1n16x5 FILLER_261_2084 ();
 b15zdnd11an1n08x5 FILLER_261_2100 ();
 b15zdnd11an1n04x5 FILLER_261_2108 ();
 b15zdnd11an1n16x5 FILLER_261_2122 ();
 b15zdnd00an1n02x5 FILLER_261_2138 ();
 b15zdnd11an1n04x5 FILLER_261_2144 ();
 b15zdnd11an1n64x5 FILLER_261_2159 ();
 b15zdnd11an1n32x5 FILLER_261_2223 ();
 b15zdnd11an1n16x5 FILLER_261_2255 ();
 b15zdnd11an1n08x5 FILLER_261_2271 ();
 b15zdnd11an1n04x5 FILLER_261_2279 ();
 b15zdnd00an1n01x5 FILLER_261_2283 ();
 b15zdnd11an1n32x5 FILLER_262_8 ();
 b15zdnd11an1n04x5 FILLER_262_40 ();
 b15zdnd00an1n02x5 FILLER_262_44 ();
 b15zdnd11an1n04x5 FILLER_262_58 ();
 b15zdnd11an1n64x5 FILLER_262_72 ();
 b15zdnd11an1n08x5 FILLER_262_136 ();
 b15zdnd11an1n04x5 FILLER_262_144 ();
 b15zdnd00an1n02x5 FILLER_262_148 ();
 b15zdnd00an1n01x5 FILLER_262_150 ();
 b15zdnd11an1n04x5 FILLER_262_172 ();
 b15zdnd00an1n02x5 FILLER_262_176 ();
 b15zdnd00an1n01x5 FILLER_262_178 ();
 b15zdnd11an1n16x5 FILLER_262_185 ();
 b15zdnd11an1n08x5 FILLER_262_201 ();
 b15zdnd11an1n32x5 FILLER_262_214 ();
 b15zdnd11an1n16x5 FILLER_262_246 ();
 b15zdnd11an1n08x5 FILLER_262_262 ();
 b15zdnd00an1n02x5 FILLER_262_270 ();
 b15zdnd00an1n01x5 FILLER_262_272 ();
 b15zdnd11an1n04x5 FILLER_262_279 ();
 b15zdnd00an1n02x5 FILLER_262_283 ();
 b15zdnd00an1n01x5 FILLER_262_285 ();
 b15zdnd11an1n64x5 FILLER_262_291 ();
 b15zdnd11an1n64x5 FILLER_262_355 ();
 b15zdnd11an1n64x5 FILLER_262_419 ();
 b15zdnd11an1n32x5 FILLER_262_483 ();
 b15zdnd11an1n04x5 FILLER_262_515 ();
 b15zdnd00an1n01x5 FILLER_262_519 ();
 b15zdnd11an1n16x5 FILLER_262_527 ();
 b15zdnd11an1n08x5 FILLER_262_543 ();
 b15zdnd00an1n02x5 FILLER_262_551 ();
 b15zdnd11an1n16x5 FILLER_262_583 ();
 b15zdnd11an1n08x5 FILLER_262_599 ();
 b15zdnd11an1n04x5 FILLER_262_607 ();
 b15zdnd00an1n02x5 FILLER_262_611 ();
 b15zdnd11an1n64x5 FILLER_262_619 ();
 b15zdnd11an1n32x5 FILLER_262_683 ();
 b15zdnd00an1n02x5 FILLER_262_715 ();
 b15zdnd00an1n01x5 FILLER_262_717 ();
 b15zdnd11an1n04x5 FILLER_262_726 ();
 b15zdnd00an1n02x5 FILLER_262_730 ();
 b15zdnd00an1n01x5 FILLER_262_732 ();
 b15zdnd11an1n64x5 FILLER_262_749 ();
 b15zdnd00an1n02x5 FILLER_262_813 ();
 b15zdnd11an1n64x5 FILLER_262_821 ();
 b15zdnd11an1n64x5 FILLER_262_885 ();
 b15zdnd11an1n32x5 FILLER_262_949 ();
 b15zdnd11an1n08x5 FILLER_262_981 ();
 b15zdnd11an1n04x5 FILLER_262_989 ();
 b15zdnd11an1n04x5 FILLER_262_999 ();
 b15zdnd00an1n02x5 FILLER_262_1003 ();
 b15zdnd11an1n32x5 FILLER_262_1011 ();
 b15zdnd11an1n08x5 FILLER_262_1043 ();
 b15zdnd00an1n01x5 FILLER_262_1051 ();
 b15zdnd11an1n32x5 FILLER_262_1057 ();
 b15zdnd11an1n04x5 FILLER_262_1089 ();
 b15zdnd00an1n01x5 FILLER_262_1093 ();
 b15zdnd11an1n32x5 FILLER_262_1100 ();
 b15zdnd11an1n16x5 FILLER_262_1132 ();
 b15zdnd00an1n02x5 FILLER_262_1148 ();
 b15zdnd00an1n01x5 FILLER_262_1150 ();
 b15zdnd11an1n16x5 FILLER_262_1158 ();
 b15zdnd00an1n02x5 FILLER_262_1174 ();
 b15zdnd00an1n01x5 FILLER_262_1176 ();
 b15zdnd11an1n04x5 FILLER_262_1189 ();
 b15zdnd11an1n64x5 FILLER_262_1197 ();
 b15zdnd00an1n02x5 FILLER_262_1261 ();
 b15zdnd11an1n04x5 FILLER_262_1277 ();
 b15zdnd11an1n08x5 FILLER_262_1286 ();
 b15zdnd00an1n02x5 FILLER_262_1294 ();
 b15zdnd00an1n01x5 FILLER_262_1296 ();
 b15zdnd11an1n04x5 FILLER_262_1323 ();
 b15zdnd11an1n04x5 FILLER_262_1336 ();
 b15zdnd11an1n64x5 FILLER_262_1350 ();
 b15zdnd11an1n64x5 FILLER_262_1414 ();
 b15zdnd11an1n16x5 FILLER_262_1478 ();
 b15zdnd11an1n04x5 FILLER_262_1494 ();
 b15zdnd00an1n01x5 FILLER_262_1498 ();
 b15zdnd11an1n16x5 FILLER_262_1506 ();
 b15zdnd11an1n08x5 FILLER_262_1522 ();
 b15zdnd11an1n04x5 FILLER_262_1530 ();
 b15zdnd11an1n16x5 FILLER_262_1544 ();
 b15zdnd00an1n02x5 FILLER_262_1560 ();
 b15zdnd11an1n16x5 FILLER_262_1568 ();
 b15zdnd11an1n08x5 FILLER_262_1584 ();
 b15zdnd11an1n04x5 FILLER_262_1592 ();
 b15zdnd11an1n16x5 FILLER_262_1609 ();
 b15zdnd00an1n01x5 FILLER_262_1625 ();
 b15zdnd11an1n32x5 FILLER_262_1636 ();
 b15zdnd11an1n08x5 FILLER_262_1668 ();
 b15zdnd00an1n02x5 FILLER_262_1676 ();
 b15zdnd11an1n04x5 FILLER_262_1686 ();
 b15zdnd11an1n16x5 FILLER_262_1711 ();
 b15zdnd11an1n08x5 FILLER_262_1727 ();
 b15zdnd11an1n04x5 FILLER_262_1735 ();
 b15zdnd00an1n02x5 FILLER_262_1739 ();
 b15zdnd11an1n04x5 FILLER_262_1747 ();
 b15zdnd11an1n04x5 FILLER_262_1760 ();
 b15zdnd00an1n02x5 FILLER_262_1764 ();
 b15zdnd00an1n01x5 FILLER_262_1766 ();
 b15zdnd11an1n16x5 FILLER_262_1781 ();
 b15zdnd00an1n01x5 FILLER_262_1797 ();
 b15zdnd11an1n64x5 FILLER_262_1806 ();
 b15zdnd11an1n08x5 FILLER_262_1870 ();
 b15zdnd11an1n04x5 FILLER_262_1878 ();
 b15zdnd00an1n02x5 FILLER_262_1882 ();
 b15zdnd00an1n01x5 FILLER_262_1884 ();
 b15zdnd11an1n16x5 FILLER_262_1889 ();
 b15zdnd00an1n02x5 FILLER_262_1905 ();
 b15zdnd11an1n04x5 FILLER_262_1913 ();
 b15zdnd11an1n04x5 FILLER_262_1921 ();
 b15zdnd00an1n02x5 FILLER_262_1925 ();
 b15zdnd00an1n01x5 FILLER_262_1927 ();
 b15zdnd11an1n64x5 FILLER_262_1935 ();
 b15zdnd11an1n04x5 FILLER_262_1999 ();
 b15zdnd00an1n01x5 FILLER_262_2003 ();
 b15zdnd11an1n64x5 FILLER_262_2011 ();
 b15zdnd11an1n08x5 FILLER_262_2082 ();
 b15zdnd11an1n04x5 FILLER_262_2090 ();
 b15zdnd00an1n01x5 FILLER_262_2094 ();
 b15zdnd11an1n04x5 FILLER_262_2100 ();
 b15zdnd00an1n02x5 FILLER_262_2104 ();
 b15zdnd00an1n01x5 FILLER_262_2106 ();
 b15zdnd11an1n04x5 FILLER_262_2113 ();
 b15zdnd11an1n16x5 FILLER_262_2124 ();
 b15zdnd11an1n04x5 FILLER_262_2140 ();
 b15zdnd00an1n02x5 FILLER_262_2144 ();
 b15zdnd00an1n02x5 FILLER_262_2151 ();
 b15zdnd00an1n01x5 FILLER_262_2153 ();
 b15zdnd11an1n16x5 FILLER_262_2162 ();
 b15zdnd11an1n08x5 FILLER_262_2178 ();
 b15zdnd11an1n04x5 FILLER_262_2186 ();
 b15zdnd00an1n01x5 FILLER_262_2190 ();
 b15zdnd11an1n08x5 FILLER_262_2196 ();
 b15zdnd11an1n04x5 FILLER_262_2204 ();
 b15zdnd00an1n01x5 FILLER_262_2208 ();
 b15zdnd11an1n08x5 FILLER_262_2216 ();
 b15zdnd11an1n04x5 FILLER_262_2224 ();
 b15zdnd00an1n02x5 FILLER_262_2228 ();
 b15zdnd00an1n01x5 FILLER_262_2230 ();
 b15zdnd11an1n32x5 FILLER_262_2237 ();
 b15zdnd11an1n04x5 FILLER_262_2269 ();
 b15zdnd00an1n02x5 FILLER_262_2273 ();
 b15zdnd00an1n01x5 FILLER_262_2275 ();
 b15zdnd11an1n64x5 FILLER_263_0 ();
 b15zdnd11an1n16x5 FILLER_263_68 ();
 b15zdnd11an1n08x5 FILLER_263_84 ();
 b15zdnd00an1n02x5 FILLER_263_92 ();
 b15zdnd00an1n01x5 FILLER_263_94 ();
 b15zdnd11an1n64x5 FILLER_263_101 ();
 b15zdnd11an1n32x5 FILLER_263_165 ();
 b15zdnd11an1n08x5 FILLER_263_197 ();
 b15zdnd11an1n04x5 FILLER_263_205 ();
 b15zdnd00an1n02x5 FILLER_263_209 ();
 b15zdnd00an1n01x5 FILLER_263_211 ();
 b15zdnd11an1n16x5 FILLER_263_218 ();
 b15zdnd11an1n08x5 FILLER_263_234 ();
 b15zdnd11an1n04x5 FILLER_263_242 ();
 b15zdnd00an1n02x5 FILLER_263_246 ();
 b15zdnd11an1n32x5 FILLER_263_253 ();
 b15zdnd11an1n04x5 FILLER_263_285 ();
 b15zdnd00an1n02x5 FILLER_263_289 ();
 b15zdnd00an1n01x5 FILLER_263_291 ();
 b15zdnd11an1n64x5 FILLER_263_301 ();
 b15zdnd11an1n64x5 FILLER_263_365 ();
 b15zdnd11an1n08x5 FILLER_263_429 ();
 b15zdnd11an1n16x5 FILLER_263_449 ();
 b15zdnd11an1n04x5 FILLER_263_473 ();
 b15zdnd11an1n64x5 FILLER_263_481 ();
 b15zdnd11an1n16x5 FILLER_263_545 ();
 b15zdnd11an1n08x5 FILLER_263_561 ();
 b15zdnd11an1n04x5 FILLER_263_569 ();
 b15zdnd11an1n32x5 FILLER_263_583 ();
 b15zdnd11an1n04x5 FILLER_263_615 ();
 b15zdnd11an1n16x5 FILLER_263_629 ();
 b15zdnd00an1n02x5 FILLER_263_645 ();
 b15zdnd11an1n08x5 FILLER_263_657 ();
 b15zdnd11an1n04x5 FILLER_263_665 ();
 b15zdnd11an1n16x5 FILLER_263_689 ();
 b15zdnd11an1n08x5 FILLER_263_705 ();
 b15zdnd00an1n02x5 FILLER_263_713 ();
 b15zdnd00an1n01x5 FILLER_263_715 ();
 b15zdnd11an1n16x5 FILLER_263_730 ();
 b15zdnd11an1n08x5 FILLER_263_746 ();
 b15zdnd11an1n04x5 FILLER_263_754 ();
 b15zdnd11an1n04x5 FILLER_263_762 ();
 b15zdnd00an1n02x5 FILLER_263_766 ();
 b15zdnd11an1n16x5 FILLER_263_783 ();
 b15zdnd11an1n08x5 FILLER_263_799 ();
 b15zdnd11an1n04x5 FILLER_263_807 ();
 b15zdnd00an1n02x5 FILLER_263_811 ();
 b15zdnd00an1n01x5 FILLER_263_813 ();
 b15zdnd11an1n64x5 FILLER_263_820 ();
 b15zdnd11an1n16x5 FILLER_263_884 ();
 b15zdnd00an1n02x5 FILLER_263_900 ();
 b15zdnd00an1n01x5 FILLER_263_902 ();
 b15zdnd11an1n32x5 FILLER_263_913 ();
 b15zdnd11an1n08x5 FILLER_263_945 ();
 b15zdnd11an1n04x5 FILLER_263_953 ();
 b15zdnd11an1n32x5 FILLER_263_975 ();
 b15zdnd11an1n08x5 FILLER_263_1007 ();
 b15zdnd00an1n01x5 FILLER_263_1015 ();
 b15zdnd11an1n32x5 FILLER_263_1021 ();
 b15zdnd11an1n08x5 FILLER_263_1053 ();
 b15zdnd11an1n04x5 FILLER_263_1061 ();
 b15zdnd00an1n02x5 FILLER_263_1065 ();
 b15zdnd11an1n16x5 FILLER_263_1073 ();
 b15zdnd11an1n04x5 FILLER_263_1089 ();
 b15zdnd00an1n01x5 FILLER_263_1093 ();
 b15zdnd11an1n32x5 FILLER_263_1100 ();
 b15zdnd00an1n02x5 FILLER_263_1132 ();
 b15zdnd11an1n08x5 FILLER_263_1140 ();
 b15zdnd00an1n01x5 FILLER_263_1148 ();
 b15zdnd11an1n16x5 FILLER_263_1165 ();
 b15zdnd11an1n08x5 FILLER_263_1181 ();
 b15zdnd11an1n04x5 FILLER_263_1189 ();
 b15zdnd00an1n02x5 FILLER_263_1193 ();
 b15zdnd11an1n04x5 FILLER_263_1207 ();
 b15zdnd00an1n01x5 FILLER_263_1211 ();
 b15zdnd11an1n16x5 FILLER_263_1217 ();
 b15zdnd11an1n08x5 FILLER_263_1233 ();
 b15zdnd00an1n02x5 FILLER_263_1241 ();
 b15zdnd00an1n01x5 FILLER_263_1243 ();
 b15zdnd11an1n04x5 FILLER_263_1251 ();
 b15zdnd11an1n04x5 FILLER_263_1272 ();
 b15zdnd00an1n02x5 FILLER_263_1276 ();
 b15zdnd11an1n32x5 FILLER_263_1290 ();
 b15zdnd11an1n08x5 FILLER_263_1322 ();
 b15zdnd00an1n02x5 FILLER_263_1330 ();
 b15zdnd00an1n01x5 FILLER_263_1332 ();
 b15zdnd11an1n04x5 FILLER_263_1342 ();
 b15zdnd00an1n01x5 FILLER_263_1346 ();
 b15zdnd11an1n04x5 FILLER_263_1355 ();
 b15zdnd11an1n64x5 FILLER_263_1368 ();
 b15zdnd11an1n04x5 FILLER_263_1432 ();
 b15zdnd00an1n01x5 FILLER_263_1436 ();
 b15zdnd11an1n04x5 FILLER_263_1453 ();
 b15zdnd11an1n04x5 FILLER_263_1482 ();
 b15zdnd11an1n16x5 FILLER_263_1491 ();
 b15zdnd11an1n04x5 FILLER_263_1507 ();
 b15zdnd11an1n04x5 FILLER_263_1532 ();
 b15zdnd11an1n16x5 FILLER_263_1541 ();
 b15zdnd00an1n02x5 FILLER_263_1557 ();
 b15zdnd11an1n32x5 FILLER_263_1565 ();
 b15zdnd00an1n02x5 FILLER_263_1597 ();
 b15zdnd11an1n64x5 FILLER_263_1614 ();
 b15zdnd11an1n64x5 FILLER_263_1678 ();
 b15zdnd11an1n32x5 FILLER_263_1742 ();
 b15zdnd11an1n16x5 FILLER_263_1774 ();
 b15zdnd11an1n08x5 FILLER_263_1790 ();
 b15zdnd11an1n32x5 FILLER_263_1811 ();
 b15zdnd11an1n16x5 FILLER_263_1843 ();
 b15zdnd11an1n08x5 FILLER_263_1859 ();
 b15zdnd11an1n04x5 FILLER_263_1867 ();
 b15zdnd00an1n02x5 FILLER_263_1871 ();
 b15zdnd11an1n04x5 FILLER_263_1882 ();
 b15zdnd11an1n16x5 FILLER_263_1892 ();
 b15zdnd11an1n08x5 FILLER_263_1908 ();
 b15zdnd00an1n01x5 FILLER_263_1916 ();
 b15zdnd11an1n64x5 FILLER_263_1933 ();
 b15zdnd00an1n02x5 FILLER_263_1997 ();
 b15zdnd00an1n01x5 FILLER_263_1999 ();
 b15zdnd11an1n16x5 FILLER_263_2014 ();
 b15zdnd11an1n04x5 FILLER_263_2030 ();
 b15zdnd00an1n01x5 FILLER_263_2034 ();
 b15zdnd11an1n16x5 FILLER_263_2041 ();
 b15zdnd11an1n08x5 FILLER_263_2057 ();
 b15zdnd11an1n04x5 FILLER_263_2065 ();
 b15zdnd11an1n08x5 FILLER_263_2079 ();
 b15zdnd11an1n64x5 FILLER_263_2102 ();
 b15zdnd11an1n16x5 FILLER_263_2166 ();
 b15zdnd00an1n02x5 FILLER_263_2182 ();
 b15zdnd00an1n01x5 FILLER_263_2184 ();
 b15zdnd11an1n32x5 FILLER_263_2191 ();
 b15zdnd00an1n02x5 FILLER_263_2223 ();
 b15zdnd11an1n32x5 FILLER_263_2233 ();
 b15zdnd11an1n16x5 FILLER_263_2265 ();
 b15zdnd00an1n02x5 FILLER_263_2281 ();
 b15zdnd00an1n01x5 FILLER_263_2283 ();
 b15zdnd11an1n64x5 FILLER_264_8 ();
 b15zdnd11an1n08x5 FILLER_264_72 ();
 b15zdnd11an1n04x5 FILLER_264_80 ();
 b15zdnd11an1n08x5 FILLER_264_96 ();
 b15zdnd00an1n02x5 FILLER_264_104 ();
 b15zdnd00an1n01x5 FILLER_264_106 ();
 b15zdnd11an1n32x5 FILLER_264_121 ();
 b15zdnd11an1n16x5 FILLER_264_153 ();
 b15zdnd00an1n02x5 FILLER_264_169 ();
 b15zdnd11an1n32x5 FILLER_264_183 ();
 b15zdnd11an1n08x5 FILLER_264_215 ();
 b15zdnd11an1n04x5 FILLER_264_223 ();
 b15zdnd11an1n04x5 FILLER_264_244 ();
 b15zdnd00an1n01x5 FILLER_264_248 ();
 b15zdnd11an1n04x5 FILLER_264_253 ();
 b15zdnd11an1n08x5 FILLER_264_261 ();
 b15zdnd11an1n04x5 FILLER_264_269 ();
 b15zdnd00an1n01x5 FILLER_264_273 ();
 b15zdnd11an1n08x5 FILLER_264_281 ();
 b15zdnd11an1n04x5 FILLER_264_289 ();
 b15zdnd00an1n02x5 FILLER_264_293 ();
 b15zdnd11an1n08x5 FILLER_264_301 ();
 b15zdnd00an1n02x5 FILLER_264_309 ();
 b15zdnd11an1n04x5 FILLER_264_317 ();
 b15zdnd11an1n08x5 FILLER_264_331 ();
 b15zdnd00an1n02x5 FILLER_264_339 ();
 b15zdnd00an1n01x5 FILLER_264_341 ();
 b15zdnd11an1n64x5 FILLER_264_348 ();
 b15zdnd11an1n64x5 FILLER_264_412 ();
 b15zdnd11an1n16x5 FILLER_264_476 ();
 b15zdnd11an1n08x5 FILLER_264_492 ();
 b15zdnd00an1n02x5 FILLER_264_500 ();
 b15zdnd00an1n01x5 FILLER_264_502 ();
 b15zdnd11an1n64x5 FILLER_264_511 ();
 b15zdnd00an1n02x5 FILLER_264_575 ();
 b15zdnd11an1n04x5 FILLER_264_581 ();
 b15zdnd00an1n02x5 FILLER_264_585 ();
 b15zdnd00an1n01x5 FILLER_264_587 ();
 b15zdnd11an1n32x5 FILLER_264_601 ();
 b15zdnd11an1n16x5 FILLER_264_633 ();
 b15zdnd11an1n04x5 FILLER_264_649 ();
 b15zdnd00an1n01x5 FILLER_264_653 ();
 b15zdnd11an1n08x5 FILLER_264_686 ();
 b15zdnd11an1n16x5 FILLER_264_701 ();
 b15zdnd00an1n01x5 FILLER_264_717 ();
 b15zdnd11an1n16x5 FILLER_264_726 ();
 b15zdnd11an1n04x5 FILLER_264_742 ();
 b15zdnd11an1n32x5 FILLER_264_751 ();
 b15zdnd11an1n16x5 FILLER_264_783 ();
 b15zdnd11an1n08x5 FILLER_264_799 ();
 b15zdnd11an1n04x5 FILLER_264_807 ();
 b15zdnd00an1n01x5 FILLER_264_811 ();
 b15zdnd11an1n64x5 FILLER_264_816 ();
 b15zdnd11an1n64x5 FILLER_264_880 ();
 b15zdnd11an1n16x5 FILLER_264_944 ();
 b15zdnd00an1n02x5 FILLER_264_960 ();
 b15zdnd00an1n01x5 FILLER_264_962 ();
 b15zdnd11an1n04x5 FILLER_264_977 ();
 b15zdnd11an1n04x5 FILLER_264_999 ();
 b15zdnd11an1n32x5 FILLER_264_1015 ();
 b15zdnd11an1n16x5 FILLER_264_1047 ();
 b15zdnd11an1n04x5 FILLER_264_1063 ();
 b15zdnd11an1n32x5 FILLER_264_1072 ();
 b15zdnd11an1n16x5 FILLER_264_1104 ();
 b15zdnd11an1n08x5 FILLER_264_1120 ();
 b15zdnd11an1n64x5 FILLER_264_1134 ();
 b15zdnd11an1n16x5 FILLER_264_1219 ();
 b15zdnd11an1n08x5 FILLER_264_1235 ();
 b15zdnd00an1n02x5 FILLER_264_1243 ();
 b15zdnd11an1n04x5 FILLER_264_1249 ();
 b15zdnd11an1n64x5 FILLER_264_1258 ();
 b15zdnd11an1n04x5 FILLER_264_1322 ();
 b15zdnd00an1n02x5 FILLER_264_1326 ();
 b15zdnd11an1n16x5 FILLER_264_1350 ();
 b15zdnd11an1n08x5 FILLER_264_1366 ();
 b15zdnd11an1n04x5 FILLER_264_1374 ();
 b15zdnd00an1n02x5 FILLER_264_1378 ();
 b15zdnd00an1n01x5 FILLER_264_1380 ();
 b15zdnd11an1n16x5 FILLER_264_1407 ();
 b15zdnd00an1n02x5 FILLER_264_1423 ();
 b15zdnd00an1n01x5 FILLER_264_1425 ();
 b15zdnd11an1n16x5 FILLER_264_1445 ();
 b15zdnd11an1n08x5 FILLER_264_1461 ();
 b15zdnd00an1n01x5 FILLER_264_1469 ();
 b15zdnd11an1n04x5 FILLER_264_1478 ();
 b15zdnd11an1n04x5 FILLER_264_1496 ();
 b15zdnd11an1n16x5 FILLER_264_1509 ();
 b15zdnd11an1n08x5 FILLER_264_1525 ();
 b15zdnd00an1n02x5 FILLER_264_1533 ();
 b15zdnd00an1n01x5 FILLER_264_1535 ();
 b15zdnd11an1n16x5 FILLER_264_1541 ();
 b15zdnd11an1n16x5 FILLER_264_1562 ();
 b15zdnd11an1n08x5 FILLER_264_1578 ();
 b15zdnd11an1n04x5 FILLER_264_1586 ();
 b15zdnd11an1n04x5 FILLER_264_1595 ();
 b15zdnd11an1n08x5 FILLER_264_1604 ();
 b15zdnd00an1n02x5 FILLER_264_1612 ();
 b15zdnd11an1n32x5 FILLER_264_1622 ();
 b15zdnd11an1n16x5 FILLER_264_1654 ();
 b15zdnd11an1n32x5 FILLER_264_1682 ();
 b15zdnd11an1n04x5 FILLER_264_1723 ();
 b15zdnd11an1n16x5 FILLER_264_1736 ();
 b15zdnd11an1n08x5 FILLER_264_1752 ();
 b15zdnd11an1n04x5 FILLER_264_1776 ();
 b15zdnd00an1n01x5 FILLER_264_1780 ();
 b15zdnd11an1n04x5 FILLER_264_1788 ();
 b15zdnd11an1n08x5 FILLER_264_1799 ();
 b15zdnd00an1n02x5 FILLER_264_1807 ();
 b15zdnd11an1n32x5 FILLER_264_1827 ();
 b15zdnd11an1n08x5 FILLER_264_1859 ();
 b15zdnd11an1n04x5 FILLER_264_1867 ();
 b15zdnd00an1n02x5 FILLER_264_1871 ();
 b15zdnd00an1n01x5 FILLER_264_1873 ();
 b15zdnd11an1n32x5 FILLER_264_1906 ();
 b15zdnd00an1n02x5 FILLER_264_1938 ();
 b15zdnd11an1n08x5 FILLER_264_1966 ();
 b15zdnd00an1n02x5 FILLER_264_1974 ();
 b15zdnd11an1n08x5 FILLER_264_1992 ();
 b15zdnd11an1n04x5 FILLER_264_2000 ();
 b15zdnd00an1n01x5 FILLER_264_2004 ();
 b15zdnd11an1n16x5 FILLER_264_2009 ();
 b15zdnd11an1n08x5 FILLER_264_2025 ();
 b15zdnd00an1n02x5 FILLER_264_2033 ();
 b15zdnd00an1n01x5 FILLER_264_2035 ();
 b15zdnd11an1n04x5 FILLER_264_2042 ();
 b15zdnd00an1n02x5 FILLER_264_2046 ();
 b15zdnd00an1n01x5 FILLER_264_2048 ();
 b15zdnd11an1n64x5 FILLER_264_2056 ();
 b15zdnd11an1n32x5 FILLER_264_2120 ();
 b15zdnd00an1n02x5 FILLER_264_2152 ();
 b15zdnd00an1n02x5 FILLER_264_2162 ();
 b15zdnd11an1n08x5 FILLER_264_2170 ();
 b15zdnd11an1n04x5 FILLER_264_2178 ();
 b15zdnd00an1n02x5 FILLER_264_2182 ();
 b15zdnd11an1n16x5 FILLER_264_2189 ();
 b15zdnd00an1n02x5 FILLER_264_2205 ();
 b15zdnd00an1n01x5 FILLER_264_2207 ();
 b15zdnd11an1n08x5 FILLER_264_2213 ();
 b15zdnd11an1n04x5 FILLER_264_2221 ();
 b15zdnd00an1n02x5 FILLER_264_2225 ();
 b15zdnd00an1n01x5 FILLER_264_2227 ();
 b15zdnd11an1n04x5 FILLER_264_2233 ();
 b15zdnd11an1n16x5 FILLER_264_2246 ();
 b15zdnd11an1n08x5 FILLER_264_2262 ();
 b15zdnd11an1n04x5 FILLER_264_2270 ();
 b15zdnd00an1n02x5 FILLER_264_2274 ();
 b15zdnd11an1n32x5 FILLER_265_0 ();
 b15zdnd11an1n16x5 FILLER_265_32 ();
 b15zdnd11an1n08x5 FILLER_265_48 ();
 b15zdnd11an1n04x5 FILLER_265_56 ();
 b15zdnd11an1n32x5 FILLER_265_69 ();
 b15zdnd11an1n08x5 FILLER_265_106 ();
 b15zdnd11an1n04x5 FILLER_265_114 ();
 b15zdnd00an1n02x5 FILLER_265_118 ();
 b15zdnd11an1n08x5 FILLER_265_125 ();
 b15zdnd00an1n02x5 FILLER_265_133 ();
 b15zdnd11an1n16x5 FILLER_265_147 ();
 b15zdnd00an1n01x5 FILLER_265_163 ();
 b15zdnd11an1n04x5 FILLER_265_168 ();
 b15zdnd11an1n32x5 FILLER_265_180 ();
 b15zdnd00an1n02x5 FILLER_265_212 ();
 b15zdnd00an1n01x5 FILLER_265_214 ();
 b15zdnd11an1n08x5 FILLER_265_220 ();
 b15zdnd11an1n04x5 FILLER_265_228 ();
 b15zdnd00an1n02x5 FILLER_265_232 ();
 b15zdnd00an1n01x5 FILLER_265_234 ();
 b15zdnd11an1n04x5 FILLER_265_247 ();
 b15zdnd11an1n32x5 FILLER_265_257 ();
 b15zdnd00an1n02x5 FILLER_265_289 ();
 b15zdnd00an1n01x5 FILLER_265_291 ();
 b15zdnd11an1n32x5 FILLER_265_297 ();
 b15zdnd11an1n08x5 FILLER_265_329 ();
 b15zdnd00an1n01x5 FILLER_265_337 ();
 b15zdnd11an1n16x5 FILLER_265_343 ();
 b15zdnd11an1n08x5 FILLER_265_359 ();
 b15zdnd00an1n01x5 FILLER_265_367 ();
 b15zdnd11an1n32x5 FILLER_265_378 ();
 b15zdnd11an1n08x5 FILLER_265_410 ();
 b15zdnd11an1n04x5 FILLER_265_418 ();
 b15zdnd00an1n02x5 FILLER_265_422 ();
 b15zdnd00an1n01x5 FILLER_265_424 ();
 b15zdnd11an1n04x5 FILLER_265_429 ();
 b15zdnd11an1n04x5 FILLER_265_447 ();
 b15zdnd11an1n08x5 FILLER_265_461 ();
 b15zdnd11an1n04x5 FILLER_265_469 ();
 b15zdnd00an1n02x5 FILLER_265_473 ();
 b15zdnd11an1n04x5 FILLER_265_487 ();
 b15zdnd11an1n08x5 FILLER_265_495 ();
 b15zdnd00an1n02x5 FILLER_265_503 ();
 b15zdnd00an1n01x5 FILLER_265_505 ();
 b15zdnd11an1n16x5 FILLER_265_511 ();
 b15zdnd11an1n08x5 FILLER_265_527 ();
 b15zdnd11an1n04x5 FILLER_265_535 ();
 b15zdnd00an1n01x5 FILLER_265_539 ();
 b15zdnd11an1n32x5 FILLER_265_545 ();
 b15zdnd11an1n16x5 FILLER_265_577 ();
 b15zdnd11an1n08x5 FILLER_265_593 ();
 b15zdnd11an1n04x5 FILLER_265_601 ();
 b15zdnd00an1n02x5 FILLER_265_605 ();
 b15zdnd00an1n01x5 FILLER_265_607 ();
 b15zdnd11an1n04x5 FILLER_265_612 ();
 b15zdnd11an1n64x5 FILLER_265_621 ();
 b15zdnd00an1n01x5 FILLER_265_685 ();
 b15zdnd11an1n64x5 FILLER_265_699 ();
 b15zdnd11an1n16x5 FILLER_265_763 ();
 b15zdnd11an1n08x5 FILLER_265_779 ();
 b15zdnd11an1n04x5 FILLER_265_787 ();
 b15zdnd11an1n32x5 FILLER_265_796 ();
 b15zdnd11an1n08x5 FILLER_265_828 ();
 b15zdnd11an1n16x5 FILLER_265_861 ();
 b15zdnd11an1n04x5 FILLER_265_877 ();
 b15zdnd00an1n01x5 FILLER_265_881 ();
 b15zdnd11an1n32x5 FILLER_265_894 ();
 b15zdnd11an1n16x5 FILLER_265_926 ();
 b15zdnd11an1n08x5 FILLER_265_942 ();
 b15zdnd11an1n04x5 FILLER_265_950 ();
 b15zdnd00an1n01x5 FILLER_265_954 ();
 b15zdnd11an1n04x5 FILLER_265_963 ();
 b15zdnd11an1n04x5 FILLER_265_976 ();
 b15zdnd11an1n32x5 FILLER_265_995 ();
 b15zdnd11an1n08x5 FILLER_265_1027 ();
 b15zdnd00an1n01x5 FILLER_265_1035 ();
 b15zdnd11an1n32x5 FILLER_265_1040 ();
 b15zdnd11an1n04x5 FILLER_265_1072 ();
 b15zdnd00an1n02x5 FILLER_265_1076 ();
 b15zdnd00an1n01x5 FILLER_265_1078 ();
 b15zdnd11an1n08x5 FILLER_265_1088 ();
 b15zdnd11an1n04x5 FILLER_265_1102 ();
 b15zdnd11an1n04x5 FILLER_265_1116 ();
 b15zdnd00an1n01x5 FILLER_265_1120 ();
 b15zdnd11an1n04x5 FILLER_265_1133 ();
 b15zdnd11an1n16x5 FILLER_265_1145 ();
 b15zdnd11an1n04x5 FILLER_265_1161 ();
 b15zdnd11an1n16x5 FILLER_265_1170 ();
 b15zdnd11an1n08x5 FILLER_265_1186 ();
 b15zdnd00an1n01x5 FILLER_265_1194 ();
 b15zdnd11an1n04x5 FILLER_265_1201 ();
 b15zdnd11an1n32x5 FILLER_265_1211 ();
 b15zdnd11an1n16x5 FILLER_265_1243 ();
 b15zdnd11an1n04x5 FILLER_265_1259 ();
 b15zdnd00an1n02x5 FILLER_265_1263 ();
 b15zdnd00an1n01x5 FILLER_265_1265 ();
 b15zdnd11an1n32x5 FILLER_265_1270 ();
 b15zdnd11an1n16x5 FILLER_265_1302 ();
 b15zdnd00an1n01x5 FILLER_265_1318 ();
 b15zdnd11an1n04x5 FILLER_265_1326 ();
 b15zdnd00an1n01x5 FILLER_265_1330 ();
 b15zdnd11an1n32x5 FILLER_265_1345 ();
 b15zdnd11an1n04x5 FILLER_265_1377 ();
 b15zdnd11an1n32x5 FILLER_265_1407 ();
 b15zdnd11an1n08x5 FILLER_265_1439 ();
 b15zdnd11an1n04x5 FILLER_265_1447 ();
 b15zdnd00an1n02x5 FILLER_265_1451 ();
 b15zdnd00an1n01x5 FILLER_265_1453 ();
 b15zdnd11an1n64x5 FILLER_265_1464 ();
 b15zdnd11an1n32x5 FILLER_265_1528 ();
 b15zdnd00an1n02x5 FILLER_265_1560 ();
 b15zdnd00an1n01x5 FILLER_265_1562 ();
 b15zdnd11an1n32x5 FILLER_265_1570 ();
 b15zdnd11an1n16x5 FILLER_265_1602 ();
 b15zdnd11an1n08x5 FILLER_265_1618 ();
 b15zdnd11an1n04x5 FILLER_265_1626 ();
 b15zdnd00an1n01x5 FILLER_265_1630 ();
 b15zdnd11an1n08x5 FILLER_265_1637 ();
 b15zdnd11an1n04x5 FILLER_265_1645 ();
 b15zdnd00an1n02x5 FILLER_265_1649 ();
 b15zdnd00an1n01x5 FILLER_265_1651 ();
 b15zdnd11an1n64x5 FILLER_265_1658 ();
 b15zdnd11an1n32x5 FILLER_265_1729 ();
 b15zdnd11an1n16x5 FILLER_265_1761 ();
 b15zdnd11an1n04x5 FILLER_265_1777 ();
 b15zdnd00an1n02x5 FILLER_265_1781 ();
 b15zdnd00an1n01x5 FILLER_265_1783 ();
 b15zdnd11an1n64x5 FILLER_265_1790 ();
 b15zdnd11an1n64x5 FILLER_265_1854 ();
 b15zdnd11an1n64x5 FILLER_265_1918 ();
 b15zdnd11an1n16x5 FILLER_265_1982 ();
 b15zdnd11an1n04x5 FILLER_265_1998 ();
 b15zdnd00an1n02x5 FILLER_265_2002 ();
 b15zdnd00an1n01x5 FILLER_265_2004 ();
 b15zdnd11an1n16x5 FILLER_265_2014 ();
 b15zdnd11an1n04x5 FILLER_265_2030 ();
 b15zdnd11an1n32x5 FILLER_265_2041 ();
 b15zdnd11an1n16x5 FILLER_265_2073 ();
 b15zdnd11an1n04x5 FILLER_265_2089 ();
 b15zdnd00an1n02x5 FILLER_265_2093 ();
 b15zdnd00an1n01x5 FILLER_265_2095 ();
 b15zdnd11an1n04x5 FILLER_265_2108 ();
 b15zdnd11an1n64x5 FILLER_265_2117 ();
 b15zdnd11an1n64x5 FILLER_265_2193 ();
 b15zdnd11an1n16x5 FILLER_265_2257 ();
 b15zdnd11an1n08x5 FILLER_265_2273 ();
 b15zdnd00an1n02x5 FILLER_265_2281 ();
 b15zdnd00an1n01x5 FILLER_265_2283 ();
 b15zdnd11an1n16x5 FILLER_266_8 ();
 b15zdnd11an1n08x5 FILLER_266_24 ();
 b15zdnd00an1n02x5 FILLER_266_32 ();
 b15zdnd11an1n16x5 FILLER_266_38 ();
 b15zdnd00an1n01x5 FILLER_266_54 ();
 b15zdnd11an1n08x5 FILLER_266_71 ();
 b15zdnd11an1n04x5 FILLER_266_79 ();
 b15zdnd00an1n02x5 FILLER_266_83 ();
 b15zdnd11an1n16x5 FILLER_266_96 ();
 b15zdnd11an1n04x5 FILLER_266_112 ();
 b15zdnd00an1n01x5 FILLER_266_116 ();
 b15zdnd11an1n64x5 FILLER_266_126 ();
 b15zdnd11an1n64x5 FILLER_266_190 ();
 b15zdnd11an1n08x5 FILLER_266_254 ();
 b15zdnd11an1n32x5 FILLER_266_280 ();
 b15zdnd11an1n16x5 FILLER_266_312 ();
 b15zdnd11an1n08x5 FILLER_266_343 ();
 b15zdnd00an1n02x5 FILLER_266_351 ();
 b15zdnd11an1n32x5 FILLER_266_374 ();
 b15zdnd11an1n16x5 FILLER_266_406 ();
 b15zdnd11an1n04x5 FILLER_266_422 ();
 b15zdnd11an1n32x5 FILLER_266_444 ();
 b15zdnd11an1n08x5 FILLER_266_476 ();
 b15zdnd11an1n04x5 FILLER_266_484 ();
 b15zdnd00an1n02x5 FILLER_266_488 ();
 b15zdnd00an1n01x5 FILLER_266_490 ();
 b15zdnd11an1n04x5 FILLER_266_505 ();
 b15zdnd00an1n01x5 FILLER_266_509 ();
 b15zdnd11an1n04x5 FILLER_266_516 ();
 b15zdnd00an1n02x5 FILLER_266_520 ();
 b15zdnd00an1n01x5 FILLER_266_522 ();
 b15zdnd11an1n08x5 FILLER_266_533 ();
 b15zdnd00an1n01x5 FILLER_266_541 ();
 b15zdnd11an1n32x5 FILLER_266_548 ();
 b15zdnd11an1n16x5 FILLER_266_580 ();
 b15zdnd11an1n08x5 FILLER_266_596 ();
 b15zdnd11an1n04x5 FILLER_266_604 ();
 b15zdnd00an1n02x5 FILLER_266_608 ();
 b15zdnd00an1n01x5 FILLER_266_610 ();
 b15zdnd11an1n32x5 FILLER_266_624 ();
 b15zdnd11an1n16x5 FILLER_266_656 ();
 b15zdnd11an1n08x5 FILLER_266_672 ();
 b15zdnd11an1n04x5 FILLER_266_680 ();
 b15zdnd00an1n02x5 FILLER_266_684 ();
 b15zdnd11an1n08x5 FILLER_266_707 ();
 b15zdnd00an1n02x5 FILLER_266_715 ();
 b15zdnd00an1n01x5 FILLER_266_717 ();
 b15zdnd11an1n08x5 FILLER_266_726 ();
 b15zdnd11an1n04x5 FILLER_266_734 ();
 b15zdnd00an1n01x5 FILLER_266_738 ();
 b15zdnd11an1n32x5 FILLER_266_754 ();
 b15zdnd11an1n16x5 FILLER_266_798 ();
 b15zdnd11an1n04x5 FILLER_266_814 ();
 b15zdnd00an1n02x5 FILLER_266_818 ();
 b15zdnd00an1n01x5 FILLER_266_820 ();
 b15zdnd11an1n04x5 FILLER_266_841 ();
 b15zdnd00an1n02x5 FILLER_266_845 ();
 b15zdnd00an1n01x5 FILLER_266_847 ();
 b15zdnd11an1n04x5 FILLER_266_879 ();
 b15zdnd11an1n64x5 FILLER_266_892 ();
 b15zdnd11an1n32x5 FILLER_266_956 ();
 b15zdnd11an1n16x5 FILLER_266_988 ();
 b15zdnd00an1n02x5 FILLER_266_1004 ();
 b15zdnd11an1n16x5 FILLER_266_1018 ();
 b15zdnd00an1n02x5 FILLER_266_1034 ();
 b15zdnd00an1n01x5 FILLER_266_1036 ();
 b15zdnd11an1n32x5 FILLER_266_1044 ();
 b15zdnd11an1n16x5 FILLER_266_1076 ();
 b15zdnd00an1n02x5 FILLER_266_1092 ();
 b15zdnd11an1n16x5 FILLER_266_1108 ();
 b15zdnd11an1n08x5 FILLER_266_1124 ();
 b15zdnd11an1n16x5 FILLER_266_1137 ();
 b15zdnd11an1n08x5 FILLER_266_1153 ();
 b15zdnd00an1n02x5 FILLER_266_1161 ();
 b15zdnd00an1n01x5 FILLER_266_1163 ();
 b15zdnd11an1n32x5 FILLER_266_1171 ();
 b15zdnd11an1n32x5 FILLER_266_1210 ();
 b15zdnd11an1n04x5 FILLER_266_1242 ();
 b15zdnd00an1n02x5 FILLER_266_1246 ();
 b15zdnd00an1n01x5 FILLER_266_1248 ();
 b15zdnd11an1n32x5 FILLER_266_1258 ();
 b15zdnd11an1n08x5 FILLER_266_1290 ();
 b15zdnd11an1n04x5 FILLER_266_1298 ();
 b15zdnd11an1n04x5 FILLER_266_1314 ();
 b15zdnd00an1n01x5 FILLER_266_1318 ();
 b15zdnd11an1n64x5 FILLER_266_1325 ();
 b15zdnd11an1n32x5 FILLER_266_1389 ();
 b15zdnd11an1n08x5 FILLER_266_1421 ();
 b15zdnd00an1n02x5 FILLER_266_1429 ();
 b15zdnd11an1n64x5 FILLER_266_1440 ();
 b15zdnd11an1n32x5 FILLER_266_1504 ();
 b15zdnd00an1n02x5 FILLER_266_1536 ();
 b15zdnd00an1n01x5 FILLER_266_1538 ();
 b15zdnd11an1n16x5 FILLER_266_1545 ();
 b15zdnd00an1n01x5 FILLER_266_1561 ();
 b15zdnd11an1n64x5 FILLER_266_1567 ();
 b15zdnd00an1n02x5 FILLER_266_1631 ();
 b15zdnd00an1n01x5 FILLER_266_1633 ();
 b15zdnd11an1n16x5 FILLER_266_1639 ();
 b15zdnd11an1n08x5 FILLER_266_1655 ();
 b15zdnd11an1n08x5 FILLER_266_1668 ();
 b15zdnd00an1n01x5 FILLER_266_1676 ();
 b15zdnd11an1n32x5 FILLER_266_1683 ();
 b15zdnd11an1n08x5 FILLER_266_1715 ();
 b15zdnd11an1n16x5 FILLER_266_1729 ();
 b15zdnd11an1n08x5 FILLER_266_1745 ();
 b15zdnd00an1n01x5 FILLER_266_1753 ();
 b15zdnd11an1n08x5 FILLER_266_1759 ();
 b15zdnd11an1n04x5 FILLER_266_1767 ();
 b15zdnd00an1n02x5 FILLER_266_1771 ();
 b15zdnd11an1n16x5 FILLER_266_1780 ();
 b15zdnd11an1n04x5 FILLER_266_1796 ();
 b15zdnd00an1n01x5 FILLER_266_1800 ();
 b15zdnd11an1n64x5 FILLER_266_1827 ();
 b15zdnd11an1n08x5 FILLER_266_1891 ();
 b15zdnd11an1n04x5 FILLER_266_1899 ();
 b15zdnd00an1n01x5 FILLER_266_1903 ();
 b15zdnd11an1n64x5 FILLER_266_1908 ();
 b15zdnd11an1n08x5 FILLER_266_1972 ();
 b15zdnd11an1n04x5 FILLER_266_1980 ();
 b15zdnd00an1n02x5 FILLER_266_1984 ();
 b15zdnd00an1n01x5 FILLER_266_1986 ();
 b15zdnd11an1n08x5 FILLER_266_1993 ();
 b15zdnd11an1n04x5 FILLER_266_2001 ();
 b15zdnd11an1n08x5 FILLER_266_2010 ();
 b15zdnd11an1n04x5 FILLER_266_2018 ();
 b15zdnd00an1n02x5 FILLER_266_2022 ();
 b15zdnd00an1n01x5 FILLER_266_2024 ();
 b15zdnd11an1n08x5 FILLER_266_2042 ();
 b15zdnd00an1n02x5 FILLER_266_2050 ();
 b15zdnd11an1n32x5 FILLER_266_2057 ();
 b15zdnd11an1n16x5 FILLER_266_2089 ();
 b15zdnd11an1n08x5 FILLER_266_2105 ();
 b15zdnd00an1n01x5 FILLER_266_2113 ();
 b15zdnd11an1n04x5 FILLER_266_2120 ();
 b15zdnd11an1n04x5 FILLER_266_2130 ();
 b15zdnd00an1n02x5 FILLER_266_2134 ();
 b15zdnd00an1n02x5 FILLER_266_2152 ();
 b15zdnd11an1n32x5 FILLER_266_2162 ();
 b15zdnd11an1n16x5 FILLER_266_2194 ();
 b15zdnd11an1n08x5 FILLER_266_2210 ();
 b15zdnd11an1n04x5 FILLER_266_2218 ();
 b15zdnd00an1n01x5 FILLER_266_2222 ();
 b15zdnd11an1n32x5 FILLER_266_2227 ();
 b15zdnd11an1n16x5 FILLER_266_2259 ();
 b15zdnd00an1n01x5 FILLER_266_2275 ();
 b15zdnd11an1n32x5 FILLER_267_0 ();
 b15zdnd11an1n04x5 FILLER_267_32 ();
 b15zdnd00an1n01x5 FILLER_267_36 ();
 b15zdnd11an1n08x5 FILLER_267_44 ();
 b15zdnd11an1n04x5 FILLER_267_52 ();
 b15zdnd00an1n02x5 FILLER_267_56 ();
 b15zdnd11an1n08x5 FILLER_267_62 ();
 b15zdnd00an1n02x5 FILLER_267_70 ();
 b15zdnd00an1n01x5 FILLER_267_72 ();
 b15zdnd11an1n04x5 FILLER_267_94 ();
 b15zdnd11an1n32x5 FILLER_267_103 ();
 b15zdnd11an1n08x5 FILLER_267_135 ();
 b15zdnd11an1n32x5 FILLER_267_150 ();
 b15zdnd00an1n01x5 FILLER_267_182 ();
 b15zdnd11an1n04x5 FILLER_267_189 ();
 b15zdnd00an1n02x5 FILLER_267_193 ();
 b15zdnd11an1n64x5 FILLER_267_205 ();
 b15zdnd11an1n64x5 FILLER_267_269 ();
 b15zdnd11an1n16x5 FILLER_267_333 ();
 b15zdnd11an1n08x5 FILLER_267_349 ();
 b15zdnd00an1n02x5 FILLER_267_357 ();
 b15zdnd00an1n01x5 FILLER_267_359 ();
 b15zdnd11an1n64x5 FILLER_267_366 ();
 b15zdnd11an1n64x5 FILLER_267_430 ();
 b15zdnd11an1n16x5 FILLER_267_494 ();
 b15zdnd00an1n02x5 FILLER_267_510 ();
 b15zdnd11an1n04x5 FILLER_267_533 ();
 b15zdnd11an1n08x5 FILLER_267_550 ();
 b15zdnd11an1n04x5 FILLER_267_558 ();
 b15zdnd00an1n02x5 FILLER_267_562 ();
 b15zdnd00an1n01x5 FILLER_267_564 ();
 b15zdnd11an1n08x5 FILLER_267_570 ();
 b15zdnd11an1n04x5 FILLER_267_578 ();
 b15zdnd00an1n02x5 FILLER_267_582 ();
 b15zdnd11an1n32x5 FILLER_267_596 ();
 b15zdnd11an1n16x5 FILLER_267_628 ();
 b15zdnd11an1n08x5 FILLER_267_644 ();
 b15zdnd00an1n02x5 FILLER_267_652 ();
 b15zdnd11an1n16x5 FILLER_267_658 ();
 b15zdnd11an1n08x5 FILLER_267_674 ();
 b15zdnd11an1n04x5 FILLER_267_682 ();
 b15zdnd00an1n02x5 FILLER_267_686 ();
 b15zdnd11an1n04x5 FILLER_267_694 ();
 b15zdnd00an1n01x5 FILLER_267_698 ();
 b15zdnd11an1n04x5 FILLER_267_704 ();
 b15zdnd11an1n04x5 FILLER_267_719 ();
 b15zdnd11an1n04x5 FILLER_267_731 ();
 b15zdnd11an1n08x5 FILLER_267_741 ();
 b15zdnd11an1n04x5 FILLER_267_749 ();
 b15zdnd00an1n01x5 FILLER_267_753 ();
 b15zdnd11an1n08x5 FILLER_267_759 ();
 b15zdnd11an1n04x5 FILLER_267_767 ();
 b15zdnd00an1n02x5 FILLER_267_771 ();
 b15zdnd11an1n08x5 FILLER_267_784 ();
 b15zdnd00an1n01x5 FILLER_267_792 ();
 b15zdnd11an1n64x5 FILLER_267_798 ();
 b15zdnd11an1n64x5 FILLER_267_862 ();
 b15zdnd11an1n64x5 FILLER_267_926 ();
 b15zdnd11an1n08x5 FILLER_267_990 ();
 b15zdnd11an1n04x5 FILLER_267_998 ();
 b15zdnd00an1n02x5 FILLER_267_1002 ();
 b15zdnd00an1n01x5 FILLER_267_1004 ();
 b15zdnd11an1n08x5 FILLER_267_1017 ();
 b15zdnd00an1n02x5 FILLER_267_1025 ();
 b15zdnd00an1n01x5 FILLER_267_1027 ();
 b15zdnd11an1n32x5 FILLER_267_1046 ();
 b15zdnd11an1n08x5 FILLER_267_1078 ();
 b15zdnd11an1n04x5 FILLER_267_1086 ();
 b15zdnd11an1n64x5 FILLER_267_1097 ();
 b15zdnd11an1n64x5 FILLER_267_1161 ();
 b15zdnd11an1n16x5 FILLER_267_1225 ();
 b15zdnd11an1n08x5 FILLER_267_1241 ();
 b15zdnd00an1n01x5 FILLER_267_1249 ();
 b15zdnd11an1n04x5 FILLER_267_1256 ();
 b15zdnd00an1n01x5 FILLER_267_1260 ();
 b15zdnd11an1n32x5 FILLER_267_1267 ();
 b15zdnd11an1n04x5 FILLER_267_1299 ();
 b15zdnd00an1n02x5 FILLER_267_1303 ();
 b15zdnd11an1n32x5 FILLER_267_1314 ();
 b15zdnd00an1n02x5 FILLER_267_1346 ();
 b15zdnd00an1n01x5 FILLER_267_1348 ();
 b15zdnd11an1n32x5 FILLER_267_1356 ();
 b15zdnd11an1n16x5 FILLER_267_1388 ();
 b15zdnd00an1n01x5 FILLER_267_1404 ();
 b15zdnd11an1n16x5 FILLER_267_1425 ();
 b15zdnd11an1n16x5 FILLER_267_1453 ();
 b15zdnd11an1n08x5 FILLER_267_1469 ();
 b15zdnd11an1n04x5 FILLER_267_1477 ();
 b15zdnd00an1n02x5 FILLER_267_1481 ();
 b15zdnd11an1n08x5 FILLER_267_1496 ();
 b15zdnd00an1n02x5 FILLER_267_1504 ();
 b15zdnd11an1n16x5 FILLER_267_1522 ();
 b15zdnd11an1n64x5 FILLER_267_1543 ();
 b15zdnd11an1n32x5 FILLER_267_1607 ();
 b15zdnd11an1n16x5 FILLER_267_1639 ();
 b15zdnd11an1n04x5 FILLER_267_1655 ();
 b15zdnd00an1n02x5 FILLER_267_1659 ();
 b15zdnd11an1n16x5 FILLER_267_1665 ();
 b15zdnd11an1n08x5 FILLER_267_1681 ();
 b15zdnd11an1n04x5 FILLER_267_1689 ();
 b15zdnd11an1n32x5 FILLER_267_1697 ();
 b15zdnd11an1n16x5 FILLER_267_1729 ();
 b15zdnd11an1n08x5 FILLER_267_1745 ();
 b15zdnd00an1n02x5 FILLER_267_1753 ();
 b15zdnd11an1n32x5 FILLER_267_1761 ();
 b15zdnd11an1n16x5 FILLER_267_1793 ();
 b15zdnd00an1n02x5 FILLER_267_1809 ();
 b15zdnd00an1n01x5 FILLER_267_1811 ();
 b15zdnd11an1n64x5 FILLER_267_1818 ();
 b15zdnd11an1n16x5 FILLER_267_1882 ();
 b15zdnd11an1n08x5 FILLER_267_1898 ();
 b15zdnd00an1n01x5 FILLER_267_1906 ();
 b15zdnd11an1n16x5 FILLER_267_1914 ();
 b15zdnd11an1n04x5 FILLER_267_1930 ();
 b15zdnd00an1n01x5 FILLER_267_1934 ();
 b15zdnd11an1n04x5 FILLER_267_1941 ();
 b15zdnd00an1n02x5 FILLER_267_1945 ();
 b15zdnd11an1n08x5 FILLER_267_1955 ();
 b15zdnd11an1n04x5 FILLER_267_1963 ();
 b15zdnd00an1n01x5 FILLER_267_1967 ();
 b15zdnd11an1n08x5 FILLER_267_1974 ();
 b15zdnd11an1n32x5 FILLER_267_1992 ();
 b15zdnd11an1n04x5 FILLER_267_2024 ();
 b15zdnd00an1n01x5 FILLER_267_2028 ();
 b15zdnd11an1n16x5 FILLER_267_2035 ();
 b15zdnd00an1n02x5 FILLER_267_2051 ();
 b15zdnd00an1n01x5 FILLER_267_2053 ();
 b15zdnd11an1n16x5 FILLER_267_2066 ();
 b15zdnd11an1n04x5 FILLER_267_2082 ();
 b15zdnd00an1n02x5 FILLER_267_2086 ();
 b15zdnd11an1n64x5 FILLER_267_2100 ();
 b15zdnd11an1n32x5 FILLER_267_2164 ();
 b15zdnd00an1n01x5 FILLER_267_2196 ();
 b15zdnd11an1n04x5 FILLER_267_2203 ();
 b15zdnd00an1n02x5 FILLER_267_2207 ();
 b15zdnd11an1n04x5 FILLER_267_2215 ();
 b15zdnd00an1n02x5 FILLER_267_2219 ();
 b15zdnd00an1n01x5 FILLER_267_2221 ();
 b15zdnd11an1n04x5 FILLER_267_2230 ();
 b15zdnd00an1n02x5 FILLER_267_2234 ();
 b15zdnd11an1n32x5 FILLER_267_2240 ();
 b15zdnd11an1n08x5 FILLER_267_2272 ();
 b15zdnd11an1n04x5 FILLER_267_2280 ();
 b15zdnd11an1n32x5 FILLER_268_8 ();
 b15zdnd11an1n08x5 FILLER_268_40 ();
 b15zdnd00an1n01x5 FILLER_268_48 ();
 b15zdnd11an1n16x5 FILLER_268_67 ();
 b15zdnd11an1n04x5 FILLER_268_83 ();
 b15zdnd00an1n01x5 FILLER_268_87 ();
 b15zdnd11an1n64x5 FILLER_268_97 ();
 b15zdnd11an1n32x5 FILLER_268_161 ();
 b15zdnd11an1n04x5 FILLER_268_193 ();
 b15zdnd11an1n08x5 FILLER_268_201 ();
 b15zdnd11an1n04x5 FILLER_268_209 ();
 b15zdnd11an1n16x5 FILLER_268_218 ();
 b15zdnd00an1n01x5 FILLER_268_234 ();
 b15zdnd11an1n32x5 FILLER_268_249 ();
 b15zdnd11an1n08x5 FILLER_268_281 ();
 b15zdnd00an1n01x5 FILLER_268_289 ();
 b15zdnd11an1n32x5 FILLER_268_305 ();
 b15zdnd11an1n16x5 FILLER_268_337 ();
 b15zdnd11an1n64x5 FILLER_268_361 ();
 b15zdnd11an1n64x5 FILLER_268_425 ();
 b15zdnd11an1n64x5 FILLER_268_489 ();
 b15zdnd11an1n16x5 FILLER_268_553 ();
 b15zdnd11an1n08x5 FILLER_268_569 ();
 b15zdnd11an1n04x5 FILLER_268_577 ();
 b15zdnd00an1n02x5 FILLER_268_581 ();
 b15zdnd00an1n01x5 FILLER_268_583 ();
 b15zdnd11an1n16x5 FILLER_268_590 ();
 b15zdnd00an1n02x5 FILLER_268_606 ();
 b15zdnd11an1n08x5 FILLER_268_614 ();
 b15zdnd11an1n04x5 FILLER_268_622 ();
 b15zdnd00an1n02x5 FILLER_268_626 ();
 b15zdnd11an1n04x5 FILLER_268_636 ();
 b15zdnd00an1n02x5 FILLER_268_640 ();
 b15zdnd00an1n01x5 FILLER_268_642 ();
 b15zdnd11an1n32x5 FILLER_268_648 ();
 b15zdnd11an1n04x5 FILLER_268_680 ();
 b15zdnd00an1n02x5 FILLER_268_684 ();
 b15zdnd00an1n01x5 FILLER_268_686 ();
 b15zdnd11an1n16x5 FILLER_268_697 ();
 b15zdnd11an1n04x5 FILLER_268_713 ();
 b15zdnd00an1n01x5 FILLER_268_717 ();
 b15zdnd11an1n04x5 FILLER_268_726 ();
 b15zdnd00an1n02x5 FILLER_268_730 ();
 b15zdnd00an1n01x5 FILLER_268_732 ();
 b15zdnd11an1n32x5 FILLER_268_739 ();
 b15zdnd11an1n04x5 FILLER_268_771 ();
 b15zdnd00an1n02x5 FILLER_268_775 ();
 b15zdnd11an1n16x5 FILLER_268_793 ();
 b15zdnd11an1n64x5 FILLER_268_813 ();
 b15zdnd11an1n08x5 FILLER_268_877 ();
 b15zdnd11an1n64x5 FILLER_268_894 ();
 b15zdnd11an1n32x5 FILLER_268_958 ();
 b15zdnd00an1n01x5 FILLER_268_990 ();
 b15zdnd11an1n64x5 FILLER_268_997 ();
 b15zdnd11an1n64x5 FILLER_268_1061 ();
 b15zdnd11an1n64x5 FILLER_268_1125 ();
 b15zdnd11an1n64x5 FILLER_268_1189 ();
 b15zdnd00an1n01x5 FILLER_268_1253 ();
 b15zdnd11an1n64x5 FILLER_268_1264 ();
 b15zdnd11an1n64x5 FILLER_268_1328 ();
 b15zdnd11an1n32x5 FILLER_268_1392 ();
 b15zdnd11an1n08x5 FILLER_268_1424 ();
 b15zdnd11an1n04x5 FILLER_268_1432 ();
 b15zdnd00an1n02x5 FILLER_268_1436 ();
 b15zdnd11an1n04x5 FILLER_268_1450 ();
 b15zdnd11an1n16x5 FILLER_268_1473 ();
 b15zdnd00an1n02x5 FILLER_268_1489 ();
 b15zdnd11an1n32x5 FILLER_268_1501 ();
 b15zdnd11an1n08x5 FILLER_268_1533 ();
 b15zdnd11an1n04x5 FILLER_268_1541 ();
 b15zdnd00an1n01x5 FILLER_268_1545 ();
 b15zdnd11an1n04x5 FILLER_268_1554 ();
 b15zdnd00an1n01x5 FILLER_268_1558 ();
 b15zdnd11an1n04x5 FILLER_268_1569 ();
 b15zdnd00an1n02x5 FILLER_268_1573 ();
 b15zdnd11an1n04x5 FILLER_268_1582 ();
 b15zdnd11an1n04x5 FILLER_268_1598 ();
 b15zdnd11an1n04x5 FILLER_268_1607 ();
 b15zdnd00an1n01x5 FILLER_268_1611 ();
 b15zdnd11an1n04x5 FILLER_268_1617 ();
 b15zdnd11an1n16x5 FILLER_268_1627 ();
 b15zdnd11an1n08x5 FILLER_268_1643 ();
 b15zdnd11an1n04x5 FILLER_268_1651 ();
 b15zdnd00an1n02x5 FILLER_268_1655 ();
 b15zdnd11an1n08x5 FILLER_268_1666 ();
 b15zdnd11an1n04x5 FILLER_268_1688 ();
 b15zdnd11an1n16x5 FILLER_268_1698 ();
 b15zdnd11an1n08x5 FILLER_268_1714 ();
 b15zdnd00an1n01x5 FILLER_268_1722 ();
 b15zdnd11an1n08x5 FILLER_268_1730 ();
 b15zdnd00an1n01x5 FILLER_268_1738 ();
 b15zdnd11an1n04x5 FILLER_268_1743 ();
 b15zdnd00an1n02x5 FILLER_268_1747 ();
 b15zdnd00an1n01x5 FILLER_268_1749 ();
 b15zdnd11an1n32x5 FILLER_268_1756 ();
 b15zdnd11an1n08x5 FILLER_268_1788 ();
 b15zdnd11an1n04x5 FILLER_268_1796 ();
 b15zdnd00an1n02x5 FILLER_268_1800 ();
 b15zdnd11an1n04x5 FILLER_268_1811 ();
 b15zdnd00an1n01x5 FILLER_268_1815 ();
 b15zdnd11an1n32x5 FILLER_268_1823 ();
 b15zdnd11an1n16x5 FILLER_268_1855 ();
 b15zdnd11an1n08x5 FILLER_268_1871 ();
 b15zdnd11an1n04x5 FILLER_268_1879 ();
 b15zdnd00an1n02x5 FILLER_268_1883 ();
 b15zdnd00an1n01x5 FILLER_268_1885 ();
 b15zdnd11an1n32x5 FILLER_268_1896 ();
 b15zdnd00an1n02x5 FILLER_268_1928 ();
 b15zdnd00an1n01x5 FILLER_268_1930 ();
 b15zdnd11an1n16x5 FILLER_268_1941 ();
 b15zdnd11an1n08x5 FILLER_268_1957 ();
 b15zdnd00an1n02x5 FILLER_268_1965 ();
 b15zdnd11an1n04x5 FILLER_268_1979 ();
 b15zdnd00an1n02x5 FILLER_268_1983 ();
 b15zdnd00an1n01x5 FILLER_268_1985 ();
 b15zdnd11an1n32x5 FILLER_268_1992 ();
 b15zdnd00an1n02x5 FILLER_268_2024 ();
 b15zdnd11an1n04x5 FILLER_268_2041 ();
 b15zdnd11an1n04x5 FILLER_268_2055 ();
 b15zdnd11an1n64x5 FILLER_268_2064 ();
 b15zdnd11an1n04x5 FILLER_268_2128 ();
 b15zdnd00an1n02x5 FILLER_268_2152 ();
 b15zdnd11an1n32x5 FILLER_268_2162 ();
 b15zdnd11an1n16x5 FILLER_268_2194 ();
 b15zdnd11an1n04x5 FILLER_268_2218 ();
 b15zdnd00an1n01x5 FILLER_268_2222 ();
 b15zdnd11an1n32x5 FILLER_268_2229 ();
 b15zdnd11an1n08x5 FILLER_268_2261 ();
 b15zdnd11an1n04x5 FILLER_268_2269 ();
 b15zdnd00an1n02x5 FILLER_268_2273 ();
 b15zdnd00an1n01x5 FILLER_268_2275 ();
 b15zdnd11an1n32x5 FILLER_269_0 ();
 b15zdnd11an1n16x5 FILLER_269_32 ();
 b15zdnd11an1n08x5 FILLER_269_48 ();
 b15zdnd11an1n04x5 FILLER_269_56 ();
 b15zdnd00an1n02x5 FILLER_269_60 ();
 b15zdnd00an1n01x5 FILLER_269_62 ();
 b15zdnd11an1n16x5 FILLER_269_68 ();
 b15zdnd11an1n04x5 FILLER_269_84 ();
 b15zdnd00an1n02x5 FILLER_269_88 ();
 b15zdnd00an1n01x5 FILLER_269_90 ();
 b15zdnd11an1n32x5 FILLER_269_98 ();
 b15zdnd11an1n16x5 FILLER_269_130 ();
 b15zdnd11an1n08x5 FILLER_269_146 ();
 b15zdnd11an1n04x5 FILLER_269_154 ();
 b15zdnd11an1n04x5 FILLER_269_163 ();
 b15zdnd11an1n04x5 FILLER_269_183 ();
 b15zdnd00an1n01x5 FILLER_269_187 ();
 b15zdnd11an1n32x5 FILLER_269_195 ();
 b15zdnd11an1n16x5 FILLER_269_227 ();
 b15zdnd11an1n04x5 FILLER_269_243 ();
 b15zdnd11an1n32x5 FILLER_269_253 ();
 b15zdnd00an1n02x5 FILLER_269_285 ();
 b15zdnd00an1n01x5 FILLER_269_287 ();
 b15zdnd11an1n08x5 FILLER_269_294 ();
 b15zdnd00an1n02x5 FILLER_269_302 ();
 b15zdnd00an1n01x5 FILLER_269_304 ();
 b15zdnd11an1n04x5 FILLER_269_318 ();
 b15zdnd11an1n04x5 FILLER_269_327 ();
 b15zdnd00an1n01x5 FILLER_269_331 ();
 b15zdnd11an1n64x5 FILLER_269_339 ();
 b15zdnd11an1n32x5 FILLER_269_403 ();
 b15zdnd11an1n16x5 FILLER_269_435 ();
 b15zdnd11an1n04x5 FILLER_269_451 ();
 b15zdnd00an1n02x5 FILLER_269_455 ();
 b15zdnd00an1n01x5 FILLER_269_457 ();
 b15zdnd11an1n32x5 FILLER_269_462 ();
 b15zdnd11an1n08x5 FILLER_269_494 ();
 b15zdnd11an1n04x5 FILLER_269_502 ();
 b15zdnd11an1n32x5 FILLER_269_524 ();
 b15zdnd11an1n04x5 FILLER_269_556 ();
 b15zdnd00an1n02x5 FILLER_269_560 ();
 b15zdnd11an1n64x5 FILLER_269_572 ();
 b15zdnd11an1n64x5 FILLER_269_636 ();
 b15zdnd11an1n64x5 FILLER_269_700 ();
 b15zdnd11an1n16x5 FILLER_269_764 ();
 b15zdnd11an1n04x5 FILLER_269_780 ();
 b15zdnd00an1n02x5 FILLER_269_784 ();
 b15zdnd11an1n04x5 FILLER_269_798 ();
 b15zdnd11an1n32x5 FILLER_269_813 ();
 b15zdnd11an1n08x5 FILLER_269_845 ();
 b15zdnd11an1n04x5 FILLER_269_871 ();
 b15zdnd11an1n04x5 FILLER_269_894 ();
 b15zdnd11an1n64x5 FILLER_269_923 ();
 b15zdnd11an1n08x5 FILLER_269_987 ();
 b15zdnd00an1n01x5 FILLER_269_995 ();
 b15zdnd11an1n32x5 FILLER_269_1002 ();
 b15zdnd00an1n02x5 FILLER_269_1034 ();
 b15zdnd11an1n08x5 FILLER_269_1051 ();
 b15zdnd11an1n04x5 FILLER_269_1059 ();
 b15zdnd00an1n01x5 FILLER_269_1063 ();
 b15zdnd11an1n08x5 FILLER_269_1084 ();
 b15zdnd11an1n32x5 FILLER_269_1098 ();
 b15zdnd11an1n08x5 FILLER_269_1130 ();
 b15zdnd00an1n01x5 FILLER_269_1138 ();
 b15zdnd11an1n32x5 FILLER_269_1144 ();
 b15zdnd11an1n16x5 FILLER_269_1176 ();
 b15zdnd11an1n08x5 FILLER_269_1192 ();
 b15zdnd11an1n32x5 FILLER_269_1205 ();
 b15zdnd11an1n08x5 FILLER_269_1237 ();
 b15zdnd00an1n02x5 FILLER_269_1245 ();
 b15zdnd00an1n01x5 FILLER_269_1247 ();
 b15zdnd11an1n04x5 FILLER_269_1253 ();
 b15zdnd00an1n02x5 FILLER_269_1257 ();
 b15zdnd11an1n08x5 FILLER_269_1263 ();
 b15zdnd00an1n02x5 FILLER_269_1271 ();
 b15zdnd00an1n01x5 FILLER_269_1273 ();
 b15zdnd11an1n16x5 FILLER_269_1284 ();
 b15zdnd11an1n32x5 FILLER_269_1306 ();
 b15zdnd11an1n16x5 FILLER_269_1338 ();
 b15zdnd00an1n02x5 FILLER_269_1354 ();
 b15zdnd00an1n01x5 FILLER_269_1356 ();
 b15zdnd11an1n04x5 FILLER_269_1363 ();
 b15zdnd00an1n01x5 FILLER_269_1367 ();
 b15zdnd11an1n64x5 FILLER_269_1374 ();
 b15zdnd11an1n32x5 FILLER_269_1438 ();
 b15zdnd11an1n04x5 FILLER_269_1470 ();
 b15zdnd11an1n04x5 FILLER_269_1478 ();
 b15zdnd00an1n02x5 FILLER_269_1482 ();
 b15zdnd11an1n04x5 FILLER_269_1490 ();
 b15zdnd11an1n16x5 FILLER_269_1500 ();
 b15zdnd11an1n04x5 FILLER_269_1516 ();
 b15zdnd00an1n01x5 FILLER_269_1520 ();
 b15zdnd11an1n08x5 FILLER_269_1527 ();
 b15zdnd00an1n02x5 FILLER_269_1535 ();
 b15zdnd00an1n01x5 FILLER_269_1537 ();
 b15zdnd11an1n08x5 FILLER_269_1548 ();
 b15zdnd00an1n01x5 FILLER_269_1556 ();
 b15zdnd11an1n32x5 FILLER_269_1589 ();
 b15zdnd11an1n04x5 FILLER_269_1626 ();
 b15zdnd11an1n04x5 FILLER_269_1635 ();
 b15zdnd00an1n02x5 FILLER_269_1639 ();
 b15zdnd11an1n32x5 FILLER_269_1649 ();
 b15zdnd11an1n08x5 FILLER_269_1681 ();
 b15zdnd11an1n16x5 FILLER_269_1699 ();
 b15zdnd11an1n04x5 FILLER_269_1715 ();
 b15zdnd00an1n01x5 FILLER_269_1719 ();
 b15zdnd11an1n16x5 FILLER_269_1736 ();
 b15zdnd11an1n04x5 FILLER_269_1752 ();
 b15zdnd00an1n01x5 FILLER_269_1756 ();
 b15zdnd11an1n04x5 FILLER_269_1773 ();
 b15zdnd11an1n64x5 FILLER_269_1782 ();
 b15zdnd11an1n32x5 FILLER_269_1846 ();
 b15zdnd11an1n08x5 FILLER_269_1878 ();
 b15zdnd00an1n01x5 FILLER_269_1886 ();
 b15zdnd11an1n16x5 FILLER_269_1897 ();
 b15zdnd11an1n04x5 FILLER_269_1913 ();
 b15zdnd00an1n01x5 FILLER_269_1917 ();
 b15zdnd11an1n04x5 FILLER_269_1930 ();
 b15zdnd11an1n08x5 FILLER_269_1939 ();
 b15zdnd00an1n01x5 FILLER_269_1947 ();
 b15zdnd11an1n64x5 FILLER_269_1969 ();
 b15zdnd11an1n16x5 FILLER_269_2033 ();
 b15zdnd00an1n01x5 FILLER_269_2049 ();
 b15zdnd11an1n32x5 FILLER_269_2062 ();
 b15zdnd00an1n02x5 FILLER_269_2094 ();
 b15zdnd00an1n01x5 FILLER_269_2096 ();
 b15zdnd11an1n32x5 FILLER_269_2103 ();
 b15zdnd00an1n01x5 FILLER_269_2135 ();
 b15zdnd11an1n64x5 FILLER_269_2150 ();
 b15zdnd11an1n64x5 FILLER_269_2214 ();
 b15zdnd11an1n04x5 FILLER_269_2278 ();
 b15zdnd00an1n02x5 FILLER_269_2282 ();
 b15zdnd11an1n64x5 FILLER_270_8 ();
 b15zdnd11an1n16x5 FILLER_270_72 ();
 b15zdnd11an1n04x5 FILLER_270_88 ();
 b15zdnd11an1n08x5 FILLER_270_102 ();
 b15zdnd11an1n04x5 FILLER_270_110 ();
 b15zdnd11an1n64x5 FILLER_270_124 ();
 b15zdnd11an1n32x5 FILLER_270_188 ();
 b15zdnd11an1n04x5 FILLER_270_220 ();
 b15zdnd00an1n02x5 FILLER_270_224 ();
 b15zdnd00an1n01x5 FILLER_270_226 ();
 b15zdnd11an1n64x5 FILLER_270_232 ();
 b15zdnd11an1n04x5 FILLER_270_302 ();
 b15zdnd11an1n16x5 FILLER_270_312 ();
 b15zdnd11an1n08x5 FILLER_270_344 ();
 b15zdnd11an1n04x5 FILLER_270_352 ();
 b15zdnd11an1n32x5 FILLER_270_366 ();
 b15zdnd11an1n16x5 FILLER_270_398 ();
 b15zdnd11an1n08x5 FILLER_270_414 ();
 b15zdnd11an1n04x5 FILLER_270_422 ();
 b15zdnd00an1n02x5 FILLER_270_426 ();
 b15zdnd00an1n01x5 FILLER_270_428 ();
 b15zdnd11an1n16x5 FILLER_270_438 ();
 b15zdnd11an1n04x5 FILLER_270_454 ();
 b15zdnd00an1n01x5 FILLER_270_458 ();
 b15zdnd11an1n08x5 FILLER_270_467 ();
 b15zdnd11an1n32x5 FILLER_270_481 ();
 b15zdnd11an1n08x5 FILLER_270_513 ();
 b15zdnd11an1n04x5 FILLER_270_521 ();
 b15zdnd00an1n01x5 FILLER_270_525 ();
 b15zdnd11an1n32x5 FILLER_270_542 ();
 b15zdnd00an1n02x5 FILLER_270_574 ();
 b15zdnd11an1n16x5 FILLER_270_581 ();
 b15zdnd11an1n08x5 FILLER_270_597 ();
 b15zdnd11an1n04x5 FILLER_270_612 ();
 b15zdnd11an1n64x5 FILLER_270_628 ();
 b15zdnd11an1n16x5 FILLER_270_692 ();
 b15zdnd11an1n08x5 FILLER_270_708 ();
 b15zdnd00an1n02x5 FILLER_270_716 ();
 b15zdnd11an1n64x5 FILLER_270_726 ();
 b15zdnd11an1n32x5 FILLER_270_790 ();
 b15zdnd00an1n02x5 FILLER_270_822 ();
 b15zdnd00an1n01x5 FILLER_270_824 ();
 b15zdnd11an1n64x5 FILLER_270_856 ();
 b15zdnd11an1n32x5 FILLER_270_920 ();
 b15zdnd11an1n16x5 FILLER_270_952 ();
 b15zdnd11an1n04x5 FILLER_270_968 ();
 b15zdnd00an1n01x5 FILLER_270_972 ();
 b15zdnd11an1n16x5 FILLER_270_978 ();
 b15zdnd00an1n02x5 FILLER_270_994 ();
 b15zdnd11an1n32x5 FILLER_270_1005 ();
 b15zdnd11an1n16x5 FILLER_270_1037 ();
 b15zdnd11an1n08x5 FILLER_270_1053 ();
 b15zdnd00an1n01x5 FILLER_270_1061 ();
 b15zdnd11an1n16x5 FILLER_270_1072 ();
 b15zdnd00an1n01x5 FILLER_270_1088 ();
 b15zdnd11an1n32x5 FILLER_270_1095 ();
 b15zdnd11an1n16x5 FILLER_270_1127 ();
 b15zdnd11an1n04x5 FILLER_270_1143 ();
 b15zdnd00an1n02x5 FILLER_270_1147 ();
 b15zdnd11an1n04x5 FILLER_270_1155 ();
 b15zdnd00an1n02x5 FILLER_270_1159 ();
 b15zdnd11an1n04x5 FILLER_270_1167 ();
 b15zdnd00an1n01x5 FILLER_270_1171 ();
 b15zdnd11an1n16x5 FILLER_270_1179 ();
 b15zdnd11an1n04x5 FILLER_270_1195 ();
 b15zdnd00an1n02x5 FILLER_270_1199 ();
 b15zdnd00an1n01x5 FILLER_270_1201 ();
 b15zdnd11an1n64x5 FILLER_270_1208 ();
 b15zdnd11an1n64x5 FILLER_270_1272 ();
 b15zdnd11an1n16x5 FILLER_270_1336 ();
 b15zdnd00an1n01x5 FILLER_270_1352 ();
 b15zdnd11an1n64x5 FILLER_270_1362 ();
 b15zdnd00an1n02x5 FILLER_270_1426 ();
 b15zdnd00an1n01x5 FILLER_270_1428 ();
 b15zdnd11an1n32x5 FILLER_270_1444 ();
 b15zdnd00an1n01x5 FILLER_270_1476 ();
 b15zdnd11an1n64x5 FILLER_270_1483 ();
 b15zdnd11an1n64x5 FILLER_270_1547 ();
 b15zdnd11an1n64x5 FILLER_270_1611 ();
 b15zdnd11an1n16x5 FILLER_270_1675 ();
 b15zdnd11an1n04x5 FILLER_270_1691 ();
 b15zdnd00an1n02x5 FILLER_270_1695 ();
 b15zdnd11an1n64x5 FILLER_270_1701 ();
 b15zdnd11an1n16x5 FILLER_270_1765 ();
 b15zdnd11an1n08x5 FILLER_270_1781 ();
 b15zdnd00an1n02x5 FILLER_270_1789 ();
 b15zdnd00an1n01x5 FILLER_270_1791 ();
 b15zdnd11an1n04x5 FILLER_270_1796 ();
 b15zdnd00an1n01x5 FILLER_270_1800 ();
 b15zdnd11an1n64x5 FILLER_270_1813 ();
 b15zdnd11an1n16x5 FILLER_270_1877 ();
 b15zdnd11an1n08x5 FILLER_270_1893 ();
 b15zdnd11an1n04x5 FILLER_270_1901 ();
 b15zdnd11an1n32x5 FILLER_270_1910 ();
 b15zdnd11an1n08x5 FILLER_270_1942 ();
 b15zdnd11an1n04x5 FILLER_270_1950 ();
 b15zdnd00an1n02x5 FILLER_270_1954 ();
 b15zdnd11an1n64x5 FILLER_270_1965 ();
 b15zdnd11an1n64x5 FILLER_270_2029 ();
 b15zdnd11an1n04x5 FILLER_270_2093 ();
 b15zdnd11an1n32x5 FILLER_270_2107 ();
 b15zdnd11an1n08x5 FILLER_270_2139 ();
 b15zdnd11an1n04x5 FILLER_270_2147 ();
 b15zdnd00an1n02x5 FILLER_270_2151 ();
 b15zdnd00an1n01x5 FILLER_270_2153 ();
 b15zdnd11an1n16x5 FILLER_270_2162 ();
 b15zdnd00an1n01x5 FILLER_270_2178 ();
 b15zdnd11an1n08x5 FILLER_270_2188 ();
 b15zdnd00an1n01x5 FILLER_270_2196 ();
 b15zdnd11an1n16x5 FILLER_270_2212 ();
 b15zdnd00an1n02x5 FILLER_270_2228 ();
 b15zdnd00an1n01x5 FILLER_270_2230 ();
 b15zdnd11an1n04x5 FILLER_270_2236 ();
 b15zdnd11an1n16x5 FILLER_270_2245 ();
 b15zdnd11an1n08x5 FILLER_270_2261 ();
 b15zdnd11an1n04x5 FILLER_270_2269 ();
 b15zdnd00an1n02x5 FILLER_270_2273 ();
 b15zdnd00an1n01x5 FILLER_270_2275 ();
 b15zdnd11an1n64x5 FILLER_271_0 ();
 b15zdnd11an1n16x5 FILLER_271_64 ();
 b15zdnd11an1n04x5 FILLER_271_80 ();
 b15zdnd00an1n02x5 FILLER_271_84 ();
 b15zdnd11an1n04x5 FILLER_271_107 ();
 b15zdnd11an1n04x5 FILLER_271_119 ();
 b15zdnd11an1n04x5 FILLER_271_136 ();
 b15zdnd11an1n64x5 FILLER_271_156 ();
 b15zdnd11an1n08x5 FILLER_271_220 ();
 b15zdnd11an1n08x5 FILLER_271_233 ();
 b15zdnd11an1n04x5 FILLER_271_241 ();
 b15zdnd00an1n01x5 FILLER_271_245 ();
 b15zdnd11an1n04x5 FILLER_271_253 ();
 b15zdnd11an1n32x5 FILLER_271_265 ();
 b15zdnd11an1n16x5 FILLER_271_297 ();
 b15zdnd11an1n08x5 FILLER_271_313 ();
 b15zdnd11an1n04x5 FILLER_271_321 ();
 b15zdnd00an1n02x5 FILLER_271_325 ();
 b15zdnd00an1n01x5 FILLER_271_327 ();
 b15zdnd11an1n16x5 FILLER_271_334 ();
 b15zdnd00an1n02x5 FILLER_271_350 ();
 b15zdnd00an1n01x5 FILLER_271_352 ();
 b15zdnd11an1n32x5 FILLER_271_369 ();
 b15zdnd11an1n16x5 FILLER_271_401 ();
 b15zdnd11an1n08x5 FILLER_271_417 ();
 b15zdnd00an1n02x5 FILLER_271_425 ();
 b15zdnd00an1n01x5 FILLER_271_427 ();
 b15zdnd11an1n16x5 FILLER_271_439 ();
 b15zdnd11an1n08x5 FILLER_271_455 ();
 b15zdnd00an1n02x5 FILLER_271_463 ();
 b15zdnd11an1n08x5 FILLER_271_479 ();
 b15zdnd00an1n02x5 FILLER_271_487 ();
 b15zdnd00an1n01x5 FILLER_271_489 ();
 b15zdnd11an1n04x5 FILLER_271_510 ();
 b15zdnd11an1n04x5 FILLER_271_519 ();
 b15zdnd11an1n08x5 FILLER_271_528 ();
 b15zdnd11an1n04x5 FILLER_271_557 ();
 b15zdnd00an1n02x5 FILLER_271_561 ();
 b15zdnd11an1n04x5 FILLER_271_571 ();
 b15zdnd11an1n32x5 FILLER_271_587 ();
 b15zdnd11an1n08x5 FILLER_271_619 ();
 b15zdnd00an1n02x5 FILLER_271_627 ();
 b15zdnd00an1n01x5 FILLER_271_629 ();
 b15zdnd11an1n16x5 FILLER_271_644 ();
 b15zdnd00an1n01x5 FILLER_271_660 ();
 b15zdnd11an1n04x5 FILLER_271_671 ();
 b15zdnd11an1n04x5 FILLER_271_695 ();
 b15zdnd11an1n16x5 FILLER_271_709 ();
 b15zdnd11an1n04x5 FILLER_271_725 ();
 b15zdnd00an1n02x5 FILLER_271_729 ();
 b15zdnd00an1n01x5 FILLER_271_731 ();
 b15zdnd11an1n04x5 FILLER_271_737 ();
 b15zdnd11an1n04x5 FILLER_271_751 ();
 b15zdnd11an1n08x5 FILLER_271_760 ();
 b15zdnd00an1n02x5 FILLER_271_768 ();
 b15zdnd00an1n01x5 FILLER_271_770 ();
 b15zdnd11an1n04x5 FILLER_271_780 ();
 b15zdnd11an1n64x5 FILLER_271_789 ();
 b15zdnd11an1n64x5 FILLER_271_853 ();
 b15zdnd11an1n32x5 FILLER_271_917 ();
 b15zdnd11an1n16x5 FILLER_271_949 ();
 b15zdnd11an1n08x5 FILLER_271_965 ();
 b15zdnd11an1n04x5 FILLER_271_973 ();
 b15zdnd00an1n01x5 FILLER_271_977 ();
 b15zdnd11an1n08x5 FILLER_271_990 ();
 b15zdnd00an1n02x5 FILLER_271_998 ();
 b15zdnd11an1n32x5 FILLER_271_1015 ();
 b15zdnd11an1n08x5 FILLER_271_1047 ();
 b15zdnd00an1n01x5 FILLER_271_1055 ();
 b15zdnd11an1n32x5 FILLER_271_1060 ();
 b15zdnd00an1n02x5 FILLER_271_1092 ();
 b15zdnd00an1n01x5 FILLER_271_1094 ();
 b15zdnd11an1n04x5 FILLER_271_1102 ();
 b15zdnd11an1n32x5 FILLER_271_1110 ();
 b15zdnd11an1n04x5 FILLER_271_1154 ();
 b15zdnd00an1n02x5 FILLER_271_1158 ();
 b15zdnd00an1n01x5 FILLER_271_1160 ();
 b15zdnd11an1n04x5 FILLER_271_1176 ();
 b15zdnd00an1n02x5 FILLER_271_1180 ();
 b15zdnd11an1n04x5 FILLER_271_1189 ();
 b15zdnd11an1n08x5 FILLER_271_1208 ();
 b15zdnd11an1n04x5 FILLER_271_1216 ();
 b15zdnd11an1n04x5 FILLER_271_1234 ();
 b15zdnd11an1n04x5 FILLER_271_1251 ();
 b15zdnd11an1n16x5 FILLER_271_1274 ();
 b15zdnd11an1n04x5 FILLER_271_1290 ();
 b15zdnd00an1n01x5 FILLER_271_1294 ();
 b15zdnd11an1n04x5 FILLER_271_1309 ();
 b15zdnd11an1n08x5 FILLER_271_1320 ();
 b15zdnd00an1n02x5 FILLER_271_1328 ();
 b15zdnd11an1n04x5 FILLER_271_1346 ();
 b15zdnd11an1n64x5 FILLER_271_1367 ();
 b15zdnd11an1n16x5 FILLER_271_1431 ();
 b15zdnd00an1n01x5 FILLER_271_1447 ();
 b15zdnd11an1n16x5 FILLER_271_1453 ();
 b15zdnd11an1n04x5 FILLER_271_1469 ();
 b15zdnd00an1n01x5 FILLER_271_1473 ();
 b15zdnd11an1n64x5 FILLER_271_1480 ();
 b15zdnd11an1n32x5 FILLER_271_1544 ();
 b15zdnd11an1n08x5 FILLER_271_1576 ();
 b15zdnd00an1n01x5 FILLER_271_1584 ();
 b15zdnd11an1n64x5 FILLER_271_1605 ();
 b15zdnd11an1n64x5 FILLER_271_1669 ();
 b15zdnd11an1n32x5 FILLER_271_1733 ();
 b15zdnd11an1n08x5 FILLER_271_1765 ();
 b15zdnd00an1n02x5 FILLER_271_1773 ();
 b15zdnd00an1n01x5 FILLER_271_1775 ();
 b15zdnd11an1n08x5 FILLER_271_1783 ();
 b15zdnd11an1n04x5 FILLER_271_1791 ();
 b15zdnd11an1n04x5 FILLER_271_1800 ();
 b15zdnd00an1n02x5 FILLER_271_1804 ();
 b15zdnd00an1n01x5 FILLER_271_1806 ();
 b15zdnd11an1n04x5 FILLER_271_1819 ();
 b15zdnd11an1n64x5 FILLER_271_1832 ();
 b15zdnd11an1n64x5 FILLER_271_1896 ();
 b15zdnd11an1n16x5 FILLER_271_1960 ();
 b15zdnd11an1n08x5 FILLER_271_1976 ();
 b15zdnd00an1n02x5 FILLER_271_1984 ();
 b15zdnd00an1n01x5 FILLER_271_1986 ();
 b15zdnd11an1n08x5 FILLER_271_1992 ();
 b15zdnd11an1n04x5 FILLER_271_2000 ();
 b15zdnd11an1n32x5 FILLER_271_2010 ();
 b15zdnd00an1n02x5 FILLER_271_2042 ();
 b15zdnd00an1n01x5 FILLER_271_2044 ();
 b15zdnd11an1n32x5 FILLER_271_2054 ();
 b15zdnd11an1n08x5 FILLER_271_2086 ();
 b15zdnd11an1n04x5 FILLER_271_2094 ();
 b15zdnd11an1n04x5 FILLER_271_2104 ();
 b15zdnd11an1n04x5 FILLER_271_2120 ();
 b15zdnd11an1n04x5 FILLER_271_2135 ();
 b15zdnd11an1n08x5 FILLER_271_2145 ();
 b15zdnd00an1n01x5 FILLER_271_2153 ();
 b15zdnd11an1n04x5 FILLER_271_2166 ();
 b15zdnd11an1n32x5 FILLER_271_2177 ();
 b15zdnd11an1n16x5 FILLER_271_2209 ();
 b15zdnd11an1n08x5 FILLER_271_2225 ();
 b15zdnd11an1n04x5 FILLER_271_2233 ();
 b15zdnd11an1n32x5 FILLER_271_2251 ();
 b15zdnd00an1n01x5 FILLER_271_2283 ();
 b15zdnd11an1n16x5 FILLER_272_8 ();
 b15zdnd11an1n08x5 FILLER_272_24 ();
 b15zdnd11an1n04x5 FILLER_272_32 ();
 b15zdnd00an1n02x5 FILLER_272_36 ();
 b15zdnd11an1n08x5 FILLER_272_43 ();
 b15zdnd11an1n04x5 FILLER_272_51 ();
 b15zdnd00an1n01x5 FILLER_272_55 ();
 b15zdnd11an1n16x5 FILLER_272_66 ();
 b15zdnd11an1n04x5 FILLER_272_88 ();
 b15zdnd11an1n32x5 FILLER_272_101 ();
 b15zdnd11an1n04x5 FILLER_272_133 ();
 b15zdnd11an1n04x5 FILLER_272_149 ();
 b15zdnd11an1n16x5 FILLER_272_169 ();
 b15zdnd00an1n02x5 FILLER_272_185 ();
 b15zdnd11an1n08x5 FILLER_272_201 ();
 b15zdnd00an1n01x5 FILLER_272_209 ();
 b15zdnd11an1n64x5 FILLER_272_219 ();
 b15zdnd11an1n32x5 FILLER_272_283 ();
 b15zdnd11an1n08x5 FILLER_272_315 ();
 b15zdnd00an1n02x5 FILLER_272_323 ();
 b15zdnd11an1n64x5 FILLER_272_336 ();
 b15zdnd11an1n16x5 FILLER_272_400 ();
 b15zdnd11an1n08x5 FILLER_272_416 ();
 b15zdnd11an1n04x5 FILLER_272_424 ();
 b15zdnd00an1n01x5 FILLER_272_428 ();
 b15zdnd11an1n04x5 FILLER_272_436 ();
 b15zdnd11an1n32x5 FILLER_272_452 ();
 b15zdnd11an1n04x5 FILLER_272_484 ();
 b15zdnd00an1n02x5 FILLER_272_488 ();
 b15zdnd00an1n01x5 FILLER_272_490 ();
 b15zdnd11an1n16x5 FILLER_272_501 ();
 b15zdnd00an1n01x5 FILLER_272_517 ();
 b15zdnd11an1n32x5 FILLER_272_528 ();
 b15zdnd11an1n08x5 FILLER_272_560 ();
 b15zdnd11an1n04x5 FILLER_272_568 ();
 b15zdnd00an1n01x5 FILLER_272_572 ();
 b15zdnd11an1n04x5 FILLER_272_585 ();
 b15zdnd11an1n32x5 FILLER_272_595 ();
 b15zdnd11an1n04x5 FILLER_272_627 ();
 b15zdnd00an1n01x5 FILLER_272_631 ();
 b15zdnd11an1n08x5 FILLER_272_645 ();
 b15zdnd00an1n02x5 FILLER_272_653 ();
 b15zdnd11an1n04x5 FILLER_272_676 ();
 b15zdnd11an1n16x5 FILLER_272_693 ();
 b15zdnd11an1n08x5 FILLER_272_709 ();
 b15zdnd00an1n01x5 FILLER_272_717 ();
 b15zdnd11an1n32x5 FILLER_272_726 ();
 b15zdnd11an1n08x5 FILLER_272_758 ();
 b15zdnd00an1n02x5 FILLER_272_766 ();
 b15zdnd11an1n32x5 FILLER_272_772 ();
 b15zdnd11an1n04x5 FILLER_272_804 ();
 b15zdnd11an1n16x5 FILLER_272_812 ();
 b15zdnd11an1n08x5 FILLER_272_828 ();
 b15zdnd11an1n04x5 FILLER_272_836 ();
 b15zdnd00an1n02x5 FILLER_272_840 ();
 b15zdnd00an1n01x5 FILLER_272_842 ();
 b15zdnd11an1n32x5 FILLER_272_855 ();
 b15zdnd11an1n16x5 FILLER_272_887 ();
 b15zdnd11an1n08x5 FILLER_272_903 ();
 b15zdnd11an1n04x5 FILLER_272_911 ();
 b15zdnd00an1n01x5 FILLER_272_915 ();
 b15zdnd11an1n64x5 FILLER_272_948 ();
 b15zdnd11an1n08x5 FILLER_272_1012 ();
 b15zdnd11an1n04x5 FILLER_272_1020 ();
 b15zdnd00an1n01x5 FILLER_272_1024 ();
 b15zdnd11an1n08x5 FILLER_272_1030 ();
 b15zdnd00an1n01x5 FILLER_272_1038 ();
 b15zdnd11an1n04x5 FILLER_272_1052 ();
 b15zdnd11an1n04x5 FILLER_272_1070 ();
 b15zdnd11an1n64x5 FILLER_272_1086 ();
 b15zdnd11an1n08x5 FILLER_272_1150 ();
 b15zdnd00an1n01x5 FILLER_272_1158 ();
 b15zdnd11an1n32x5 FILLER_272_1173 ();
 b15zdnd11an1n16x5 FILLER_272_1205 ();
 b15zdnd11an1n08x5 FILLER_272_1221 ();
 b15zdnd00an1n02x5 FILLER_272_1229 ();
 b15zdnd00an1n01x5 FILLER_272_1231 ();
 b15zdnd11an1n32x5 FILLER_272_1258 ();
 b15zdnd11an1n04x5 FILLER_272_1290 ();
 b15zdnd11an1n04x5 FILLER_272_1303 ();
 b15zdnd00an1n01x5 FILLER_272_1307 ();
 b15zdnd11an1n04x5 FILLER_272_1314 ();
 b15zdnd00an1n02x5 FILLER_272_1318 ();
 b15zdnd11an1n04x5 FILLER_272_1340 ();
 b15zdnd00an1n02x5 FILLER_272_1344 ();
 b15zdnd11an1n04x5 FILLER_272_1350 ();
 b15zdnd00an1n02x5 FILLER_272_1354 ();
 b15zdnd00an1n01x5 FILLER_272_1356 ();
 b15zdnd11an1n64x5 FILLER_272_1363 ();
 b15zdnd11an1n08x5 FILLER_272_1427 ();
 b15zdnd00an1n02x5 FILLER_272_1435 ();
 b15zdnd00an1n01x5 FILLER_272_1437 ();
 b15zdnd11an1n16x5 FILLER_272_1452 ();
 b15zdnd11an1n04x5 FILLER_272_1468 ();
 b15zdnd11an1n16x5 FILLER_272_1486 ();
 b15zdnd11an1n08x5 FILLER_272_1502 ();
 b15zdnd11an1n04x5 FILLER_272_1510 ();
 b15zdnd11an1n32x5 FILLER_272_1520 ();
 b15zdnd11an1n08x5 FILLER_272_1552 ();
 b15zdnd00an1n01x5 FILLER_272_1560 ();
 b15zdnd11an1n16x5 FILLER_272_1567 ();
 b15zdnd11an1n04x5 FILLER_272_1583 ();
 b15zdnd00an1n02x5 FILLER_272_1587 ();
 b15zdnd00an1n01x5 FILLER_272_1589 ();
 b15zdnd11an1n04x5 FILLER_272_1596 ();
 b15zdnd11an1n32x5 FILLER_272_1611 ();
 b15zdnd11an1n16x5 FILLER_272_1643 ();
 b15zdnd11an1n04x5 FILLER_272_1659 ();
 b15zdnd00an1n01x5 FILLER_272_1663 ();
 b15zdnd11an1n64x5 FILLER_272_1670 ();
 b15zdnd11an1n04x5 FILLER_272_1734 ();
 b15zdnd11an1n32x5 FILLER_272_1756 ();
 b15zdnd11an1n64x5 FILLER_272_1801 ();
 b15zdnd11an1n16x5 FILLER_272_1865 ();
 b15zdnd11an1n04x5 FILLER_272_1881 ();
 b15zdnd00an1n02x5 FILLER_272_1885 ();
 b15zdnd00an1n01x5 FILLER_272_1887 ();
 b15zdnd11an1n32x5 FILLER_272_1896 ();
 b15zdnd11an1n16x5 FILLER_272_1928 ();
 b15zdnd11an1n04x5 FILLER_272_1944 ();
 b15zdnd00an1n01x5 FILLER_272_1948 ();
 b15zdnd11an1n08x5 FILLER_272_1961 ();
 b15zdnd11an1n04x5 FILLER_272_1969 ();
 b15zdnd00an1n02x5 FILLER_272_1973 ();
 b15zdnd00an1n01x5 FILLER_272_1975 ();
 b15zdnd11an1n32x5 FILLER_272_1991 ();
 b15zdnd11an1n08x5 FILLER_272_2023 ();
 b15zdnd00an1n01x5 FILLER_272_2031 ();
 b15zdnd11an1n04x5 FILLER_272_2040 ();
 b15zdnd11an1n04x5 FILLER_272_2057 ();
 b15zdnd11an1n04x5 FILLER_272_2068 ();
 b15zdnd11an1n64x5 FILLER_272_2076 ();
 b15zdnd11an1n08x5 FILLER_272_2140 ();
 b15zdnd11an1n04x5 FILLER_272_2148 ();
 b15zdnd00an1n02x5 FILLER_272_2152 ();
 b15zdnd11an1n04x5 FILLER_272_2162 ();
 b15zdnd00an1n02x5 FILLER_272_2166 ();
 b15zdnd00an1n01x5 FILLER_272_2168 ();
 b15zdnd11an1n04x5 FILLER_272_2176 ();
 b15zdnd00an1n01x5 FILLER_272_2180 ();
 b15zdnd11an1n04x5 FILLER_272_2185 ();
 b15zdnd11an1n04x5 FILLER_272_2205 ();
 b15zdnd11an1n32x5 FILLER_272_2221 ();
 b15zdnd11an1n16x5 FILLER_272_2253 ();
 b15zdnd11an1n04x5 FILLER_272_2269 ();
 b15zdnd00an1n02x5 FILLER_272_2273 ();
 b15zdnd00an1n01x5 FILLER_272_2275 ();
 b15zdnd11an1n32x5 FILLER_273_0 ();
 b15zdnd11an1n08x5 FILLER_273_32 ();
 b15zdnd11an1n04x5 FILLER_273_50 ();
 b15zdnd00an1n01x5 FILLER_273_54 ();
 b15zdnd11an1n64x5 FILLER_273_69 ();
 b15zdnd11an1n16x5 FILLER_273_133 ();
 b15zdnd11an1n08x5 FILLER_273_158 ();
 b15zdnd00an1n01x5 FILLER_273_166 ();
 b15zdnd11an1n04x5 FILLER_273_180 ();
 b15zdnd11an1n04x5 FILLER_273_191 ();
 b15zdnd00an1n01x5 FILLER_273_195 ();
 b15zdnd11an1n16x5 FILLER_273_212 ();
 b15zdnd00an1n01x5 FILLER_273_228 ();
 b15zdnd11an1n16x5 FILLER_273_245 ();
 b15zdnd11an1n04x5 FILLER_273_261 ();
 b15zdnd11an1n64x5 FILLER_273_277 ();
 b15zdnd11an1n64x5 FILLER_273_341 ();
 b15zdnd11an1n64x5 FILLER_273_405 ();
 b15zdnd00an1n01x5 FILLER_273_469 ();
 b15zdnd11an1n64x5 FILLER_273_498 ();
 b15zdnd11an1n16x5 FILLER_273_562 ();
 b15zdnd11an1n08x5 FILLER_273_578 ();
 b15zdnd00an1n01x5 FILLER_273_586 ();
 b15zdnd11an1n04x5 FILLER_273_603 ();
 b15zdnd11an1n16x5 FILLER_273_613 ();
 b15zdnd11an1n08x5 FILLER_273_629 ();
 b15zdnd00an1n02x5 FILLER_273_637 ();
 b15zdnd00an1n01x5 FILLER_273_639 ();
 b15zdnd11an1n04x5 FILLER_273_647 ();
 b15zdnd00an1n02x5 FILLER_273_651 ();
 b15zdnd11an1n04x5 FILLER_273_662 ();
 b15zdnd11an1n32x5 FILLER_273_677 ();
 b15zdnd11an1n08x5 FILLER_273_709 ();
 b15zdnd00an1n01x5 FILLER_273_717 ();
 b15zdnd11an1n04x5 FILLER_273_722 ();
 b15zdnd11an1n08x5 FILLER_273_740 ();
 b15zdnd00an1n02x5 FILLER_273_748 ();
 b15zdnd11an1n08x5 FILLER_273_755 ();
 b15zdnd00an1n02x5 FILLER_273_763 ();
 b15zdnd11an1n04x5 FILLER_273_775 ();
 b15zdnd11an1n64x5 FILLER_273_783 ();
 b15zdnd11an1n64x5 FILLER_273_847 ();
 b15zdnd11an1n32x5 FILLER_273_911 ();
 b15zdnd11an1n08x5 FILLER_273_943 ();
 b15zdnd00an1n02x5 FILLER_273_951 ();
 b15zdnd00an1n01x5 FILLER_273_953 ();
 b15zdnd11an1n64x5 FILLER_273_962 ();
 b15zdnd11an1n64x5 FILLER_273_1026 ();
 b15zdnd00an1n01x5 FILLER_273_1090 ();
 b15zdnd11an1n04x5 FILLER_273_1095 ();
 b15zdnd11an1n64x5 FILLER_273_1109 ();
 b15zdnd11an1n64x5 FILLER_273_1173 ();
 b15zdnd11an1n64x5 FILLER_273_1237 ();
 b15zdnd11an1n32x5 FILLER_273_1301 ();
 b15zdnd11an1n16x5 FILLER_273_1333 ();
 b15zdnd11an1n08x5 FILLER_273_1349 ();
 b15zdnd11an1n04x5 FILLER_273_1357 ();
 b15zdnd11an1n32x5 FILLER_273_1366 ();
 b15zdnd11an1n16x5 FILLER_273_1398 ();
 b15zdnd11an1n08x5 FILLER_273_1414 ();
 b15zdnd00an1n02x5 FILLER_273_1422 ();
 b15zdnd00an1n01x5 FILLER_273_1424 ();
 b15zdnd11an1n04x5 FILLER_273_1429 ();
 b15zdnd11an1n16x5 FILLER_273_1445 ();
 b15zdnd00an1n02x5 FILLER_273_1461 ();
 b15zdnd11an1n16x5 FILLER_273_1479 ();
 b15zdnd11an1n08x5 FILLER_273_1495 ();
 b15zdnd00an1n02x5 FILLER_273_1503 ();
 b15zdnd00an1n01x5 FILLER_273_1505 ();
 b15zdnd11an1n08x5 FILLER_273_1513 ();
 b15zdnd00an1n02x5 FILLER_273_1521 ();
 b15zdnd11an1n04x5 FILLER_273_1527 ();
 b15zdnd11an1n04x5 FILLER_273_1547 ();
 b15zdnd11an1n32x5 FILLER_273_1556 ();
 b15zdnd11an1n04x5 FILLER_273_1588 ();
 b15zdnd00an1n02x5 FILLER_273_1592 ();
 b15zdnd00an1n01x5 FILLER_273_1594 ();
 b15zdnd11an1n04x5 FILLER_273_1621 ();
 b15zdnd11an1n04x5 FILLER_273_1632 ();
 b15zdnd00an1n02x5 FILLER_273_1636 ();
 b15zdnd11an1n04x5 FILLER_273_1658 ();
 b15zdnd00an1n02x5 FILLER_273_1662 ();
 b15zdnd00an1n01x5 FILLER_273_1664 ();
 b15zdnd11an1n64x5 FILLER_273_1675 ();
 b15zdnd11an1n64x5 FILLER_273_1739 ();
 b15zdnd11an1n64x5 FILLER_273_1803 ();
 b15zdnd11an1n16x5 FILLER_273_1867 ();
 b15zdnd11an1n08x5 FILLER_273_1883 ();
 b15zdnd11an1n04x5 FILLER_273_1891 ();
 b15zdnd00an1n02x5 FILLER_273_1895 ();
 b15zdnd11an1n08x5 FILLER_273_1903 ();
 b15zdnd11an1n04x5 FILLER_273_1911 ();
 b15zdnd11an1n16x5 FILLER_273_1919 ();
 b15zdnd11an1n08x5 FILLER_273_1935 ();
 b15zdnd11an1n04x5 FILLER_273_1943 ();
 b15zdnd00an1n02x5 FILLER_273_1947 ();
 b15zdnd11an1n16x5 FILLER_273_1958 ();
 b15zdnd11an1n04x5 FILLER_273_1974 ();
 b15zdnd00an1n02x5 FILLER_273_1978 ();
 b15zdnd00an1n01x5 FILLER_273_1980 ();
 b15zdnd11an1n32x5 FILLER_273_1985 ();
 b15zdnd11an1n08x5 FILLER_273_2017 ();
 b15zdnd11an1n04x5 FILLER_273_2025 ();
 b15zdnd00an1n02x5 FILLER_273_2029 ();
 b15zdnd00an1n01x5 FILLER_273_2031 ();
 b15zdnd11an1n32x5 FILLER_273_2042 ();
 b15zdnd11an1n08x5 FILLER_273_2074 ();
 b15zdnd11an1n04x5 FILLER_273_2082 ();
 b15zdnd00an1n01x5 FILLER_273_2086 ();
 b15zdnd11an1n64x5 FILLER_273_2097 ();
 b15zdnd11an1n32x5 FILLER_273_2161 ();
 b15zdnd11an1n16x5 FILLER_273_2193 ();
 b15zdnd11an1n08x5 FILLER_273_2209 ();
 b15zdnd11an1n04x5 FILLER_273_2217 ();
 b15zdnd11an1n32x5 FILLER_273_2225 ();
 b15zdnd11an1n16x5 FILLER_273_2257 ();
 b15zdnd11an1n08x5 FILLER_273_2273 ();
 b15zdnd00an1n02x5 FILLER_273_2281 ();
 b15zdnd00an1n01x5 FILLER_273_2283 ();
 b15zdnd11an1n32x5 FILLER_274_8 ();
 b15zdnd11an1n04x5 FILLER_274_40 ();
 b15zdnd11an1n16x5 FILLER_274_51 ();
 b15zdnd00an1n02x5 FILLER_274_67 ();
 b15zdnd00an1n01x5 FILLER_274_69 ();
 b15zdnd11an1n08x5 FILLER_274_75 ();
 b15zdnd11an1n04x5 FILLER_274_83 ();
 b15zdnd00an1n02x5 FILLER_274_87 ();
 b15zdnd00an1n01x5 FILLER_274_89 ();
 b15zdnd11an1n16x5 FILLER_274_95 ();
 b15zdnd11an1n08x5 FILLER_274_111 ();
 b15zdnd11an1n32x5 FILLER_274_132 ();
 b15zdnd11an1n16x5 FILLER_274_169 ();
 b15zdnd11an1n04x5 FILLER_274_185 ();
 b15zdnd00an1n01x5 FILLER_274_189 ();
 b15zdnd11an1n32x5 FILLER_274_194 ();
 b15zdnd11an1n08x5 FILLER_274_226 ();
 b15zdnd00an1n02x5 FILLER_274_234 ();
 b15zdnd00an1n01x5 FILLER_274_236 ();
 b15zdnd11an1n16x5 FILLER_274_255 ();
 b15zdnd11an1n04x5 FILLER_274_271 ();
 b15zdnd00an1n02x5 FILLER_274_275 ();
 b15zdnd11an1n16x5 FILLER_274_287 ();
 b15zdnd11an1n08x5 FILLER_274_303 ();
 b15zdnd00an1n01x5 FILLER_274_311 ();
 b15zdnd11an1n64x5 FILLER_274_320 ();
 b15zdnd11an1n32x5 FILLER_274_384 ();
 b15zdnd11an1n16x5 FILLER_274_416 ();
 b15zdnd11an1n08x5 FILLER_274_432 ();
 b15zdnd11an1n04x5 FILLER_274_440 ();
 b15zdnd00an1n02x5 FILLER_274_444 ();
 b15zdnd00an1n01x5 FILLER_274_446 ();
 b15zdnd11an1n16x5 FILLER_274_463 ();
 b15zdnd11an1n32x5 FILLER_274_483 ();
 b15zdnd11an1n16x5 FILLER_274_515 ();
 b15zdnd11an1n08x5 FILLER_274_541 ();
 b15zdnd11an1n04x5 FILLER_274_549 ();
 b15zdnd00an1n02x5 FILLER_274_553 ();
 b15zdnd11an1n64x5 FILLER_274_559 ();
 b15zdnd11an1n32x5 FILLER_274_623 ();
 b15zdnd11an1n16x5 FILLER_274_655 ();
 b15zdnd11an1n08x5 FILLER_274_671 ();
 b15zdnd11an1n04x5 FILLER_274_679 ();
 b15zdnd00an1n02x5 FILLER_274_683 ();
 b15zdnd11an1n16x5 FILLER_274_690 ();
 b15zdnd11an1n08x5 FILLER_274_706 ();
 b15zdnd11an1n04x5 FILLER_274_714 ();
 b15zdnd11an1n64x5 FILLER_274_726 ();
 b15zdnd11an1n16x5 FILLER_274_790 ();
 b15zdnd00an1n01x5 FILLER_274_806 ();
 b15zdnd11an1n32x5 FILLER_274_813 ();
 b15zdnd11an1n08x5 FILLER_274_845 ();
 b15zdnd11an1n04x5 FILLER_274_853 ();
 b15zdnd11an1n04x5 FILLER_274_888 ();
 b15zdnd11an1n64x5 FILLER_274_917 ();
 b15zdnd11an1n64x5 FILLER_274_989 ();
 b15zdnd11an1n64x5 FILLER_274_1053 ();
 b15zdnd11an1n32x5 FILLER_274_1117 ();
 b15zdnd11an1n04x5 FILLER_274_1149 ();
 b15zdnd00an1n02x5 FILLER_274_1153 ();
 b15zdnd11an1n16x5 FILLER_274_1167 ();
 b15zdnd11an1n08x5 FILLER_274_1183 ();
 b15zdnd00an1n01x5 FILLER_274_1191 ();
 b15zdnd11an1n32x5 FILLER_274_1198 ();
 b15zdnd11an1n08x5 FILLER_274_1230 ();
 b15zdnd11an1n04x5 FILLER_274_1238 ();
 b15zdnd11an1n08x5 FILLER_274_1247 ();
 b15zdnd11an1n04x5 FILLER_274_1255 ();
 b15zdnd00an1n02x5 FILLER_274_1259 ();
 b15zdnd11an1n64x5 FILLER_274_1270 ();
 b15zdnd11an1n04x5 FILLER_274_1334 ();
 b15zdnd00an1n02x5 FILLER_274_1338 ();
 b15zdnd11an1n64x5 FILLER_274_1346 ();
 b15zdnd11an1n64x5 FILLER_274_1410 ();
 b15zdnd11an1n16x5 FILLER_274_1474 ();
 b15zdnd11an1n08x5 FILLER_274_1490 ();
 b15zdnd11an1n04x5 FILLER_274_1498 ();
 b15zdnd00an1n02x5 FILLER_274_1502 ();
 b15zdnd11an1n32x5 FILLER_274_1511 ();
 b15zdnd11an1n16x5 FILLER_274_1543 ();
 b15zdnd11an1n08x5 FILLER_274_1559 ();
 b15zdnd11an1n08x5 FILLER_274_1574 ();
 b15zdnd00an1n02x5 FILLER_274_1582 ();
 b15zdnd11an1n08x5 FILLER_274_1600 ();
 b15zdnd11an1n04x5 FILLER_274_1608 ();
 b15zdnd00an1n01x5 FILLER_274_1612 ();
 b15zdnd11an1n08x5 FILLER_274_1617 ();
 b15zdnd11an1n04x5 FILLER_274_1625 ();
 b15zdnd00an1n02x5 FILLER_274_1629 ();
 b15zdnd00an1n01x5 FILLER_274_1631 ();
 b15zdnd11an1n32x5 FILLER_274_1639 ();
 b15zdnd11an1n16x5 FILLER_274_1671 ();
 b15zdnd11an1n08x5 FILLER_274_1687 ();
 b15zdnd11an1n04x5 FILLER_274_1695 ();
 b15zdnd11an1n16x5 FILLER_274_1711 ();
 b15zdnd11an1n08x5 FILLER_274_1727 ();
 b15zdnd00an1n02x5 FILLER_274_1735 ();
 b15zdnd00an1n01x5 FILLER_274_1737 ();
 b15zdnd11an1n64x5 FILLER_274_1764 ();
 b15zdnd11an1n64x5 FILLER_274_1828 ();
 b15zdnd00an1n01x5 FILLER_274_1892 ();
 b15zdnd11an1n16x5 FILLER_274_1897 ();
 b15zdnd11an1n08x5 FILLER_274_1913 ();
 b15zdnd00an1n02x5 FILLER_274_1921 ();
 b15zdnd11an1n08x5 FILLER_274_1936 ();
 b15zdnd11an1n04x5 FILLER_274_1944 ();
 b15zdnd00an1n01x5 FILLER_274_1948 ();
 b15zdnd11an1n64x5 FILLER_274_1971 ();
 b15zdnd11an1n04x5 FILLER_274_2035 ();
 b15zdnd00an1n01x5 FILLER_274_2039 ();
 b15zdnd11an1n04x5 FILLER_274_2048 ();
 b15zdnd11an1n32x5 FILLER_274_2056 ();
 b15zdnd00an1n01x5 FILLER_274_2088 ();
 b15zdnd11an1n16x5 FILLER_274_2094 ();
 b15zdnd11an1n04x5 FILLER_274_2110 ();
 b15zdnd00an1n02x5 FILLER_274_2114 ();
 b15zdnd11an1n08x5 FILLER_274_2127 ();
 b15zdnd00an1n02x5 FILLER_274_2135 ();
 b15zdnd00an1n01x5 FILLER_274_2137 ();
 b15zdnd11an1n04x5 FILLER_274_2148 ();
 b15zdnd00an1n02x5 FILLER_274_2152 ();
 b15zdnd11an1n64x5 FILLER_274_2162 ();
 b15zdnd11an1n32x5 FILLER_274_2226 ();
 b15zdnd11an1n16x5 FILLER_274_2258 ();
 b15zdnd00an1n02x5 FILLER_274_2274 ();
 b15zdnd11an1n32x5 FILLER_275_0 ();
 b15zdnd11an1n04x5 FILLER_275_32 ();
 b15zdnd00an1n02x5 FILLER_275_36 ();
 b15zdnd11an1n64x5 FILLER_275_46 ();
 b15zdnd00an1n01x5 FILLER_275_110 ();
 b15zdnd11an1n64x5 FILLER_275_126 ();
 b15zdnd11an1n16x5 FILLER_275_190 ();
 b15zdnd11an1n08x5 FILLER_275_206 ();
 b15zdnd11an1n04x5 FILLER_275_214 ();
 b15zdnd11an1n08x5 FILLER_275_230 ();
 b15zdnd11an1n32x5 FILLER_275_261 ();
 b15zdnd11an1n16x5 FILLER_275_293 ();
 b15zdnd00an1n02x5 FILLER_275_309 ();
 b15zdnd00an1n01x5 FILLER_275_311 ();
 b15zdnd11an1n04x5 FILLER_275_324 ();
 b15zdnd00an1n02x5 FILLER_275_328 ();
 b15zdnd00an1n01x5 FILLER_275_330 ();
 b15zdnd11an1n64x5 FILLER_275_352 ();
 b15zdnd11an1n16x5 FILLER_275_416 ();
 b15zdnd00an1n02x5 FILLER_275_432 ();
 b15zdnd11an1n08x5 FILLER_275_446 ();
 b15zdnd11an1n04x5 FILLER_275_454 ();
 b15zdnd00an1n02x5 FILLER_275_458 ();
 b15zdnd00an1n01x5 FILLER_275_460 ();
 b15zdnd11an1n64x5 FILLER_275_466 ();
 b15zdnd00an1n02x5 FILLER_275_530 ();
 b15zdnd11an1n08x5 FILLER_275_538 ();
 b15zdnd11an1n04x5 FILLER_275_546 ();
 b15zdnd00an1n02x5 FILLER_275_550 ();
 b15zdnd00an1n01x5 FILLER_275_552 ();
 b15zdnd11an1n32x5 FILLER_275_559 ();
 b15zdnd11an1n08x5 FILLER_275_591 ();
 b15zdnd11an1n04x5 FILLER_275_599 ();
 b15zdnd00an1n01x5 FILLER_275_603 ();
 b15zdnd11an1n32x5 FILLER_275_636 ();
 b15zdnd11an1n16x5 FILLER_275_668 ();
 b15zdnd00an1n01x5 FILLER_275_684 ();
 b15zdnd11an1n32x5 FILLER_275_690 ();
 b15zdnd11an1n16x5 FILLER_275_722 ();
 b15zdnd11an1n08x5 FILLER_275_738 ();
 b15zdnd00an1n02x5 FILLER_275_746 ();
 b15zdnd11an1n32x5 FILLER_275_752 ();
 b15zdnd11an1n08x5 FILLER_275_784 ();
 b15zdnd11an1n04x5 FILLER_275_792 ();
 b15zdnd00an1n02x5 FILLER_275_796 ();
 b15zdnd11an1n64x5 FILLER_275_814 ();
 b15zdnd11an1n08x5 FILLER_275_878 ();
 b15zdnd11an1n04x5 FILLER_275_886 ();
 b15zdnd00an1n01x5 FILLER_275_890 ();
 b15zdnd11an1n32x5 FILLER_275_922 ();
 b15zdnd11an1n16x5 FILLER_275_954 ();
 b15zdnd11an1n04x5 FILLER_275_970 ();
 b15zdnd11an1n08x5 FILLER_275_982 ();
 b15zdnd11an1n64x5 FILLER_275_1000 ();
 b15zdnd11an1n08x5 FILLER_275_1064 ();
 b15zdnd00an1n01x5 FILLER_275_1072 ();
 b15zdnd11an1n04x5 FILLER_275_1088 ();
 b15zdnd11an1n16x5 FILLER_275_1098 ();
 b15zdnd11an1n04x5 FILLER_275_1114 ();
 b15zdnd00an1n02x5 FILLER_275_1118 ();
 b15zdnd00an1n01x5 FILLER_275_1120 ();
 b15zdnd11an1n04x5 FILLER_275_1141 ();
 b15zdnd11an1n32x5 FILLER_275_1149 ();
 b15zdnd11an1n08x5 FILLER_275_1181 ();
 b15zdnd00an1n02x5 FILLER_275_1189 ();
 b15zdnd11an1n32x5 FILLER_275_1198 ();
 b15zdnd11an1n16x5 FILLER_275_1234 ();
 b15zdnd11an1n08x5 FILLER_275_1250 ();
 b15zdnd11an1n04x5 FILLER_275_1258 ();
 b15zdnd00an1n02x5 FILLER_275_1262 ();
 b15zdnd00an1n01x5 FILLER_275_1264 ();
 b15zdnd11an1n64x5 FILLER_275_1269 ();
 b15zdnd11an1n04x5 FILLER_275_1333 ();
 b15zdnd11an1n08x5 FILLER_275_1346 ();
 b15zdnd11an1n64x5 FILLER_275_1363 ();
 b15zdnd00an1n02x5 FILLER_275_1427 ();
 b15zdnd00an1n01x5 FILLER_275_1429 ();
 b15zdnd11an1n04x5 FILLER_275_1435 ();
 b15zdnd11an1n04x5 FILLER_275_1453 ();
 b15zdnd00an1n02x5 FILLER_275_1457 ();
 b15zdnd11an1n08x5 FILLER_275_1468 ();
 b15zdnd11an1n04x5 FILLER_275_1476 ();
 b15zdnd00an1n01x5 FILLER_275_1480 ();
 b15zdnd11an1n04x5 FILLER_275_1501 ();
 b15zdnd11an1n32x5 FILLER_275_1515 ();
 b15zdnd11an1n16x5 FILLER_275_1547 ();
 b15zdnd11an1n04x5 FILLER_275_1563 ();
 b15zdnd11an1n32x5 FILLER_275_1576 ();
 b15zdnd00an1n01x5 FILLER_275_1608 ();
 b15zdnd11an1n04x5 FILLER_275_1614 ();
 b15zdnd00an1n02x5 FILLER_275_1618 ();
 b15zdnd11an1n04x5 FILLER_275_1626 ();
 b15zdnd11an1n08x5 FILLER_275_1639 ();
 b15zdnd11an1n16x5 FILLER_275_1662 ();
 b15zdnd11an1n04x5 FILLER_275_1686 ();
 b15zdnd00an1n02x5 FILLER_275_1690 ();
 b15zdnd00an1n01x5 FILLER_275_1692 ();
 b15zdnd11an1n16x5 FILLER_275_1706 ();
 b15zdnd11an1n04x5 FILLER_275_1722 ();
 b15zdnd00an1n01x5 FILLER_275_1726 ();
 b15zdnd11an1n04x5 FILLER_275_1748 ();
 b15zdnd11an1n08x5 FILLER_275_1760 ();
 b15zdnd11an1n04x5 FILLER_275_1768 ();
 b15zdnd00an1n02x5 FILLER_275_1772 ();
 b15zdnd00an1n01x5 FILLER_275_1774 ();
 b15zdnd11an1n04x5 FILLER_275_1795 ();
 b15zdnd11an1n04x5 FILLER_275_1811 ();
 b15zdnd11an1n64x5 FILLER_275_1824 ();
 b15zdnd11an1n64x5 FILLER_275_1888 ();
 b15zdnd11an1n64x5 FILLER_275_1952 ();
 b15zdnd11an1n32x5 FILLER_275_2016 ();
 b15zdnd00an1n02x5 FILLER_275_2048 ();
 b15zdnd00an1n01x5 FILLER_275_2050 ();
 b15zdnd11an1n16x5 FILLER_275_2057 ();
 b15zdnd11an1n08x5 FILLER_275_2073 ();
 b15zdnd11an1n04x5 FILLER_275_2081 ();
 b15zdnd00an1n02x5 FILLER_275_2085 ();
 b15zdnd11an1n64x5 FILLER_275_2092 ();
 b15zdnd11an1n04x5 FILLER_275_2156 ();
 b15zdnd00an1n02x5 FILLER_275_2160 ();
 b15zdnd11an1n08x5 FILLER_275_2174 ();
 b15zdnd11an1n04x5 FILLER_275_2182 ();
 b15zdnd00an1n01x5 FILLER_275_2186 ();
 b15zdnd11an1n04x5 FILLER_275_2202 ();
 b15zdnd11an1n16x5 FILLER_275_2213 ();
 b15zdnd00an1n02x5 FILLER_275_2229 ();
 b15zdnd11an1n32x5 FILLER_275_2240 ();
 b15zdnd11an1n08x5 FILLER_275_2272 ();
 b15zdnd11an1n04x5 FILLER_275_2280 ();
 b15zdnd11an1n64x5 FILLER_276_8 ();
 b15zdnd11an1n64x5 FILLER_276_72 ();
 b15zdnd00an1n02x5 FILLER_276_136 ();
 b15zdnd11an1n64x5 FILLER_276_145 ();
 b15zdnd11an1n08x5 FILLER_276_209 ();
 b15zdnd11an1n04x5 FILLER_276_217 ();
 b15zdnd11an1n08x5 FILLER_276_228 ();
 b15zdnd11an1n04x5 FILLER_276_236 ();
 b15zdnd00an1n02x5 FILLER_276_240 ();
 b15zdnd00an1n01x5 FILLER_276_242 ();
 b15zdnd11an1n32x5 FILLER_276_255 ();
 b15zdnd11an1n16x5 FILLER_276_287 ();
 b15zdnd11an1n04x5 FILLER_276_303 ();
 b15zdnd00an1n02x5 FILLER_276_307 ();
 b15zdnd00an1n01x5 FILLER_276_309 ();
 b15zdnd11an1n16x5 FILLER_276_321 ();
 b15zdnd11an1n08x5 FILLER_276_337 ();
 b15zdnd11an1n04x5 FILLER_276_345 ();
 b15zdnd00an1n02x5 FILLER_276_349 ();
 b15zdnd00an1n01x5 FILLER_276_351 ();
 b15zdnd11an1n08x5 FILLER_276_360 ();
 b15zdnd11an1n04x5 FILLER_276_368 ();
 b15zdnd00an1n02x5 FILLER_276_372 ();
 b15zdnd00an1n01x5 FILLER_276_374 ();
 b15zdnd11an1n32x5 FILLER_276_380 ();
 b15zdnd11an1n16x5 FILLER_276_412 ();
 b15zdnd11an1n08x5 FILLER_276_428 ();
 b15zdnd00an1n02x5 FILLER_276_436 ();
 b15zdnd00an1n01x5 FILLER_276_438 ();
 b15zdnd11an1n08x5 FILLER_276_454 ();
 b15zdnd11an1n04x5 FILLER_276_462 ();
 b15zdnd11an1n32x5 FILLER_276_478 ();
 b15zdnd11an1n08x5 FILLER_276_510 ();
 b15zdnd00an1n02x5 FILLER_276_518 ();
 b15zdnd00an1n01x5 FILLER_276_520 ();
 b15zdnd11an1n32x5 FILLER_276_526 ();
 b15zdnd11an1n16x5 FILLER_276_558 ();
 b15zdnd11an1n08x5 FILLER_276_574 ();
 b15zdnd11an1n16x5 FILLER_276_590 ();
 b15zdnd00an1n02x5 FILLER_276_606 ();
 b15zdnd11an1n32x5 FILLER_276_614 ();
 b15zdnd11an1n16x5 FILLER_276_646 ();
 b15zdnd11an1n08x5 FILLER_276_662 ();
 b15zdnd00an1n01x5 FILLER_276_670 ();
 b15zdnd11an1n32x5 FILLER_276_675 ();
 b15zdnd11an1n08x5 FILLER_276_707 ();
 b15zdnd00an1n02x5 FILLER_276_715 ();
 b15zdnd00an1n01x5 FILLER_276_717 ();
 b15zdnd11an1n16x5 FILLER_276_726 ();
 b15zdnd11an1n04x5 FILLER_276_742 ();
 b15zdnd00an1n02x5 FILLER_276_746 ();
 b15zdnd00an1n01x5 FILLER_276_748 ();
 b15zdnd11an1n16x5 FILLER_276_758 ();
 b15zdnd11an1n08x5 FILLER_276_774 ();
 b15zdnd11an1n64x5 FILLER_276_788 ();
 b15zdnd11an1n16x5 FILLER_276_852 ();
 b15zdnd11an1n08x5 FILLER_276_868 ();
 b15zdnd11an1n04x5 FILLER_276_876 ();
 b15zdnd00an1n02x5 FILLER_276_880 ();
 b15zdnd00an1n01x5 FILLER_276_882 ();
 b15zdnd11an1n08x5 FILLER_276_901 ();
 b15zdnd11an1n04x5 FILLER_276_909 ();
 b15zdnd11an1n32x5 FILLER_276_938 ();
 b15zdnd11an1n16x5 FILLER_276_970 ();
 b15zdnd11an1n04x5 FILLER_276_986 ();
 b15zdnd00an1n01x5 FILLER_276_990 ();
 b15zdnd11an1n08x5 FILLER_276_1011 ();
 b15zdnd11an1n04x5 FILLER_276_1019 ();
 b15zdnd11an1n04x5 FILLER_276_1028 ();
 b15zdnd11an1n16x5 FILLER_276_1042 ();
 b15zdnd11an1n04x5 FILLER_276_1058 ();
 b15zdnd00an1n01x5 FILLER_276_1062 ();
 b15zdnd11an1n04x5 FILLER_276_1095 ();
 b15zdnd11an1n16x5 FILLER_276_1103 ();
 b15zdnd11an1n08x5 FILLER_276_1119 ();
 b15zdnd11an1n64x5 FILLER_276_1137 ();
 b15zdnd11an1n08x5 FILLER_276_1201 ();
 b15zdnd11an1n04x5 FILLER_276_1209 ();
 b15zdnd00an1n02x5 FILLER_276_1213 ();
 b15zdnd11an1n16x5 FILLER_276_1227 ();
 b15zdnd00an1n01x5 FILLER_276_1243 ();
 b15zdnd11an1n32x5 FILLER_276_1253 ();
 b15zdnd11an1n08x5 FILLER_276_1285 ();
 b15zdnd11an1n04x5 FILLER_276_1293 ();
 b15zdnd00an1n02x5 FILLER_276_1297 ();
 b15zdnd00an1n01x5 FILLER_276_1299 ();
 b15zdnd11an1n04x5 FILLER_276_1306 ();
 b15zdnd00an1n01x5 FILLER_276_1310 ();
 b15zdnd11an1n64x5 FILLER_276_1327 ();
 b15zdnd11an1n64x5 FILLER_276_1391 ();
 b15zdnd00an1n01x5 FILLER_276_1455 ();
 b15zdnd11an1n64x5 FILLER_276_1461 ();
 b15zdnd11an1n08x5 FILLER_276_1525 ();
 b15zdnd00an1n02x5 FILLER_276_1533 ();
 b15zdnd11an1n64x5 FILLER_276_1547 ();
 b15zdnd11an1n32x5 FILLER_276_1611 ();
 b15zdnd11an1n16x5 FILLER_276_1643 ();
 b15zdnd11an1n08x5 FILLER_276_1659 ();
 b15zdnd00an1n02x5 FILLER_276_1667 ();
 b15zdnd00an1n01x5 FILLER_276_1669 ();
 b15zdnd11an1n04x5 FILLER_276_1685 ();
 b15zdnd11an1n08x5 FILLER_276_1701 ();
 b15zdnd00an1n02x5 FILLER_276_1709 ();
 b15zdnd00an1n01x5 FILLER_276_1711 ();
 b15zdnd11an1n32x5 FILLER_276_1718 ();
 b15zdnd11an1n16x5 FILLER_276_1750 ();
 b15zdnd11an1n08x5 FILLER_276_1766 ();
 b15zdnd11an1n08x5 FILLER_276_1781 ();
 b15zdnd00an1n01x5 FILLER_276_1789 ();
 b15zdnd11an1n32x5 FILLER_276_1795 ();
 b15zdnd11an1n16x5 FILLER_276_1827 ();
 b15zdnd11an1n32x5 FILLER_276_1854 ();
 b15zdnd11an1n16x5 FILLER_276_1886 ();
 b15zdnd11an1n08x5 FILLER_276_1902 ();
 b15zdnd11an1n04x5 FILLER_276_1910 ();
 b15zdnd11an1n16x5 FILLER_276_1938 ();
 b15zdnd11an1n16x5 FILLER_276_1959 ();
 b15zdnd11an1n04x5 FILLER_276_1975 ();
 b15zdnd00an1n02x5 FILLER_276_1979 ();
 b15zdnd11an1n32x5 FILLER_276_1993 ();
 b15zdnd11an1n16x5 FILLER_276_2025 ();
 b15zdnd11an1n08x5 FILLER_276_2041 ();
 b15zdnd00an1n02x5 FILLER_276_2049 ();
 b15zdnd11an1n32x5 FILLER_276_2058 ();
 b15zdnd11an1n16x5 FILLER_276_2090 ();
 b15zdnd11an1n04x5 FILLER_276_2106 ();
 b15zdnd00an1n01x5 FILLER_276_2110 ();
 b15zdnd11an1n32x5 FILLER_276_2116 ();
 b15zdnd11an1n04x5 FILLER_276_2148 ();
 b15zdnd00an1n02x5 FILLER_276_2152 ();
 b15zdnd11an1n32x5 FILLER_276_2162 ();
 b15zdnd11an1n08x5 FILLER_276_2215 ();
 b15zdnd11an1n04x5 FILLER_276_2223 ();
 b15zdnd00an1n02x5 FILLER_276_2227 ();
 b15zdnd00an1n01x5 FILLER_276_2229 ();
 b15zdnd11an1n04x5 FILLER_276_2239 ();
 b15zdnd11an1n04x5 FILLER_276_2250 ();
 b15zdnd11an1n08x5 FILLER_276_2268 ();
 b15zdnd11an1n64x5 FILLER_277_0 ();
 b15zdnd11an1n04x5 FILLER_277_64 ();
 b15zdnd00an1n02x5 FILLER_277_68 ();
 b15zdnd11an1n08x5 FILLER_277_88 ();
 b15zdnd11an1n04x5 FILLER_277_96 ();
 b15zdnd11an1n04x5 FILLER_277_114 ();
 b15zdnd00an1n01x5 FILLER_277_118 ();
 b15zdnd11an1n64x5 FILLER_277_132 ();
 b15zdnd11an1n64x5 FILLER_277_196 ();
 b15zdnd00an1n01x5 FILLER_277_260 ();
 b15zdnd11an1n32x5 FILLER_277_265 ();
 b15zdnd11an1n16x5 FILLER_277_297 ();
 b15zdnd11an1n08x5 FILLER_277_313 ();
 b15zdnd00an1n02x5 FILLER_277_321 ();
 b15zdnd11an1n16x5 FILLER_277_329 ();
 b15zdnd11an1n04x5 FILLER_277_345 ();
 b15zdnd00an1n02x5 FILLER_277_349 ();
 b15zdnd00an1n01x5 FILLER_277_351 ();
 b15zdnd11an1n04x5 FILLER_277_359 ();
 b15zdnd11an1n04x5 FILLER_277_370 ();
 b15zdnd11an1n32x5 FILLER_277_380 ();
 b15zdnd11an1n16x5 FILLER_277_412 ();
 b15zdnd00an1n01x5 FILLER_277_428 ();
 b15zdnd11an1n64x5 FILLER_277_436 ();
 b15zdnd11an1n04x5 FILLER_277_500 ();
 b15zdnd00an1n02x5 FILLER_277_504 ();
 b15zdnd11an1n04x5 FILLER_277_511 ();
 b15zdnd00an1n02x5 FILLER_277_515 ();
 b15zdnd00an1n01x5 FILLER_277_517 ();
 b15zdnd11an1n04x5 FILLER_277_524 ();
 b15zdnd11an1n64x5 FILLER_277_548 ();
 b15zdnd11an1n32x5 FILLER_277_612 ();
 b15zdnd00an1n02x5 FILLER_277_644 ();
 b15zdnd11an1n16x5 FILLER_277_652 ();
 b15zdnd00an1n02x5 FILLER_277_668 ();
 b15zdnd00an1n01x5 FILLER_277_670 ();
 b15zdnd11an1n16x5 FILLER_277_692 ();
 b15zdnd11an1n08x5 FILLER_277_708 ();
 b15zdnd00an1n02x5 FILLER_277_716 ();
 b15zdnd11an1n32x5 FILLER_277_749 ();
 b15zdnd11an1n16x5 FILLER_277_781 ();
 b15zdnd11an1n08x5 FILLER_277_797 ();
 b15zdnd00an1n01x5 FILLER_277_805 ();
 b15zdnd11an1n08x5 FILLER_277_837 ();
 b15zdnd11an1n04x5 FILLER_277_845 ();
 b15zdnd00an1n01x5 FILLER_277_849 ();
 b15zdnd11an1n04x5 FILLER_277_876 ();
 b15zdnd11an1n32x5 FILLER_277_892 ();
 b15zdnd00an1n01x5 FILLER_277_924 ();
 b15zdnd11an1n16x5 FILLER_277_956 ();
 b15zdnd11an1n08x5 FILLER_277_972 ();
 b15zdnd00an1n01x5 FILLER_277_980 ();
 b15zdnd11an1n08x5 FILLER_277_996 ();
 b15zdnd00an1n02x5 FILLER_277_1004 ();
 b15zdnd00an1n01x5 FILLER_277_1006 ();
 b15zdnd11an1n16x5 FILLER_277_1011 ();
 b15zdnd11an1n08x5 FILLER_277_1027 ();
 b15zdnd00an1n02x5 FILLER_277_1035 ();
 b15zdnd11an1n04x5 FILLER_277_1041 ();
 b15zdnd11an1n32x5 FILLER_277_1060 ();
 b15zdnd11an1n08x5 FILLER_277_1092 ();
 b15zdnd11an1n08x5 FILLER_277_1117 ();
 b15zdnd00an1n01x5 FILLER_277_1125 ();
 b15zdnd11an1n16x5 FILLER_277_1138 ();
 b15zdnd00an1n02x5 FILLER_277_1154 ();
 b15zdnd00an1n01x5 FILLER_277_1156 ();
 b15zdnd11an1n04x5 FILLER_277_1161 ();
 b15zdnd11an1n16x5 FILLER_277_1182 ();
 b15zdnd00an1n02x5 FILLER_277_1198 ();
 b15zdnd11an1n16x5 FILLER_277_1205 ();
 b15zdnd11an1n08x5 FILLER_277_1221 ();
 b15zdnd00an1n01x5 FILLER_277_1229 ();
 b15zdnd11an1n16x5 FILLER_277_1235 ();
 b15zdnd00an1n01x5 FILLER_277_1251 ();
 b15zdnd11an1n32x5 FILLER_277_1262 ();
 b15zdnd11an1n16x5 FILLER_277_1309 ();
 b15zdnd11an1n08x5 FILLER_277_1325 ();
 b15zdnd11an1n04x5 FILLER_277_1333 ();
 b15zdnd00an1n02x5 FILLER_277_1337 ();
 b15zdnd00an1n01x5 FILLER_277_1339 ();
 b15zdnd11an1n16x5 FILLER_277_1345 ();
 b15zdnd11an1n04x5 FILLER_277_1365 ();
 b15zdnd11an1n64x5 FILLER_277_1376 ();
 b15zdnd11an1n32x5 FILLER_277_1440 ();
 b15zdnd11an1n04x5 FILLER_277_1472 ();
 b15zdnd00an1n02x5 FILLER_277_1476 ();
 b15zdnd11an1n64x5 FILLER_277_1492 ();
 b15zdnd11an1n16x5 FILLER_277_1556 ();
 b15zdnd11an1n04x5 FILLER_277_1572 ();
 b15zdnd11an1n64x5 FILLER_277_1593 ();
 b15zdnd00an1n01x5 FILLER_277_1657 ();
 b15zdnd11an1n32x5 FILLER_277_1670 ();
 b15zdnd11an1n08x5 FILLER_277_1702 ();
 b15zdnd11an1n04x5 FILLER_277_1720 ();
 b15zdnd00an1n02x5 FILLER_277_1724 ();
 b15zdnd00an1n01x5 FILLER_277_1726 ();
 b15zdnd11an1n04x5 FILLER_277_1743 ();
 b15zdnd11an1n16x5 FILLER_277_1752 ();
 b15zdnd11an1n04x5 FILLER_277_1768 ();
 b15zdnd11an1n64x5 FILLER_277_1777 ();
 b15zdnd11an1n04x5 FILLER_277_1841 ();
 b15zdnd00an1n02x5 FILLER_277_1845 ();
 b15zdnd11an1n04x5 FILLER_277_1856 ();
 b15zdnd11an1n64x5 FILLER_277_1880 ();
 b15zdnd11an1n08x5 FILLER_277_1944 ();
 b15zdnd11an1n04x5 FILLER_277_1952 ();
 b15zdnd00an1n01x5 FILLER_277_1956 ();
 b15zdnd11an1n04x5 FILLER_277_1969 ();
 b15zdnd11an1n04x5 FILLER_277_1978 ();
 b15zdnd11an1n08x5 FILLER_277_1986 ();
 b15zdnd00an1n02x5 FILLER_277_1994 ();
 b15zdnd11an1n64x5 FILLER_277_2009 ();
 b15zdnd11an1n64x5 FILLER_277_2073 ();
 b15zdnd11an1n08x5 FILLER_277_2137 ();
 b15zdnd00an1n02x5 FILLER_277_2145 ();
 b15zdnd11an1n08x5 FILLER_277_2159 ();
 b15zdnd11an1n04x5 FILLER_277_2167 ();
 b15zdnd00an1n02x5 FILLER_277_2171 ();
 b15zdnd00an1n01x5 FILLER_277_2173 ();
 b15zdnd11an1n04x5 FILLER_277_2194 ();
 b15zdnd00an1n01x5 FILLER_277_2198 ();
 b15zdnd11an1n08x5 FILLER_277_2213 ();
 b15zdnd00an1n01x5 FILLER_277_2221 ();
 b15zdnd11an1n32x5 FILLER_277_2237 ();
 b15zdnd11an1n08x5 FILLER_277_2269 ();
 b15zdnd11an1n04x5 FILLER_277_2277 ();
 b15zdnd00an1n02x5 FILLER_277_2281 ();
 b15zdnd00an1n01x5 FILLER_277_2283 ();
 b15zdnd11an1n32x5 FILLER_278_8 ();
 b15zdnd11an1n08x5 FILLER_278_40 ();
 b15zdnd00an1n02x5 FILLER_278_48 ();
 b15zdnd00an1n01x5 FILLER_278_50 ();
 b15zdnd11an1n16x5 FILLER_278_60 ();
 b15zdnd11an1n08x5 FILLER_278_76 ();
 b15zdnd11an1n04x5 FILLER_278_84 ();
 b15zdnd11an1n16x5 FILLER_278_92 ();
 b15zdnd11an1n04x5 FILLER_278_108 ();
 b15zdnd00an1n02x5 FILLER_278_112 ();
 b15zdnd11an1n04x5 FILLER_278_123 ();
 b15zdnd00an1n01x5 FILLER_278_127 ();
 b15zdnd11an1n04x5 FILLER_278_140 ();
 b15zdnd00an1n01x5 FILLER_278_144 ();
 b15zdnd11an1n04x5 FILLER_278_152 ();
 b15zdnd11an1n16x5 FILLER_278_163 ();
 b15zdnd00an1n02x5 FILLER_278_179 ();
 b15zdnd11an1n16x5 FILLER_278_187 ();
 b15zdnd11an1n04x5 FILLER_278_203 ();
 b15zdnd11an1n32x5 FILLER_278_214 ();
 b15zdnd11an1n16x5 FILLER_278_246 ();
 b15zdnd00an1n01x5 FILLER_278_262 ();
 b15zdnd11an1n16x5 FILLER_278_269 ();
 b15zdnd11an1n08x5 FILLER_278_285 ();
 b15zdnd00an1n01x5 FILLER_278_293 ();
 b15zdnd11an1n64x5 FILLER_278_301 ();
 b15zdnd11an1n64x5 FILLER_278_365 ();
 b15zdnd11an1n32x5 FILLER_278_429 ();
 b15zdnd11an1n08x5 FILLER_278_468 ();
 b15zdnd11an1n04x5 FILLER_278_476 ();
 b15zdnd00an1n01x5 FILLER_278_480 ();
 b15zdnd11an1n64x5 FILLER_278_489 ();
 b15zdnd11an1n08x5 FILLER_278_553 ();
 b15zdnd11an1n04x5 FILLER_278_561 ();
 b15zdnd00an1n01x5 FILLER_278_565 ();
 b15zdnd11an1n08x5 FILLER_278_572 ();
 b15zdnd11an1n04x5 FILLER_278_580 ();
 b15zdnd00an1n02x5 FILLER_278_584 ();
 b15zdnd00an1n01x5 FILLER_278_586 ();
 b15zdnd11an1n32x5 FILLER_278_599 ();
 b15zdnd11an1n08x5 FILLER_278_631 ();
 b15zdnd11an1n04x5 FILLER_278_639 ();
 b15zdnd00an1n02x5 FILLER_278_643 ();
 b15zdnd00an1n01x5 FILLER_278_645 ();
 b15zdnd11an1n04x5 FILLER_278_650 ();
 b15zdnd00an1n01x5 FILLER_278_654 ();
 b15zdnd11an1n32x5 FILLER_278_668 ();
 b15zdnd11an1n16x5 FILLER_278_700 ();
 b15zdnd00an1n02x5 FILLER_278_716 ();
 b15zdnd11an1n16x5 FILLER_278_726 ();
 b15zdnd11an1n08x5 FILLER_278_742 ();
 b15zdnd11an1n16x5 FILLER_278_756 ();
 b15zdnd11an1n08x5 FILLER_278_772 ();
 b15zdnd11an1n64x5 FILLER_278_784 ();
 b15zdnd11an1n04x5 FILLER_278_848 ();
 b15zdnd00an1n02x5 FILLER_278_852 ();
 b15zdnd00an1n01x5 FILLER_278_854 ();
 b15zdnd11an1n32x5 FILLER_278_880 ();
 b15zdnd11an1n04x5 FILLER_278_912 ();
 b15zdnd00an1n02x5 FILLER_278_916 ();
 b15zdnd00an1n01x5 FILLER_278_918 ();
 b15zdnd11an1n16x5 FILLER_278_950 ();
 b15zdnd11an1n08x5 FILLER_278_966 ();
 b15zdnd11an1n04x5 FILLER_278_974 ();
 b15zdnd11an1n16x5 FILLER_278_985 ();
 b15zdnd11an1n08x5 FILLER_278_1001 ();
 b15zdnd00an1n02x5 FILLER_278_1009 ();
 b15zdnd00an1n01x5 FILLER_278_1011 ();
 b15zdnd11an1n16x5 FILLER_278_1016 ();
 b15zdnd00an1n02x5 FILLER_278_1032 ();
 b15zdnd11an1n32x5 FILLER_278_1038 ();
 b15zdnd11an1n16x5 FILLER_278_1070 ();
 b15zdnd11an1n08x5 FILLER_278_1086 ();
 b15zdnd00an1n01x5 FILLER_278_1094 ();
 b15zdnd11an1n32x5 FILLER_278_1103 ();
 b15zdnd11an1n16x5 FILLER_278_1135 ();
 b15zdnd11an1n04x5 FILLER_278_1151 ();
 b15zdnd00an1n02x5 FILLER_278_1155 ();
 b15zdnd11an1n08x5 FILLER_278_1166 ();
 b15zdnd00an1n02x5 FILLER_278_1174 ();
 b15zdnd11an1n04x5 FILLER_278_1194 ();
 b15zdnd11an1n16x5 FILLER_278_1203 ();
 b15zdnd11an1n08x5 FILLER_278_1219 ();
 b15zdnd00an1n02x5 FILLER_278_1227 ();
 b15zdnd11an1n08x5 FILLER_278_1234 ();
 b15zdnd11an1n04x5 FILLER_278_1242 ();
 b15zdnd00an1n02x5 FILLER_278_1246 ();
 b15zdnd00an1n01x5 FILLER_278_1248 ();
 b15zdnd11an1n16x5 FILLER_278_1256 ();
 b15zdnd00an1n02x5 FILLER_278_1272 ();
 b15zdnd11an1n16x5 FILLER_278_1278 ();
 b15zdnd11an1n04x5 FILLER_278_1294 ();
 b15zdnd00an1n02x5 FILLER_278_1298 ();
 b15zdnd11an1n32x5 FILLER_278_1311 ();
 b15zdnd11an1n04x5 FILLER_278_1343 ();
 b15zdnd00an1n01x5 FILLER_278_1347 ();
 b15zdnd11an1n04x5 FILLER_278_1358 ();
 b15zdnd11an1n32x5 FILLER_278_1377 ();
 b15zdnd11an1n16x5 FILLER_278_1409 ();
 b15zdnd11an1n08x5 FILLER_278_1425 ();
 b15zdnd11an1n16x5 FILLER_278_1445 ();
 b15zdnd11an1n04x5 FILLER_278_1461 ();
 b15zdnd11an1n04x5 FILLER_278_1471 ();
 b15zdnd11an1n08x5 FILLER_278_1480 ();
 b15zdnd00an1n01x5 FILLER_278_1488 ();
 b15zdnd11an1n08x5 FILLER_278_1500 ();
 b15zdnd11an1n04x5 FILLER_278_1508 ();
 b15zdnd00an1n01x5 FILLER_278_1512 ();
 b15zdnd11an1n04x5 FILLER_278_1525 ();
 b15zdnd00an1n01x5 FILLER_278_1529 ();
 b15zdnd11an1n04x5 FILLER_278_1535 ();
 b15zdnd00an1n02x5 FILLER_278_1539 ();
 b15zdnd11an1n04x5 FILLER_278_1547 ();
 b15zdnd00an1n02x5 FILLER_278_1551 ();
 b15zdnd11an1n04x5 FILLER_278_1560 ();
 b15zdnd11an1n64x5 FILLER_278_1570 ();
 b15zdnd11an1n16x5 FILLER_278_1634 ();
 b15zdnd00an1n01x5 FILLER_278_1650 ();
 b15zdnd11an1n08x5 FILLER_278_1660 ();
 b15zdnd00an1n01x5 FILLER_278_1668 ();
 b15zdnd11an1n64x5 FILLER_278_1680 ();
 b15zdnd00an1n02x5 FILLER_278_1744 ();
 b15zdnd00an1n01x5 FILLER_278_1746 ();
 b15zdnd11an1n08x5 FILLER_278_1756 ();
 b15zdnd11an1n04x5 FILLER_278_1764 ();
 b15zdnd11an1n04x5 FILLER_278_1777 ();
 b15zdnd00an1n02x5 FILLER_278_1781 ();
 b15zdnd00an1n01x5 FILLER_278_1783 ();
 b15zdnd11an1n64x5 FILLER_278_1797 ();
 b15zdnd11an1n32x5 FILLER_278_1861 ();
 b15zdnd11an1n04x5 FILLER_278_1893 ();
 b15zdnd00an1n02x5 FILLER_278_1897 ();
 b15zdnd00an1n01x5 FILLER_278_1899 ();
 b15zdnd11an1n16x5 FILLER_278_1926 ();
 b15zdnd11an1n64x5 FILLER_278_1954 ();
 b15zdnd11an1n64x5 FILLER_278_2018 ();
 b15zdnd11an1n32x5 FILLER_278_2082 ();
 b15zdnd00an1n02x5 FILLER_278_2114 ();
 b15zdnd00an1n01x5 FILLER_278_2116 ();
 b15zdnd11an1n16x5 FILLER_278_2122 ();
 b15zdnd11an1n04x5 FILLER_278_2138 ();
 b15zdnd11an1n04x5 FILLER_278_2148 ();
 b15zdnd00an1n02x5 FILLER_278_2152 ();
 b15zdnd11an1n64x5 FILLER_278_2162 ();
 b15zdnd11an1n32x5 FILLER_278_2226 ();
 b15zdnd11an1n16x5 FILLER_278_2258 ();
 b15zdnd00an1n02x5 FILLER_278_2274 ();
 b15zdnd11an1n32x5 FILLER_279_0 ();
 b15zdnd11an1n16x5 FILLER_279_32 ();
 b15zdnd00an1n02x5 FILLER_279_48 ();
 b15zdnd11an1n16x5 FILLER_279_56 ();
 b15zdnd11an1n08x5 FILLER_279_72 ();
 b15zdnd11an1n04x5 FILLER_279_80 ();
 b15zdnd11an1n16x5 FILLER_279_100 ();
 b15zdnd11an1n04x5 FILLER_279_116 ();
 b15zdnd00an1n01x5 FILLER_279_120 ();
 b15zdnd11an1n08x5 FILLER_279_137 ();
 b15zdnd11an1n16x5 FILLER_279_155 ();
 b15zdnd00an1n02x5 FILLER_279_171 ();
 b15zdnd11an1n16x5 FILLER_279_189 ();
 b15zdnd00an1n01x5 FILLER_279_205 ();
 b15zdnd11an1n32x5 FILLER_279_211 ();
 b15zdnd11an1n16x5 FILLER_279_243 ();
 b15zdnd00an1n02x5 FILLER_279_259 ();
 b15zdnd11an1n16x5 FILLER_279_266 ();
 b15zdnd11an1n04x5 FILLER_279_282 ();
 b15zdnd00an1n02x5 FILLER_279_286 ();
 b15zdnd00an1n01x5 FILLER_279_288 ();
 b15zdnd11an1n64x5 FILLER_279_321 ();
 b15zdnd11an1n64x5 FILLER_279_385 ();
 b15zdnd11an1n16x5 FILLER_279_449 ();
 b15zdnd11an1n04x5 FILLER_279_465 ();
 b15zdnd00an1n02x5 FILLER_279_469 ();
 b15zdnd11an1n04x5 FILLER_279_477 ();
 b15zdnd11an1n32x5 FILLER_279_486 ();
 b15zdnd11an1n04x5 FILLER_279_518 ();
 b15zdnd11an1n16x5 FILLER_279_534 ();
 b15zdnd11an1n08x5 FILLER_279_550 ();
 b15zdnd00an1n02x5 FILLER_279_558 ();
 b15zdnd11an1n04x5 FILLER_279_567 ();
 b15zdnd11an1n16x5 FILLER_279_576 ();
 b15zdnd11an1n04x5 FILLER_279_592 ();
 b15zdnd11an1n08x5 FILLER_279_611 ();
 b15zdnd00an1n02x5 FILLER_279_619 ();
 b15zdnd11an1n64x5 FILLER_279_625 ();
 b15zdnd11an1n32x5 FILLER_279_689 ();
 b15zdnd11an1n16x5 FILLER_279_721 ();
 b15zdnd11an1n08x5 FILLER_279_737 ();
 b15zdnd11an1n04x5 FILLER_279_745 ();
 b15zdnd11an1n16x5 FILLER_279_759 ();
 b15zdnd11an1n08x5 FILLER_279_775 ();
 b15zdnd11an1n04x5 FILLER_279_783 ();
 b15zdnd00an1n02x5 FILLER_279_787 ();
 b15zdnd11an1n16x5 FILLER_279_801 ();
 b15zdnd00an1n02x5 FILLER_279_817 ();
 b15zdnd11an1n04x5 FILLER_279_850 ();
 b15zdnd11an1n64x5 FILLER_279_885 ();
 b15zdnd11an1n16x5 FILLER_279_949 ();
 b15zdnd11an1n08x5 FILLER_279_965 ();
 b15zdnd00an1n01x5 FILLER_279_973 ();
 b15zdnd11an1n16x5 FILLER_279_984 ();
 b15zdnd11an1n04x5 FILLER_279_1000 ();
 b15zdnd11an1n64x5 FILLER_279_1011 ();
 b15zdnd11an1n64x5 FILLER_279_1075 ();
 b15zdnd11an1n04x5 FILLER_279_1139 ();
 b15zdnd00an1n02x5 FILLER_279_1143 ();
 b15zdnd00an1n01x5 FILLER_279_1145 ();
 b15zdnd11an1n32x5 FILLER_279_1162 ();
 b15zdnd11an1n04x5 FILLER_279_1194 ();
 b15zdnd00an1n01x5 FILLER_279_1198 ();
 b15zdnd11an1n32x5 FILLER_279_1210 ();
 b15zdnd11an1n16x5 FILLER_279_1242 ();
 b15zdnd11an1n08x5 FILLER_279_1258 ();
 b15zdnd00an1n01x5 FILLER_279_1266 ();
 b15zdnd11an1n08x5 FILLER_279_1283 ();
 b15zdnd00an1n02x5 FILLER_279_1291 ();
 b15zdnd00an1n01x5 FILLER_279_1293 ();
 b15zdnd11an1n08x5 FILLER_279_1306 ();
 b15zdnd11an1n04x5 FILLER_279_1314 ();
 b15zdnd00an1n02x5 FILLER_279_1318 ();
 b15zdnd11an1n64x5 FILLER_279_1328 ();
 b15zdnd11an1n32x5 FILLER_279_1392 ();
 b15zdnd11an1n08x5 FILLER_279_1424 ();
 b15zdnd00an1n02x5 FILLER_279_1432 ();
 b15zdnd00an1n01x5 FILLER_279_1434 ();
 b15zdnd11an1n08x5 FILLER_279_1455 ();
 b15zdnd11an1n04x5 FILLER_279_1463 ();
 b15zdnd00an1n02x5 FILLER_279_1467 ();
 b15zdnd11an1n04x5 FILLER_279_1479 ();
 b15zdnd11an1n04x5 FILLER_279_1489 ();
 b15zdnd11an1n16x5 FILLER_279_1504 ();
 b15zdnd11an1n04x5 FILLER_279_1520 ();
 b15zdnd11an1n16x5 FILLER_279_1532 ();
 b15zdnd11an1n08x5 FILLER_279_1548 ();
 b15zdnd11an1n32x5 FILLER_279_1562 ();
 b15zdnd11an1n16x5 FILLER_279_1594 ();
 b15zdnd11an1n04x5 FILLER_279_1610 ();
 b15zdnd00an1n02x5 FILLER_279_1614 ();
 b15zdnd11an1n04x5 FILLER_279_1622 ();
 b15zdnd11an1n04x5 FILLER_279_1630 ();
 b15zdnd11an1n32x5 FILLER_279_1644 ();
 b15zdnd11an1n16x5 FILLER_279_1676 ();
 b15zdnd11an1n04x5 FILLER_279_1692 ();
 b15zdnd11an1n16x5 FILLER_279_1703 ();
 b15zdnd11an1n08x5 FILLER_279_1719 ();
 b15zdnd11an1n04x5 FILLER_279_1727 ();
 b15zdnd00an1n02x5 FILLER_279_1731 ();
 b15zdnd11an1n16x5 FILLER_279_1742 ();
 b15zdnd11an1n08x5 FILLER_279_1758 ();
 b15zdnd00an1n01x5 FILLER_279_1766 ();
 b15zdnd11an1n08x5 FILLER_279_1773 ();
 b15zdnd11an1n04x5 FILLER_279_1781 ();
 b15zdnd11an1n64x5 FILLER_279_1790 ();
 b15zdnd11an1n64x5 FILLER_279_1854 ();
 b15zdnd11an1n32x5 FILLER_279_1918 ();
 b15zdnd11an1n16x5 FILLER_279_1950 ();
 b15zdnd00an1n02x5 FILLER_279_1966 ();
 b15zdnd11an1n16x5 FILLER_279_1973 ();
 b15zdnd11an1n08x5 FILLER_279_1989 ();
 b15zdnd00an1n02x5 FILLER_279_1997 ();
 b15zdnd11an1n16x5 FILLER_279_2014 ();
 b15zdnd11an1n16x5 FILLER_279_2037 ();
 b15zdnd11an1n08x5 FILLER_279_2065 ();
 b15zdnd00an1n02x5 FILLER_279_2073 ();
 b15zdnd11an1n04x5 FILLER_279_2080 ();
 b15zdnd11an1n04x5 FILLER_279_2090 ();
 b15zdnd00an1n02x5 FILLER_279_2094 ();
 b15zdnd00an1n01x5 FILLER_279_2096 ();
 b15zdnd11an1n08x5 FILLER_279_2103 ();
 b15zdnd11an1n04x5 FILLER_279_2111 ();
 b15zdnd00an1n02x5 FILLER_279_2115 ();
 b15zdnd11an1n04x5 FILLER_279_2124 ();
 b15zdnd00an1n02x5 FILLER_279_2128 ();
 b15zdnd00an1n01x5 FILLER_279_2130 ();
 b15zdnd11an1n04x5 FILLER_279_2137 ();
 b15zdnd11an1n64x5 FILLER_279_2151 ();
 b15zdnd11an1n08x5 FILLER_279_2215 ();
 b15zdnd11an1n04x5 FILLER_279_2223 ();
 b15zdnd11an1n32x5 FILLER_279_2239 ();
 b15zdnd11an1n08x5 FILLER_279_2271 ();
 b15zdnd11an1n04x5 FILLER_279_2279 ();
 b15zdnd00an1n01x5 FILLER_279_2283 ();
 b15zdnd11an1n32x5 FILLER_280_8 ();
 b15zdnd11an1n08x5 FILLER_280_40 ();
 b15zdnd11an1n08x5 FILLER_280_53 ();
 b15zdnd11an1n04x5 FILLER_280_61 ();
 b15zdnd11an1n64x5 FILLER_280_81 ();
 b15zdnd11an1n16x5 FILLER_280_145 ();
 b15zdnd11an1n08x5 FILLER_280_161 ();
 b15zdnd11an1n04x5 FILLER_280_169 ();
 b15zdnd00an1n02x5 FILLER_280_173 ();
 b15zdnd11an1n04x5 FILLER_280_182 ();
 b15zdnd11an1n08x5 FILLER_280_191 ();
 b15zdnd00an1n02x5 FILLER_280_199 ();
 b15zdnd11an1n08x5 FILLER_280_210 ();
 b15zdnd11an1n04x5 FILLER_280_218 ();
 b15zdnd00an1n02x5 FILLER_280_222 ();
 b15zdnd00an1n01x5 FILLER_280_224 ();
 b15zdnd11an1n16x5 FILLER_280_231 ();
 b15zdnd00an1n01x5 FILLER_280_247 ();
 b15zdnd11an1n16x5 FILLER_280_252 ();
 b15zdnd11an1n08x5 FILLER_280_268 ();
 b15zdnd11an1n04x5 FILLER_280_276 ();
 b15zdnd00an1n01x5 FILLER_280_280 ();
 b15zdnd11an1n04x5 FILLER_280_288 ();
 b15zdnd11an1n64x5 FILLER_280_307 ();
 b15zdnd11an1n64x5 FILLER_280_371 ();
 b15zdnd11an1n32x5 FILLER_280_435 ();
 b15zdnd11an1n04x5 FILLER_280_467 ();
 b15zdnd00an1n02x5 FILLER_280_471 ();
 b15zdnd11an1n16x5 FILLER_280_478 ();
 b15zdnd11an1n08x5 FILLER_280_494 ();
 b15zdnd00an1n02x5 FILLER_280_502 ();
 b15zdnd11an1n04x5 FILLER_280_514 ();
 b15zdnd00an1n02x5 FILLER_280_518 ();
 b15zdnd11an1n16x5 FILLER_280_540 ();
 b15zdnd11an1n16x5 FILLER_280_563 ();
 b15zdnd11an1n08x5 FILLER_280_579 ();
 b15zdnd11an1n04x5 FILLER_280_587 ();
 b15zdnd00an1n02x5 FILLER_280_591 ();
 b15zdnd11an1n04x5 FILLER_280_600 ();
 b15zdnd11an1n64x5 FILLER_280_618 ();
 b15zdnd11an1n16x5 FILLER_280_682 ();
 b15zdnd11an1n04x5 FILLER_280_698 ();
 b15zdnd00an1n02x5 FILLER_280_716 ();
 b15zdnd11an1n32x5 FILLER_280_726 ();
 b15zdnd11an1n16x5 FILLER_280_758 ();
 b15zdnd00an1n02x5 FILLER_280_774 ();
 b15zdnd11an1n64x5 FILLER_280_808 ();
 b15zdnd11an1n64x5 FILLER_280_872 ();
 b15zdnd11an1n32x5 FILLER_280_936 ();
 b15zdnd11an1n04x5 FILLER_280_968 ();
 b15zdnd11an1n16x5 FILLER_280_982 ();
 b15zdnd11an1n08x5 FILLER_280_998 ();
 b15zdnd11an1n04x5 FILLER_280_1006 ();
 b15zdnd00an1n02x5 FILLER_280_1010 ();
 b15zdnd11an1n32x5 FILLER_280_1018 ();
 b15zdnd11an1n16x5 FILLER_280_1050 ();
 b15zdnd11an1n08x5 FILLER_280_1066 ();
 b15zdnd11an1n04x5 FILLER_280_1074 ();
 b15zdnd00an1n02x5 FILLER_280_1078 ();
 b15zdnd11an1n04x5 FILLER_280_1090 ();
 b15zdnd11an1n32x5 FILLER_280_1099 ();
 b15zdnd11an1n16x5 FILLER_280_1131 ();
 b15zdnd00an1n02x5 FILLER_280_1147 ();
 b15zdnd11an1n64x5 FILLER_280_1159 ();
 b15zdnd11an1n64x5 FILLER_280_1223 ();
 b15zdnd11an1n32x5 FILLER_280_1287 ();
 b15zdnd00an1n02x5 FILLER_280_1319 ();
 b15zdnd11an1n04x5 FILLER_280_1330 ();
 b15zdnd11an1n64x5 FILLER_280_1347 ();
 b15zdnd11an1n16x5 FILLER_280_1411 ();
 b15zdnd11an1n04x5 FILLER_280_1427 ();
 b15zdnd00an1n01x5 FILLER_280_1431 ();
 b15zdnd11an1n32x5 FILLER_280_1457 ();
 b15zdnd11an1n08x5 FILLER_280_1489 ();
 b15zdnd11an1n04x5 FILLER_280_1497 ();
 b15zdnd00an1n02x5 FILLER_280_1501 ();
 b15zdnd11an1n64x5 FILLER_280_1514 ();
 b15zdnd11an1n16x5 FILLER_280_1578 ();
 b15zdnd00an1n02x5 FILLER_280_1594 ();
 b15zdnd11an1n04x5 FILLER_280_1602 ();
 b15zdnd00an1n02x5 FILLER_280_1606 ();
 b15zdnd11an1n04x5 FILLER_280_1620 ();
 b15zdnd11an1n32x5 FILLER_280_1628 ();
 b15zdnd11an1n04x5 FILLER_280_1660 ();
 b15zdnd00an1n01x5 FILLER_280_1664 ();
 b15zdnd11an1n16x5 FILLER_280_1670 ();
 b15zdnd00an1n02x5 FILLER_280_1686 ();
 b15zdnd00an1n01x5 FILLER_280_1688 ();
 b15zdnd11an1n16x5 FILLER_280_1695 ();
 b15zdnd00an1n02x5 FILLER_280_1711 ();
 b15zdnd00an1n01x5 FILLER_280_1713 ();
 b15zdnd11an1n32x5 FILLER_280_1719 ();
 b15zdnd11an1n04x5 FILLER_280_1751 ();
 b15zdnd00an1n02x5 FILLER_280_1755 ();
 b15zdnd00an1n01x5 FILLER_280_1757 ();
 b15zdnd11an1n16x5 FILLER_280_1778 ();
 b15zdnd11an1n04x5 FILLER_280_1794 ();
 b15zdnd00an1n02x5 FILLER_280_1798 ();
 b15zdnd11an1n64x5 FILLER_280_1807 ();
 b15zdnd11an1n04x5 FILLER_280_1871 ();
 b15zdnd11an1n04x5 FILLER_280_1893 ();
 b15zdnd11an1n16x5 FILLER_280_1903 ();
 b15zdnd11an1n04x5 FILLER_280_1919 ();
 b15zdnd00an1n02x5 FILLER_280_1923 ();
 b15zdnd11an1n64x5 FILLER_280_1934 ();
 b15zdnd11an1n16x5 FILLER_280_2002 ();
 b15zdnd11an1n08x5 FILLER_280_2018 ();
 b15zdnd00an1n02x5 FILLER_280_2026 ();
 b15zdnd00an1n01x5 FILLER_280_2028 ();
 b15zdnd11an1n04x5 FILLER_280_2060 ();
 b15zdnd11an1n04x5 FILLER_280_2076 ();
 b15zdnd00an1n02x5 FILLER_280_2080 ();
 b15zdnd00an1n01x5 FILLER_280_2082 ();
 b15zdnd11an1n32x5 FILLER_280_2094 ();
 b15zdnd11an1n16x5 FILLER_280_2126 ();
 b15zdnd11an1n08x5 FILLER_280_2142 ();
 b15zdnd11an1n04x5 FILLER_280_2150 ();
 b15zdnd11an1n08x5 FILLER_280_2162 ();
 b15zdnd11an1n04x5 FILLER_280_2170 ();
 b15zdnd00an1n01x5 FILLER_280_2174 ();
 b15zdnd11an1n08x5 FILLER_280_2187 ();
 b15zdnd11an1n04x5 FILLER_280_2195 ();
 b15zdnd00an1n02x5 FILLER_280_2199 ();
 b15zdnd11an1n16x5 FILLER_280_2208 ();
 b15zdnd11an1n08x5 FILLER_280_2224 ();
 b15zdnd11an1n04x5 FILLER_280_2232 ();
 b15zdnd00an1n01x5 FILLER_280_2236 ();
 b15zdnd11an1n32x5 FILLER_280_2242 ();
 b15zdnd00an1n02x5 FILLER_280_2274 ();
 b15zdnd11an1n32x5 FILLER_281_0 ();
 b15zdnd11an1n08x5 FILLER_281_32 ();
 b15zdnd00an1n02x5 FILLER_281_40 ();
 b15zdnd11an1n08x5 FILLER_281_60 ();
 b15zdnd11an1n04x5 FILLER_281_68 ();
 b15zdnd00an1n02x5 FILLER_281_72 ();
 b15zdnd00an1n01x5 FILLER_281_74 ();
 b15zdnd11an1n16x5 FILLER_281_84 ();
 b15zdnd11an1n04x5 FILLER_281_100 ();
 b15zdnd00an1n01x5 FILLER_281_104 ();
 b15zdnd11an1n64x5 FILLER_281_116 ();
 b15zdnd11an1n64x5 FILLER_281_180 ();
 b15zdnd11an1n04x5 FILLER_281_244 ();
 b15zdnd00an1n02x5 FILLER_281_248 ();
 b15zdnd11an1n04x5 FILLER_281_255 ();
 b15zdnd11an1n16x5 FILLER_281_271 ();
 b15zdnd11an1n04x5 FILLER_281_287 ();
 b15zdnd00an1n01x5 FILLER_281_291 ();
 b15zdnd11an1n16x5 FILLER_281_298 ();
 b15zdnd00an1n01x5 FILLER_281_314 ();
 b15zdnd11an1n04x5 FILLER_281_320 ();
 b15zdnd00an1n01x5 FILLER_281_324 ();
 b15zdnd11an1n04x5 FILLER_281_329 ();
 b15zdnd00an1n02x5 FILLER_281_333 ();
 b15zdnd00an1n01x5 FILLER_281_335 ();
 b15zdnd11an1n08x5 FILLER_281_341 ();
 b15zdnd00an1n02x5 FILLER_281_349 ();
 b15zdnd11an1n64x5 FILLER_281_361 ();
 b15zdnd11an1n08x5 FILLER_281_425 ();
 b15zdnd11an1n04x5 FILLER_281_433 ();
 b15zdnd00an1n02x5 FILLER_281_437 ();
 b15zdnd11an1n32x5 FILLER_281_449 ();
 b15zdnd11an1n16x5 FILLER_281_481 ();
 b15zdnd11an1n08x5 FILLER_281_497 ();
 b15zdnd00an1n02x5 FILLER_281_505 ();
 b15zdnd11an1n04x5 FILLER_281_525 ();
 b15zdnd00an1n02x5 FILLER_281_529 ();
 b15zdnd11an1n64x5 FILLER_281_539 ();
 b15zdnd11an1n08x5 FILLER_281_603 ();
 b15zdnd00an1n01x5 FILLER_281_611 ();
 b15zdnd11an1n64x5 FILLER_281_618 ();
 b15zdnd11an1n16x5 FILLER_281_682 ();
 b15zdnd11an1n08x5 FILLER_281_698 ();
 b15zdnd11an1n04x5 FILLER_281_706 ();
 b15zdnd11an1n08x5 FILLER_281_732 ();
 b15zdnd11an1n04x5 FILLER_281_740 ();
 b15zdnd11an1n32x5 FILLER_281_756 ();
 b15zdnd11an1n04x5 FILLER_281_788 ();
 b15zdnd00an1n01x5 FILLER_281_792 ();
 b15zdnd11an1n64x5 FILLER_281_798 ();
 b15zdnd11an1n16x5 FILLER_281_862 ();
 b15zdnd11an1n08x5 FILLER_281_878 ();
 b15zdnd00an1n02x5 FILLER_281_886 ();
 b15zdnd11an1n04x5 FILLER_281_903 ();
 b15zdnd11an1n32x5 FILLER_281_933 ();
 b15zdnd11an1n16x5 FILLER_281_965 ();
 b15zdnd00an1n01x5 FILLER_281_981 ();
 b15zdnd11an1n64x5 FILLER_281_994 ();
 b15zdnd11an1n32x5 FILLER_281_1058 ();
 b15zdnd11an1n04x5 FILLER_281_1090 ();
 b15zdnd11an1n04x5 FILLER_281_1103 ();
 b15zdnd11an1n08x5 FILLER_281_1115 ();
 b15zdnd00an1n02x5 FILLER_281_1123 ();
 b15zdnd00an1n01x5 FILLER_281_1125 ();
 b15zdnd11an1n64x5 FILLER_281_1134 ();
 b15zdnd11an1n08x5 FILLER_281_1198 ();
 b15zdnd00an1n02x5 FILLER_281_1206 ();
 b15zdnd00an1n01x5 FILLER_281_1208 ();
 b15zdnd11an1n16x5 FILLER_281_1214 ();
 b15zdnd11an1n08x5 FILLER_281_1230 ();
 b15zdnd11an1n04x5 FILLER_281_1238 ();
 b15zdnd00an1n02x5 FILLER_281_1242 ();
 b15zdnd00an1n01x5 FILLER_281_1244 ();
 b15zdnd11an1n64x5 FILLER_281_1251 ();
 b15zdnd11an1n08x5 FILLER_281_1315 ();
 b15zdnd11an1n04x5 FILLER_281_1323 ();
 b15zdnd11an1n16x5 FILLER_281_1334 ();
 b15zdnd11an1n04x5 FILLER_281_1350 ();
 b15zdnd00an1n01x5 FILLER_281_1354 ();
 b15zdnd11an1n64x5 FILLER_281_1376 ();
 b15zdnd11an1n64x5 FILLER_281_1440 ();
 b15zdnd11an1n64x5 FILLER_281_1504 ();
 b15zdnd11an1n08x5 FILLER_281_1568 ();
 b15zdnd11an1n04x5 FILLER_281_1576 ();
 b15zdnd00an1n02x5 FILLER_281_1580 ();
 b15zdnd11an1n32x5 FILLER_281_1588 ();
 b15zdnd00an1n01x5 FILLER_281_1620 ();
 b15zdnd11an1n32x5 FILLER_281_1629 ();
 b15zdnd00an1n01x5 FILLER_281_1661 ();
 b15zdnd11an1n16x5 FILLER_281_1668 ();
 b15zdnd00an1n01x5 FILLER_281_1684 ();
 b15zdnd11an1n64x5 FILLER_281_1695 ();
 b15zdnd11an1n16x5 FILLER_281_1759 ();
 b15zdnd11an1n08x5 FILLER_281_1775 ();
 b15zdnd00an1n02x5 FILLER_281_1783 ();
 b15zdnd00an1n01x5 FILLER_281_1785 ();
 b15zdnd11an1n04x5 FILLER_281_1791 ();
 b15zdnd00an1n02x5 FILLER_281_1795 ();
 b15zdnd00an1n01x5 FILLER_281_1797 ();
 b15zdnd11an1n64x5 FILLER_281_1804 ();
 b15zdnd11an1n16x5 FILLER_281_1868 ();
 b15zdnd11an1n04x5 FILLER_281_1884 ();
 b15zdnd00an1n02x5 FILLER_281_1888 ();
 b15zdnd11an1n16x5 FILLER_281_1908 ();
 b15zdnd11an1n08x5 FILLER_281_1924 ();
 b15zdnd11an1n04x5 FILLER_281_1938 ();
 b15zdnd11an1n04x5 FILLER_281_1951 ();
 b15zdnd11an1n04x5 FILLER_281_1961 ();
 b15zdnd11an1n64x5 FILLER_281_1971 ();
 b15zdnd11an1n04x5 FILLER_281_2035 ();
 b15zdnd00an1n02x5 FILLER_281_2039 ();
 b15zdnd00an1n01x5 FILLER_281_2041 ();
 b15zdnd11an1n04x5 FILLER_281_2047 ();
 b15zdnd00an1n01x5 FILLER_281_2051 ();
 b15zdnd11an1n16x5 FILLER_281_2058 ();
 b15zdnd00an1n01x5 FILLER_281_2074 ();
 b15zdnd11an1n64x5 FILLER_281_2081 ();
 b15zdnd11an1n08x5 FILLER_281_2145 ();
 b15zdnd00an1n02x5 FILLER_281_2153 ();
 b15zdnd00an1n01x5 FILLER_281_2155 ();
 b15zdnd11an1n08x5 FILLER_281_2166 ();
 b15zdnd11an1n04x5 FILLER_281_2174 ();
 b15zdnd11an1n64x5 FILLER_281_2183 ();
 b15zdnd11an1n32x5 FILLER_281_2247 ();
 b15zdnd11an1n04x5 FILLER_281_2279 ();
 b15zdnd00an1n01x5 FILLER_281_2283 ();
 b15zdnd11an1n64x5 FILLER_282_8 ();
 b15zdnd11an1n04x5 FILLER_282_72 ();
 b15zdnd00an1n01x5 FILLER_282_76 ();
 b15zdnd11an1n32x5 FILLER_282_82 ();
 b15zdnd00an1n02x5 FILLER_282_114 ();
 b15zdnd11an1n16x5 FILLER_282_120 ();
 b15zdnd11an1n32x5 FILLER_282_145 ();
 b15zdnd11an1n16x5 FILLER_282_177 ();
 b15zdnd11an1n08x5 FILLER_282_193 ();
 b15zdnd00an1n02x5 FILLER_282_201 ();
 b15zdnd00an1n01x5 FILLER_282_203 ();
 b15zdnd11an1n64x5 FILLER_282_212 ();
 b15zdnd11an1n16x5 FILLER_282_276 ();
 b15zdnd11an1n04x5 FILLER_282_292 ();
 b15zdnd11an1n32x5 FILLER_282_302 ();
 b15zdnd11an1n04x5 FILLER_282_334 ();
 b15zdnd11an1n64x5 FILLER_282_342 ();
 b15zdnd11an1n32x5 FILLER_282_406 ();
 b15zdnd11an1n04x5 FILLER_282_438 ();
 b15zdnd00an1n02x5 FILLER_282_442 ();
 b15zdnd00an1n01x5 FILLER_282_444 ();
 b15zdnd11an1n64x5 FILLER_282_455 ();
 b15zdnd11an1n16x5 FILLER_282_550 ();
 b15zdnd00an1n01x5 FILLER_282_566 ();
 b15zdnd11an1n32x5 FILLER_282_574 ();
 b15zdnd11an1n16x5 FILLER_282_606 ();
 b15zdnd11an1n08x5 FILLER_282_622 ();
 b15zdnd11an1n04x5 FILLER_282_630 ();
 b15zdnd00an1n02x5 FILLER_282_634 ();
 b15zdnd00an1n01x5 FILLER_282_636 ();
 b15zdnd11an1n16x5 FILLER_282_646 ();
 b15zdnd11an1n08x5 FILLER_282_662 ();
 b15zdnd11an1n04x5 FILLER_282_676 ();
 b15zdnd11an1n08x5 FILLER_282_692 ();
 b15zdnd00an1n02x5 FILLER_282_700 ();
 b15zdnd11an1n04x5 FILLER_282_711 ();
 b15zdnd00an1n02x5 FILLER_282_715 ();
 b15zdnd00an1n01x5 FILLER_282_717 ();
 b15zdnd11an1n08x5 FILLER_282_726 ();
 b15zdnd00an1n02x5 FILLER_282_734 ();
 b15zdnd00an1n01x5 FILLER_282_736 ();
 b15zdnd11an1n04x5 FILLER_282_742 ();
 b15zdnd11an1n32x5 FILLER_282_753 ();
 b15zdnd11an1n04x5 FILLER_282_785 ();
 b15zdnd11an1n64x5 FILLER_282_797 ();
 b15zdnd11an1n08x5 FILLER_282_861 ();
 b15zdnd00an1n02x5 FILLER_282_869 ();
 b15zdnd11an1n64x5 FILLER_282_880 ();
 b15zdnd11an1n16x5 FILLER_282_944 ();
 b15zdnd11an1n08x5 FILLER_282_960 ();
 b15zdnd11an1n04x5 FILLER_282_968 ();
 b15zdnd00an1n02x5 FILLER_282_972 ();
 b15zdnd00an1n01x5 FILLER_282_974 ();
 b15zdnd11an1n64x5 FILLER_282_982 ();
 b15zdnd11an1n16x5 FILLER_282_1046 ();
 b15zdnd11an1n08x5 FILLER_282_1062 ();
 b15zdnd11an1n04x5 FILLER_282_1070 ();
 b15zdnd00an1n02x5 FILLER_282_1074 ();
 b15zdnd00an1n01x5 FILLER_282_1076 ();
 b15zdnd11an1n04x5 FILLER_282_1082 ();
 b15zdnd00an1n02x5 FILLER_282_1086 ();
 b15zdnd00an1n01x5 FILLER_282_1088 ();
 b15zdnd11an1n32x5 FILLER_282_1095 ();
 b15zdnd11an1n08x5 FILLER_282_1127 ();
 b15zdnd11an1n04x5 FILLER_282_1135 ();
 b15zdnd11an1n08x5 FILLER_282_1151 ();
 b15zdnd11an1n04x5 FILLER_282_1159 ();
 b15zdnd11an1n32x5 FILLER_282_1169 ();
 b15zdnd11an1n08x5 FILLER_282_1201 ();
 b15zdnd00an1n01x5 FILLER_282_1209 ();
 b15zdnd11an1n16x5 FILLER_282_1215 ();
 b15zdnd11an1n04x5 FILLER_282_1231 ();
 b15zdnd11an1n16x5 FILLER_282_1244 ();
 b15zdnd11an1n04x5 FILLER_282_1260 ();
 b15zdnd00an1n02x5 FILLER_282_1264 ();
 b15zdnd00an1n01x5 FILLER_282_1266 ();
 b15zdnd11an1n32x5 FILLER_282_1275 ();
 b15zdnd11an1n16x5 FILLER_282_1307 ();
 b15zdnd00an1n02x5 FILLER_282_1323 ();
 b15zdnd00an1n01x5 FILLER_282_1325 ();
 b15zdnd11an1n16x5 FILLER_282_1331 ();
 b15zdnd11an1n08x5 FILLER_282_1347 ();
 b15zdnd11an1n04x5 FILLER_282_1355 ();
 b15zdnd00an1n02x5 FILLER_282_1359 ();
 b15zdnd00an1n01x5 FILLER_282_1361 ();
 b15zdnd11an1n64x5 FILLER_282_1366 ();
 b15zdnd11an1n32x5 FILLER_282_1430 ();
 b15zdnd11an1n16x5 FILLER_282_1462 ();
 b15zdnd11an1n32x5 FILLER_282_1486 ();
 b15zdnd11an1n16x5 FILLER_282_1518 ();
 b15zdnd11an1n04x5 FILLER_282_1534 ();
 b15zdnd00an1n01x5 FILLER_282_1538 ();
 b15zdnd11an1n08x5 FILLER_282_1545 ();
 b15zdnd00an1n02x5 FILLER_282_1553 ();
 b15zdnd11an1n04x5 FILLER_282_1563 ();
 b15zdnd11an1n64x5 FILLER_282_1573 ();
 b15zdnd11an1n16x5 FILLER_282_1637 ();
 b15zdnd11an1n08x5 FILLER_282_1653 ();
 b15zdnd00an1n01x5 FILLER_282_1661 ();
 b15zdnd11an1n64x5 FILLER_282_1670 ();
 b15zdnd11an1n64x5 FILLER_282_1734 ();
 b15zdnd11an1n64x5 FILLER_282_1798 ();
 b15zdnd11an1n16x5 FILLER_282_1862 ();
 b15zdnd11an1n04x5 FILLER_282_1878 ();
 b15zdnd00an1n01x5 FILLER_282_1882 ();
 b15zdnd11an1n04x5 FILLER_282_1914 ();
 b15zdnd11an1n04x5 FILLER_282_1944 ();
 b15zdnd00an1n02x5 FILLER_282_1948 ();
 b15zdnd11an1n04x5 FILLER_282_1956 ();
 b15zdnd11an1n16x5 FILLER_282_1972 ();
 b15zdnd11an1n08x5 FILLER_282_1988 ();
 b15zdnd11an1n64x5 FILLER_282_2006 ();
 b15zdnd11an1n32x5 FILLER_282_2070 ();
 b15zdnd11an1n16x5 FILLER_282_2102 ();
 b15zdnd11an1n04x5 FILLER_282_2118 ();
 b15zdnd11an1n04x5 FILLER_282_2136 ();
 b15zdnd00an1n01x5 FILLER_282_2140 ();
 b15zdnd11an1n04x5 FILLER_282_2148 ();
 b15zdnd00an1n02x5 FILLER_282_2152 ();
 b15zdnd11an1n16x5 FILLER_282_2162 ();
 b15zdnd11an1n04x5 FILLER_282_2178 ();
 b15zdnd00an1n02x5 FILLER_282_2182 ();
 b15zdnd00an1n01x5 FILLER_282_2184 ();
 b15zdnd11an1n04x5 FILLER_282_2199 ();
 b15zdnd11an1n04x5 FILLER_282_2212 ();
 b15zdnd11an1n08x5 FILLER_282_2226 ();
 b15zdnd00an1n01x5 FILLER_282_2234 ();
 b15zdnd11an1n32x5 FILLER_282_2241 ();
 b15zdnd00an1n02x5 FILLER_282_2273 ();
 b15zdnd00an1n01x5 FILLER_282_2275 ();
 b15zdnd11an1n32x5 FILLER_283_0 ();
 b15zdnd11an1n08x5 FILLER_283_32 ();
 b15zdnd11an1n16x5 FILLER_283_58 ();
 b15zdnd11an1n08x5 FILLER_283_74 ();
 b15zdnd11an1n08x5 FILLER_283_92 ();
 b15zdnd00an1n01x5 FILLER_283_100 ();
 b15zdnd11an1n32x5 FILLER_283_111 ();
 b15zdnd00an1n01x5 FILLER_283_143 ();
 b15zdnd11an1n32x5 FILLER_283_156 ();
 b15zdnd11an1n08x5 FILLER_283_188 ();
 b15zdnd11an1n04x5 FILLER_283_196 ();
 b15zdnd00an1n02x5 FILLER_283_200 ();
 b15zdnd11an1n04x5 FILLER_283_212 ();
 b15zdnd11an1n64x5 FILLER_283_220 ();
 b15zdnd11an1n32x5 FILLER_283_284 ();
 b15zdnd11an1n08x5 FILLER_283_316 ();
 b15zdnd00an1n01x5 FILLER_283_324 ();
 b15zdnd11an1n16x5 FILLER_283_331 ();
 b15zdnd11an1n08x5 FILLER_283_347 ();
 b15zdnd11an1n64x5 FILLER_283_360 ();
 b15zdnd00an1n02x5 FILLER_283_424 ();
 b15zdnd00an1n01x5 FILLER_283_426 ();
 b15zdnd11an1n04x5 FILLER_283_436 ();
 b15zdnd11an1n64x5 FILLER_283_448 ();
 b15zdnd11an1n16x5 FILLER_283_512 ();
 b15zdnd11an1n04x5 FILLER_283_528 ();
 b15zdnd00an1n02x5 FILLER_283_532 ();
 b15zdnd11an1n04x5 FILLER_283_547 ();
 b15zdnd00an1n01x5 FILLER_283_551 ();
 b15zdnd11an1n04x5 FILLER_283_558 ();
 b15zdnd11an1n32x5 FILLER_283_569 ();
 b15zdnd11an1n08x5 FILLER_283_601 ();
 b15zdnd11an1n32x5 FILLER_283_619 ();
 b15zdnd11an1n16x5 FILLER_283_651 ();
 b15zdnd11an1n04x5 FILLER_283_667 ();
 b15zdnd11an1n16x5 FILLER_283_685 ();
 b15zdnd11an1n04x5 FILLER_283_701 ();
 b15zdnd00an1n02x5 FILLER_283_705 ();
 b15zdnd11an1n04x5 FILLER_283_727 ();
 b15zdnd11an1n32x5 FILLER_283_737 ();
 b15zdnd00an1n02x5 FILLER_283_769 ();
 b15zdnd11an1n16x5 FILLER_283_781 ();
 b15zdnd11an1n08x5 FILLER_283_797 ();
 b15zdnd00an1n02x5 FILLER_283_805 ();
 b15zdnd11an1n16x5 FILLER_283_814 ();
 b15zdnd00an1n01x5 FILLER_283_830 ();
 b15zdnd11an1n16x5 FILLER_283_846 ();
 b15zdnd11an1n08x5 FILLER_283_862 ();
 b15zdnd11an1n04x5 FILLER_283_870 ();
 b15zdnd11an1n64x5 FILLER_283_889 ();
 b15zdnd11an1n32x5 FILLER_283_953 ();
 b15zdnd11an1n16x5 FILLER_283_985 ();
 b15zdnd00an1n02x5 FILLER_283_1001 ();
 b15zdnd11an1n08x5 FILLER_283_1009 ();
 b15zdnd11an1n04x5 FILLER_283_1017 ();
 b15zdnd00an1n02x5 FILLER_283_1021 ();
 b15zdnd11an1n04x5 FILLER_283_1028 ();
 b15zdnd11an1n04x5 FILLER_283_1036 ();
 b15zdnd00an1n01x5 FILLER_283_1040 ();
 b15zdnd11an1n16x5 FILLER_283_1053 ();
 b15zdnd11an1n08x5 FILLER_283_1069 ();
 b15zdnd11an1n04x5 FILLER_283_1077 ();
 b15zdnd00an1n02x5 FILLER_283_1081 ();
 b15zdnd11an1n32x5 FILLER_283_1093 ();
 b15zdnd11an1n04x5 FILLER_283_1125 ();
 b15zdnd00an1n02x5 FILLER_283_1129 ();
 b15zdnd00an1n01x5 FILLER_283_1131 ();
 b15zdnd11an1n04x5 FILLER_283_1146 ();
 b15zdnd00an1n02x5 FILLER_283_1150 ();
 b15zdnd11an1n04x5 FILLER_283_1157 ();
 b15zdnd11an1n04x5 FILLER_283_1167 ();
 b15zdnd11an1n16x5 FILLER_283_1179 ();
 b15zdnd11an1n08x5 FILLER_283_1195 ();
 b15zdnd11an1n04x5 FILLER_283_1203 ();
 b15zdnd00an1n02x5 FILLER_283_1207 ();
 b15zdnd00an1n01x5 FILLER_283_1209 ();
 b15zdnd11an1n16x5 FILLER_283_1214 ();
 b15zdnd11an1n04x5 FILLER_283_1230 ();
 b15zdnd00an1n02x5 FILLER_283_1234 ();
 b15zdnd00an1n01x5 FILLER_283_1236 ();
 b15zdnd11an1n08x5 FILLER_283_1249 ();
 b15zdnd11an1n16x5 FILLER_283_1273 ();
 b15zdnd11an1n08x5 FILLER_283_1289 ();
 b15zdnd00an1n01x5 FILLER_283_1297 ();
 b15zdnd11an1n64x5 FILLER_283_1310 ();
 b15zdnd11an1n16x5 FILLER_283_1374 ();
 b15zdnd11an1n04x5 FILLER_283_1390 ();
 b15zdnd00an1n02x5 FILLER_283_1394 ();
 b15zdnd00an1n01x5 FILLER_283_1396 ();
 b15zdnd11an1n08x5 FILLER_283_1417 ();
 b15zdnd11an1n04x5 FILLER_283_1425 ();
 b15zdnd00an1n01x5 FILLER_283_1429 ();
 b15zdnd11an1n04x5 FILLER_283_1446 ();
 b15zdnd11an1n04x5 FILLER_283_1455 ();
 b15zdnd11an1n64x5 FILLER_283_1483 ();
 b15zdnd11an1n16x5 FILLER_283_1547 ();
 b15zdnd00an1n01x5 FILLER_283_1563 ();
 b15zdnd11an1n08x5 FILLER_283_1570 ();
 b15zdnd11an1n04x5 FILLER_283_1589 ();
 b15zdnd11an1n64x5 FILLER_283_1603 ();
 b15zdnd11an1n32x5 FILLER_283_1667 ();
 b15zdnd11an1n08x5 FILLER_283_1699 ();
 b15zdnd11an1n04x5 FILLER_283_1707 ();
 b15zdnd00an1n02x5 FILLER_283_1711 ();
 b15zdnd00an1n01x5 FILLER_283_1713 ();
 b15zdnd11an1n04x5 FILLER_283_1721 ();
 b15zdnd11an1n32x5 FILLER_283_1730 ();
 b15zdnd00an1n01x5 FILLER_283_1762 ();
 b15zdnd11an1n04x5 FILLER_283_1773 ();
 b15zdnd11an1n16x5 FILLER_283_1787 ();
 b15zdnd11an1n64x5 FILLER_283_1807 ();
 b15zdnd11an1n64x5 FILLER_283_1871 ();
 b15zdnd11an1n04x5 FILLER_283_1947 ();
 b15zdnd11an1n32x5 FILLER_283_1956 ();
 b15zdnd11an1n08x5 FILLER_283_1988 ();
 b15zdnd00an1n01x5 FILLER_283_1996 ();
 b15zdnd11an1n04x5 FILLER_283_2009 ();
 b15zdnd00an1n02x5 FILLER_283_2013 ();
 b15zdnd00an1n01x5 FILLER_283_2015 ();
 b15zdnd11an1n08x5 FILLER_283_2025 ();
 b15zdnd11an1n64x5 FILLER_283_2039 ();
 b15zdnd11an1n04x5 FILLER_283_2103 ();
 b15zdnd00an1n02x5 FILLER_283_2107 ();
 b15zdnd00an1n01x5 FILLER_283_2109 ();
 b15zdnd11an1n16x5 FILLER_283_2114 ();
 b15zdnd11an1n08x5 FILLER_283_2130 ();
 b15zdnd11an1n04x5 FILLER_283_2138 ();
 b15zdnd00an1n02x5 FILLER_283_2142 ();
 b15zdnd11an1n32x5 FILLER_283_2162 ();
 b15zdnd11an1n08x5 FILLER_283_2194 ();
 b15zdnd11an1n04x5 FILLER_283_2202 ();
 b15zdnd00an1n02x5 FILLER_283_2206 ();
 b15zdnd00an1n01x5 FILLER_283_2208 ();
 b15zdnd11an1n16x5 FILLER_283_2215 ();
 b15zdnd00an1n01x5 FILLER_283_2231 ();
 b15zdnd11an1n32x5 FILLER_283_2238 ();
 b15zdnd11an1n08x5 FILLER_283_2270 ();
 b15zdnd11an1n04x5 FILLER_283_2278 ();
 b15zdnd00an1n02x5 FILLER_283_2282 ();
 b15zdnd11an1n64x5 FILLER_284_8 ();
 b15zdnd11an1n08x5 FILLER_284_72 ();
 b15zdnd11an1n04x5 FILLER_284_80 ();
 b15zdnd11an1n08x5 FILLER_284_90 ();
 b15zdnd11an1n04x5 FILLER_284_98 ();
 b15zdnd00an1n02x5 FILLER_284_102 ();
 b15zdnd11an1n32x5 FILLER_284_110 ();
 b15zdnd11an1n04x5 FILLER_284_142 ();
 b15zdnd00an1n02x5 FILLER_284_146 ();
 b15zdnd11an1n04x5 FILLER_284_160 ();
 b15zdnd11an1n04x5 FILLER_284_172 ();
 b15zdnd11an1n32x5 FILLER_284_181 ();
 b15zdnd11an1n08x5 FILLER_284_213 ();
 b15zdnd11an1n04x5 FILLER_284_221 ();
 b15zdnd00an1n02x5 FILLER_284_225 ();
 b15zdnd00an1n01x5 FILLER_284_227 ();
 b15zdnd11an1n04x5 FILLER_284_235 ();
 b15zdnd11an1n64x5 FILLER_284_248 ();
 b15zdnd11an1n32x5 FILLER_284_312 ();
 b15zdnd11an1n08x5 FILLER_284_344 ();
 b15zdnd00an1n01x5 FILLER_284_352 ();
 b15zdnd11an1n64x5 FILLER_284_363 ();
 b15zdnd11an1n08x5 FILLER_284_427 ();
 b15zdnd00an1n01x5 FILLER_284_435 ();
 b15zdnd11an1n16x5 FILLER_284_450 ();
 b15zdnd00an1n02x5 FILLER_284_466 ();
 b15zdnd11an1n04x5 FILLER_284_474 ();
 b15zdnd11an1n32x5 FILLER_284_483 ();
 b15zdnd11an1n16x5 FILLER_284_515 ();
 b15zdnd11an1n08x5 FILLER_284_531 ();
 b15zdnd00an1n02x5 FILLER_284_539 ();
 b15zdnd00an1n01x5 FILLER_284_541 ();
 b15zdnd11an1n64x5 FILLER_284_557 ();
 b15zdnd11an1n08x5 FILLER_284_621 ();
 b15zdnd11an1n04x5 FILLER_284_629 ();
 b15zdnd00an1n02x5 FILLER_284_633 ();
 b15zdnd11an1n32x5 FILLER_284_642 ();
 b15zdnd11an1n16x5 FILLER_284_674 ();
 b15zdnd11an1n08x5 FILLER_284_690 ();
 b15zdnd11an1n04x5 FILLER_284_698 ();
 b15zdnd00an1n01x5 FILLER_284_702 ();
 b15zdnd00an1n02x5 FILLER_284_716 ();
 b15zdnd11an1n32x5 FILLER_284_726 ();
 b15zdnd11an1n16x5 FILLER_284_758 ();
 b15zdnd11an1n04x5 FILLER_284_774 ();
 b15zdnd11an1n04x5 FILLER_284_794 ();
 b15zdnd11an1n32x5 FILLER_284_802 ();
 b15zdnd11an1n04x5 FILLER_284_834 ();
 b15zdnd00an1n01x5 FILLER_284_838 ();
 b15zdnd11an1n04x5 FILLER_284_870 ();
 b15zdnd11an1n16x5 FILLER_284_889 ();
 b15zdnd00an1n01x5 FILLER_284_905 ();
 b15zdnd11an1n04x5 FILLER_284_916 ();
 b15zdnd11an1n64x5 FILLER_284_929 ();
 b15zdnd11an1n08x5 FILLER_284_993 ();
 b15zdnd11an1n64x5 FILLER_284_1011 ();
 b15zdnd11an1n08x5 FILLER_284_1075 ();
 b15zdnd11an1n04x5 FILLER_284_1083 ();
 b15zdnd00an1n01x5 FILLER_284_1087 ();
 b15zdnd11an1n04x5 FILLER_284_1102 ();
 b15zdnd00an1n02x5 FILLER_284_1106 ();
 b15zdnd11an1n16x5 FILLER_284_1117 ();
 b15zdnd11an1n08x5 FILLER_284_1133 ();
 b15zdnd00an1n02x5 FILLER_284_1141 ();
 b15zdnd00an1n01x5 FILLER_284_1143 ();
 b15zdnd11an1n16x5 FILLER_284_1160 ();
 b15zdnd00an1n01x5 FILLER_284_1176 ();
 b15zdnd11an1n08x5 FILLER_284_1182 ();
 b15zdnd11an1n64x5 FILLER_284_1198 ();
 b15zdnd11an1n32x5 FILLER_284_1262 ();
 b15zdnd11an1n04x5 FILLER_284_1294 ();
 b15zdnd00an1n02x5 FILLER_284_1298 ();
 b15zdnd00an1n01x5 FILLER_284_1300 ();
 b15zdnd11an1n04x5 FILLER_284_1321 ();
 b15zdnd11an1n16x5 FILLER_284_1335 ();
 b15zdnd00an1n01x5 FILLER_284_1351 ();
 b15zdnd11an1n64x5 FILLER_284_1371 ();
 b15zdnd11an1n32x5 FILLER_284_1435 ();
 b15zdnd11an1n08x5 FILLER_284_1467 ();
 b15zdnd00an1n02x5 FILLER_284_1475 ();
 b15zdnd11an1n32x5 FILLER_284_1481 ();
 b15zdnd11an1n16x5 FILLER_284_1513 ();
 b15zdnd11an1n04x5 FILLER_284_1529 ();
 b15zdnd00an1n01x5 FILLER_284_1533 ();
 b15zdnd11an1n64x5 FILLER_284_1541 ();
 b15zdnd11an1n08x5 FILLER_284_1605 ();
 b15zdnd11an1n04x5 FILLER_284_1613 ();
 b15zdnd00an1n02x5 FILLER_284_1617 ();
 b15zdnd11an1n32x5 FILLER_284_1625 ();
 b15zdnd11an1n16x5 FILLER_284_1657 ();
 b15zdnd11an1n08x5 FILLER_284_1673 ();
 b15zdnd11an1n04x5 FILLER_284_1681 ();
 b15zdnd00an1n01x5 FILLER_284_1685 ();
 b15zdnd11an1n32x5 FILLER_284_1696 ();
 b15zdnd11an1n08x5 FILLER_284_1728 ();
 b15zdnd11an1n04x5 FILLER_284_1736 ();
 b15zdnd00an1n02x5 FILLER_284_1740 ();
 b15zdnd11an1n08x5 FILLER_284_1748 ();
 b15zdnd11an1n04x5 FILLER_284_1756 ();
 b15zdnd00an1n02x5 FILLER_284_1760 ();
 b15zdnd11an1n08x5 FILLER_284_1774 ();
 b15zdnd11an1n04x5 FILLER_284_1793 ();
 b15zdnd00an1n02x5 FILLER_284_1797 ();
 b15zdnd11an1n64x5 FILLER_284_1812 ();
 b15zdnd11an1n64x5 FILLER_284_1876 ();
 b15zdnd00an1n01x5 FILLER_284_1940 ();
 b15zdnd11an1n04x5 FILLER_284_1951 ();
 b15zdnd11an1n32x5 FILLER_284_1963 ();
 b15zdnd11an1n16x5 FILLER_284_1995 ();
 b15zdnd00an1n02x5 FILLER_284_2011 ();
 b15zdnd11an1n64x5 FILLER_284_2023 ();
 b15zdnd11an1n16x5 FILLER_284_2087 ();
 b15zdnd11an1n08x5 FILLER_284_2103 ();
 b15zdnd11an1n04x5 FILLER_284_2111 ();
 b15zdnd11an1n04x5 FILLER_284_2127 ();
 b15zdnd11an1n04x5 FILLER_284_2147 ();
 b15zdnd00an1n02x5 FILLER_284_2151 ();
 b15zdnd00an1n01x5 FILLER_284_2153 ();
 b15zdnd11an1n08x5 FILLER_284_2162 ();
 b15zdnd11an1n04x5 FILLER_284_2176 ();
 b15zdnd11an1n32x5 FILLER_284_2186 ();
 b15zdnd00an1n02x5 FILLER_284_2218 ();
 b15zdnd00an1n01x5 FILLER_284_2220 ();
 b15zdnd11an1n04x5 FILLER_284_2233 ();
 b15zdnd11an1n16x5 FILLER_284_2253 ();
 b15zdnd11an1n04x5 FILLER_284_2269 ();
 b15zdnd00an1n02x5 FILLER_284_2273 ();
 b15zdnd00an1n01x5 FILLER_284_2275 ();
 b15zdnd11an1n32x5 FILLER_285_0 ();
 b15zdnd11an1n04x5 FILLER_285_32 ();
 b15zdnd11an1n08x5 FILLER_285_56 ();
 b15zdnd11an1n08x5 FILLER_285_82 ();
 b15zdnd11an1n04x5 FILLER_285_90 ();
 b15zdnd00an1n01x5 FILLER_285_94 ();
 b15zdnd11an1n32x5 FILLER_285_111 ();
 b15zdnd11an1n16x5 FILLER_285_143 ();
 b15zdnd00an1n01x5 FILLER_285_159 ();
 b15zdnd11an1n04x5 FILLER_285_172 ();
 b15zdnd11an1n04x5 FILLER_285_180 ();
 b15zdnd00an1n02x5 FILLER_285_184 ();
 b15zdnd11an1n32x5 FILLER_285_192 ();
 b15zdnd11an1n16x5 FILLER_285_224 ();
 b15zdnd11an1n16x5 FILLER_285_245 ();
 b15zdnd11an1n04x5 FILLER_285_274 ();
 b15zdnd11an1n04x5 FILLER_285_282 ();
 b15zdnd00an1n01x5 FILLER_285_286 ();
 b15zdnd11an1n32x5 FILLER_285_296 ();
 b15zdnd11an1n16x5 FILLER_285_328 ();
 b15zdnd11an1n08x5 FILLER_285_344 ();
 b15zdnd11an1n04x5 FILLER_285_352 ();
 b15zdnd00an1n02x5 FILLER_285_356 ();
 b15zdnd11an1n64x5 FILLER_285_368 ();
 b15zdnd11an1n16x5 FILLER_285_432 ();
 b15zdnd00an1n01x5 FILLER_285_448 ();
 b15zdnd11an1n08x5 FILLER_285_460 ();
 b15zdnd11an1n04x5 FILLER_285_484 ();
 b15zdnd11an1n08x5 FILLER_285_494 ();
 b15zdnd00an1n02x5 FILLER_285_502 ();
 b15zdnd00an1n01x5 FILLER_285_504 ();
 b15zdnd11an1n04x5 FILLER_285_511 ();
 b15zdnd11an1n32x5 FILLER_285_527 ();
 b15zdnd11an1n08x5 FILLER_285_559 ();
 b15zdnd11an1n04x5 FILLER_285_567 ();
 b15zdnd00an1n02x5 FILLER_285_571 ();
 b15zdnd11an1n04x5 FILLER_285_580 ();
 b15zdnd11an1n04x5 FILLER_285_591 ();
 b15zdnd00an1n02x5 FILLER_285_595 ();
 b15zdnd00an1n01x5 FILLER_285_597 ();
 b15zdnd11an1n04x5 FILLER_285_610 ();
 b15zdnd11an1n08x5 FILLER_285_624 ();
 b15zdnd11an1n04x5 FILLER_285_632 ();
 b15zdnd11an1n32x5 FILLER_285_641 ();
 b15zdnd11an1n04x5 FILLER_285_673 ();
 b15zdnd00an1n02x5 FILLER_285_677 ();
 b15zdnd00an1n01x5 FILLER_285_679 ();
 b15zdnd11an1n16x5 FILLER_285_685 ();
 b15zdnd11an1n08x5 FILLER_285_701 ();
 b15zdnd00an1n02x5 FILLER_285_709 ();
 b15zdnd11an1n32x5 FILLER_285_716 ();
 b15zdnd11an1n16x5 FILLER_285_748 ();
 b15zdnd11an1n08x5 FILLER_285_764 ();
 b15zdnd11an1n04x5 FILLER_285_772 ();
 b15zdnd11an1n04x5 FILLER_285_781 ();
 b15zdnd11an1n04x5 FILLER_285_790 ();
 b15zdnd00an1n01x5 FILLER_285_794 ();
 b15zdnd11an1n32x5 FILLER_285_827 ();
 b15zdnd11an1n16x5 FILLER_285_859 ();
 b15zdnd11an1n04x5 FILLER_285_875 ();
 b15zdnd00an1n01x5 FILLER_285_879 ();
 b15zdnd11an1n04x5 FILLER_285_906 ();
 b15zdnd11an1n64x5 FILLER_285_920 ();
 b15zdnd11an1n16x5 FILLER_285_984 ();
 b15zdnd11an1n08x5 FILLER_285_1000 ();
 b15zdnd11an1n08x5 FILLER_285_1020 ();
 b15zdnd11an1n64x5 FILLER_285_1034 ();
 b15zdnd11an1n32x5 FILLER_285_1098 ();
 b15zdnd11an1n08x5 FILLER_285_1130 ();
 b15zdnd11an1n04x5 FILLER_285_1138 ();
 b15zdnd00an1n01x5 FILLER_285_1142 ();
 b15zdnd11an1n64x5 FILLER_285_1152 ();
 b15zdnd11an1n04x5 FILLER_285_1216 ();
 b15zdnd00an1n01x5 FILLER_285_1220 ();
 b15zdnd11an1n04x5 FILLER_285_1233 ();
 b15zdnd11an1n08x5 FILLER_285_1242 ();
 b15zdnd11an1n04x5 FILLER_285_1250 ();
 b15zdnd00an1n02x5 FILLER_285_1254 ();
 b15zdnd11an1n16x5 FILLER_285_1261 ();
 b15zdnd11an1n04x5 FILLER_285_1277 ();
 b15zdnd00an1n02x5 FILLER_285_1281 ();
 b15zdnd00an1n01x5 FILLER_285_1283 ();
 b15zdnd11an1n08x5 FILLER_285_1293 ();
 b15zdnd11an1n16x5 FILLER_285_1305 ();
 b15zdnd00an1n01x5 FILLER_285_1321 ();
 b15zdnd11an1n64x5 FILLER_285_1333 ();
 b15zdnd11an1n32x5 FILLER_285_1397 ();
 b15zdnd11an1n08x5 FILLER_285_1429 ();
 b15zdnd00an1n02x5 FILLER_285_1437 ();
 b15zdnd11an1n16x5 FILLER_285_1445 ();
 b15zdnd11an1n04x5 FILLER_285_1461 ();
 b15zdnd11an1n04x5 FILLER_285_1470 ();
 b15zdnd11an1n32x5 FILLER_285_1486 ();
 b15zdnd11an1n04x5 FILLER_285_1522 ();
 b15zdnd00an1n02x5 FILLER_285_1526 ();
 b15zdnd00an1n01x5 FILLER_285_1528 ();
 b15zdnd11an1n04x5 FILLER_285_1537 ();
 b15zdnd11an1n04x5 FILLER_285_1546 ();
 b15zdnd11an1n16x5 FILLER_285_1558 ();
 b15zdnd11an1n04x5 FILLER_285_1574 ();
 b15zdnd00an1n02x5 FILLER_285_1578 ();
 b15zdnd11an1n16x5 FILLER_285_1587 ();
 b15zdnd00an1n02x5 FILLER_285_1603 ();
 b15zdnd00an1n01x5 FILLER_285_1605 ();
 b15zdnd11an1n04x5 FILLER_285_1615 ();
 b15zdnd11an1n16x5 FILLER_285_1632 ();
 b15zdnd11an1n04x5 FILLER_285_1648 ();
 b15zdnd00an1n01x5 FILLER_285_1652 ();
 b15zdnd11an1n32x5 FILLER_285_1665 ();
 b15zdnd11an1n16x5 FILLER_285_1697 ();
 b15zdnd00an1n01x5 FILLER_285_1713 ();
 b15zdnd11an1n32x5 FILLER_285_1721 ();
 b15zdnd11an1n16x5 FILLER_285_1753 ();
 b15zdnd11an1n08x5 FILLER_285_1769 ();
 b15zdnd00an1n02x5 FILLER_285_1777 ();
 b15zdnd11an1n16x5 FILLER_285_1785 ();
 b15zdnd11an1n08x5 FILLER_285_1801 ();
 b15zdnd11an1n04x5 FILLER_285_1809 ();
 b15zdnd00an1n02x5 FILLER_285_1813 ();
 b15zdnd11an1n32x5 FILLER_285_1819 ();
 b15zdnd11an1n16x5 FILLER_285_1851 ();
 b15zdnd11an1n04x5 FILLER_285_1867 ();
 b15zdnd11an1n04x5 FILLER_285_1878 ();
 b15zdnd11an1n04x5 FILLER_285_1891 ();
 b15zdnd11an1n08x5 FILLER_285_1900 ();
 b15zdnd00an1n02x5 FILLER_285_1908 ();
 b15zdnd11an1n08x5 FILLER_285_1918 ();
 b15zdnd11an1n04x5 FILLER_285_1926 ();
 b15zdnd00an1n02x5 FILLER_285_1930 ();
 b15zdnd00an1n01x5 FILLER_285_1932 ();
 b15zdnd11an1n04x5 FILLER_285_1946 ();
 b15zdnd00an1n01x5 FILLER_285_1950 ();
 b15zdnd11an1n32x5 FILLER_285_1956 ();
 b15zdnd11an1n04x5 FILLER_285_1988 ();
 b15zdnd00an1n01x5 FILLER_285_1992 ();
 b15zdnd11an1n16x5 FILLER_285_1997 ();
 b15zdnd11an1n04x5 FILLER_285_2013 ();
 b15zdnd00an1n02x5 FILLER_285_2017 ();
 b15zdnd00an1n01x5 FILLER_285_2019 ();
 b15zdnd11an1n04x5 FILLER_285_2040 ();
 b15zdnd00an1n02x5 FILLER_285_2044 ();
 b15zdnd11an1n04x5 FILLER_285_2053 ();
 b15zdnd11an1n16x5 FILLER_285_2062 ();
 b15zdnd00an1n02x5 FILLER_285_2078 ();
 b15zdnd00an1n01x5 FILLER_285_2080 ();
 b15zdnd11an1n04x5 FILLER_285_2087 ();
 b15zdnd11an1n04x5 FILLER_285_2096 ();
 b15zdnd11an1n64x5 FILLER_285_2106 ();
 b15zdnd11an1n64x5 FILLER_285_2170 ();
 b15zdnd11an1n32x5 FILLER_285_2234 ();
 b15zdnd11an1n16x5 FILLER_285_2266 ();
 b15zdnd00an1n02x5 FILLER_285_2282 ();
 b15zdnd11an1n16x5 FILLER_286_8 ();
 b15zdnd11an1n08x5 FILLER_286_24 ();
 b15zdnd00an1n02x5 FILLER_286_32 ();
 b15zdnd00an1n01x5 FILLER_286_34 ();
 b15zdnd11an1n32x5 FILLER_286_58 ();
 b15zdnd11an1n08x5 FILLER_286_90 ();
 b15zdnd11an1n04x5 FILLER_286_98 ();
 b15zdnd00an1n02x5 FILLER_286_102 ();
 b15zdnd11an1n16x5 FILLER_286_110 ();
 b15zdnd00an1n02x5 FILLER_286_126 ();
 b15zdnd11an1n32x5 FILLER_286_149 ();
 b15zdnd11an1n04x5 FILLER_286_181 ();
 b15zdnd00an1n01x5 FILLER_286_185 ();
 b15zdnd11an1n16x5 FILLER_286_192 ();
 b15zdnd11an1n08x5 FILLER_286_208 ();
 b15zdnd11an1n16x5 FILLER_286_232 ();
 b15zdnd11an1n04x5 FILLER_286_248 ();
 b15zdnd00an1n01x5 FILLER_286_252 ();
 b15zdnd11an1n08x5 FILLER_286_260 ();
 b15zdnd11an1n04x5 FILLER_286_273 ();
 b15zdnd00an1n02x5 FILLER_286_277 ();
 b15zdnd00an1n01x5 FILLER_286_279 ();
 b15zdnd11an1n04x5 FILLER_286_286 ();
 b15zdnd11an1n32x5 FILLER_286_303 ();
 b15zdnd11an1n04x5 FILLER_286_335 ();
 b15zdnd11an1n04x5 FILLER_286_351 ();
 b15zdnd11an1n64x5 FILLER_286_364 ();
 b15zdnd11an1n64x5 FILLER_286_428 ();
 b15zdnd11an1n08x5 FILLER_286_492 ();
 b15zdnd00an1n02x5 FILLER_286_500 ();
 b15zdnd11an1n32x5 FILLER_286_508 ();
 b15zdnd11an1n16x5 FILLER_286_540 ();
 b15zdnd11an1n64x5 FILLER_286_566 ();
 b15zdnd11an1n08x5 FILLER_286_630 ();
 b15zdnd00an1n01x5 FILLER_286_638 ();
 b15zdnd11an1n16x5 FILLER_286_646 ();
 b15zdnd11an1n08x5 FILLER_286_662 ();
 b15zdnd11an1n04x5 FILLER_286_670 ();
 b15zdnd00an1n01x5 FILLER_286_674 ();
 b15zdnd11an1n32x5 FILLER_286_684 ();
 b15zdnd00an1n02x5 FILLER_286_716 ();
 b15zdnd11an1n04x5 FILLER_286_726 ();
 b15zdnd00an1n01x5 FILLER_286_730 ();
 b15zdnd11an1n64x5 FILLER_286_735 ();
 b15zdnd11an1n16x5 FILLER_286_799 ();
 b15zdnd00an1n02x5 FILLER_286_815 ();
 b15zdnd11an1n64x5 FILLER_286_842 ();
 b15zdnd11an1n32x5 FILLER_286_906 ();
 b15zdnd11an1n16x5 FILLER_286_938 ();
 b15zdnd00an1n02x5 FILLER_286_954 ();
 b15zdnd11an1n04x5 FILLER_286_962 ();
 b15zdnd11an1n16x5 FILLER_286_978 ();
 b15zdnd00an1n01x5 FILLER_286_994 ();
 b15zdnd11an1n08x5 FILLER_286_1021 ();
 b15zdnd00an1n02x5 FILLER_286_1029 ();
 b15zdnd00an1n01x5 FILLER_286_1031 ();
 b15zdnd11an1n08x5 FILLER_286_1038 ();
 b15zdnd11an1n04x5 FILLER_286_1046 ();
 b15zdnd00an1n01x5 FILLER_286_1050 ();
 b15zdnd11an1n32x5 FILLER_286_1055 ();
 b15zdnd11an1n16x5 FILLER_286_1087 ();
 b15zdnd11an1n04x5 FILLER_286_1103 ();
 b15zdnd00an1n02x5 FILLER_286_1107 ();
 b15zdnd11an1n64x5 FILLER_286_1116 ();
 b15zdnd11an1n64x5 FILLER_286_1180 ();
 b15zdnd11an1n08x5 FILLER_286_1244 ();
 b15zdnd00an1n02x5 FILLER_286_1252 ();
 b15zdnd11an1n08x5 FILLER_286_1270 ();
 b15zdnd11an1n04x5 FILLER_286_1278 ();
 b15zdnd00an1n01x5 FILLER_286_1282 ();
 b15zdnd11an1n08x5 FILLER_286_1288 ();
 b15zdnd11an1n04x5 FILLER_286_1310 ();
 b15zdnd11an1n04x5 FILLER_286_1340 ();
 b15zdnd11an1n08x5 FILLER_286_1360 ();
 b15zdnd00an1n01x5 FILLER_286_1368 ();
 b15zdnd11an1n32x5 FILLER_286_1382 ();
 b15zdnd11an1n16x5 FILLER_286_1414 ();
 b15zdnd11an1n08x5 FILLER_286_1430 ();
 b15zdnd00an1n02x5 FILLER_286_1438 ();
 b15zdnd11an1n08x5 FILLER_286_1448 ();
 b15zdnd00an1n02x5 FILLER_286_1456 ();
 b15zdnd11an1n64x5 FILLER_286_1471 ();
 b15zdnd11an1n08x5 FILLER_286_1535 ();
 b15zdnd11an1n16x5 FILLER_286_1548 ();
 b15zdnd11an1n04x5 FILLER_286_1564 ();
 b15zdnd00an1n02x5 FILLER_286_1568 ();
 b15zdnd00an1n01x5 FILLER_286_1570 ();
 b15zdnd11an1n32x5 FILLER_286_1578 ();
 b15zdnd11an1n08x5 FILLER_286_1610 ();
 b15zdnd00an1n01x5 FILLER_286_1618 ();
 b15zdnd11an1n08x5 FILLER_286_1630 ();
 b15zdnd00an1n02x5 FILLER_286_1638 ();
 b15zdnd11an1n04x5 FILLER_286_1645 ();
 b15zdnd11an1n32x5 FILLER_286_1655 ();
 b15zdnd11an1n16x5 FILLER_286_1687 ();
 b15zdnd11an1n08x5 FILLER_286_1703 ();
 b15zdnd11an1n04x5 FILLER_286_1711 ();
 b15zdnd11an1n08x5 FILLER_286_1730 ();
 b15zdnd11an1n04x5 FILLER_286_1744 ();
 b15zdnd00an1n02x5 FILLER_286_1748 ();
 b15zdnd00an1n01x5 FILLER_286_1750 ();
 b15zdnd11an1n08x5 FILLER_286_1762 ();
 b15zdnd00an1n02x5 FILLER_286_1770 ();
 b15zdnd00an1n01x5 FILLER_286_1772 ();
 b15zdnd11an1n32x5 FILLER_286_1780 ();
 b15zdnd00an1n01x5 FILLER_286_1812 ();
 b15zdnd11an1n32x5 FILLER_286_1835 ();
 b15zdnd11an1n32x5 FILLER_286_1887 ();
 b15zdnd11an1n16x5 FILLER_286_1919 ();
 b15zdnd00an1n02x5 FILLER_286_1935 ();
 b15zdnd11an1n04x5 FILLER_286_1957 ();
 b15zdnd00an1n02x5 FILLER_286_1961 ();
 b15zdnd11an1n08x5 FILLER_286_1973 ();
 b15zdnd11an1n04x5 FILLER_286_1981 ();
 b15zdnd00an1n01x5 FILLER_286_1985 ();
 b15zdnd11an1n08x5 FILLER_286_1995 ();
 b15zdnd11an1n04x5 FILLER_286_2003 ();
 b15zdnd00an1n02x5 FILLER_286_2007 ();
 b15zdnd11an1n04x5 FILLER_286_2013 ();
 b15zdnd11an1n16x5 FILLER_286_2024 ();
 b15zdnd11an1n04x5 FILLER_286_2040 ();
 b15zdnd00an1n01x5 FILLER_286_2044 ();
 b15zdnd11an1n16x5 FILLER_286_2051 ();
 b15zdnd11an1n08x5 FILLER_286_2067 ();
 b15zdnd11an1n04x5 FILLER_286_2075 ();
 b15zdnd00an1n02x5 FILLER_286_2079 ();
 b15zdnd11an1n08x5 FILLER_286_2087 ();
 b15zdnd11an1n16x5 FILLER_286_2107 ();
 b15zdnd00an1n02x5 FILLER_286_2123 ();
 b15zdnd00an1n01x5 FILLER_286_2125 ();
 b15zdnd00an1n02x5 FILLER_286_2152 ();
 b15zdnd00an1n02x5 FILLER_286_2162 ();
 b15zdnd00an1n01x5 FILLER_286_2164 ();
 b15zdnd11an1n32x5 FILLER_286_2177 ();
 b15zdnd11an1n16x5 FILLER_286_2209 ();
 b15zdnd00an1n01x5 FILLER_286_2225 ();
 b15zdnd11an1n32x5 FILLER_286_2240 ();
 b15zdnd11an1n04x5 FILLER_286_2272 ();
 b15zdnd11an1n32x5 FILLER_287_0 ();
 b15zdnd11an1n16x5 FILLER_287_32 ();
 b15zdnd11an1n04x5 FILLER_287_48 ();
 b15zdnd00an1n02x5 FILLER_287_52 ();
 b15zdnd11an1n04x5 FILLER_287_63 ();
 b15zdnd00an1n02x5 FILLER_287_67 ();
 b15zdnd11an1n64x5 FILLER_287_74 ();
 b15zdnd11an1n64x5 FILLER_287_138 ();
 b15zdnd11an1n64x5 FILLER_287_202 ();
 b15zdnd11an1n04x5 FILLER_287_266 ();
 b15zdnd00an1n02x5 FILLER_287_270 ();
 b15zdnd00an1n01x5 FILLER_287_272 ();
 b15zdnd11an1n32x5 FILLER_287_282 ();
 b15zdnd11an1n08x5 FILLER_287_314 ();
 b15zdnd00an1n02x5 FILLER_287_322 ();
 b15zdnd00an1n01x5 FILLER_287_324 ();
 b15zdnd11an1n04x5 FILLER_287_330 ();
 b15zdnd11an1n08x5 FILLER_287_349 ();
 b15zdnd11an1n04x5 FILLER_287_357 ();
 b15zdnd00an1n02x5 FILLER_287_361 ();
 b15zdnd11an1n32x5 FILLER_287_371 ();
 b15zdnd11an1n16x5 FILLER_287_403 ();
 b15zdnd00an1n02x5 FILLER_287_419 ();
 b15zdnd11an1n16x5 FILLER_287_437 ();
 b15zdnd11an1n32x5 FILLER_287_463 ();
 b15zdnd11an1n16x5 FILLER_287_495 ();
 b15zdnd11an1n04x5 FILLER_287_511 ();
 b15zdnd00an1n01x5 FILLER_287_515 ();
 b15zdnd11an1n32x5 FILLER_287_526 ();
 b15zdnd11an1n16x5 FILLER_287_558 ();
 b15zdnd11an1n04x5 FILLER_287_574 ();
 b15zdnd00an1n02x5 FILLER_287_578 ();
 b15zdnd11an1n32x5 FILLER_287_592 ();
 b15zdnd11an1n08x5 FILLER_287_624 ();
 b15zdnd11an1n04x5 FILLER_287_632 ();
 b15zdnd00an1n02x5 FILLER_287_636 ();
 b15zdnd11an1n64x5 FILLER_287_652 ();
 b15zdnd11an1n08x5 FILLER_287_716 ();
 b15zdnd00an1n02x5 FILLER_287_724 ();
 b15zdnd00an1n01x5 FILLER_287_726 ();
 b15zdnd11an1n32x5 FILLER_287_739 ();
 b15zdnd11an1n16x5 FILLER_287_771 ();
 b15zdnd11an1n04x5 FILLER_287_787 ();
 b15zdnd00an1n01x5 FILLER_287_791 ();
 b15zdnd11an1n16x5 FILLER_287_812 ();
 b15zdnd00an1n02x5 FILLER_287_828 ();
 b15zdnd11an1n16x5 FILLER_287_855 ();
 b15zdnd11an1n08x5 FILLER_287_871 ();
 b15zdnd00an1n02x5 FILLER_287_879 ();
 b15zdnd11an1n32x5 FILLER_287_906 ();
 b15zdnd11an1n16x5 FILLER_287_938 ();
 b15zdnd11an1n08x5 FILLER_287_954 ();
 b15zdnd00an1n02x5 FILLER_287_962 ();
 b15zdnd00an1n01x5 FILLER_287_964 ();
 b15zdnd11an1n16x5 FILLER_287_971 ();
 b15zdnd11an1n08x5 FILLER_287_987 ();
 b15zdnd11an1n04x5 FILLER_287_995 ();
 b15zdnd00an1n02x5 FILLER_287_999 ();
 b15zdnd00an1n01x5 FILLER_287_1001 ();
 b15zdnd11an1n32x5 FILLER_287_1012 ();
 b15zdnd11an1n16x5 FILLER_287_1044 ();
 b15zdnd11an1n04x5 FILLER_287_1060 ();
 b15zdnd00an1n01x5 FILLER_287_1064 ();
 b15zdnd11an1n04x5 FILLER_287_1079 ();
 b15zdnd11an1n64x5 FILLER_287_1092 ();
 b15zdnd11an1n16x5 FILLER_287_1156 ();
 b15zdnd11an1n08x5 FILLER_287_1172 ();
 b15zdnd00an1n02x5 FILLER_287_1180 ();
 b15zdnd11an1n04x5 FILLER_287_1188 ();
 b15zdnd11an1n08x5 FILLER_287_1198 ();
 b15zdnd11an1n04x5 FILLER_287_1206 ();
 b15zdnd00an1n02x5 FILLER_287_1210 ();
 b15zdnd00an1n01x5 FILLER_287_1212 ();
 b15zdnd11an1n04x5 FILLER_287_1229 ();
 b15zdnd11an1n64x5 FILLER_287_1238 ();
 b15zdnd11an1n64x5 FILLER_287_1302 ();
 b15zdnd11an1n32x5 FILLER_287_1366 ();
 b15zdnd11an1n16x5 FILLER_287_1398 ();
 b15zdnd11an1n08x5 FILLER_287_1414 ();
 b15zdnd11an1n04x5 FILLER_287_1422 ();
 b15zdnd00an1n02x5 FILLER_287_1426 ();
 b15zdnd00an1n01x5 FILLER_287_1428 ();
 b15zdnd11an1n16x5 FILLER_287_1436 ();
 b15zdnd11an1n08x5 FILLER_287_1452 ();
 b15zdnd00an1n02x5 FILLER_287_1460 ();
 b15zdnd11an1n64x5 FILLER_287_1476 ();
 b15zdnd11an1n16x5 FILLER_287_1540 ();
 b15zdnd11an1n08x5 FILLER_287_1556 ();
 b15zdnd00an1n01x5 FILLER_287_1564 ();
 b15zdnd11an1n04x5 FILLER_287_1570 ();
 b15zdnd11an1n08x5 FILLER_287_1605 ();
 b15zdnd11an1n04x5 FILLER_287_1629 ();
 b15zdnd00an1n02x5 FILLER_287_1633 ();
 b15zdnd00an1n01x5 FILLER_287_1635 ();
 b15zdnd11an1n08x5 FILLER_287_1641 ();
 b15zdnd00an1n01x5 FILLER_287_1649 ();
 b15zdnd11an1n08x5 FILLER_287_1656 ();
 b15zdnd00an1n01x5 FILLER_287_1664 ();
 b15zdnd11an1n04x5 FILLER_287_1670 ();
 b15zdnd00an1n02x5 FILLER_287_1674 ();
 b15zdnd11an1n04x5 FILLER_287_1687 ();
 b15zdnd11an1n16x5 FILLER_287_1703 ();
 b15zdnd11an1n08x5 FILLER_287_1725 ();
 b15zdnd11an1n64x5 FILLER_287_1744 ();
 b15zdnd11an1n08x5 FILLER_287_1808 ();
 b15zdnd00an1n02x5 FILLER_287_1816 ();
 b15zdnd11an1n64x5 FILLER_287_1830 ();
 b15zdnd11an1n32x5 FILLER_287_1894 ();
 b15zdnd11an1n04x5 FILLER_287_1926 ();
 b15zdnd00an1n02x5 FILLER_287_1930 ();
 b15zdnd00an1n01x5 FILLER_287_1932 ();
 b15zdnd11an1n16x5 FILLER_287_1949 ();
 b15zdnd11an1n08x5 FILLER_287_1965 ();
 b15zdnd11an1n04x5 FILLER_287_1973 ();
 b15zdnd11an1n04x5 FILLER_287_1986 ();
 b15zdnd11an1n08x5 FILLER_287_2004 ();
 b15zdnd11an1n04x5 FILLER_287_2012 ();
 b15zdnd00an1n01x5 FILLER_287_2016 ();
 b15zdnd11an1n16x5 FILLER_287_2023 ();
 b15zdnd11an1n08x5 FILLER_287_2039 ();
 b15zdnd11an1n04x5 FILLER_287_2067 ();
 b15zdnd00an1n02x5 FILLER_287_2071 ();
 b15zdnd11an1n04x5 FILLER_287_2093 ();
 b15zdnd11an1n04x5 FILLER_287_2105 ();
 b15zdnd11an1n08x5 FILLER_287_2121 ();
 b15zdnd11an1n04x5 FILLER_287_2129 ();
 b15zdnd00an1n02x5 FILLER_287_2133 ();
 b15zdnd00an1n01x5 FILLER_287_2135 ();
 b15zdnd11an1n08x5 FILLER_287_2140 ();
 b15zdnd00an1n02x5 FILLER_287_2148 ();
 b15zdnd11an1n16x5 FILLER_287_2164 ();
 b15zdnd11an1n04x5 FILLER_287_2180 ();
 b15zdnd00an1n02x5 FILLER_287_2184 ();
 b15zdnd11an1n04x5 FILLER_287_2197 ();
 b15zdnd11an1n64x5 FILLER_287_2205 ();
 b15zdnd11an1n08x5 FILLER_287_2269 ();
 b15zdnd11an1n04x5 FILLER_287_2277 ();
 b15zdnd00an1n02x5 FILLER_287_2281 ();
 b15zdnd00an1n01x5 FILLER_287_2283 ();
 b15zdnd11an1n32x5 FILLER_288_8 ();
 b15zdnd11an1n16x5 FILLER_288_40 ();
 b15zdnd11an1n08x5 FILLER_288_56 ();
 b15zdnd11an1n04x5 FILLER_288_64 ();
 b15zdnd00an1n02x5 FILLER_288_68 ();
 b15zdnd11an1n64x5 FILLER_288_83 ();
 b15zdnd11an1n04x5 FILLER_288_147 ();
 b15zdnd00an1n02x5 FILLER_288_151 ();
 b15zdnd11an1n64x5 FILLER_288_158 ();
 b15zdnd11an1n64x5 FILLER_288_222 ();
 b15zdnd11an1n32x5 FILLER_288_286 ();
 b15zdnd11an1n16x5 FILLER_288_318 ();
 b15zdnd11an1n04x5 FILLER_288_334 ();
 b15zdnd00an1n01x5 FILLER_288_338 ();
 b15zdnd11an1n08x5 FILLER_288_343 ();
 b15zdnd11an1n04x5 FILLER_288_351 ();
 b15zdnd11an1n32x5 FILLER_288_371 ();
 b15zdnd11an1n16x5 FILLER_288_403 ();
 b15zdnd00an1n02x5 FILLER_288_419 ();
 b15zdnd11an1n16x5 FILLER_288_437 ();
 b15zdnd00an1n02x5 FILLER_288_453 ();
 b15zdnd11an1n32x5 FILLER_288_473 ();
 b15zdnd11an1n08x5 FILLER_288_505 ();
 b15zdnd11an1n04x5 FILLER_288_513 ();
 b15zdnd11an1n04x5 FILLER_288_525 ();
 b15zdnd11an1n08x5 FILLER_288_534 ();
 b15zdnd11an1n04x5 FILLER_288_542 ();
 b15zdnd00an1n02x5 FILLER_288_546 ();
 b15zdnd11an1n04x5 FILLER_288_554 ();
 b15zdnd11an1n32x5 FILLER_288_564 ();
 b15zdnd11an1n16x5 FILLER_288_596 ();
 b15zdnd11an1n04x5 FILLER_288_612 ();
 b15zdnd00an1n01x5 FILLER_288_616 ();
 b15zdnd11an1n32x5 FILLER_288_627 ();
 b15zdnd11an1n16x5 FILLER_288_659 ();
 b15zdnd11an1n04x5 FILLER_288_675 ();
 b15zdnd11an1n08x5 FILLER_288_691 ();
 b15zdnd11an1n04x5 FILLER_288_699 ();
 b15zdnd00an1n02x5 FILLER_288_703 ();
 b15zdnd00an1n01x5 FILLER_288_705 ();
 b15zdnd00an1n02x5 FILLER_288_716 ();
 b15zdnd00an1n02x5 FILLER_288_726 ();
 b15zdnd11an1n16x5 FILLER_288_744 ();
 b15zdnd11an1n08x5 FILLER_288_760 ();
 b15zdnd11an1n04x5 FILLER_288_768 ();
 b15zdnd00an1n02x5 FILLER_288_772 ();
 b15zdnd00an1n01x5 FILLER_288_774 ();
 b15zdnd11an1n04x5 FILLER_288_781 ();
 b15zdnd00an1n01x5 FILLER_288_785 ();
 b15zdnd11an1n64x5 FILLER_288_792 ();
 b15zdnd11an1n64x5 FILLER_288_856 ();
 b15zdnd11an1n64x5 FILLER_288_920 ();
 b15zdnd11an1n32x5 FILLER_288_984 ();
 b15zdnd11an1n04x5 FILLER_288_1016 ();
 b15zdnd11an1n04x5 FILLER_288_1024 ();
 b15zdnd11an1n32x5 FILLER_288_1034 ();
 b15zdnd11an1n08x5 FILLER_288_1066 ();
 b15zdnd00an1n01x5 FILLER_288_1074 ();
 b15zdnd11an1n16x5 FILLER_288_1085 ();
 b15zdnd11an1n04x5 FILLER_288_1101 ();
 b15zdnd00an1n01x5 FILLER_288_1105 ();
 b15zdnd11an1n04x5 FILLER_288_1111 ();
 b15zdnd00an1n02x5 FILLER_288_1115 ();
 b15zdnd00an1n01x5 FILLER_288_1117 ();
 b15zdnd11an1n04x5 FILLER_288_1127 ();
 b15zdnd11an1n04x5 FILLER_288_1151 ();
 b15zdnd00an1n02x5 FILLER_288_1155 ();
 b15zdnd11an1n64x5 FILLER_288_1163 ();
 b15zdnd11an1n64x5 FILLER_288_1227 ();
 b15zdnd11an1n04x5 FILLER_288_1291 ();
 b15zdnd11an1n16x5 FILLER_288_1313 ();
 b15zdnd00an1n02x5 FILLER_288_1329 ();
 b15zdnd00an1n01x5 FILLER_288_1331 ();
 b15zdnd11an1n64x5 FILLER_288_1344 ();
 b15zdnd11an1n16x5 FILLER_288_1408 ();
 b15zdnd00an1n02x5 FILLER_288_1424 ();
 b15zdnd11an1n04x5 FILLER_288_1430 ();
 b15zdnd11an1n16x5 FILLER_288_1442 ();
 b15zdnd11an1n08x5 FILLER_288_1458 ();
 b15zdnd11an1n04x5 FILLER_288_1466 ();
 b15zdnd00an1n02x5 FILLER_288_1470 ();
 b15zdnd00an1n01x5 FILLER_288_1472 ();
 b15zdnd11an1n64x5 FILLER_288_1482 ();
 b15zdnd11an1n16x5 FILLER_288_1546 ();
 b15zdnd11an1n08x5 FILLER_288_1562 ();
 b15zdnd11an1n04x5 FILLER_288_1570 ();
 b15zdnd00an1n02x5 FILLER_288_1574 ();
 b15zdnd00an1n01x5 FILLER_288_1576 ();
 b15zdnd11an1n64x5 FILLER_288_1594 ();
 b15zdnd11an1n16x5 FILLER_288_1658 ();
 b15zdnd11an1n04x5 FILLER_288_1674 ();
 b15zdnd00an1n02x5 FILLER_288_1678 ();
 b15zdnd11an1n32x5 FILLER_288_1686 ();
 b15zdnd11an1n16x5 FILLER_288_1718 ();
 b15zdnd00an1n02x5 FILLER_288_1734 ();
 b15zdnd00an1n01x5 FILLER_288_1736 ();
 b15zdnd11an1n32x5 FILLER_288_1749 ();
 b15zdnd11an1n04x5 FILLER_288_1781 ();
 b15zdnd00an1n01x5 FILLER_288_1785 ();
 b15zdnd11an1n08x5 FILLER_288_1802 ();
 b15zdnd00an1n02x5 FILLER_288_1810 ();
 b15zdnd11an1n64x5 FILLER_288_1819 ();
 b15zdnd11an1n64x5 FILLER_288_1883 ();
 b15zdnd11an1n32x5 FILLER_288_1947 ();
 b15zdnd11an1n08x5 FILLER_288_1979 ();
 b15zdnd11an1n64x5 FILLER_288_1992 ();
 b15zdnd11an1n64x5 FILLER_288_2056 ();
 b15zdnd11an1n32x5 FILLER_288_2120 ();
 b15zdnd00an1n02x5 FILLER_288_2152 ();
 b15zdnd11an1n32x5 FILLER_288_2162 ();
 b15zdnd00an1n01x5 FILLER_288_2194 ();
 b15zdnd11an1n64x5 FILLER_288_2202 ();
 b15zdnd11an1n08x5 FILLER_288_2266 ();
 b15zdnd00an1n02x5 FILLER_288_2274 ();
 b15zdnd11an1n32x5 FILLER_289_0 ();
 b15zdnd11an1n08x5 FILLER_289_32 ();
 b15zdnd11an1n04x5 FILLER_289_40 ();
 b15zdnd00an1n02x5 FILLER_289_44 ();
 b15zdnd00an1n01x5 FILLER_289_46 ();
 b15zdnd11an1n08x5 FILLER_289_63 ();
 b15zdnd00an1n02x5 FILLER_289_71 ();
 b15zdnd11an1n08x5 FILLER_289_80 ();
 b15zdnd11an1n04x5 FILLER_289_88 ();
 b15zdnd00an1n02x5 FILLER_289_92 ();
 b15zdnd11an1n04x5 FILLER_289_100 ();
 b15zdnd11an1n04x5 FILLER_289_110 ();
 b15zdnd11an1n08x5 FILLER_289_138 ();
 b15zdnd11an1n04x5 FILLER_289_146 ();
 b15zdnd11an1n08x5 FILLER_289_159 ();
 b15zdnd11an1n04x5 FILLER_289_167 ();
 b15zdnd11an1n32x5 FILLER_289_178 ();
 b15zdnd11an1n08x5 FILLER_289_210 ();
 b15zdnd11an1n04x5 FILLER_289_218 ();
 b15zdnd00an1n02x5 FILLER_289_222 ();
 b15zdnd11an1n04x5 FILLER_289_236 ();
 b15zdnd11an1n64x5 FILLER_289_245 ();
 b15zdnd11an1n64x5 FILLER_289_309 ();
 b15zdnd11an1n32x5 FILLER_289_373 ();
 b15zdnd11an1n16x5 FILLER_289_405 ();
 b15zdnd11an1n04x5 FILLER_289_421 ();
 b15zdnd00an1n02x5 FILLER_289_425 ();
 b15zdnd00an1n01x5 FILLER_289_427 ();
 b15zdnd11an1n04x5 FILLER_289_435 ();
 b15zdnd11an1n64x5 FILLER_289_449 ();
 b15zdnd11an1n64x5 FILLER_289_513 ();
 b15zdnd11an1n04x5 FILLER_289_577 ();
 b15zdnd00an1n02x5 FILLER_289_581 ();
 b15zdnd11an1n08x5 FILLER_289_592 ();
 b15zdnd00an1n02x5 FILLER_289_600 ();
 b15zdnd00an1n01x5 FILLER_289_602 ();
 b15zdnd11an1n16x5 FILLER_289_611 ();
 b15zdnd00an1n01x5 FILLER_289_627 ();
 b15zdnd11an1n08x5 FILLER_289_638 ();
 b15zdnd00an1n01x5 FILLER_289_646 ();
 b15zdnd11an1n08x5 FILLER_289_667 ();
 b15zdnd00an1n01x5 FILLER_289_675 ();
 b15zdnd11an1n32x5 FILLER_289_688 ();
 b15zdnd11an1n16x5 FILLER_289_720 ();
 b15zdnd11an1n04x5 FILLER_289_736 ();
 b15zdnd00an1n02x5 FILLER_289_740 ();
 b15zdnd11an1n04x5 FILLER_289_746 ();
 b15zdnd11an1n04x5 FILLER_289_773 ();
 b15zdnd00an1n01x5 FILLER_289_777 ();
 b15zdnd11an1n04x5 FILLER_289_785 ();
 b15zdnd00an1n01x5 FILLER_289_789 ();
 b15zdnd11an1n64x5 FILLER_289_797 ();
 b15zdnd11an1n64x5 FILLER_289_861 ();
 b15zdnd11an1n32x5 FILLER_289_925 ();
 b15zdnd11an1n16x5 FILLER_289_957 ();
 b15zdnd11an1n08x5 FILLER_289_973 ();
 b15zdnd11an1n04x5 FILLER_289_981 ();
 b15zdnd00an1n02x5 FILLER_289_985 ();
 b15zdnd11an1n04x5 FILLER_289_995 ();
 b15zdnd11an1n16x5 FILLER_289_1009 ();
 b15zdnd11an1n32x5 FILLER_289_1035 ();
 b15zdnd00an1n01x5 FILLER_289_1067 ();
 b15zdnd11an1n08x5 FILLER_289_1082 ();
 b15zdnd00an1n01x5 FILLER_289_1090 ();
 b15zdnd11an1n08x5 FILLER_289_1101 ();
 b15zdnd00an1n01x5 FILLER_289_1109 ();
 b15zdnd11an1n08x5 FILLER_289_1116 ();
 b15zdnd11an1n16x5 FILLER_289_1129 ();
 b15zdnd11an1n08x5 FILLER_289_1145 ();
 b15zdnd00an1n02x5 FILLER_289_1153 ();
 b15zdnd11an1n64x5 FILLER_289_1160 ();
 b15zdnd11an1n64x5 FILLER_289_1224 ();
 b15zdnd11an1n16x5 FILLER_289_1288 ();
 b15zdnd11an1n08x5 FILLER_289_1304 ();
 b15zdnd00an1n01x5 FILLER_289_1312 ();
 b15zdnd11an1n08x5 FILLER_289_1322 ();
 b15zdnd00an1n01x5 FILLER_289_1330 ();
 b15zdnd11an1n04x5 FILLER_289_1335 ();
 b15zdnd00an1n02x5 FILLER_289_1339 ();
 b15zdnd00an1n01x5 FILLER_289_1341 ();
 b15zdnd11an1n64x5 FILLER_289_1366 ();
 b15zdnd11an1n32x5 FILLER_289_1430 ();
 b15zdnd11an1n08x5 FILLER_289_1462 ();
 b15zdnd00an1n02x5 FILLER_289_1470 ();
 b15zdnd11an1n32x5 FILLER_289_1486 ();
 b15zdnd00an1n02x5 FILLER_289_1518 ();
 b15zdnd00an1n01x5 FILLER_289_1520 ();
 b15zdnd11an1n16x5 FILLER_289_1533 ();
 b15zdnd11an1n08x5 FILLER_289_1549 ();
 b15zdnd00an1n02x5 FILLER_289_1557 ();
 b15zdnd00an1n01x5 FILLER_289_1559 ();
 b15zdnd11an1n08x5 FILLER_289_1566 ();
 b15zdnd11an1n04x5 FILLER_289_1574 ();
 b15zdnd00an1n02x5 FILLER_289_1578 ();
 b15zdnd11an1n64x5 FILLER_289_1592 ();
 b15zdnd11an1n64x5 FILLER_289_1656 ();
 b15zdnd11an1n32x5 FILLER_289_1720 ();
 b15zdnd11an1n16x5 FILLER_289_1752 ();
 b15zdnd11an1n08x5 FILLER_289_1768 ();
 b15zdnd11an1n04x5 FILLER_289_1776 ();
 b15zdnd11an1n64x5 FILLER_289_1790 ();
 b15zdnd11an1n32x5 FILLER_289_1854 ();
 b15zdnd00an1n02x5 FILLER_289_1886 ();
 b15zdnd00an1n01x5 FILLER_289_1888 ();
 b15zdnd11an1n04x5 FILLER_289_1921 ();
 b15zdnd00an1n02x5 FILLER_289_1925 ();
 b15zdnd11an1n04x5 FILLER_289_1939 ();
 b15zdnd11an1n64x5 FILLER_289_1960 ();
 b15zdnd11an1n32x5 FILLER_289_2024 ();
 b15zdnd11an1n08x5 FILLER_289_2056 ();
 b15zdnd00an1n02x5 FILLER_289_2064 ();
 b15zdnd11an1n64x5 FILLER_289_2078 ();
 b15zdnd11an1n32x5 FILLER_289_2142 ();
 b15zdnd11an1n16x5 FILLER_289_2174 ();
 b15zdnd11an1n16x5 FILLER_289_2195 ();
 b15zdnd11an1n08x5 FILLER_289_2211 ();
 b15zdnd00an1n01x5 FILLER_289_2219 ();
 b15zdnd11an1n08x5 FILLER_289_2226 ();
 b15zdnd11an1n04x5 FILLER_289_2240 ();
 b15zdnd11an1n32x5 FILLER_289_2248 ();
 b15zdnd11an1n04x5 FILLER_289_2280 ();
 b15zdnd11an1n32x5 FILLER_290_8 ();
 b15zdnd11an1n16x5 FILLER_290_40 ();
 b15zdnd11an1n08x5 FILLER_290_56 ();
 b15zdnd00an1n02x5 FILLER_290_64 ();
 b15zdnd11an1n64x5 FILLER_290_75 ();
 b15zdnd11an1n04x5 FILLER_290_139 ();
 b15zdnd00an1n01x5 FILLER_290_143 ();
 b15zdnd11an1n08x5 FILLER_290_154 ();
 b15zdnd11an1n16x5 FILLER_290_181 ();
 b15zdnd11an1n04x5 FILLER_290_197 ();
 b15zdnd11an1n04x5 FILLER_290_213 ();
 b15zdnd11an1n08x5 FILLER_290_229 ();
 b15zdnd11an1n04x5 FILLER_290_237 ();
 b15zdnd00an1n02x5 FILLER_290_241 ();
 b15zdnd11an1n08x5 FILLER_290_250 ();
 b15zdnd00an1n02x5 FILLER_290_258 ();
 b15zdnd00an1n01x5 FILLER_290_260 ();
 b15zdnd11an1n04x5 FILLER_290_269 ();
 b15zdnd00an1n02x5 FILLER_290_273 ();
 b15zdnd00an1n01x5 FILLER_290_275 ();
 b15zdnd11an1n16x5 FILLER_290_281 ();
 b15zdnd00an1n02x5 FILLER_290_297 ();
 b15zdnd11an1n04x5 FILLER_290_305 ();
 b15zdnd00an1n02x5 FILLER_290_309 ();
 b15zdnd11an1n32x5 FILLER_290_322 ();
 b15zdnd11an1n04x5 FILLER_290_354 ();
 b15zdnd11an1n64x5 FILLER_290_377 ();
 b15zdnd11an1n16x5 FILLER_290_441 ();
 b15zdnd11an1n08x5 FILLER_290_457 ();
 b15zdnd11an1n16x5 FILLER_290_474 ();
 b15zdnd11an1n04x5 FILLER_290_490 ();
 b15zdnd00an1n02x5 FILLER_290_494 ();
 b15zdnd11an1n04x5 FILLER_290_506 ();
 b15zdnd11an1n32x5 FILLER_290_515 ();
 b15zdnd11an1n16x5 FILLER_290_547 ();
 b15zdnd00an1n01x5 FILLER_290_563 ();
 b15zdnd11an1n08x5 FILLER_290_570 ();
 b15zdnd11an1n16x5 FILLER_290_599 ();
 b15zdnd00an1n02x5 FILLER_290_615 ();
 b15zdnd00an1n01x5 FILLER_290_617 ();
 b15zdnd11an1n16x5 FILLER_290_632 ();
 b15zdnd11an1n08x5 FILLER_290_648 ();
 b15zdnd11an1n08x5 FILLER_290_664 ();
 b15zdnd11an1n04x5 FILLER_290_672 ();
 b15zdnd00an1n02x5 FILLER_290_676 ();
 b15zdnd11an1n08x5 FILLER_290_688 ();
 b15zdnd00an1n01x5 FILLER_290_696 ();
 b15zdnd00an1n02x5 FILLER_290_716 ();
 b15zdnd11an1n64x5 FILLER_290_726 ();
 b15zdnd11an1n64x5 FILLER_290_790 ();
 b15zdnd11an1n04x5 FILLER_290_854 ();
 b15zdnd11an1n04x5 FILLER_290_884 ();
 b15zdnd11an1n64x5 FILLER_290_945 ();
 b15zdnd11an1n64x5 FILLER_290_1009 ();
 b15zdnd11an1n32x5 FILLER_290_1073 ();
 b15zdnd11an1n16x5 FILLER_290_1105 ();
 b15zdnd11an1n04x5 FILLER_290_1128 ();
 b15zdnd00an1n01x5 FILLER_290_1132 ();
 b15zdnd11an1n04x5 FILLER_290_1137 ();
 b15zdnd00an1n01x5 FILLER_290_1141 ();
 b15zdnd11an1n08x5 FILLER_290_1168 ();
 b15zdnd11an1n04x5 FILLER_290_1183 ();
 b15zdnd00an1n02x5 FILLER_290_1187 ();
 b15zdnd11an1n16x5 FILLER_290_1201 ();
 b15zdnd11an1n04x5 FILLER_290_1217 ();
 b15zdnd00an1n01x5 FILLER_290_1221 ();
 b15zdnd11an1n04x5 FILLER_290_1229 ();
 b15zdnd11an1n04x5 FILLER_290_1237 ();
 b15zdnd11an1n04x5 FILLER_290_1256 ();
 b15zdnd00an1n01x5 FILLER_290_1260 ();
 b15zdnd11an1n64x5 FILLER_290_1272 ();
 b15zdnd11an1n16x5 FILLER_290_1336 ();
 b15zdnd11an1n08x5 FILLER_290_1352 ();
 b15zdnd00an1n02x5 FILLER_290_1360 ();
 b15zdnd11an1n08x5 FILLER_290_1366 ();
 b15zdnd11an1n04x5 FILLER_290_1374 ();
 b15zdnd11an1n32x5 FILLER_290_1393 ();
 b15zdnd11an1n08x5 FILLER_290_1425 ();
 b15zdnd11an1n04x5 FILLER_290_1433 ();
 b15zdnd00an1n02x5 FILLER_290_1437 ();
 b15zdnd00an1n01x5 FILLER_290_1439 ();
 b15zdnd11an1n16x5 FILLER_290_1449 ();
 b15zdnd11an1n08x5 FILLER_290_1485 ();
 b15zdnd11an1n16x5 FILLER_290_1499 ();
 b15zdnd11an1n04x5 FILLER_290_1515 ();
 b15zdnd11an1n04x5 FILLER_290_1524 ();
 b15zdnd00an1n02x5 FILLER_290_1528 ();
 b15zdnd11an1n08x5 FILLER_290_1546 ();
 b15zdnd11an1n64x5 FILLER_290_1567 ();
 b15zdnd11an1n32x5 FILLER_290_1631 ();
 b15zdnd11an1n16x5 FILLER_290_1663 ();
 b15zdnd11an1n04x5 FILLER_290_1679 ();
 b15zdnd00an1n01x5 FILLER_290_1683 ();
 b15zdnd11an1n04x5 FILLER_290_1696 ();
 b15zdnd11an1n32x5 FILLER_290_1706 ();
 b15zdnd11an1n16x5 FILLER_290_1738 ();
 b15zdnd11an1n08x5 FILLER_290_1754 ();
 b15zdnd00an1n01x5 FILLER_290_1762 ();
 b15zdnd11an1n04x5 FILLER_290_1768 ();
 b15zdnd11an1n32x5 FILLER_290_1776 ();
 b15zdnd11an1n04x5 FILLER_290_1808 ();
 b15zdnd11an1n64x5 FILLER_290_1817 ();
 b15zdnd11an1n32x5 FILLER_290_1881 ();
 b15zdnd00an1n02x5 FILLER_290_1913 ();
 b15zdnd11an1n08x5 FILLER_290_1933 ();
 b15zdnd11an1n04x5 FILLER_290_1941 ();
 b15zdnd00an1n01x5 FILLER_290_1945 ();
 b15zdnd11an1n08x5 FILLER_290_1950 ();
 b15zdnd11an1n04x5 FILLER_290_1958 ();
 b15zdnd00an1n01x5 FILLER_290_1962 ();
 b15zdnd11an1n08x5 FILLER_290_1969 ();
 b15zdnd11an1n04x5 FILLER_290_1977 ();
 b15zdnd00an1n01x5 FILLER_290_1981 ();
 b15zdnd11an1n64x5 FILLER_290_1987 ();
 b15zdnd00an1n02x5 FILLER_290_2051 ();
 b15zdnd00an1n01x5 FILLER_290_2053 ();
 b15zdnd11an1n32x5 FILLER_290_2059 ();
 b15zdnd11an1n08x5 FILLER_290_2091 ();
 b15zdnd11an1n04x5 FILLER_290_2099 ();
 b15zdnd00an1n02x5 FILLER_290_2103 ();
 b15zdnd00an1n01x5 FILLER_290_2105 ();
 b15zdnd11an1n04x5 FILLER_290_2112 ();
 b15zdnd00an1n01x5 FILLER_290_2116 ();
 b15zdnd11an1n16x5 FILLER_290_2123 ();
 b15zdnd11an1n08x5 FILLER_290_2139 ();
 b15zdnd11an1n04x5 FILLER_290_2147 ();
 b15zdnd00an1n02x5 FILLER_290_2151 ();
 b15zdnd00an1n01x5 FILLER_290_2153 ();
 b15zdnd11an1n32x5 FILLER_290_2162 ();
 b15zdnd11an1n08x5 FILLER_290_2194 ();
 b15zdnd00an1n01x5 FILLER_290_2202 ();
 b15zdnd11an1n08x5 FILLER_290_2208 ();
 b15zdnd11an1n04x5 FILLER_290_2216 ();
 b15zdnd00an1n01x5 FILLER_290_2220 ();
 b15zdnd11an1n04x5 FILLER_290_2230 ();
 b15zdnd11an1n08x5 FILLER_290_2239 ();
 b15zdnd11an1n04x5 FILLER_290_2247 ();
 b15zdnd00an1n02x5 FILLER_290_2251 ();
 b15zdnd11an1n16x5 FILLER_290_2260 ();
 b15zdnd11an1n32x5 FILLER_291_0 ();
 b15zdnd11an1n04x5 FILLER_291_32 ();
 b15zdnd00an1n01x5 FILLER_291_36 ();
 b15zdnd11an1n08x5 FILLER_291_55 ();
 b15zdnd11an1n04x5 FILLER_291_63 ();
 b15zdnd00an1n02x5 FILLER_291_67 ();
 b15zdnd00an1n01x5 FILLER_291_69 ();
 b15zdnd11an1n32x5 FILLER_291_76 ();
 b15zdnd11an1n08x5 FILLER_291_108 ();
 b15zdnd11an1n04x5 FILLER_291_116 ();
 b15zdnd11an1n64x5 FILLER_291_124 ();
 b15zdnd11an1n32x5 FILLER_291_188 ();
 b15zdnd11an1n32x5 FILLER_291_227 ();
 b15zdnd11an1n08x5 FILLER_291_259 ();
 b15zdnd11an1n04x5 FILLER_291_267 ();
 b15zdnd00an1n02x5 FILLER_291_271 ();
 b15zdnd11an1n04x5 FILLER_291_280 ();
 b15zdnd11an1n04x5 FILLER_291_288 ();
 b15zdnd00an1n01x5 FILLER_291_292 ();
 b15zdnd11an1n08x5 FILLER_291_307 ();
 b15zdnd11an1n04x5 FILLER_291_315 ();
 b15zdnd11an1n04x5 FILLER_291_335 ();
 b15zdnd11an1n16x5 FILLER_291_344 ();
 b15zdnd00an1n02x5 FILLER_291_360 ();
 b15zdnd00an1n01x5 FILLER_291_362 ();
 b15zdnd11an1n64x5 FILLER_291_383 ();
 b15zdnd11an1n32x5 FILLER_291_447 ();
 b15zdnd00an1n02x5 FILLER_291_479 ();
 b15zdnd11an1n16x5 FILLER_291_497 ();
 b15zdnd11an1n04x5 FILLER_291_513 ();
 b15zdnd00an1n01x5 FILLER_291_517 ();
 b15zdnd11an1n16x5 FILLER_291_524 ();
 b15zdnd11an1n08x5 FILLER_291_540 ();
 b15zdnd00an1n02x5 FILLER_291_548 ();
 b15zdnd00an1n01x5 FILLER_291_550 ();
 b15zdnd11an1n16x5 FILLER_291_558 ();
 b15zdnd00an1n01x5 FILLER_291_574 ();
 b15zdnd11an1n32x5 FILLER_291_587 ();
 b15zdnd11an1n16x5 FILLER_291_619 ();
 b15zdnd11an1n04x5 FILLER_291_635 ();
 b15zdnd00an1n02x5 FILLER_291_639 ();
 b15zdnd00an1n01x5 FILLER_291_641 ();
 b15zdnd11an1n16x5 FILLER_291_654 ();
 b15zdnd11an1n08x5 FILLER_291_670 ();
 b15zdnd00an1n02x5 FILLER_291_678 ();
 b15zdnd11an1n64x5 FILLER_291_685 ();
 b15zdnd11an1n32x5 FILLER_291_749 ();
 b15zdnd11an1n04x5 FILLER_291_781 ();
 b15zdnd00an1n02x5 FILLER_291_785 ();
 b15zdnd11an1n64x5 FILLER_291_808 ();
 b15zdnd11an1n08x5 FILLER_291_872 ();
 b15zdnd11an1n04x5 FILLER_291_880 ();
 b15zdnd00an1n02x5 FILLER_291_884 ();
 b15zdnd00an1n01x5 FILLER_291_886 ();
 b15zdnd11an1n64x5 FILLER_291_899 ();
 b15zdnd11an1n08x5 FILLER_291_963 ();
 b15zdnd11an1n04x5 FILLER_291_971 ();
 b15zdnd00an1n01x5 FILLER_291_975 ();
 b15zdnd11an1n04x5 FILLER_291_989 ();
 b15zdnd00an1n02x5 FILLER_291_993 ();
 b15zdnd00an1n01x5 FILLER_291_995 ();
 b15zdnd11an1n32x5 FILLER_291_1002 ();
 b15zdnd11an1n08x5 FILLER_291_1034 ();
 b15zdnd11an1n04x5 FILLER_291_1042 ();
 b15zdnd00an1n02x5 FILLER_291_1046 ();
 b15zdnd11an1n64x5 FILLER_291_1057 ();
 b15zdnd11an1n16x5 FILLER_291_1121 ();
 b15zdnd11an1n08x5 FILLER_291_1137 ();
 b15zdnd00an1n01x5 FILLER_291_1145 ();
 b15zdnd11an1n32x5 FILLER_291_1157 ();
 b15zdnd11an1n16x5 FILLER_291_1189 ();
 b15zdnd11an1n08x5 FILLER_291_1205 ();
 b15zdnd11an1n04x5 FILLER_291_1213 ();
 b15zdnd00an1n02x5 FILLER_291_1217 ();
 b15zdnd00an1n01x5 FILLER_291_1219 ();
 b15zdnd11an1n08x5 FILLER_291_1231 ();
 b15zdnd00an1n01x5 FILLER_291_1239 ();
 b15zdnd11an1n16x5 FILLER_291_1248 ();
 b15zdnd11an1n08x5 FILLER_291_1264 ();
 b15zdnd11an1n04x5 FILLER_291_1272 ();
 b15zdnd00an1n02x5 FILLER_291_1276 ();
 b15zdnd00an1n01x5 FILLER_291_1278 ();
 b15zdnd11an1n04x5 FILLER_291_1285 ();
 b15zdnd11an1n32x5 FILLER_291_1297 ();
 b15zdnd00an1n02x5 FILLER_291_1329 ();
 b15zdnd00an1n01x5 FILLER_291_1331 ();
 b15zdnd11an1n64x5 FILLER_291_1344 ();
 b15zdnd11an1n32x5 FILLER_291_1408 ();
 b15zdnd11an1n08x5 FILLER_291_1440 ();
 b15zdnd00an1n01x5 FILLER_291_1448 ();
 b15zdnd11an1n16x5 FILLER_291_1463 ();
 b15zdnd11an1n08x5 FILLER_291_1479 ();
 b15zdnd11an1n04x5 FILLER_291_1487 ();
 b15zdnd00an1n02x5 FILLER_291_1491 ();
 b15zdnd00an1n01x5 FILLER_291_1493 ();
 b15zdnd11an1n04x5 FILLER_291_1501 ();
 b15zdnd00an1n01x5 FILLER_291_1505 ();
 b15zdnd11an1n04x5 FILLER_291_1532 ();
 b15zdnd11an1n04x5 FILLER_291_1548 ();
 b15zdnd11an1n04x5 FILLER_291_1573 ();
 b15zdnd11an1n32x5 FILLER_291_1586 ();
 b15zdnd00an1n02x5 FILLER_291_1618 ();
 b15zdnd00an1n01x5 FILLER_291_1620 ();
 b15zdnd11an1n32x5 FILLER_291_1635 ();
 b15zdnd11an1n16x5 FILLER_291_1667 ();
 b15zdnd00an1n02x5 FILLER_291_1683 ();
 b15zdnd11an1n16x5 FILLER_291_1690 ();
 b15zdnd11an1n08x5 FILLER_291_1711 ();
 b15zdnd11an1n04x5 FILLER_291_1719 ();
 b15zdnd11an1n04x5 FILLER_291_1731 ();
 b15zdnd11an1n32x5 FILLER_291_1740 ();
 b15zdnd11an1n04x5 FILLER_291_1779 ();
 b15zdnd11an1n16x5 FILLER_291_1787 ();
 b15zdnd11an1n08x5 FILLER_291_1803 ();
 b15zdnd00an1n02x5 FILLER_291_1811 ();
 b15zdnd11an1n64x5 FILLER_291_1822 ();
 b15zdnd11an1n64x5 FILLER_291_1886 ();
 b15zdnd11an1n16x5 FILLER_291_1950 ();
 b15zdnd11an1n08x5 FILLER_291_1973 ();
 b15zdnd11an1n16x5 FILLER_291_1995 ();
 b15zdnd00an1n01x5 FILLER_291_2011 ();
 b15zdnd11an1n16x5 FILLER_291_2033 ();
 b15zdnd11an1n04x5 FILLER_291_2049 ();
 b15zdnd00an1n02x5 FILLER_291_2053 ();
 b15zdnd00an1n01x5 FILLER_291_2055 ();
 b15zdnd11an1n04x5 FILLER_291_2061 ();
 b15zdnd00an1n02x5 FILLER_291_2065 ();
 b15zdnd00an1n01x5 FILLER_291_2067 ();
 b15zdnd11an1n08x5 FILLER_291_2075 ();
 b15zdnd00an1n02x5 FILLER_291_2083 ();
 b15zdnd11an1n04x5 FILLER_291_2095 ();
 b15zdnd00an1n02x5 FILLER_291_2099 ();
 b15zdnd00an1n01x5 FILLER_291_2101 ();
 b15zdnd11an1n08x5 FILLER_291_2109 ();
 b15zdnd00an1n02x5 FILLER_291_2117 ();
 b15zdnd11an1n16x5 FILLER_291_2123 ();
 b15zdnd00an1n02x5 FILLER_291_2139 ();
 b15zdnd11an1n16x5 FILLER_291_2145 ();
 b15zdnd00an1n02x5 FILLER_291_2161 ();
 b15zdnd00an1n01x5 FILLER_291_2163 ();
 b15zdnd11an1n32x5 FILLER_291_2182 ();
 b15zdnd11an1n16x5 FILLER_291_2214 ();
 b15zdnd11an1n32x5 FILLER_291_2240 ();
 b15zdnd11an1n08x5 FILLER_291_2272 ();
 b15zdnd11an1n04x5 FILLER_291_2280 ();
 b15zdnd11an1n32x5 FILLER_292_8 ();
 b15zdnd11an1n04x5 FILLER_292_40 ();
 b15zdnd00an1n01x5 FILLER_292_44 ();
 b15zdnd11an1n16x5 FILLER_292_63 ();
 b15zdnd11an1n08x5 FILLER_292_79 ();
 b15zdnd11an1n04x5 FILLER_292_87 ();
 b15zdnd11an1n64x5 FILLER_292_104 ();
 b15zdnd11an1n08x5 FILLER_292_168 ();
 b15zdnd11an1n04x5 FILLER_292_176 ();
 b15zdnd00an1n02x5 FILLER_292_180 ();
 b15zdnd11an1n16x5 FILLER_292_197 ();
 b15zdnd11an1n04x5 FILLER_292_213 ();
 b15zdnd00an1n01x5 FILLER_292_217 ();
 b15zdnd11an1n32x5 FILLER_292_224 ();
 b15zdnd11an1n16x5 FILLER_292_256 ();
 b15zdnd11an1n04x5 FILLER_292_272 ();
 b15zdnd11an1n08x5 FILLER_292_284 ();
 b15zdnd11an1n16x5 FILLER_292_296 ();
 b15zdnd11an1n08x5 FILLER_292_312 ();
 b15zdnd00an1n01x5 FILLER_292_320 ();
 b15zdnd11an1n64x5 FILLER_292_337 ();
 b15zdnd11an1n16x5 FILLER_292_401 ();
 b15zdnd11an1n08x5 FILLER_292_417 ();
 b15zdnd11an1n04x5 FILLER_292_425 ();
 b15zdnd00an1n02x5 FILLER_292_429 ();
 b15zdnd00an1n01x5 FILLER_292_431 ();
 b15zdnd11an1n16x5 FILLER_292_448 ();
 b15zdnd00an1n01x5 FILLER_292_464 ();
 b15zdnd11an1n16x5 FILLER_292_475 ();
 b15zdnd11an1n08x5 FILLER_292_497 ();
 b15zdnd11an1n04x5 FILLER_292_505 ();
 b15zdnd00an1n01x5 FILLER_292_509 ();
 b15zdnd11an1n04x5 FILLER_292_515 ();
 b15zdnd00an1n01x5 FILLER_292_519 ();
 b15zdnd11an1n64x5 FILLER_292_530 ();
 b15zdnd11an1n64x5 FILLER_292_594 ();
 b15zdnd11an1n32x5 FILLER_292_658 ();
 b15zdnd11an1n04x5 FILLER_292_690 ();
 b15zdnd00an1n02x5 FILLER_292_694 ();
 b15zdnd11an1n04x5 FILLER_292_714 ();
 b15zdnd00an1n02x5 FILLER_292_726 ();
 b15zdnd00an1n01x5 FILLER_292_728 ();
 b15zdnd11an1n04x5 FILLER_292_754 ();
 b15zdnd11an1n64x5 FILLER_292_762 ();
 b15zdnd11an1n08x5 FILLER_292_826 ();
 b15zdnd11an1n16x5 FILLER_292_844 ();
 b15zdnd11an1n08x5 FILLER_292_860 ();
 b15zdnd11an1n04x5 FILLER_292_893 ();
 b15zdnd11an1n16x5 FILLER_292_912 ();
 b15zdnd11an1n32x5 FILLER_292_952 ();
 b15zdnd11an1n04x5 FILLER_292_984 ();
 b15zdnd00an1n02x5 FILLER_292_988 ();
 b15zdnd00an1n01x5 FILLER_292_990 ();
 b15zdnd11an1n08x5 FILLER_292_1007 ();
 b15zdnd00an1n02x5 FILLER_292_1015 ();
 b15zdnd00an1n01x5 FILLER_292_1017 ();
 b15zdnd11an1n08x5 FILLER_292_1022 ();
 b15zdnd00an1n01x5 FILLER_292_1030 ();
 b15zdnd11an1n16x5 FILLER_292_1037 ();
 b15zdnd11an1n08x5 FILLER_292_1053 ();
 b15zdnd11an1n04x5 FILLER_292_1061 ();
 b15zdnd00an1n01x5 FILLER_292_1065 ();
 b15zdnd11an1n04x5 FILLER_292_1082 ();
 b15zdnd11an1n16x5 FILLER_292_1092 ();
 b15zdnd00an1n01x5 FILLER_292_1108 ();
 b15zdnd11an1n32x5 FILLER_292_1117 ();
 b15zdnd11an1n16x5 FILLER_292_1149 ();
 b15zdnd11an1n04x5 FILLER_292_1165 ();
 b15zdnd00an1n01x5 FILLER_292_1169 ();
 b15zdnd11an1n64x5 FILLER_292_1177 ();
 b15zdnd11an1n32x5 FILLER_292_1241 ();
 b15zdnd11an1n04x5 FILLER_292_1273 ();
 b15zdnd11an1n04x5 FILLER_292_1284 ();
 b15zdnd11an1n04x5 FILLER_292_1295 ();
 b15zdnd11an1n16x5 FILLER_292_1308 ();
 b15zdnd00an1n01x5 FILLER_292_1324 ();
 b15zdnd11an1n16x5 FILLER_292_1330 ();
 b15zdnd11an1n08x5 FILLER_292_1346 ();
 b15zdnd11an1n04x5 FILLER_292_1354 ();
 b15zdnd11an1n32x5 FILLER_292_1378 ();
 b15zdnd11an1n16x5 FILLER_292_1410 ();
 b15zdnd11an1n04x5 FILLER_292_1426 ();
 b15zdnd00an1n02x5 FILLER_292_1430 ();
 b15zdnd00an1n01x5 FILLER_292_1432 ();
 b15zdnd11an1n04x5 FILLER_292_1457 ();
 b15zdnd11an1n32x5 FILLER_292_1473 ();
 b15zdnd11an1n32x5 FILLER_292_1509 ();
 b15zdnd11an1n16x5 FILLER_292_1541 ();
 b15zdnd00an1n02x5 FILLER_292_1557 ();
 b15zdnd00an1n01x5 FILLER_292_1559 ();
 b15zdnd11an1n04x5 FILLER_292_1581 ();
 b15zdnd11an1n16x5 FILLER_292_1592 ();
 b15zdnd11an1n08x5 FILLER_292_1608 ();
 b15zdnd11an1n04x5 FILLER_292_1616 ();
 b15zdnd00an1n02x5 FILLER_292_1620 ();
 b15zdnd00an1n01x5 FILLER_292_1622 ();
 b15zdnd11an1n08x5 FILLER_292_1643 ();
 b15zdnd11an1n04x5 FILLER_292_1651 ();
 b15zdnd00an1n02x5 FILLER_292_1655 ();
 b15zdnd11an1n08x5 FILLER_292_1669 ();
 b15zdnd00an1n02x5 FILLER_292_1677 ();
 b15zdnd11an1n16x5 FILLER_292_1689 ();
 b15zdnd11an1n04x5 FILLER_292_1705 ();
 b15zdnd00an1n02x5 FILLER_292_1709 ();
 b15zdnd11an1n08x5 FILLER_292_1718 ();
 b15zdnd11an1n04x5 FILLER_292_1726 ();
 b15zdnd00an1n02x5 FILLER_292_1730 ();
 b15zdnd11an1n32x5 FILLER_292_1737 ();
 b15zdnd11an1n08x5 FILLER_292_1769 ();
 b15zdnd00an1n02x5 FILLER_292_1777 ();
 b15zdnd00an1n01x5 FILLER_292_1779 ();
 b15zdnd11an1n08x5 FILLER_292_1789 ();
 b15zdnd11an1n04x5 FILLER_292_1803 ();
 b15zdnd11an1n08x5 FILLER_292_1812 ();
 b15zdnd11an1n64x5 FILLER_292_1825 ();
 b15zdnd11an1n32x5 FILLER_292_1920 ();
 b15zdnd11an1n08x5 FILLER_292_1952 ();
 b15zdnd11an1n04x5 FILLER_292_1960 ();
 b15zdnd00an1n01x5 FILLER_292_1964 ();
 b15zdnd11an1n16x5 FILLER_292_1970 ();
 b15zdnd11an1n64x5 FILLER_292_2006 ();
 b15zdnd11an1n08x5 FILLER_292_2070 ();
 b15zdnd00an1n02x5 FILLER_292_2078 ();
 b15zdnd11an1n04x5 FILLER_292_2085 ();
 b15zdnd11an1n04x5 FILLER_292_2093 ();
 b15zdnd11an1n32x5 FILLER_292_2103 ();
 b15zdnd11an1n04x5 FILLER_292_2135 ();
 b15zdnd00an1n02x5 FILLER_292_2151 ();
 b15zdnd00an1n01x5 FILLER_292_2153 ();
 b15zdnd11an1n64x5 FILLER_292_2162 ();
 b15zdnd11an1n32x5 FILLER_292_2226 ();
 b15zdnd11an1n16x5 FILLER_292_2258 ();
 b15zdnd00an1n02x5 FILLER_292_2274 ();
 b15zdnd11an1n64x5 FILLER_293_0 ();
 b15zdnd11an1n08x5 FILLER_293_64 ();
 b15zdnd00an1n01x5 FILLER_293_72 ();
 b15zdnd11an1n04x5 FILLER_293_78 ();
 b15zdnd00an1n01x5 FILLER_293_82 ();
 b15zdnd11an1n32x5 FILLER_293_92 ();
 b15zdnd11an1n16x5 FILLER_293_124 ();
 b15zdnd11an1n04x5 FILLER_293_140 ();
 b15zdnd11an1n04x5 FILLER_293_149 ();
 b15zdnd00an1n01x5 FILLER_293_153 ();
 b15zdnd11an1n04x5 FILLER_293_168 ();
 b15zdnd11an1n64x5 FILLER_293_184 ();
 b15zdnd11an1n08x5 FILLER_293_248 ();
 b15zdnd00an1n01x5 FILLER_293_256 ();
 b15zdnd11an1n16x5 FILLER_293_271 ();
 b15zdnd00an1n01x5 FILLER_293_287 ();
 b15zdnd11an1n64x5 FILLER_293_300 ();
 b15zdnd11an1n64x5 FILLER_293_364 ();
 b15zdnd11an1n32x5 FILLER_293_428 ();
 b15zdnd00an1n02x5 FILLER_293_460 ();
 b15zdnd00an1n01x5 FILLER_293_462 ();
 b15zdnd11an1n16x5 FILLER_293_482 ();
 b15zdnd11an1n04x5 FILLER_293_498 ();
 b15zdnd00an1n02x5 FILLER_293_502 ();
 b15zdnd11an1n32x5 FILLER_293_508 ();
 b15zdnd11an1n08x5 FILLER_293_540 ();
 b15zdnd00an1n01x5 FILLER_293_548 ();
 b15zdnd11an1n08x5 FILLER_293_557 ();
 b15zdnd11an1n04x5 FILLER_293_565 ();
 b15zdnd00an1n01x5 FILLER_293_569 ();
 b15zdnd11an1n64x5 FILLER_293_584 ();
 b15zdnd11an1n32x5 FILLER_293_648 ();
 b15zdnd11an1n16x5 FILLER_293_680 ();
 b15zdnd00an1n02x5 FILLER_293_696 ();
 b15zdnd00an1n01x5 FILLER_293_698 ();
 b15zdnd11an1n16x5 FILLER_293_703 ();
 b15zdnd11an1n04x5 FILLER_293_719 ();
 b15zdnd00an1n02x5 FILLER_293_723 ();
 b15zdnd11an1n16x5 FILLER_293_729 ();
 b15zdnd11an1n04x5 FILLER_293_745 ();
 b15zdnd00an1n02x5 FILLER_293_749 ();
 b15zdnd00an1n01x5 FILLER_293_751 ();
 b15zdnd11an1n08x5 FILLER_293_764 ();
 b15zdnd11an1n32x5 FILLER_293_784 ();
 b15zdnd11an1n16x5 FILLER_293_816 ();
 b15zdnd11an1n04x5 FILLER_293_832 ();
 b15zdnd11an1n64x5 FILLER_293_847 ();
 b15zdnd11an1n32x5 FILLER_293_911 ();
 b15zdnd00an1n02x5 FILLER_293_943 ();
 b15zdnd11an1n08x5 FILLER_293_970 ();
 b15zdnd11an1n04x5 FILLER_293_978 ();
 b15zdnd00an1n01x5 FILLER_293_982 ();
 b15zdnd11an1n16x5 FILLER_293_992 ();
 b15zdnd11an1n08x5 FILLER_293_1008 ();
 b15zdnd11an1n04x5 FILLER_293_1016 ();
 b15zdnd00an1n02x5 FILLER_293_1020 ();
 b15zdnd00an1n01x5 FILLER_293_1022 ();
 b15zdnd11an1n04x5 FILLER_293_1030 ();
 b15zdnd11an1n32x5 FILLER_293_1048 ();
 b15zdnd00an1n02x5 FILLER_293_1080 ();
 b15zdnd00an1n01x5 FILLER_293_1082 ();
 b15zdnd11an1n08x5 FILLER_293_1089 ();
 b15zdnd00an1n02x5 FILLER_293_1097 ();
 b15zdnd00an1n01x5 FILLER_293_1099 ();
 b15zdnd11an1n04x5 FILLER_293_1111 ();
 b15zdnd11an1n32x5 FILLER_293_1119 ();
 b15zdnd11an1n16x5 FILLER_293_1151 ();
 b15zdnd11an1n04x5 FILLER_293_1167 ();
 b15zdnd00an1n02x5 FILLER_293_1171 ();
 b15zdnd00an1n01x5 FILLER_293_1173 ();
 b15zdnd11an1n04x5 FILLER_293_1189 ();
 b15zdnd11an1n64x5 FILLER_293_1199 ();
 b15zdnd11an1n04x5 FILLER_293_1263 ();
 b15zdnd00an1n02x5 FILLER_293_1267 ();
 b15zdnd00an1n01x5 FILLER_293_1269 ();
 b15zdnd11an1n16x5 FILLER_293_1296 ();
 b15zdnd00an1n01x5 FILLER_293_1312 ();
 b15zdnd11an1n08x5 FILLER_293_1325 ();
 b15zdnd00an1n01x5 FILLER_293_1333 ();
 b15zdnd11an1n64x5 FILLER_293_1355 ();
 b15zdnd11an1n16x5 FILLER_293_1419 ();
 b15zdnd11an1n04x5 FILLER_293_1451 ();
 b15zdnd00an1n02x5 FILLER_293_1455 ();
 b15zdnd11an1n04x5 FILLER_293_1463 ();
 b15zdnd11an1n08x5 FILLER_293_1472 ();
 b15zdnd11an1n04x5 FILLER_293_1480 ();
 b15zdnd00an1n02x5 FILLER_293_1484 ();
 b15zdnd11an1n64x5 FILLER_293_1502 ();
 b15zdnd11an1n08x5 FILLER_293_1566 ();
 b15zdnd11an1n04x5 FILLER_293_1574 ();
 b15zdnd00an1n01x5 FILLER_293_1578 ();
 b15zdnd11an1n16x5 FILLER_293_1585 ();
 b15zdnd00an1n02x5 FILLER_293_1601 ();
 b15zdnd11an1n08x5 FILLER_293_1609 ();
 b15zdnd00an1n02x5 FILLER_293_1617 ();
 b15zdnd11an1n16x5 FILLER_293_1631 ();
 b15zdnd11an1n08x5 FILLER_293_1647 ();
 b15zdnd00an1n01x5 FILLER_293_1655 ();
 b15zdnd11an1n08x5 FILLER_293_1664 ();
 b15zdnd11an1n04x5 FILLER_293_1672 ();
 b15zdnd00an1n01x5 FILLER_293_1676 ();
 b15zdnd11an1n64x5 FILLER_293_1684 ();
 b15zdnd11an1n32x5 FILLER_293_1748 ();
 b15zdnd11an1n04x5 FILLER_293_1780 ();
 b15zdnd11an1n64x5 FILLER_293_1796 ();
 b15zdnd11an1n32x5 FILLER_293_1860 ();
 b15zdnd11an1n16x5 FILLER_293_1892 ();
 b15zdnd11an1n08x5 FILLER_293_1908 ();
 b15zdnd00an1n01x5 FILLER_293_1916 ();
 b15zdnd11an1n32x5 FILLER_293_1929 ();
 b15zdnd11an1n16x5 FILLER_293_1961 ();
 b15zdnd11an1n08x5 FILLER_293_1977 ();
 b15zdnd11an1n04x5 FILLER_293_1985 ();
 b15zdnd00an1n02x5 FILLER_293_1989 ();
 b15zdnd11an1n04x5 FILLER_293_2003 ();
 b15zdnd11an1n64x5 FILLER_293_2021 ();
 b15zdnd11an1n32x5 FILLER_293_2085 ();
 b15zdnd11an1n08x5 FILLER_293_2117 ();
 b15zdnd11an1n04x5 FILLER_293_2156 ();
 b15zdnd00an1n02x5 FILLER_293_2160 ();
 b15zdnd00an1n01x5 FILLER_293_2162 ();
 b15zdnd11an1n16x5 FILLER_293_2169 ();
 b15zdnd11an1n08x5 FILLER_293_2185 ();
 b15zdnd00an1n02x5 FILLER_293_2193 ();
 b15zdnd00an1n01x5 FILLER_293_2195 ();
 b15zdnd11an1n64x5 FILLER_293_2208 ();
 b15zdnd11an1n08x5 FILLER_293_2272 ();
 b15zdnd11an1n04x5 FILLER_293_2280 ();
 b15zdnd11an1n32x5 FILLER_294_8 ();
 b15zdnd00an1n02x5 FILLER_294_40 ();
 b15zdnd00an1n01x5 FILLER_294_42 ();
 b15zdnd11an1n32x5 FILLER_294_57 ();
 b15zdnd11an1n04x5 FILLER_294_89 ();
 b15zdnd00an1n02x5 FILLER_294_93 ();
 b15zdnd11an1n04x5 FILLER_294_101 ();
 b15zdnd11an1n32x5 FILLER_294_121 ();
 b15zdnd11an1n16x5 FILLER_294_153 ();
 b15zdnd11an1n08x5 FILLER_294_169 ();
 b15zdnd00an1n02x5 FILLER_294_177 ();
 b15zdnd00an1n01x5 FILLER_294_179 ();
 b15zdnd11an1n16x5 FILLER_294_200 ();
 b15zdnd11an1n08x5 FILLER_294_216 ();
 b15zdnd00an1n01x5 FILLER_294_224 ();
 b15zdnd11an1n64x5 FILLER_294_256 ();
 b15zdnd11an1n16x5 FILLER_294_320 ();
 b15zdnd11an1n08x5 FILLER_294_336 ();
 b15zdnd00an1n01x5 FILLER_294_344 ();
 b15zdnd11an1n64x5 FILLER_294_366 ();
 b15zdnd11an1n08x5 FILLER_294_430 ();
 b15zdnd00an1n01x5 FILLER_294_438 ();
 b15zdnd11an1n64x5 FILLER_294_449 ();
 b15zdnd11an1n08x5 FILLER_294_513 ();
 b15zdnd11an1n04x5 FILLER_294_521 ();
 b15zdnd00an1n02x5 FILLER_294_525 ();
 b15zdnd11an1n08x5 FILLER_294_531 ();
 b15zdnd00an1n01x5 FILLER_294_539 ();
 b15zdnd11an1n16x5 FILLER_294_558 ();
 b15zdnd11an1n04x5 FILLER_294_574 ();
 b15zdnd00an1n02x5 FILLER_294_578 ();
 b15zdnd00an1n01x5 FILLER_294_580 ();
 b15zdnd11an1n32x5 FILLER_294_586 ();
 b15zdnd11an1n08x5 FILLER_294_618 ();
 b15zdnd11an1n64x5 FILLER_294_639 ();
 b15zdnd11an1n08x5 FILLER_294_703 ();
 b15zdnd11an1n04x5 FILLER_294_711 ();
 b15zdnd00an1n02x5 FILLER_294_715 ();
 b15zdnd00an1n01x5 FILLER_294_717 ();
 b15zdnd11an1n16x5 FILLER_294_726 ();
 b15zdnd00an1n02x5 FILLER_294_742 ();
 b15zdnd00an1n01x5 FILLER_294_744 ();
 b15zdnd11an1n16x5 FILLER_294_750 ();
 b15zdnd11an1n04x5 FILLER_294_766 ();
 b15zdnd11an1n64x5 FILLER_294_778 ();
 b15zdnd11an1n32x5 FILLER_294_842 ();
 b15zdnd11an1n16x5 FILLER_294_874 ();
 b15zdnd11an1n04x5 FILLER_294_890 ();
 b15zdnd00an1n02x5 FILLER_294_894 ();
 b15zdnd11an1n64x5 FILLER_294_913 ();
 b15zdnd11an1n32x5 FILLER_294_977 ();
 b15zdnd11an1n08x5 FILLER_294_1009 ();
 b15zdnd11an1n04x5 FILLER_294_1017 ();
 b15zdnd00an1n02x5 FILLER_294_1021 ();
 b15zdnd00an1n01x5 FILLER_294_1023 ();
 b15zdnd11an1n32x5 FILLER_294_1040 ();
 b15zdnd11an1n16x5 FILLER_294_1072 ();
 b15zdnd11an1n04x5 FILLER_294_1088 ();
 b15zdnd00an1n02x5 FILLER_294_1092 ();
 b15zdnd00an1n01x5 FILLER_294_1094 ();
 b15zdnd11an1n16x5 FILLER_294_1108 ();
 b15zdnd11an1n04x5 FILLER_294_1124 ();
 b15zdnd11an1n16x5 FILLER_294_1132 ();
 b15zdnd11an1n04x5 FILLER_294_1148 ();
 b15zdnd00an1n02x5 FILLER_294_1152 ();
 b15zdnd11an1n08x5 FILLER_294_1163 ();
 b15zdnd11an1n04x5 FILLER_294_1171 ();
 b15zdnd00an1n02x5 FILLER_294_1175 ();
 b15zdnd00an1n01x5 FILLER_294_1177 ();
 b15zdnd11an1n64x5 FILLER_294_1184 ();
 b15zdnd11an1n16x5 FILLER_294_1248 ();
 b15zdnd11an1n04x5 FILLER_294_1264 ();
 b15zdnd00an1n01x5 FILLER_294_1268 ();
 b15zdnd11an1n32x5 FILLER_294_1275 ();
 b15zdnd00an1n02x5 FILLER_294_1307 ();
 b15zdnd00an1n01x5 FILLER_294_1309 ();
 b15zdnd11an1n16x5 FILLER_294_1323 ();
 b15zdnd11an1n04x5 FILLER_294_1344 ();
 b15zdnd11an1n64x5 FILLER_294_1353 ();
 b15zdnd11an1n64x5 FILLER_294_1417 ();
 b15zdnd11an1n04x5 FILLER_294_1481 ();
 b15zdnd00an1n02x5 FILLER_294_1485 ();
 b15zdnd00an1n01x5 FILLER_294_1487 ();
 b15zdnd11an1n16x5 FILLER_294_1508 ();
 b15zdnd11an1n08x5 FILLER_294_1524 ();
 b15zdnd11an1n04x5 FILLER_294_1532 ();
 b15zdnd00an1n02x5 FILLER_294_1536 ();
 b15zdnd00an1n01x5 FILLER_294_1538 ();
 b15zdnd11an1n64x5 FILLER_294_1545 ();
 b15zdnd11an1n16x5 FILLER_294_1609 ();
 b15zdnd11an1n08x5 FILLER_294_1625 ();
 b15zdnd11an1n04x5 FILLER_294_1633 ();
 b15zdnd00an1n02x5 FILLER_294_1637 ();
 b15zdnd00an1n01x5 FILLER_294_1639 ();
 b15zdnd11an1n64x5 FILLER_294_1651 ();
 b15zdnd11an1n32x5 FILLER_294_1715 ();
 b15zdnd11an1n16x5 FILLER_294_1747 ();
 b15zdnd00an1n01x5 FILLER_294_1763 ();
 b15zdnd11an1n64x5 FILLER_294_1768 ();
 b15zdnd11an1n64x5 FILLER_294_1832 ();
 b15zdnd11an1n04x5 FILLER_294_1896 ();
 b15zdnd00an1n02x5 FILLER_294_1900 ();
 b15zdnd11an1n32x5 FILLER_294_1923 ();
 b15zdnd11an1n16x5 FILLER_294_1955 ();
 b15zdnd11an1n08x5 FILLER_294_1971 ();
 b15zdnd00an1n01x5 FILLER_294_1979 ();
 b15zdnd11an1n16x5 FILLER_294_1986 ();
 b15zdnd11an1n08x5 FILLER_294_2002 ();
 b15zdnd11an1n04x5 FILLER_294_2010 ();
 b15zdnd00an1n02x5 FILLER_294_2014 ();
 b15zdnd00an1n01x5 FILLER_294_2016 ();
 b15zdnd11an1n04x5 FILLER_294_2032 ();
 b15zdnd11an1n08x5 FILLER_294_2043 ();
 b15zdnd00an1n02x5 FILLER_294_2051 ();
 b15zdnd11an1n64x5 FILLER_294_2066 ();
 b15zdnd11an1n16x5 FILLER_294_2130 ();
 b15zdnd11an1n08x5 FILLER_294_2146 ();
 b15zdnd11an1n04x5 FILLER_294_2162 ();
 b15zdnd11an1n16x5 FILLER_294_2171 ();
 b15zdnd11an1n08x5 FILLER_294_2187 ();
 b15zdnd11an1n04x5 FILLER_294_2195 ();
 b15zdnd00an1n01x5 FILLER_294_2199 ();
 b15zdnd11an1n04x5 FILLER_294_2206 ();
 b15zdnd00an1n01x5 FILLER_294_2210 ();
 b15zdnd11an1n04x5 FILLER_294_2227 ();
 b15zdnd00an1n02x5 FILLER_294_2231 ();
 b15zdnd00an1n01x5 FILLER_294_2233 ();
 b15zdnd11an1n16x5 FILLER_294_2249 ();
 b15zdnd11an1n08x5 FILLER_294_2265 ();
 b15zdnd00an1n02x5 FILLER_294_2273 ();
 b15zdnd00an1n01x5 FILLER_294_2275 ();
 b15zdnd11an1n32x5 FILLER_295_0 ();
 b15zdnd11an1n08x5 FILLER_295_32 ();
 b15zdnd00an1n02x5 FILLER_295_40 ();
 b15zdnd00an1n01x5 FILLER_295_42 ();
 b15zdnd11an1n04x5 FILLER_295_74 ();
 b15zdnd00an1n01x5 FILLER_295_78 ();
 b15zdnd11an1n64x5 FILLER_295_110 ();
 b15zdnd11an1n08x5 FILLER_295_174 ();
 b15zdnd00an1n02x5 FILLER_295_182 ();
 b15zdnd00an1n01x5 FILLER_295_184 ();
 b15zdnd11an1n32x5 FILLER_295_189 ();
 b15zdnd11an1n16x5 FILLER_295_221 ();
 b15zdnd11an1n04x5 FILLER_295_237 ();
 b15zdnd00an1n01x5 FILLER_295_241 ();
 b15zdnd11an1n64x5 FILLER_295_263 ();
 b15zdnd11an1n64x5 FILLER_295_327 ();
 b15zdnd11an1n32x5 FILLER_295_391 ();
 b15zdnd11an1n08x5 FILLER_295_423 ();
 b15zdnd00an1n02x5 FILLER_295_431 ();
 b15zdnd00an1n01x5 FILLER_295_433 ();
 b15zdnd11an1n08x5 FILLER_295_439 ();
 b15zdnd11an1n04x5 FILLER_295_447 ();
 b15zdnd00an1n02x5 FILLER_295_451 ();
 b15zdnd00an1n01x5 FILLER_295_453 ();
 b15zdnd11an1n04x5 FILLER_295_470 ();
 b15zdnd11an1n32x5 FILLER_295_492 ();
 b15zdnd11an1n16x5 FILLER_295_524 ();
 b15zdnd11an1n08x5 FILLER_295_540 ();
 b15zdnd11an1n04x5 FILLER_295_548 ();
 b15zdnd00an1n02x5 FILLER_295_552 ();
 b15zdnd11an1n32x5 FILLER_295_560 ();
 b15zdnd11an1n16x5 FILLER_295_592 ();
 b15zdnd11an1n08x5 FILLER_295_608 ();
 b15zdnd11an1n04x5 FILLER_295_647 ();
 b15zdnd11an1n08x5 FILLER_295_657 ();
 b15zdnd00an1n02x5 FILLER_295_665 ();
 b15zdnd00an1n01x5 FILLER_295_667 ();
 b15zdnd11an1n04x5 FILLER_295_672 ();
 b15zdnd11an1n32x5 FILLER_295_681 ();
 b15zdnd11an1n16x5 FILLER_295_713 ();
 b15zdnd11an1n08x5 FILLER_295_729 ();
 b15zdnd11an1n04x5 FILLER_295_737 ();
 b15zdnd00an1n02x5 FILLER_295_741 ();
 b15zdnd11an1n04x5 FILLER_295_766 ();
 b15zdnd11an1n64x5 FILLER_295_777 ();
 b15zdnd11an1n32x5 FILLER_295_841 ();
 b15zdnd11an1n16x5 FILLER_295_873 ();
 b15zdnd11an1n08x5 FILLER_295_889 ();
 b15zdnd00an1n02x5 FILLER_295_897 ();
 b15zdnd00an1n01x5 FILLER_295_899 ();
 b15zdnd11an1n64x5 FILLER_295_925 ();
 b15zdnd11an1n64x5 FILLER_295_989 ();
 b15zdnd11an1n04x5 FILLER_295_1053 ();
 b15zdnd00an1n02x5 FILLER_295_1057 ();
 b15zdnd11an1n64x5 FILLER_295_1066 ();
 b15zdnd11an1n16x5 FILLER_295_1130 ();
 b15zdnd11an1n08x5 FILLER_295_1146 ();
 b15zdnd00an1n01x5 FILLER_295_1154 ();
 b15zdnd11an1n16x5 FILLER_295_1167 ();
 b15zdnd11an1n04x5 FILLER_295_1183 ();
 b15zdnd11an1n04x5 FILLER_295_1193 ();
 b15zdnd11an1n16x5 FILLER_295_1203 ();
 b15zdnd11an1n08x5 FILLER_295_1219 ();
 b15zdnd00an1n01x5 FILLER_295_1227 ();
 b15zdnd11an1n32x5 FILLER_295_1234 ();
 b15zdnd00an1n02x5 FILLER_295_1266 ();
 b15zdnd00an1n01x5 FILLER_295_1268 ();
 b15zdnd11an1n04x5 FILLER_295_1285 ();
 b15zdnd11an1n08x5 FILLER_295_1294 ();
 b15zdnd00an1n01x5 FILLER_295_1302 ();
 b15zdnd11an1n64x5 FILLER_295_1326 ();
 b15zdnd11an1n64x5 FILLER_295_1390 ();
 b15zdnd11an1n32x5 FILLER_295_1454 ();
 b15zdnd11an1n16x5 FILLER_295_1486 ();
 b15zdnd00an1n02x5 FILLER_295_1502 ();
 b15zdnd11an1n64x5 FILLER_295_1514 ();
 b15zdnd11an1n64x5 FILLER_295_1578 ();
 b15zdnd11an1n32x5 FILLER_295_1642 ();
 b15zdnd11an1n16x5 FILLER_295_1674 ();
 b15zdnd11an1n08x5 FILLER_295_1690 ();
 b15zdnd11an1n04x5 FILLER_295_1698 ();
 b15zdnd11an1n32x5 FILLER_295_1709 ();
 b15zdnd11an1n08x5 FILLER_295_1741 ();
 b15zdnd11an1n04x5 FILLER_295_1749 ();
 b15zdnd11an1n08x5 FILLER_295_1764 ();
 b15zdnd00an1n02x5 FILLER_295_1772 ();
 b15zdnd11an1n64x5 FILLER_295_1790 ();
 b15zdnd11an1n16x5 FILLER_295_1854 ();
 b15zdnd11an1n04x5 FILLER_295_1870 ();
 b15zdnd11an1n04x5 FILLER_295_1906 ();
 b15zdnd11an1n08x5 FILLER_295_1916 ();
 b15zdnd11an1n16x5 FILLER_295_1944 ();
 b15zdnd11an1n04x5 FILLER_295_1960 ();
 b15zdnd00an1n02x5 FILLER_295_1964 ();
 b15zdnd11an1n04x5 FILLER_295_1979 ();
 b15zdnd11an1n64x5 FILLER_295_1989 ();
 b15zdnd11an1n32x5 FILLER_295_2053 ();
 b15zdnd11an1n08x5 FILLER_295_2085 ();
 b15zdnd00an1n01x5 FILLER_295_2093 ();
 b15zdnd11an1n32x5 FILLER_295_2108 ();
 b15zdnd11an1n16x5 FILLER_295_2140 ();
 b15zdnd11an1n04x5 FILLER_295_2156 ();
 b15zdnd00an1n02x5 FILLER_295_2160 ();
 b15zdnd11an1n04x5 FILLER_295_2176 ();
 b15zdnd11an1n08x5 FILLER_295_2193 ();
 b15zdnd00an1n02x5 FILLER_295_2201 ();
 b15zdnd00an1n01x5 FILLER_295_2203 ();
 b15zdnd11an1n08x5 FILLER_295_2220 ();
 b15zdnd00an1n02x5 FILLER_295_2228 ();
 b15zdnd11an1n32x5 FILLER_295_2248 ();
 b15zdnd11an1n04x5 FILLER_295_2280 ();
 b15zdnd11an1n16x5 FILLER_296_8 ();
 b15zdnd11an1n08x5 FILLER_296_24 ();
 b15zdnd00an1n02x5 FILLER_296_32 ();
 b15zdnd11an1n08x5 FILLER_296_65 ();
 b15zdnd00an1n02x5 FILLER_296_73 ();
 b15zdnd00an1n01x5 FILLER_296_75 ();
 b15zdnd11an1n16x5 FILLER_296_108 ();
 b15zdnd11an1n04x5 FILLER_296_124 ();
 b15zdnd00an1n02x5 FILLER_296_128 ();
 b15zdnd11an1n04x5 FILLER_296_138 ();
 b15zdnd11an1n32x5 FILLER_296_154 ();
 b15zdnd11an1n16x5 FILLER_296_186 ();
 b15zdnd11an1n04x5 FILLER_296_202 ();
 b15zdnd00an1n02x5 FILLER_296_206 ();
 b15zdnd11an1n04x5 FILLER_296_212 ();
 b15zdnd00an1n02x5 FILLER_296_216 ();
 b15zdnd00an1n01x5 FILLER_296_218 ();
 b15zdnd11an1n04x5 FILLER_296_235 ();
 b15zdnd00an1n02x5 FILLER_296_239 ();
 b15zdnd00an1n01x5 FILLER_296_241 ();
 b15zdnd11an1n32x5 FILLER_296_256 ();
 b15zdnd11an1n16x5 FILLER_296_288 ();
 b15zdnd11an1n08x5 FILLER_296_304 ();
 b15zdnd00an1n02x5 FILLER_296_312 ();
 b15zdnd00an1n01x5 FILLER_296_314 ();
 b15zdnd11an1n16x5 FILLER_296_347 ();
 b15zdnd11an1n04x5 FILLER_296_363 ();
 b15zdnd00an1n02x5 FILLER_296_367 ();
 b15zdnd11an1n64x5 FILLER_296_401 ();
 b15zdnd11an1n04x5 FILLER_296_465 ();
 b15zdnd00an1n01x5 FILLER_296_469 ();
 b15zdnd11an1n16x5 FILLER_296_488 ();
 b15zdnd11an1n08x5 FILLER_296_504 ();
 b15zdnd11an1n04x5 FILLER_296_512 ();
 b15zdnd00an1n01x5 FILLER_296_516 ();
 b15zdnd11an1n16x5 FILLER_296_533 ();
 b15zdnd00an1n02x5 FILLER_296_549 ();
 b15zdnd11an1n08x5 FILLER_296_559 ();
 b15zdnd00an1n01x5 FILLER_296_567 ();
 b15zdnd11an1n32x5 FILLER_296_576 ();
 b15zdnd11an1n16x5 FILLER_296_608 ();
 b15zdnd11an1n08x5 FILLER_296_624 ();
 b15zdnd11an1n04x5 FILLER_296_632 ();
 b15zdnd00an1n01x5 FILLER_296_636 ();
 b15zdnd11an1n04x5 FILLER_296_644 ();
 b15zdnd00an1n01x5 FILLER_296_648 ();
 b15zdnd11an1n08x5 FILLER_296_661 ();
 b15zdnd11an1n04x5 FILLER_296_669 ();
 b15zdnd00an1n02x5 FILLER_296_673 ();
 b15zdnd00an1n01x5 FILLER_296_675 ();
 b15zdnd11an1n16x5 FILLER_296_685 ();
 b15zdnd00an1n01x5 FILLER_296_701 ();
 b15zdnd00an1n02x5 FILLER_296_716 ();
 b15zdnd11an1n16x5 FILLER_296_726 ();
 b15zdnd11an1n32x5 FILLER_296_758 ();
 b15zdnd00an1n02x5 FILLER_296_790 ();
 b15zdnd11an1n04x5 FILLER_296_823 ();
 b15zdnd11an1n32x5 FILLER_296_836 ();
 b15zdnd11an1n04x5 FILLER_296_868 ();
 b15zdnd00an1n02x5 FILLER_296_872 ();
 b15zdnd00an1n01x5 FILLER_296_874 ();
 b15zdnd11an1n04x5 FILLER_296_906 ();
 b15zdnd11an1n04x5 FILLER_296_941 ();
 b15zdnd11an1n64x5 FILLER_296_970 ();
 b15zdnd11an1n08x5 FILLER_296_1034 ();
 b15zdnd11an1n04x5 FILLER_296_1042 ();
 b15zdnd00an1n02x5 FILLER_296_1046 ();
 b15zdnd00an1n01x5 FILLER_296_1048 ();
 b15zdnd11an1n04x5 FILLER_296_1056 ();
 b15zdnd11an1n08x5 FILLER_296_1079 ();
 b15zdnd00an1n01x5 FILLER_296_1087 ();
 b15zdnd11an1n04x5 FILLER_296_1100 ();
 b15zdnd11an1n08x5 FILLER_296_1111 ();
 b15zdnd11an1n04x5 FILLER_296_1119 ();
 b15zdnd00an1n02x5 FILLER_296_1123 ();
 b15zdnd00an1n01x5 FILLER_296_1125 ();
 b15zdnd11an1n64x5 FILLER_296_1132 ();
 b15zdnd11an1n04x5 FILLER_296_1196 ();
 b15zdnd00an1n02x5 FILLER_296_1200 ();
 b15zdnd11an1n04x5 FILLER_296_1226 ();
 b15zdnd11an1n16x5 FILLER_296_1244 ();
 b15zdnd11an1n08x5 FILLER_296_1260 ();
 b15zdnd00an1n02x5 FILLER_296_1268 ();
 b15zdnd11an1n16x5 FILLER_296_1275 ();
 b15zdnd11an1n08x5 FILLER_296_1291 ();
 b15zdnd00an1n02x5 FILLER_296_1299 ();
 b15zdnd11an1n08x5 FILLER_296_1317 ();
 b15zdnd11an1n04x5 FILLER_296_1325 ();
 b15zdnd00an1n02x5 FILLER_296_1329 ();
 b15zdnd11an1n64x5 FILLER_296_1342 ();
 b15zdnd00an1n01x5 FILLER_296_1406 ();
 b15zdnd11an1n64x5 FILLER_296_1427 ();
 b15zdnd11an1n04x5 FILLER_296_1491 ();
 b15zdnd00an1n02x5 FILLER_296_1495 ();
 b15zdnd11an1n04x5 FILLER_296_1504 ();
 b15zdnd11an1n04x5 FILLER_296_1536 ();
 b15zdnd00an1n02x5 FILLER_296_1540 ();
 b15zdnd11an1n16x5 FILLER_296_1555 ();
 b15zdnd11an1n04x5 FILLER_296_1571 ();
 b15zdnd11an1n08x5 FILLER_296_1583 ();
 b15zdnd11an1n04x5 FILLER_296_1591 ();
 b15zdnd00an1n02x5 FILLER_296_1595 ();
 b15zdnd00an1n01x5 FILLER_296_1597 ();
 b15zdnd11an1n64x5 FILLER_296_1604 ();
 b15zdnd11an1n32x5 FILLER_296_1668 ();
 b15zdnd11an1n08x5 FILLER_296_1700 ();
 b15zdnd11an1n04x5 FILLER_296_1708 ();
 b15zdnd00an1n02x5 FILLER_296_1712 ();
 b15zdnd11an1n08x5 FILLER_296_1723 ();
 b15zdnd00an1n01x5 FILLER_296_1731 ();
 b15zdnd11an1n08x5 FILLER_296_1748 ();
 b15zdnd11an1n04x5 FILLER_296_1756 ();
 b15zdnd00an1n01x5 FILLER_296_1760 ();
 b15zdnd11an1n04x5 FILLER_296_1768 ();
 b15zdnd11an1n64x5 FILLER_296_1777 ();
 b15zdnd11an1n32x5 FILLER_296_1841 ();
 b15zdnd11an1n16x5 FILLER_296_1873 ();
 b15zdnd11an1n08x5 FILLER_296_1889 ();
 b15zdnd11an1n04x5 FILLER_296_1897 ();
 b15zdnd11an1n16x5 FILLER_296_1932 ();
 b15zdnd00an1n02x5 FILLER_296_1948 ();
 b15zdnd11an1n08x5 FILLER_296_1968 ();
 b15zdnd00an1n02x5 FILLER_296_1976 ();
 b15zdnd00an1n01x5 FILLER_296_1978 ();
 b15zdnd11an1n32x5 FILLER_296_1989 ();
 b15zdnd11an1n16x5 FILLER_296_2021 ();
 b15zdnd11an1n08x5 FILLER_296_2037 ();
 b15zdnd11an1n04x5 FILLER_296_2045 ();
 b15zdnd00an1n02x5 FILLER_296_2049 ();
 b15zdnd00an1n01x5 FILLER_296_2051 ();
 b15zdnd11an1n64x5 FILLER_296_2059 ();
 b15zdnd11an1n16x5 FILLER_296_2123 ();
 b15zdnd11an1n08x5 FILLER_296_2139 ();
 b15zdnd11an1n04x5 FILLER_296_2147 ();
 b15zdnd00an1n02x5 FILLER_296_2151 ();
 b15zdnd00an1n01x5 FILLER_296_2153 ();
 b15zdnd11an1n04x5 FILLER_296_2162 ();
 b15zdnd00an1n01x5 FILLER_296_2166 ();
 b15zdnd11an1n08x5 FILLER_296_2187 ();
 b15zdnd11an1n04x5 FILLER_296_2195 ();
 b15zdnd11an1n16x5 FILLER_296_2205 ();
 b15zdnd11an1n08x5 FILLER_296_2221 ();
 b15zdnd11an1n04x5 FILLER_296_2229 ();
 b15zdnd00an1n01x5 FILLER_296_2233 ();
 b15zdnd11an1n32x5 FILLER_296_2243 ();
 b15zdnd00an1n01x5 FILLER_296_2275 ();
 b15zdnd11an1n32x5 FILLER_297_0 ();
 b15zdnd11an1n08x5 FILLER_297_32 ();
 b15zdnd00an1n02x5 FILLER_297_40 ();
 b15zdnd00an1n01x5 FILLER_297_42 ();
 b15zdnd11an1n16x5 FILLER_297_59 ();
 b15zdnd11an1n04x5 FILLER_297_89 ();
 b15zdnd11an1n16x5 FILLER_297_98 ();
 b15zdnd11an1n08x5 FILLER_297_114 ();
 b15zdnd11an1n04x5 FILLER_297_122 ();
 b15zdnd11an1n04x5 FILLER_297_130 ();
 b15zdnd11an1n08x5 FILLER_297_141 ();
 b15zdnd11an1n04x5 FILLER_297_149 ();
 b15zdnd00an1n02x5 FILLER_297_153 ();
 b15zdnd00an1n01x5 FILLER_297_155 ();
 b15zdnd11an1n64x5 FILLER_297_159 ();
 b15zdnd11an1n08x5 FILLER_297_223 ();
 b15zdnd11an1n04x5 FILLER_297_231 ();
 b15zdnd00an1n01x5 FILLER_297_235 ();
 b15zdnd11an1n32x5 FILLER_297_241 ();
 b15zdnd11an1n16x5 FILLER_297_273 ();
 b15zdnd11an1n08x5 FILLER_297_289 ();
 b15zdnd11an1n04x5 FILLER_297_297 ();
 b15zdnd00an1n02x5 FILLER_297_301 ();
 b15zdnd11an1n08x5 FILLER_297_316 ();
 b15zdnd00an1n02x5 FILLER_297_324 ();
 b15zdnd11an1n64x5 FILLER_297_357 ();
 b15zdnd11an1n16x5 FILLER_297_421 ();
 b15zdnd00an1n01x5 FILLER_297_437 ();
 b15zdnd11an1n16x5 FILLER_297_461 ();
 b15zdnd11an1n08x5 FILLER_297_477 ();
 b15zdnd11an1n04x5 FILLER_297_485 ();
 b15zdnd00an1n01x5 FILLER_297_489 ();
 b15zdnd11an1n16x5 FILLER_297_503 ();
 b15zdnd11an1n08x5 FILLER_297_519 ();
 b15zdnd11an1n08x5 FILLER_297_539 ();
 b15zdnd11an1n04x5 FILLER_297_547 ();
 b15zdnd00an1n01x5 FILLER_297_551 ();
 b15zdnd11an1n64x5 FILLER_297_558 ();
 b15zdnd11an1n64x5 FILLER_297_622 ();
 b15zdnd11an1n16x5 FILLER_297_686 ();
 b15zdnd00an1n01x5 FILLER_297_702 ();
 b15zdnd11an1n64x5 FILLER_297_712 ();
 b15zdnd11an1n32x5 FILLER_297_776 ();
 b15zdnd11an1n08x5 FILLER_297_808 ();
 b15zdnd11an1n04x5 FILLER_297_816 ();
 b15zdnd00an1n02x5 FILLER_297_820 ();
 b15zdnd00an1n01x5 FILLER_297_822 ();
 b15zdnd11an1n64x5 FILLER_297_832 ();
 b15zdnd11an1n64x5 FILLER_297_896 ();
 b15zdnd11an1n04x5 FILLER_297_960 ();
 b15zdnd00an1n02x5 FILLER_297_964 ();
 b15zdnd00an1n01x5 FILLER_297_966 ();
 b15zdnd11an1n32x5 FILLER_297_976 ();
 b15zdnd11an1n04x5 FILLER_297_1008 ();
 b15zdnd11an1n08x5 FILLER_297_1028 ();
 b15zdnd00an1n02x5 FILLER_297_1036 ();
 b15zdnd11an1n04x5 FILLER_297_1050 ();
 b15zdnd11an1n16x5 FILLER_297_1063 ();
 b15zdnd00an1n02x5 FILLER_297_1079 ();
 b15zdnd00an1n01x5 FILLER_297_1081 ();
 b15zdnd11an1n04x5 FILLER_297_1086 ();
 b15zdnd11an1n16x5 FILLER_297_1110 ();
 b15zdnd00an1n02x5 FILLER_297_1126 ();
 b15zdnd11an1n04x5 FILLER_297_1138 ();
 b15zdnd11an1n64x5 FILLER_297_1156 ();
 b15zdnd11an1n08x5 FILLER_297_1220 ();
 b15zdnd00an1n02x5 FILLER_297_1228 ();
 b15zdnd11an1n04x5 FILLER_297_1236 ();
 b15zdnd00an1n01x5 FILLER_297_1240 ();
 b15zdnd11an1n64x5 FILLER_297_1248 ();
 b15zdnd11an1n32x5 FILLER_297_1312 ();
 b15zdnd11an1n04x5 FILLER_297_1344 ();
 b15zdnd00an1n02x5 FILLER_297_1348 ();
 b15zdnd11an1n16x5 FILLER_297_1381 ();
 b15zdnd00an1n01x5 FILLER_297_1397 ();
 b15zdnd11an1n16x5 FILLER_297_1407 ();
 b15zdnd11an1n04x5 FILLER_297_1423 ();
 b15zdnd00an1n02x5 FILLER_297_1427 ();
 b15zdnd11an1n04x5 FILLER_297_1447 ();
 b15zdnd11an1n16x5 FILLER_297_1476 ();
 b15zdnd00an1n02x5 FILLER_297_1492 ();
 b15zdnd11an1n04x5 FILLER_297_1499 ();
 b15zdnd11an1n64x5 FILLER_297_1517 ();
 b15zdnd11an1n16x5 FILLER_297_1581 ();
 b15zdnd00an1n02x5 FILLER_297_1597 ();
 b15zdnd00an1n01x5 FILLER_297_1599 ();
 b15zdnd11an1n08x5 FILLER_297_1606 ();
 b15zdnd00an1n02x5 FILLER_297_1614 ();
 b15zdnd11an1n08x5 FILLER_297_1621 ();
 b15zdnd00an1n02x5 FILLER_297_1629 ();
 b15zdnd11an1n04x5 FILLER_297_1635 ();
 b15zdnd00an1n02x5 FILLER_297_1639 ();
 b15zdnd11an1n08x5 FILLER_297_1649 ();
 b15zdnd00an1n01x5 FILLER_297_1657 ();
 b15zdnd11an1n04x5 FILLER_297_1667 ();
 b15zdnd00an1n02x5 FILLER_297_1671 ();
 b15zdnd11an1n04x5 FILLER_297_1683 ();
 b15zdnd11an1n32x5 FILLER_297_1694 ();
 b15zdnd11an1n04x5 FILLER_297_1726 ();
 b15zdnd00an1n01x5 FILLER_297_1730 ();
 b15zdnd11an1n32x5 FILLER_297_1736 ();
 b15zdnd00an1n02x5 FILLER_297_1768 ();
 b15zdnd00an1n01x5 FILLER_297_1770 ();
 b15zdnd11an1n32x5 FILLER_297_1776 ();
 b15zdnd11an1n16x5 FILLER_297_1808 ();
 b15zdnd00an1n01x5 FILLER_297_1824 ();
 b15zdnd11an1n64x5 FILLER_297_1833 ();
 b15zdnd11an1n04x5 FILLER_297_1897 ();
 b15zdnd00an1n02x5 FILLER_297_1901 ();
 b15zdnd00an1n01x5 FILLER_297_1903 ();
 b15zdnd11an1n64x5 FILLER_297_1922 ();
 b15zdnd11an1n08x5 FILLER_297_1986 ();
 b15zdnd00an1n02x5 FILLER_297_1994 ();
 b15zdnd00an1n01x5 FILLER_297_1996 ();
 b15zdnd11an1n32x5 FILLER_297_2003 ();
 b15zdnd11an1n04x5 FILLER_297_2035 ();
 b15zdnd00an1n02x5 FILLER_297_2039 ();
 b15zdnd11an1n04x5 FILLER_297_2054 ();
 b15zdnd11an1n16x5 FILLER_297_2073 ();
 b15zdnd11an1n04x5 FILLER_297_2089 ();
 b15zdnd00an1n02x5 FILLER_297_2093 ();
 b15zdnd00an1n01x5 FILLER_297_2095 ();
 b15zdnd11an1n32x5 FILLER_297_2102 ();
 b15zdnd11an1n16x5 FILLER_297_2134 ();
 b15zdnd11an1n08x5 FILLER_297_2150 ();
 b15zdnd11an1n04x5 FILLER_297_2158 ();
 b15zdnd00an1n01x5 FILLER_297_2162 ();
 b15zdnd11an1n64x5 FILLER_297_2167 ();
 b15zdnd00an1n01x5 FILLER_297_2231 ();
 b15zdnd11an1n32x5 FILLER_297_2240 ();
 b15zdnd11an1n08x5 FILLER_297_2272 ();
 b15zdnd11an1n04x5 FILLER_297_2280 ();
 b15zdnd11an1n32x5 FILLER_298_8 ();
 b15zdnd11an1n16x5 FILLER_298_40 ();
 b15zdnd11an1n64x5 FILLER_298_74 ();
 b15zdnd11an1n16x5 FILLER_298_138 ();
 b15zdnd11an1n04x5 FILLER_298_175 ();
 b15zdnd11an1n04x5 FILLER_298_184 ();
 b15zdnd00an1n02x5 FILLER_298_188 ();
 b15zdnd11an1n04x5 FILLER_298_195 ();
 b15zdnd11an1n16x5 FILLER_298_211 ();
 b15zdnd11an1n08x5 FILLER_298_227 ();
 b15zdnd11an1n04x5 FILLER_298_235 ();
 b15zdnd11an1n04x5 FILLER_298_249 ();
 b15zdnd00an1n02x5 FILLER_298_253 ();
 b15zdnd11an1n04x5 FILLER_298_268 ();
 b15zdnd11an1n16x5 FILLER_298_276 ();
 b15zdnd11an1n04x5 FILLER_298_300 ();
 b15zdnd00an1n02x5 FILLER_298_304 ();
 b15zdnd11an1n08x5 FILLER_298_315 ();
 b15zdnd11an1n04x5 FILLER_298_323 ();
 b15zdnd00an1n02x5 FILLER_298_327 ();
 b15zdnd11an1n64x5 FILLER_298_339 ();
 b15zdnd11an1n64x5 FILLER_298_403 ();
 b15zdnd11an1n08x5 FILLER_298_467 ();
 b15zdnd00an1n02x5 FILLER_298_475 ();
 b15zdnd00an1n01x5 FILLER_298_477 ();
 b15zdnd11an1n04x5 FILLER_298_490 ();
 b15zdnd00an1n01x5 FILLER_298_494 ();
 b15zdnd11an1n32x5 FILLER_298_509 ();
 b15zdnd11an1n08x5 FILLER_298_541 ();
 b15zdnd00an1n02x5 FILLER_298_549 ();
 b15zdnd11an1n32x5 FILLER_298_555 ();
 b15zdnd11an1n08x5 FILLER_298_587 ();
 b15zdnd11an1n04x5 FILLER_298_595 ();
 b15zdnd00an1n02x5 FILLER_298_599 ();
 b15zdnd11an1n08x5 FILLER_298_610 ();
 b15zdnd00an1n02x5 FILLER_298_618 ();
 b15zdnd11an1n16x5 FILLER_298_624 ();
 b15zdnd11an1n08x5 FILLER_298_640 ();
 b15zdnd11an1n32x5 FILLER_298_655 ();
 b15zdnd11an1n16x5 FILLER_298_687 ();
 b15zdnd11an1n04x5 FILLER_298_703 ();
 b15zdnd00an1n02x5 FILLER_298_707 ();
 b15zdnd11an1n04x5 FILLER_298_713 ();
 b15zdnd00an1n01x5 FILLER_298_717 ();
 b15zdnd11an1n32x5 FILLER_298_726 ();
 b15zdnd00an1n01x5 FILLER_298_758 ();
 b15zdnd11an1n64x5 FILLER_298_777 ();
 b15zdnd11an1n08x5 FILLER_298_841 ();
 b15zdnd11an1n04x5 FILLER_298_849 ();
 b15zdnd00an1n02x5 FILLER_298_853 ();
 b15zdnd11an1n04x5 FILLER_298_880 ();
 b15zdnd11an1n64x5 FILLER_298_912 ();
 b15zdnd11an1n16x5 FILLER_298_976 ();
 b15zdnd11an1n04x5 FILLER_298_992 ();
 b15zdnd00an1n01x5 FILLER_298_996 ();
 b15zdnd11an1n32x5 FILLER_298_1013 ();
 b15zdnd11an1n08x5 FILLER_298_1045 ();
 b15zdnd00an1n02x5 FILLER_298_1053 ();
 b15zdnd00an1n01x5 FILLER_298_1055 ();
 b15zdnd11an1n64x5 FILLER_298_1063 ();
 b15zdnd11an1n32x5 FILLER_298_1127 ();
 b15zdnd11an1n08x5 FILLER_298_1159 ();
 b15zdnd11an1n04x5 FILLER_298_1167 ();
 b15zdnd11an1n64x5 FILLER_298_1176 ();
 b15zdnd11an1n16x5 FILLER_298_1240 ();
 b15zdnd11an1n08x5 FILLER_298_1256 ();
 b15zdnd11an1n04x5 FILLER_298_1264 ();
 b15zdnd00an1n02x5 FILLER_298_1268 ();
 b15zdnd00an1n01x5 FILLER_298_1270 ();
 b15zdnd11an1n64x5 FILLER_298_1277 ();
 b15zdnd11an1n64x5 FILLER_298_1341 ();
 b15zdnd11an1n16x5 FILLER_298_1405 ();
 b15zdnd11an1n08x5 FILLER_298_1421 ();
 b15zdnd00an1n02x5 FILLER_298_1429 ();
 b15zdnd00an1n01x5 FILLER_298_1431 ();
 b15zdnd11an1n08x5 FILLER_298_1457 ();
 b15zdnd11an1n04x5 FILLER_298_1465 ();
 b15zdnd00an1n02x5 FILLER_298_1469 ();
 b15zdnd00an1n01x5 FILLER_298_1471 ();
 b15zdnd11an1n08x5 FILLER_298_1479 ();
 b15zdnd11an1n04x5 FILLER_298_1487 ();
 b15zdnd00an1n02x5 FILLER_298_1491 ();
 b15zdnd00an1n01x5 FILLER_298_1493 ();
 b15zdnd11an1n32x5 FILLER_298_1504 ();
 b15zdnd11an1n16x5 FILLER_298_1536 ();
 b15zdnd00an1n02x5 FILLER_298_1552 ();
 b15zdnd00an1n01x5 FILLER_298_1554 ();
 b15zdnd11an1n32x5 FILLER_298_1560 ();
 b15zdnd11an1n08x5 FILLER_298_1592 ();
 b15zdnd11an1n32x5 FILLER_298_1606 ();
 b15zdnd11an1n08x5 FILLER_298_1638 ();
 b15zdnd00an1n02x5 FILLER_298_1646 ();
 b15zdnd00an1n01x5 FILLER_298_1648 ();
 b15zdnd11an1n04x5 FILLER_298_1655 ();
 b15zdnd00an1n02x5 FILLER_298_1659 ();
 b15zdnd11an1n08x5 FILLER_298_1681 ();
 b15zdnd00an1n02x5 FILLER_298_1689 ();
 b15zdnd11an1n04x5 FILLER_298_1701 ();
 b15zdnd11an1n16x5 FILLER_298_1717 ();
 b15zdnd00an1n02x5 FILLER_298_1733 ();
 b15zdnd00an1n01x5 FILLER_298_1735 ();
 b15zdnd11an1n32x5 FILLER_298_1757 ();
 b15zdnd11an1n16x5 FILLER_298_1789 ();
 b15zdnd11an1n08x5 FILLER_298_1805 ();
 b15zdnd11an1n04x5 FILLER_298_1813 ();
 b15zdnd11an1n04x5 FILLER_298_1826 ();
 b15zdnd11an1n04x5 FILLER_298_1842 ();
 b15zdnd11an1n04x5 FILLER_298_1866 ();
 b15zdnd11an1n64x5 FILLER_298_1896 ();
 b15zdnd11an1n16x5 FILLER_298_1960 ();
 b15zdnd11an1n04x5 FILLER_298_1976 ();
 b15zdnd11an1n04x5 FILLER_298_1994 ();
 b15zdnd11an1n08x5 FILLER_298_2016 ();
 b15zdnd11an1n04x5 FILLER_298_2024 ();
 b15zdnd00an1n02x5 FILLER_298_2028 ();
 b15zdnd00an1n01x5 FILLER_298_2030 ();
 b15zdnd11an1n16x5 FILLER_298_2045 ();
 b15zdnd00an1n02x5 FILLER_298_2061 ();
 b15zdnd11an1n04x5 FILLER_298_2068 ();
 b15zdnd11an1n04x5 FILLER_298_2078 ();
 b15zdnd11an1n16x5 FILLER_298_2102 ();
 b15zdnd11an1n08x5 FILLER_298_2118 ();
 b15zdnd11an1n04x5 FILLER_298_2126 ();
 b15zdnd00an1n02x5 FILLER_298_2130 ();
 b15zdnd11an1n04x5 FILLER_298_2138 ();
 b15zdnd00an1n02x5 FILLER_298_2152 ();
 b15zdnd11an1n32x5 FILLER_298_2162 ();
 b15zdnd11an1n08x5 FILLER_298_2194 ();
 b15zdnd11an1n64x5 FILLER_298_2210 ();
 b15zdnd00an1n02x5 FILLER_298_2274 ();
 b15zdnd11an1n64x5 FILLER_299_0 ();
 b15zdnd11an1n08x5 FILLER_299_64 ();
 b15zdnd11an1n04x5 FILLER_299_90 ();
 b15zdnd11an1n04x5 FILLER_299_112 ();
 b15zdnd00an1n02x5 FILLER_299_116 ();
 b15zdnd11an1n16x5 FILLER_299_130 ();
 b15zdnd11an1n08x5 FILLER_299_146 ();
 b15zdnd11an1n04x5 FILLER_299_166 ();
 b15zdnd11an1n04x5 FILLER_299_186 ();
 b15zdnd11an1n08x5 FILLER_299_195 ();
 b15zdnd00an1n02x5 FILLER_299_203 ();
 b15zdnd11an1n16x5 FILLER_299_221 ();
 b15zdnd11an1n04x5 FILLER_299_246 ();
 b15zdnd00an1n02x5 FILLER_299_250 ();
 b15zdnd11an1n04x5 FILLER_299_258 ();
 b15zdnd11an1n08x5 FILLER_299_269 ();
 b15zdnd00an1n02x5 FILLER_299_277 ();
 b15zdnd00an1n01x5 FILLER_299_279 ();
 b15zdnd11an1n16x5 FILLER_299_289 ();
 b15zdnd11an1n04x5 FILLER_299_312 ();
 b15zdnd11an1n64x5 FILLER_299_320 ();
 b15zdnd11an1n32x5 FILLER_299_384 ();
 b15zdnd11an1n08x5 FILLER_299_416 ();
 b15zdnd00an1n01x5 FILLER_299_424 ();
 b15zdnd11an1n08x5 FILLER_299_456 ();
 b15zdnd11an1n04x5 FILLER_299_464 ();
 b15zdnd00an1n02x5 FILLER_299_468 ();
 b15zdnd11an1n08x5 FILLER_299_478 ();
 b15zdnd00an1n01x5 FILLER_299_486 ();
 b15zdnd11an1n08x5 FILLER_299_505 ();
 b15zdnd11an1n04x5 FILLER_299_513 ();
 b15zdnd00an1n02x5 FILLER_299_517 ();
 b15zdnd00an1n01x5 FILLER_299_519 ();
 b15zdnd11an1n64x5 FILLER_299_532 ();
 b15zdnd00an1n01x5 FILLER_299_596 ();
 b15zdnd11an1n08x5 FILLER_299_604 ();
 b15zdnd00an1n02x5 FILLER_299_612 ();
 b15zdnd11an1n04x5 FILLER_299_620 ();
 b15zdnd11an1n04x5 FILLER_299_642 ();
 b15zdnd00an1n01x5 FILLER_299_646 ();
 b15zdnd11an1n32x5 FILLER_299_651 ();
 b15zdnd11an1n08x5 FILLER_299_683 ();
 b15zdnd11an1n04x5 FILLER_299_691 ();
 b15zdnd00an1n02x5 FILLER_299_695 ();
 b15zdnd00an1n01x5 FILLER_299_697 ();
 b15zdnd11an1n16x5 FILLER_299_705 ();
 b15zdnd11an1n04x5 FILLER_299_721 ();
 b15zdnd00an1n01x5 FILLER_299_725 ();
 b15zdnd11an1n64x5 FILLER_299_758 ();
 b15zdnd11an1n16x5 FILLER_299_822 ();
 b15zdnd11an1n04x5 FILLER_299_869 ();
 b15zdnd11an1n32x5 FILLER_299_898 ();
 b15zdnd11an1n16x5 FILLER_299_930 ();
 b15zdnd11an1n08x5 FILLER_299_946 ();
 b15zdnd11an1n04x5 FILLER_299_954 ();
 b15zdnd00an1n02x5 FILLER_299_958 ();
 b15zdnd11an1n64x5 FILLER_299_985 ();
 b15zdnd11an1n64x5 FILLER_299_1049 ();
 b15zdnd11an1n16x5 FILLER_299_1113 ();
 b15zdnd11an1n04x5 FILLER_299_1129 ();
 b15zdnd00an1n01x5 FILLER_299_1133 ();
 b15zdnd11an1n08x5 FILLER_299_1142 ();
 b15zdnd00an1n02x5 FILLER_299_1150 ();
 b15zdnd00an1n01x5 FILLER_299_1152 ();
 b15zdnd11an1n64x5 FILLER_299_1159 ();
 b15zdnd11an1n32x5 FILLER_299_1223 ();
 b15zdnd11an1n08x5 FILLER_299_1255 ();
 b15zdnd11an1n04x5 FILLER_299_1263 ();
 b15zdnd00an1n01x5 FILLER_299_1267 ();
 b15zdnd11an1n08x5 FILLER_299_1278 ();
 b15zdnd00an1n01x5 FILLER_299_1286 ();
 b15zdnd11an1n04x5 FILLER_299_1290 ();
 b15zdnd11an1n04x5 FILLER_299_1305 ();
 b15zdnd11an1n64x5 FILLER_299_1325 ();
 b15zdnd11an1n32x5 FILLER_299_1389 ();
 b15zdnd11an1n04x5 FILLER_299_1421 ();
 b15zdnd00an1n02x5 FILLER_299_1425 ();
 b15zdnd00an1n01x5 FILLER_299_1427 ();
 b15zdnd11an1n04x5 FILLER_299_1433 ();
 b15zdnd11an1n16x5 FILLER_299_1446 ();
 b15zdnd11an1n08x5 FILLER_299_1462 ();
 b15zdnd00an1n02x5 FILLER_299_1470 ();
 b15zdnd11an1n16x5 FILLER_299_1484 ();
 b15zdnd11an1n08x5 FILLER_299_1500 ();
 b15zdnd11an1n04x5 FILLER_299_1508 ();
 b15zdnd11an1n08x5 FILLER_299_1524 ();
 b15zdnd11an1n04x5 FILLER_299_1532 ();
 b15zdnd11an1n04x5 FILLER_299_1552 ();
 b15zdnd11an1n64x5 FILLER_299_1565 ();
 b15zdnd11an1n16x5 FILLER_299_1629 ();
 b15zdnd00an1n02x5 FILLER_299_1645 ();
 b15zdnd00an1n01x5 FILLER_299_1647 ();
 b15zdnd11an1n04x5 FILLER_299_1652 ();
 b15zdnd11an1n64x5 FILLER_299_1662 ();
 b15zdnd11an1n64x5 FILLER_299_1726 ();
 b15zdnd11an1n32x5 FILLER_299_1790 ();
 b15zdnd00an1n01x5 FILLER_299_1822 ();
 b15zdnd11an1n64x5 FILLER_299_1830 ();
 b15zdnd11an1n08x5 FILLER_299_1894 ();
 b15zdnd00an1n02x5 FILLER_299_1902 ();
 b15zdnd11an1n32x5 FILLER_299_1924 ();
 b15zdnd11an1n08x5 FILLER_299_1956 ();
 b15zdnd00an1n02x5 FILLER_299_1964 ();
 b15zdnd00an1n01x5 FILLER_299_1966 ();
 b15zdnd11an1n04x5 FILLER_299_1975 ();
 b15zdnd11an1n32x5 FILLER_299_2005 ();
 b15zdnd00an1n01x5 FILLER_299_2037 ();
 b15zdnd11an1n16x5 FILLER_299_2044 ();
 b15zdnd11an1n08x5 FILLER_299_2060 ();
 b15zdnd11an1n04x5 FILLER_299_2068 ();
 b15zdnd11an1n04x5 FILLER_299_2092 ();
 b15zdnd00an1n02x5 FILLER_299_2096 ();
 b15zdnd11an1n04x5 FILLER_299_2103 ();
 b15zdnd00an1n01x5 FILLER_299_2107 ();
 b15zdnd11an1n04x5 FILLER_299_2124 ();
 b15zdnd11an1n04x5 FILLER_299_2137 ();
 b15zdnd11an1n32x5 FILLER_299_2150 ();
 b15zdnd11an1n08x5 FILLER_299_2182 ();
 b15zdnd11an1n04x5 FILLER_299_2190 ();
 b15zdnd00an1n02x5 FILLER_299_2194 ();
 b15zdnd00an1n01x5 FILLER_299_2196 ();
 b15zdnd11an1n08x5 FILLER_299_2213 ();
 b15zdnd11an1n04x5 FILLER_299_2221 ();
 b15zdnd11an1n32x5 FILLER_299_2239 ();
 b15zdnd11an1n08x5 FILLER_299_2271 ();
 b15zdnd11an1n04x5 FILLER_299_2279 ();
 b15zdnd00an1n01x5 FILLER_299_2283 ();
 b15zdnd11an1n64x5 FILLER_300_8 ();
 b15zdnd11an1n64x5 FILLER_300_72 ();
 b15zdnd11an1n64x5 FILLER_300_136 ();
 b15zdnd11an1n64x5 FILLER_300_200 ();
 b15zdnd11an1n64x5 FILLER_300_264 ();
 b15zdnd11an1n64x5 FILLER_300_328 ();
 b15zdnd11an1n64x5 FILLER_300_392 ();
 b15zdnd11an1n16x5 FILLER_300_456 ();
 b15zdnd11an1n08x5 FILLER_300_472 ();
 b15zdnd11an1n04x5 FILLER_300_480 ();
 b15zdnd11an1n08x5 FILLER_300_510 ();
 b15zdnd11an1n04x5 FILLER_300_518 ();
 b15zdnd00an1n01x5 FILLER_300_522 ();
 b15zdnd11an1n04x5 FILLER_300_529 ();
 b15zdnd11an1n64x5 FILLER_300_542 ();
 b15zdnd00an1n02x5 FILLER_300_606 ();
 b15zdnd00an1n01x5 FILLER_300_608 ();
 b15zdnd11an1n64x5 FILLER_300_618 ();
 b15zdnd00an1n02x5 FILLER_300_682 ();
 b15zdnd11an1n04x5 FILLER_300_690 ();
 b15zdnd11an1n04x5 FILLER_300_714 ();
 b15zdnd11an1n08x5 FILLER_300_726 ();
 b15zdnd00an1n02x5 FILLER_300_734 ();
 b15zdnd00an1n01x5 FILLER_300_736 ();
 b15zdnd11an1n32x5 FILLER_300_769 ();
 b15zdnd00an1n02x5 FILLER_300_801 ();
 b15zdnd00an1n01x5 FILLER_300_803 ();
 b15zdnd11an1n64x5 FILLER_300_822 ();
 b15zdnd11an1n08x5 FILLER_300_886 ();
 b15zdnd00an1n01x5 FILLER_300_894 ();
 b15zdnd11an1n32x5 FILLER_300_898 ();
 b15zdnd00an1n02x5 FILLER_300_930 ();
 b15zdnd00an1n01x5 FILLER_300_932 ();
 b15zdnd11an1n04x5 FILLER_300_964 ();
 b15zdnd11an1n32x5 FILLER_300_988 ();
 b15zdnd00an1n02x5 FILLER_300_1020 ();
 b15zdnd00an1n01x5 FILLER_300_1022 ();
 b15zdnd11an1n32x5 FILLER_300_1033 ();
 b15zdnd11an1n16x5 FILLER_300_1065 ();
 b15zdnd11an1n04x5 FILLER_300_1081 ();
 b15zdnd00an1n02x5 FILLER_300_1085 ();
 b15zdnd00an1n01x5 FILLER_300_1087 ();
 b15zdnd11an1n16x5 FILLER_300_1106 ();
 b15zdnd00an1n01x5 FILLER_300_1122 ();
 b15zdnd11an1n04x5 FILLER_300_1149 ();
 b15zdnd00an1n02x5 FILLER_300_1153 ();
 b15zdnd11an1n08x5 FILLER_300_1162 ();
 b15zdnd00an1n02x5 FILLER_300_1170 ();
 b15zdnd11an1n04x5 FILLER_300_1188 ();
 b15zdnd11an1n32x5 FILLER_300_1198 ();
 b15zdnd11an1n16x5 FILLER_300_1230 ();
 b15zdnd11an1n08x5 FILLER_300_1246 ();
 b15zdnd00an1n02x5 FILLER_300_1254 ();
 b15zdnd11an1n32x5 FILLER_300_1267 ();
 b15zdnd11an1n04x5 FILLER_300_1311 ();
 b15zdnd11an1n04x5 FILLER_300_1329 ();
 b15zdnd00an1n02x5 FILLER_300_1333 ();
 b15zdnd11an1n08x5 FILLER_300_1358 ();
 b15zdnd00an1n01x5 FILLER_300_1366 ();
 b15zdnd11an1n64x5 FILLER_300_1381 ();
 b15zdnd11an1n16x5 FILLER_300_1445 ();
 b15zdnd11an1n08x5 FILLER_300_1461 ();
 b15zdnd11an1n04x5 FILLER_300_1469 ();
 b15zdnd00an1n02x5 FILLER_300_1473 ();
 b15zdnd00an1n01x5 FILLER_300_1475 ();
 b15zdnd11an1n32x5 FILLER_300_1482 ();
 b15zdnd11an1n04x5 FILLER_300_1514 ();
 b15zdnd00an1n02x5 FILLER_300_1518 ();
 b15zdnd11an1n04x5 FILLER_300_1525 ();
 b15zdnd00an1n02x5 FILLER_300_1529 ();
 b15zdnd00an1n01x5 FILLER_300_1531 ();
 b15zdnd11an1n08x5 FILLER_300_1544 ();
 b15zdnd11an1n04x5 FILLER_300_1552 ();
 b15zdnd00an1n02x5 FILLER_300_1556 ();
 b15zdnd00an1n01x5 FILLER_300_1558 ();
 b15zdnd11an1n16x5 FILLER_300_1565 ();
 b15zdnd11an1n04x5 FILLER_300_1581 ();
 b15zdnd00an1n02x5 FILLER_300_1585 ();
 b15zdnd11an1n32x5 FILLER_300_1594 ();
 b15zdnd11an1n16x5 FILLER_300_1626 ();
 b15zdnd00an1n02x5 FILLER_300_1642 ();
 b15zdnd00an1n01x5 FILLER_300_1644 ();
 b15zdnd11an1n32x5 FILLER_300_1659 ();
 b15zdnd11an1n16x5 FILLER_300_1691 ();
 b15zdnd11an1n04x5 FILLER_300_1707 ();
 b15zdnd00an1n01x5 FILLER_300_1711 ();
 b15zdnd11an1n16x5 FILLER_300_1722 ();
 b15zdnd00an1n02x5 FILLER_300_1738 ();
 b15zdnd11an1n08x5 FILLER_300_1748 ();
 b15zdnd00an1n01x5 FILLER_300_1756 ();
 b15zdnd11an1n08x5 FILLER_300_1763 ();
 b15zdnd11an1n04x5 FILLER_300_1771 ();
 b15zdnd00an1n02x5 FILLER_300_1775 ();
 b15zdnd11an1n08x5 FILLER_300_1781 ();
 b15zdnd11an1n04x5 FILLER_300_1789 ();
 b15zdnd11an1n08x5 FILLER_300_1811 ();
 b15zdnd11an1n04x5 FILLER_300_1819 ();
 b15zdnd00an1n02x5 FILLER_300_1823 ();
 b15zdnd11an1n32x5 FILLER_300_1834 ();
 b15zdnd11an1n16x5 FILLER_300_1866 ();
 b15zdnd00an1n01x5 FILLER_300_1882 ();
 b15zdnd11an1n04x5 FILLER_300_1897 ();
 b15zdnd11an1n04x5 FILLER_300_1927 ();
 b15zdnd11an1n16x5 FILLER_300_1944 ();
 b15zdnd00an1n02x5 FILLER_300_1960 ();
 b15zdnd11an1n16x5 FILLER_300_1969 ();
 b15zdnd00an1n02x5 FILLER_300_1985 ();
 b15zdnd11an1n32x5 FILLER_300_1997 ();
 b15zdnd11an1n08x5 FILLER_300_2029 ();
 b15zdnd00an1n02x5 FILLER_300_2037 ();
 b15zdnd00an1n01x5 FILLER_300_2039 ();
 b15zdnd11an1n08x5 FILLER_300_2058 ();
 b15zdnd11an1n04x5 FILLER_300_2066 ();
 b15zdnd00an1n02x5 FILLER_300_2070 ();
 b15zdnd11an1n32x5 FILLER_300_2092 ();
 b15zdnd00an1n02x5 FILLER_300_2124 ();
 b15zdnd00an1n01x5 FILLER_300_2126 ();
 b15zdnd11an1n16x5 FILLER_300_2131 ();
 b15zdnd11an1n04x5 FILLER_300_2147 ();
 b15zdnd00an1n02x5 FILLER_300_2151 ();
 b15zdnd00an1n01x5 FILLER_300_2153 ();
 b15zdnd11an1n08x5 FILLER_300_2162 ();
 b15zdnd00an1n02x5 FILLER_300_2170 ();
 b15zdnd11an1n32x5 FILLER_300_2177 ();
 b15zdnd11an1n16x5 FILLER_300_2209 ();
 b15zdnd11an1n08x5 FILLER_300_2225 ();
 b15zdnd00an1n01x5 FILLER_300_2233 ();
 b15zdnd11an1n16x5 FILLER_300_2252 ();
 b15zdnd11an1n08x5 FILLER_300_2268 ();
 b15zdnd11an1n64x5 FILLER_301_0 ();
 b15zdnd11an1n64x5 FILLER_301_64 ();
 b15zdnd11an1n64x5 FILLER_301_128 ();
 b15zdnd11an1n64x5 FILLER_301_192 ();
 b15zdnd11an1n64x5 FILLER_301_256 ();
 b15zdnd11an1n64x5 FILLER_301_320 ();
 b15zdnd11an1n64x5 FILLER_301_384 ();
 b15zdnd11an1n04x5 FILLER_301_448 ();
 b15zdnd00an1n02x5 FILLER_301_452 ();
 b15zdnd11an1n16x5 FILLER_301_470 ();
 b15zdnd11an1n08x5 FILLER_301_486 ();
 b15zdnd11an1n04x5 FILLER_301_494 ();
 b15zdnd11an1n08x5 FILLER_301_510 ();
 b15zdnd00an1n02x5 FILLER_301_518 ();
 b15zdnd11an1n16x5 FILLER_301_531 ();
 b15zdnd11an1n16x5 FILLER_301_571 ();
 b15zdnd11an1n08x5 FILLER_301_596 ();
 b15zdnd11an1n04x5 FILLER_301_604 ();
 b15zdnd11an1n04x5 FILLER_301_614 ();
 b15zdnd11an1n32x5 FILLER_301_622 ();
 b15zdnd11an1n04x5 FILLER_301_654 ();
 b15zdnd00an1n02x5 FILLER_301_658 ();
 b15zdnd00an1n01x5 FILLER_301_660 ();
 b15zdnd11an1n16x5 FILLER_301_670 ();
 b15zdnd11an1n08x5 FILLER_301_686 ();
 b15zdnd00an1n01x5 FILLER_301_694 ();
 b15zdnd11an1n04x5 FILLER_301_699 ();
 b15zdnd11an1n08x5 FILLER_301_717 ();
 b15zdnd11an1n32x5 FILLER_301_741 ();
 b15zdnd11an1n04x5 FILLER_301_773 ();
 b15zdnd00an1n02x5 FILLER_301_777 ();
 b15zdnd11an1n04x5 FILLER_301_793 ();
 b15zdnd11an1n08x5 FILLER_301_809 ();
 b15zdnd11an1n32x5 FILLER_301_832 ();
 b15zdnd11an1n16x5 FILLER_301_864 ();
 b15zdnd11an1n08x5 FILLER_301_880 ();
 b15zdnd00an1n01x5 FILLER_301_888 ();
 b15zdnd11an1n16x5 FILLER_301_909 ();
 b15zdnd00an1n02x5 FILLER_301_925 ();
 b15zdnd11an1n32x5 FILLER_301_942 ();
 b15zdnd11an1n16x5 FILLER_301_974 ();
 b15zdnd11an1n08x5 FILLER_301_990 ();
 b15zdnd11an1n04x5 FILLER_301_998 ();
 b15zdnd00an1n02x5 FILLER_301_1002 ();
 b15zdnd00an1n01x5 FILLER_301_1004 ();
 b15zdnd11an1n16x5 FILLER_301_1021 ();
 b15zdnd11an1n08x5 FILLER_301_1037 ();
 b15zdnd00an1n01x5 FILLER_301_1045 ();
 b15zdnd11an1n32x5 FILLER_301_1052 ();
 b15zdnd11an1n08x5 FILLER_301_1084 ();
 b15zdnd11an1n04x5 FILLER_301_1092 ();
 b15zdnd00an1n01x5 FILLER_301_1096 ();
 b15zdnd11an1n04x5 FILLER_301_1103 ();
 b15zdnd11an1n04x5 FILLER_301_1115 ();
 b15zdnd11an1n08x5 FILLER_301_1126 ();
 b15zdnd11an1n04x5 FILLER_301_1134 ();
 b15zdnd11an1n32x5 FILLER_301_1144 ();
 b15zdnd11an1n16x5 FILLER_301_1176 ();
 b15zdnd11an1n04x5 FILLER_301_1197 ();
 b15zdnd00an1n02x5 FILLER_301_1201 ();
 b15zdnd11an1n16x5 FILLER_301_1209 ();
 b15zdnd11an1n04x5 FILLER_301_1229 ();
 b15zdnd11an1n16x5 FILLER_301_1239 ();
 b15zdnd11an1n08x5 FILLER_301_1263 ();
 b15zdnd00an1n02x5 FILLER_301_1271 ();
 b15zdnd11an1n04x5 FILLER_301_1296 ();
 b15zdnd11an1n64x5 FILLER_301_1326 ();
 b15zdnd11an1n64x5 FILLER_301_1390 ();
 b15zdnd11an1n32x5 FILLER_301_1454 ();
 b15zdnd11an1n04x5 FILLER_301_1486 ();
 b15zdnd00an1n02x5 FILLER_301_1490 ();
 b15zdnd00an1n01x5 FILLER_301_1492 ();
 b15zdnd11an1n64x5 FILLER_301_1509 ();
 b15zdnd11an1n08x5 FILLER_301_1573 ();
 b15zdnd11an1n04x5 FILLER_301_1581 ();
 b15zdnd00an1n02x5 FILLER_301_1585 ();
 b15zdnd11an1n32x5 FILLER_301_1595 ();
 b15zdnd11an1n16x5 FILLER_301_1627 ();
 b15zdnd11an1n08x5 FILLER_301_1643 ();
 b15zdnd11an1n04x5 FILLER_301_1651 ();
 b15zdnd00an1n02x5 FILLER_301_1655 ();
 b15zdnd11an1n04x5 FILLER_301_1666 ();
 b15zdnd00an1n02x5 FILLER_301_1670 ();
 b15zdnd11an1n04x5 FILLER_301_1688 ();
 b15zdnd11an1n08x5 FILLER_301_1700 ();
 b15zdnd00an1n02x5 FILLER_301_1708 ();
 b15zdnd11an1n16x5 FILLER_301_1730 ();
 b15zdnd11an1n08x5 FILLER_301_1746 ();
 b15zdnd00an1n02x5 FILLER_301_1754 ();
 b15zdnd00an1n01x5 FILLER_301_1756 ();
 b15zdnd11an1n08x5 FILLER_301_1763 ();
 b15zdnd11an1n04x5 FILLER_301_1771 ();
 b15zdnd11an1n64x5 FILLER_301_1786 ();
 b15zdnd11an1n32x5 FILLER_301_1850 ();
 b15zdnd11an1n16x5 FILLER_301_1882 ();
 b15zdnd00an1n02x5 FILLER_301_1898 ();
 b15zdnd00an1n01x5 FILLER_301_1900 ();
 b15zdnd11an1n32x5 FILLER_301_1927 ();
 b15zdnd11an1n64x5 FILLER_301_1985 ();
 b15zdnd11an1n32x5 FILLER_301_2049 ();
 b15zdnd11an1n08x5 FILLER_301_2081 ();
 b15zdnd11an1n04x5 FILLER_301_2089 ();
 b15zdnd11an1n32x5 FILLER_301_2105 ();
 b15zdnd11an1n16x5 FILLER_301_2137 ();
 b15zdnd11an1n04x5 FILLER_301_2153 ();
 b15zdnd00an1n01x5 FILLER_301_2157 ();
 b15zdnd11an1n08x5 FILLER_301_2164 ();
 b15zdnd11an1n64x5 FILLER_301_2177 ();
 b15zdnd11an1n32x5 FILLER_301_2241 ();
 b15zdnd11an1n08x5 FILLER_301_2273 ();
 b15zdnd00an1n02x5 FILLER_301_2281 ();
 b15zdnd00an1n01x5 FILLER_301_2283 ();
 b15zdnd11an1n64x5 FILLER_302_8 ();
 b15zdnd11an1n64x5 FILLER_302_72 ();
 b15zdnd11an1n64x5 FILLER_302_136 ();
 b15zdnd11an1n64x5 FILLER_302_200 ();
 b15zdnd11an1n64x5 FILLER_302_264 ();
 b15zdnd11an1n64x5 FILLER_302_328 ();
 b15zdnd11an1n64x5 FILLER_302_392 ();
 b15zdnd11an1n64x5 FILLER_302_456 ();
 b15zdnd11an1n04x5 FILLER_302_520 ();
 b15zdnd00an1n02x5 FILLER_302_524 ();
 b15zdnd00an1n01x5 FILLER_302_526 ();
 b15zdnd11an1n08x5 FILLER_302_536 ();
 b15zdnd11an1n04x5 FILLER_302_544 ();
 b15zdnd00an1n02x5 FILLER_302_548 ();
 b15zdnd11an1n64x5 FILLER_302_554 ();
 b15zdnd11an1n64x5 FILLER_302_618 ();
 b15zdnd11an1n32x5 FILLER_302_682 ();
 b15zdnd11an1n04x5 FILLER_302_714 ();
 b15zdnd11an1n64x5 FILLER_302_726 ();
 b15zdnd11an1n16x5 FILLER_302_790 ();
 b15zdnd00an1n01x5 FILLER_302_806 ();
 b15zdnd11an1n32x5 FILLER_302_822 ();
 b15zdnd11an1n08x5 FILLER_302_854 ();
 b15zdnd11an1n04x5 FILLER_302_862 ();
 b15zdnd00an1n01x5 FILLER_302_866 ();
 b15zdnd11an1n04x5 FILLER_302_892 ();
 b15zdnd11an1n64x5 FILLER_302_901 ();
 b15zdnd11an1n64x5 FILLER_302_965 ();
 b15zdnd11an1n16x5 FILLER_302_1029 ();
 b15zdnd00an1n02x5 FILLER_302_1045 ();
 b15zdnd00an1n01x5 FILLER_302_1047 ();
 b15zdnd11an1n08x5 FILLER_302_1055 ();
 b15zdnd00an1n02x5 FILLER_302_1063 ();
 b15zdnd11an1n32x5 FILLER_302_1069 ();
 b15zdnd11an1n16x5 FILLER_302_1101 ();
 b15zdnd11an1n08x5 FILLER_302_1117 ();
 b15zdnd00an1n02x5 FILLER_302_1125 ();
 b15zdnd11an1n32x5 FILLER_302_1139 ();
 b15zdnd11an1n16x5 FILLER_302_1171 ();
 b15zdnd11an1n08x5 FILLER_302_1187 ();
 b15zdnd00an1n02x5 FILLER_302_1195 ();
 b15zdnd00an1n01x5 FILLER_302_1197 ();
 b15zdnd11an1n08x5 FILLER_302_1211 ();
 b15zdnd11an1n04x5 FILLER_302_1219 ();
 b15zdnd11an1n04x5 FILLER_302_1228 ();
 b15zdnd11an1n04x5 FILLER_302_1236 ();
 b15zdnd00an1n02x5 FILLER_302_1240 ();
 b15zdnd11an1n32x5 FILLER_302_1246 ();
 b15zdnd11an1n08x5 FILLER_302_1278 ();
 b15zdnd11an1n16x5 FILLER_302_1298 ();
 b15zdnd11an1n08x5 FILLER_302_1314 ();
 b15zdnd00an1n02x5 FILLER_302_1322 ();
 b15zdnd11an1n04x5 FILLER_302_1337 ();
 b15zdnd11an1n32x5 FILLER_302_1362 ();
 b15zdnd11an1n04x5 FILLER_302_1394 ();
 b15zdnd11an1n04x5 FILLER_302_1418 ();
 b15zdnd11an1n32x5 FILLER_302_1454 ();
 b15zdnd11an1n04x5 FILLER_302_1486 ();
 b15zdnd00an1n01x5 FILLER_302_1490 ();
 b15zdnd11an1n04x5 FILLER_302_1498 ();
 b15zdnd11an1n64x5 FILLER_302_1508 ();
 b15zdnd11an1n32x5 FILLER_302_1572 ();
 b15zdnd11an1n16x5 FILLER_302_1604 ();
 b15zdnd00an1n02x5 FILLER_302_1620 ();
 b15zdnd00an1n01x5 FILLER_302_1622 ();
 b15zdnd11an1n08x5 FILLER_302_1628 ();
 b15zdnd00an1n01x5 FILLER_302_1636 ();
 b15zdnd11an1n16x5 FILLER_302_1642 ();
 b15zdnd11an1n04x5 FILLER_302_1658 ();
 b15zdnd00an1n01x5 FILLER_302_1662 ();
 b15zdnd11an1n04x5 FILLER_302_1679 ();
 b15zdnd11an1n04x5 FILLER_302_1703 ();
 b15zdnd11an1n64x5 FILLER_302_1717 ();
 b15zdnd11an1n64x5 FILLER_302_1781 ();
 b15zdnd11an1n08x5 FILLER_302_1845 ();
 b15zdnd11an1n04x5 FILLER_302_1853 ();
 b15zdnd00an1n02x5 FILLER_302_1857 ();
 b15zdnd00an1n01x5 FILLER_302_1859 ();
 b15zdnd11an1n16x5 FILLER_302_1886 ();
 b15zdnd00an1n02x5 FILLER_302_1902 ();
 b15zdnd00an1n01x5 FILLER_302_1904 ();
 b15zdnd11an1n04x5 FILLER_302_1921 ();
 b15zdnd11an1n64x5 FILLER_302_1941 ();
 b15zdnd11an1n64x5 FILLER_302_2005 ();
 b15zdnd11an1n16x5 FILLER_302_2069 ();
 b15zdnd00an1n01x5 FILLER_302_2085 ();
 b15zdnd11an1n16x5 FILLER_302_2112 ();
 b15zdnd00an1n01x5 FILLER_302_2128 ();
 b15zdnd11an1n08x5 FILLER_302_2145 ();
 b15zdnd00an1n01x5 FILLER_302_2153 ();
 b15zdnd00an1n02x5 FILLER_302_2162 ();
 b15zdnd11an1n04x5 FILLER_302_2176 ();
 b15zdnd11an1n64x5 FILLER_302_2196 ();
 b15zdnd11an1n16x5 FILLER_302_2260 ();
 b15zdnd11an1n64x5 FILLER_303_0 ();
 b15zdnd11an1n64x5 FILLER_303_64 ();
 b15zdnd11an1n64x5 FILLER_303_128 ();
 b15zdnd11an1n64x5 FILLER_303_192 ();
 b15zdnd11an1n64x5 FILLER_303_256 ();
 b15zdnd11an1n64x5 FILLER_303_320 ();
 b15zdnd11an1n64x5 FILLER_303_384 ();
 b15zdnd11an1n64x5 FILLER_303_448 ();
 b15zdnd11an1n32x5 FILLER_303_512 ();
 b15zdnd11an1n04x5 FILLER_303_544 ();
 b15zdnd00an1n01x5 FILLER_303_548 ();
 b15zdnd11an1n64x5 FILLER_303_555 ();
 b15zdnd11an1n64x5 FILLER_303_619 ();
 b15zdnd11an1n16x5 FILLER_303_683 ();
 b15zdnd11an1n08x5 FILLER_303_699 ();
 b15zdnd00an1n02x5 FILLER_303_707 ();
 b15zdnd11an1n32x5 FILLER_303_727 ();
 b15zdnd11an1n16x5 FILLER_303_759 ();
 b15zdnd11an1n32x5 FILLER_303_807 ();
 b15zdnd11an1n16x5 FILLER_303_839 ();
 b15zdnd11an1n04x5 FILLER_303_855 ();
 b15zdnd00an1n02x5 FILLER_303_859 ();
 b15zdnd11an1n32x5 FILLER_303_892 ();
 b15zdnd11an1n04x5 FILLER_303_924 ();
 b15zdnd00an1n01x5 FILLER_303_928 ();
 b15zdnd11an1n64x5 FILLER_303_933 ();
 b15zdnd11an1n32x5 FILLER_303_997 ();
 b15zdnd11an1n16x5 FILLER_303_1029 ();
 b15zdnd00an1n02x5 FILLER_303_1045 ();
 b15zdnd11an1n08x5 FILLER_303_1052 ();
 b15zdnd11an1n04x5 FILLER_303_1060 ();
 b15zdnd11an1n64x5 FILLER_303_1078 ();
 b15zdnd11an1n64x5 FILLER_303_1142 ();
 b15zdnd11an1n64x5 FILLER_303_1206 ();
 b15zdnd11an1n32x5 FILLER_303_1270 ();
 b15zdnd11an1n04x5 FILLER_303_1302 ();
 b15zdnd00an1n01x5 FILLER_303_1306 ();
 b15zdnd11an1n08x5 FILLER_303_1321 ();
 b15zdnd00an1n02x5 FILLER_303_1329 ();
 b15zdnd00an1n01x5 FILLER_303_1331 ();
 b15zdnd11an1n64x5 FILLER_303_1358 ();
 b15zdnd11an1n16x5 FILLER_303_1422 ();
 b15zdnd11an1n08x5 FILLER_303_1438 ();
 b15zdnd11an1n16x5 FILLER_303_1462 ();
 b15zdnd11an1n08x5 FILLER_303_1478 ();
 b15zdnd11an1n16x5 FILLER_303_1494 ();
 b15zdnd11an1n08x5 FILLER_303_1510 ();
 b15zdnd11an1n04x5 FILLER_303_1518 ();
 b15zdnd00an1n02x5 FILLER_303_1522 ();
 b15zdnd11an1n16x5 FILLER_303_1530 ();
 b15zdnd11an1n08x5 FILLER_303_1546 ();
 b15zdnd11an1n04x5 FILLER_303_1554 ();
 b15zdnd11an1n08x5 FILLER_303_1564 ();
 b15zdnd11an1n32x5 FILLER_303_1576 ();
 b15zdnd00an1n02x5 FILLER_303_1608 ();
 b15zdnd11an1n16x5 FILLER_303_1615 ();
 b15zdnd00an1n02x5 FILLER_303_1631 ();
 b15zdnd00an1n01x5 FILLER_303_1633 ();
 b15zdnd11an1n08x5 FILLER_303_1638 ();
 b15zdnd00an1n02x5 FILLER_303_1646 ();
 b15zdnd11an1n04x5 FILLER_303_1661 ();
 b15zdnd11an1n16x5 FILLER_303_1680 ();
 b15zdnd11an1n04x5 FILLER_303_1696 ();
 b15zdnd11an1n64x5 FILLER_303_1710 ();
 b15zdnd00an1n02x5 FILLER_303_1774 ();
 b15zdnd11an1n32x5 FILLER_303_1799 ();
 b15zdnd11an1n32x5 FILLER_303_1841 ();
 b15zdnd11an1n08x5 FILLER_303_1873 ();
 b15zdnd11an1n04x5 FILLER_303_1881 ();
 b15zdnd00an1n02x5 FILLER_303_1885 ();
 b15zdnd11an1n08x5 FILLER_303_1910 ();
 b15zdnd11an1n04x5 FILLER_303_1918 ();
 b15zdnd00an1n02x5 FILLER_303_1922 ();
 b15zdnd00an1n01x5 FILLER_303_1924 ();
 b15zdnd11an1n32x5 FILLER_303_1938 ();
 b15zdnd11an1n04x5 FILLER_303_1970 ();
 b15zdnd11an1n04x5 FILLER_303_1984 ();
 b15zdnd00an1n01x5 FILLER_303_1988 ();
 b15zdnd11an1n08x5 FILLER_303_1993 ();
 b15zdnd00an1n01x5 FILLER_303_2001 ();
 b15zdnd11an1n08x5 FILLER_303_2009 ();
 b15zdnd00an1n01x5 FILLER_303_2017 ();
 b15zdnd11an1n08x5 FILLER_303_2024 ();
 b15zdnd11an1n04x5 FILLER_303_2032 ();
 b15zdnd00an1n01x5 FILLER_303_2036 ();
 b15zdnd11an1n16x5 FILLER_303_2050 ();
 b15zdnd00an1n01x5 FILLER_303_2066 ();
 b15zdnd11an1n04x5 FILLER_303_2071 ();
 b15zdnd00an1n02x5 FILLER_303_2075 ();
 b15zdnd00an1n01x5 FILLER_303_2077 ();
 b15zdnd11an1n08x5 FILLER_303_2083 ();
 b15zdnd11an1n04x5 FILLER_303_2091 ();
 b15zdnd00an1n01x5 FILLER_303_2095 ();
 b15zdnd11an1n04x5 FILLER_303_2104 ();
 b15zdnd11an1n08x5 FILLER_303_2112 ();
 b15zdnd00an1n01x5 FILLER_303_2120 ();
 b15zdnd11an1n08x5 FILLER_303_2141 ();
 b15zdnd11an1n04x5 FILLER_303_2149 ();
 b15zdnd00an1n01x5 FILLER_303_2153 ();
 b15zdnd11an1n04x5 FILLER_303_2170 ();
 b15zdnd11an1n16x5 FILLER_303_2181 ();
 b15zdnd11an1n08x5 FILLER_303_2197 ();
 b15zdnd00an1n02x5 FILLER_303_2205 ();
 b15zdnd00an1n01x5 FILLER_303_2207 ();
 b15zdnd11an1n16x5 FILLER_303_2217 ();
 b15zdnd11an1n04x5 FILLER_303_2233 ();
 b15zdnd11an1n32x5 FILLER_303_2251 ();
 b15zdnd00an1n01x5 FILLER_303_2283 ();
 b15zdnd11an1n64x5 FILLER_304_8 ();
 b15zdnd11an1n64x5 FILLER_304_72 ();
 b15zdnd11an1n64x5 FILLER_304_136 ();
 b15zdnd11an1n64x5 FILLER_304_200 ();
 b15zdnd11an1n64x5 FILLER_304_264 ();
 b15zdnd11an1n64x5 FILLER_304_328 ();
 b15zdnd11an1n08x5 FILLER_304_392 ();
 b15zdnd00an1n01x5 FILLER_304_400 ();
 b15zdnd11an1n04x5 FILLER_304_408 ();
 b15zdnd11an1n64x5 FILLER_304_418 ();
 b15zdnd11an1n32x5 FILLER_304_482 ();
 b15zdnd00an1n02x5 FILLER_304_514 ();
 b15zdnd00an1n01x5 FILLER_304_516 ();
 b15zdnd11an1n08x5 FILLER_304_535 ();
 b15zdnd00an1n02x5 FILLER_304_543 ();
 b15zdnd00an1n01x5 FILLER_304_545 ();
 b15zdnd11an1n32x5 FILLER_304_554 ();
 b15zdnd11an1n04x5 FILLER_304_586 ();
 b15zdnd00an1n02x5 FILLER_304_590 ();
 b15zdnd11an1n08x5 FILLER_304_602 ();
 b15zdnd00an1n01x5 FILLER_304_610 ();
 b15zdnd11an1n16x5 FILLER_304_616 ();
 b15zdnd00an1n02x5 FILLER_304_632 ();
 b15zdnd00an1n01x5 FILLER_304_634 ();
 b15zdnd11an1n08x5 FILLER_304_644 ();
 b15zdnd11an1n04x5 FILLER_304_657 ();
 b15zdnd11an1n32x5 FILLER_304_667 ();
 b15zdnd11an1n16x5 FILLER_304_699 ();
 b15zdnd00an1n02x5 FILLER_304_715 ();
 b15zdnd00an1n01x5 FILLER_304_717 ();
 b15zdnd11an1n64x5 FILLER_304_726 ();
 b15zdnd11an1n32x5 FILLER_304_790 ();
 b15zdnd11an1n16x5 FILLER_304_822 ();
 b15zdnd11an1n08x5 FILLER_304_838 ();
 b15zdnd11an1n04x5 FILLER_304_846 ();
 b15zdnd11an1n32x5 FILLER_304_868 ();
 b15zdnd11an1n08x5 FILLER_304_900 ();
 b15zdnd11an1n04x5 FILLER_304_908 ();
 b15zdnd11an1n04x5 FILLER_304_919 ();
 b15zdnd00an1n02x5 FILLER_304_923 ();
 b15zdnd11an1n04x5 FILLER_304_956 ();
 b15zdnd11an1n16x5 FILLER_304_984 ();
 b15zdnd11an1n08x5 FILLER_304_1000 ();
 b15zdnd00an1n01x5 FILLER_304_1008 ();
 b15zdnd11an1n08x5 FILLER_304_1032 ();
 b15zdnd11an1n04x5 FILLER_304_1040 ();
 b15zdnd00an1n02x5 FILLER_304_1044 ();
 b15zdnd00an1n01x5 FILLER_304_1046 ();
 b15zdnd11an1n16x5 FILLER_304_1054 ();
 b15zdnd11an1n08x5 FILLER_304_1070 ();
 b15zdnd11an1n04x5 FILLER_304_1078 ();
 b15zdnd00an1n01x5 FILLER_304_1082 ();
 b15zdnd11an1n32x5 FILLER_304_1091 ();
 b15zdnd11an1n04x5 FILLER_304_1123 ();
 b15zdnd00an1n01x5 FILLER_304_1127 ();
 b15zdnd11an1n08x5 FILLER_304_1147 ();
 b15zdnd11an1n04x5 FILLER_304_1155 ();
 b15zdnd00an1n02x5 FILLER_304_1159 ();
 b15zdnd00an1n01x5 FILLER_304_1161 ();
 b15zdnd11an1n04x5 FILLER_304_1168 ();
 b15zdnd00an1n02x5 FILLER_304_1172 ();
 b15zdnd00an1n01x5 FILLER_304_1174 ();
 b15zdnd11an1n64x5 FILLER_304_1181 ();
 b15zdnd11an1n16x5 FILLER_304_1245 ();
 b15zdnd11an1n08x5 FILLER_304_1261 ();
 b15zdnd00an1n02x5 FILLER_304_1269 ();
 b15zdnd00an1n01x5 FILLER_304_1271 ();
 b15zdnd11an1n16x5 FILLER_304_1284 ();
 b15zdnd11an1n08x5 FILLER_304_1300 ();
 b15zdnd11an1n64x5 FILLER_304_1324 ();
 b15zdnd11an1n08x5 FILLER_304_1388 ();
 b15zdnd11an1n04x5 FILLER_304_1396 ();
 b15zdnd00an1n02x5 FILLER_304_1400 ();
 b15zdnd00an1n01x5 FILLER_304_1402 ();
 b15zdnd11an1n16x5 FILLER_304_1407 ();
 b15zdnd11an1n04x5 FILLER_304_1423 ();
 b15zdnd00an1n02x5 FILLER_304_1427 ();
 b15zdnd00an1n01x5 FILLER_304_1429 ();
 b15zdnd11an1n32x5 FILLER_304_1448 ();
 b15zdnd11an1n04x5 FILLER_304_1480 ();
 b15zdnd11an1n16x5 FILLER_304_1504 ();
 b15zdnd11an1n04x5 FILLER_304_1520 ();
 b15zdnd11an1n08x5 FILLER_304_1534 ();
 b15zdnd00an1n01x5 FILLER_304_1542 ();
 b15zdnd11an1n04x5 FILLER_304_1560 ();
 b15zdnd11an1n04x5 FILLER_304_1570 ();
 b15zdnd11an1n64x5 FILLER_304_1581 ();
 b15zdnd11an1n32x5 FILLER_304_1645 ();
 b15zdnd11an1n08x5 FILLER_304_1677 ();
 b15zdnd11an1n04x5 FILLER_304_1685 ();
 b15zdnd00an1n01x5 FILLER_304_1689 ();
 b15zdnd11an1n04x5 FILLER_304_1716 ();
 b15zdnd11an1n04x5 FILLER_304_1741 ();
 b15zdnd11an1n04x5 FILLER_304_1751 ();
 b15zdnd11an1n32x5 FILLER_304_1770 ();
 b15zdnd11an1n16x5 FILLER_304_1802 ();
 b15zdnd00an1n01x5 FILLER_304_1818 ();
 b15zdnd11an1n04x5 FILLER_304_1826 ();
 b15zdnd00an1n02x5 FILLER_304_1830 ();
 b15zdnd00an1n01x5 FILLER_304_1832 ();
 b15zdnd11an1n32x5 FILLER_304_1842 ();
 b15zdnd11an1n16x5 FILLER_304_1874 ();
 b15zdnd11an1n08x5 FILLER_304_1890 ();
 b15zdnd11an1n04x5 FILLER_304_1916 ();
 b15zdnd11an1n04x5 FILLER_304_1929 ();
 b15zdnd11an1n32x5 FILLER_304_1945 ();
 b15zdnd11an1n08x5 FILLER_304_1977 ();
 b15zdnd11an1n04x5 FILLER_304_1985 ();
 b15zdnd00an1n02x5 FILLER_304_1989 ();
 b15zdnd11an1n04x5 FILLER_304_1997 ();
 b15zdnd11an1n04x5 FILLER_304_2009 ();
 b15zdnd00an1n02x5 FILLER_304_2013 ();
 b15zdnd11an1n08x5 FILLER_304_2025 ();
 b15zdnd00an1n02x5 FILLER_304_2033 ();
 b15zdnd00an1n01x5 FILLER_304_2035 ();
 b15zdnd11an1n16x5 FILLER_304_2056 ();
 b15zdnd11an1n08x5 FILLER_304_2072 ();
 b15zdnd11an1n04x5 FILLER_304_2080 ();
 b15zdnd11an1n04x5 FILLER_304_2088 ();
 b15zdnd11an1n16x5 FILLER_304_2100 ();
 b15zdnd11an1n08x5 FILLER_304_2116 ();
 b15zdnd11an1n04x5 FILLER_304_2124 ();
 b15zdnd00an1n02x5 FILLER_304_2128 ();
 b15zdnd11an1n04x5 FILLER_304_2136 ();
 b15zdnd00an1n02x5 FILLER_304_2152 ();
 b15zdnd11an1n08x5 FILLER_304_2162 ();
 b15zdnd11an1n04x5 FILLER_304_2170 ();
 b15zdnd00an1n02x5 FILLER_304_2174 ();
 b15zdnd11an1n04x5 FILLER_304_2197 ();
 b15zdnd11an1n16x5 FILLER_304_2207 ();
 b15zdnd11an1n04x5 FILLER_304_2223 ();
 b15zdnd11an1n16x5 FILLER_304_2245 ();
 b15zdnd11an1n08x5 FILLER_304_2261 ();
 b15zdnd11an1n04x5 FILLER_304_2269 ();
 b15zdnd00an1n02x5 FILLER_304_2273 ();
 b15zdnd00an1n01x5 FILLER_304_2275 ();
 b15zdnd11an1n64x5 FILLER_305_0 ();
 b15zdnd11an1n64x5 FILLER_305_64 ();
 b15zdnd11an1n64x5 FILLER_305_128 ();
 b15zdnd11an1n64x5 FILLER_305_192 ();
 b15zdnd11an1n32x5 FILLER_305_256 ();
 b15zdnd11an1n16x5 FILLER_305_288 ();
 b15zdnd11an1n08x5 FILLER_305_304 ();
 b15zdnd00an1n02x5 FILLER_305_312 ();
 b15zdnd11an1n08x5 FILLER_305_320 ();
 b15zdnd00an1n02x5 FILLER_305_328 ();
 b15zdnd11an1n04x5 FILLER_305_337 ();
 b15zdnd11an1n04x5 FILLER_305_344 ();
 b15zdnd00an1n01x5 FILLER_305_348 ();
 b15zdnd11an1n16x5 FILLER_305_356 ();
 b15zdnd11an1n08x5 FILLER_305_372 ();
 b15zdnd00an1n02x5 FILLER_305_380 ();
 b15zdnd11an1n04x5 FILLER_305_393 ();
 b15zdnd00an1n02x5 FILLER_305_397 ();
 b15zdnd11an1n08x5 FILLER_305_403 ();
 b15zdnd00an1n02x5 FILLER_305_411 ();
 b15zdnd00an1n01x5 FILLER_305_413 ();
 b15zdnd11an1n08x5 FILLER_305_419 ();
 b15zdnd11an1n04x5 FILLER_305_427 ();
 b15zdnd00an1n02x5 FILLER_305_431 ();
 b15zdnd11an1n16x5 FILLER_305_439 ();
 b15zdnd11an1n04x5 FILLER_305_455 ();
 b15zdnd11an1n64x5 FILLER_305_471 ();
 b15zdnd11an1n16x5 FILLER_305_535 ();
 b15zdnd11an1n08x5 FILLER_305_551 ();
 b15zdnd00an1n02x5 FILLER_305_559 ();
 b15zdnd00an1n01x5 FILLER_305_561 ();
 b15zdnd11an1n04x5 FILLER_305_567 ();
 b15zdnd11an1n04x5 FILLER_305_583 ();
 b15zdnd11an1n08x5 FILLER_305_598 ();
 b15zdnd11an1n04x5 FILLER_305_606 ();
 b15zdnd11an1n16x5 FILLER_305_617 ();
 b15zdnd11an1n08x5 FILLER_305_633 ();
 b15zdnd11an1n04x5 FILLER_305_641 ();
 b15zdnd00an1n01x5 FILLER_305_645 ();
 b15zdnd11an1n64x5 FILLER_305_652 ();
 b15zdnd11an1n16x5 FILLER_305_716 ();
 b15zdnd11an1n04x5 FILLER_305_732 ();
 b15zdnd11an1n08x5 FILLER_305_742 ();
 b15zdnd11an1n04x5 FILLER_305_750 ();
 b15zdnd00an1n01x5 FILLER_305_754 ();
 b15zdnd11an1n16x5 FILLER_305_760 ();
 b15zdnd11an1n08x5 FILLER_305_776 ();
 b15zdnd11an1n04x5 FILLER_305_784 ();
 b15zdnd00an1n01x5 FILLER_305_788 ();
 b15zdnd11an1n64x5 FILLER_305_820 ();
 b15zdnd11an1n32x5 FILLER_305_884 ();
 b15zdnd00an1n01x5 FILLER_305_916 ();
 b15zdnd11an1n16x5 FILLER_305_935 ();
 b15zdnd11an1n04x5 FILLER_305_951 ();
 b15zdnd00an1n01x5 FILLER_305_955 ();
 b15zdnd11an1n08x5 FILLER_305_966 ();
 b15zdnd00an1n02x5 FILLER_305_974 ();
 b15zdnd00an1n01x5 FILLER_305_976 ();
 b15zdnd11an1n04x5 FILLER_305_1003 ();
 b15zdnd11an1n64x5 FILLER_305_1019 ();
 b15zdnd00an1n02x5 FILLER_305_1083 ();
 b15zdnd00an1n01x5 FILLER_305_1085 ();
 b15zdnd11an1n16x5 FILLER_305_1098 ();
 b15zdnd11an1n08x5 FILLER_305_1114 ();
 b15zdnd11an1n08x5 FILLER_305_1129 ();
 b15zdnd00an1n01x5 FILLER_305_1137 ();
 b15zdnd11an1n08x5 FILLER_305_1158 ();
 b15zdnd11an1n16x5 FILLER_305_1173 ();
 b15zdnd11an1n08x5 FILLER_305_1189 ();
 b15zdnd11an1n04x5 FILLER_305_1197 ();
 b15zdnd00an1n02x5 FILLER_305_1201 ();
 b15zdnd00an1n01x5 FILLER_305_1203 ();
 b15zdnd11an1n32x5 FILLER_305_1212 ();
 b15zdnd11an1n16x5 FILLER_305_1244 ();
 b15zdnd11an1n04x5 FILLER_305_1260 ();
 b15zdnd00an1n01x5 FILLER_305_1264 ();
 b15zdnd11an1n08x5 FILLER_305_1277 ();
 b15zdnd00an1n01x5 FILLER_305_1285 ();
 b15zdnd11an1n04x5 FILLER_305_1292 ();
 b15zdnd11an1n64x5 FILLER_305_1312 ();
 b15zdnd11an1n08x5 FILLER_305_1376 ();
 b15zdnd00an1n01x5 FILLER_305_1384 ();
 b15zdnd11an1n64x5 FILLER_305_1405 ();
 b15zdnd11an1n32x5 FILLER_305_1469 ();
 b15zdnd11an1n08x5 FILLER_305_1501 ();
 b15zdnd00an1n02x5 FILLER_305_1509 ();
 b15zdnd00an1n01x5 FILLER_305_1511 ();
 b15zdnd11an1n16x5 FILLER_305_1526 ();
 b15zdnd00an1n01x5 FILLER_305_1542 ();
 b15zdnd11an1n08x5 FILLER_305_1554 ();
 b15zdnd00an1n02x5 FILLER_305_1562 ();
 b15zdnd11an1n32x5 FILLER_305_1570 ();
 b15zdnd11an1n04x5 FILLER_305_1602 ();
 b15zdnd00an1n02x5 FILLER_305_1606 ();
 b15zdnd00an1n01x5 FILLER_305_1608 ();
 b15zdnd11an1n64x5 FILLER_305_1617 ();
 b15zdnd11an1n04x5 FILLER_305_1681 ();
 b15zdnd11an1n32x5 FILLER_305_1691 ();
 b15zdnd11an1n08x5 FILLER_305_1723 ();
 b15zdnd11an1n04x5 FILLER_305_1731 ();
 b15zdnd00an1n02x5 FILLER_305_1735 ();
 b15zdnd00an1n01x5 FILLER_305_1737 ();
 b15zdnd11an1n04x5 FILLER_305_1749 ();
 b15zdnd11an1n16x5 FILLER_305_1773 ();
 b15zdnd11an1n08x5 FILLER_305_1789 ();
 b15zdnd11an1n04x5 FILLER_305_1797 ();
 b15zdnd00an1n01x5 FILLER_305_1801 ();
 b15zdnd11an1n08x5 FILLER_305_1820 ();
 b15zdnd00an1n02x5 FILLER_305_1828 ();
 b15zdnd00an1n01x5 FILLER_305_1830 ();
 b15zdnd11an1n64x5 FILLER_305_1838 ();
 b15zdnd11an1n08x5 FILLER_305_1902 ();
 b15zdnd00an1n02x5 FILLER_305_1910 ();
 b15zdnd00an1n01x5 FILLER_305_1912 ();
 b15zdnd11an1n08x5 FILLER_305_1933 ();
 b15zdnd00an1n02x5 FILLER_305_1941 ();
 b15zdnd11an1n08x5 FILLER_305_1955 ();
 b15zdnd11an1n04x5 FILLER_305_1969 ();
 b15zdnd11an1n32x5 FILLER_305_1978 ();
 b15zdnd11an1n16x5 FILLER_305_2010 ();
 b15zdnd11an1n08x5 FILLER_305_2026 ();
 b15zdnd11an1n04x5 FILLER_305_2034 ();
 b15zdnd00an1n01x5 FILLER_305_2038 ();
 b15zdnd11an1n04x5 FILLER_305_2044 ();
 b15zdnd11an1n08x5 FILLER_305_2052 ();
 b15zdnd11an1n04x5 FILLER_305_2060 ();
 b15zdnd00an1n02x5 FILLER_305_2064 ();
 b15zdnd11an1n04x5 FILLER_305_2078 ();
 b15zdnd11an1n64x5 FILLER_305_2094 ();
 b15zdnd11an1n32x5 FILLER_305_2158 ();
 b15zdnd11an1n08x5 FILLER_305_2190 ();
 b15zdnd11an1n04x5 FILLER_305_2198 ();
 b15zdnd00an1n01x5 FILLER_305_2202 ();
 b15zdnd11an1n16x5 FILLER_305_2212 ();
 b15zdnd00an1n02x5 FILLER_305_2228 ();
 b15zdnd11an1n32x5 FILLER_305_2248 ();
 b15zdnd11an1n04x5 FILLER_305_2280 ();
 b15zdnd11an1n64x5 FILLER_306_8 ();
 b15zdnd11an1n64x5 FILLER_306_72 ();
 b15zdnd11an1n64x5 FILLER_306_136 ();
 b15zdnd11an1n16x5 FILLER_306_200 ();
 b15zdnd00an1n02x5 FILLER_306_216 ();
 b15zdnd11an1n64x5 FILLER_306_234 ();
 b15zdnd11an1n16x5 FILLER_306_298 ();
 b15zdnd00an1n02x5 FILLER_306_314 ();
 b15zdnd11an1n04x5 FILLER_306_334 ();
 b15zdnd11an1n32x5 FILLER_306_369 ();
 b15zdnd11an1n16x5 FILLER_306_401 ();
 b15zdnd00an1n01x5 FILLER_306_417 ();
 b15zdnd11an1n08x5 FILLER_306_423 ();
 b15zdnd11an1n04x5 FILLER_306_431 ();
 b15zdnd00an1n01x5 FILLER_306_435 ();
 b15zdnd11an1n64x5 FILLER_306_443 ();
 b15zdnd11an1n64x5 FILLER_306_507 ();
 b15zdnd11an1n32x5 FILLER_306_571 ();
 b15zdnd00an1n02x5 FILLER_306_603 ();
 b15zdnd11an1n32x5 FILLER_306_620 ();
 b15zdnd11an1n16x5 FILLER_306_658 ();
 b15zdnd11an1n08x5 FILLER_306_674 ();
 b15zdnd00an1n01x5 FILLER_306_682 ();
 b15zdnd11an1n08x5 FILLER_306_703 ();
 b15zdnd11an1n04x5 FILLER_306_711 ();
 b15zdnd00an1n02x5 FILLER_306_715 ();
 b15zdnd00an1n01x5 FILLER_306_717 ();
 b15zdnd11an1n08x5 FILLER_306_726 ();
 b15zdnd11an1n04x5 FILLER_306_734 ();
 b15zdnd00an1n01x5 FILLER_306_738 ();
 b15zdnd11an1n16x5 FILLER_306_759 ();
 b15zdnd11an1n08x5 FILLER_306_775 ();
 b15zdnd11an1n04x5 FILLER_306_783 ();
 b15zdnd00an1n02x5 FILLER_306_787 ();
 b15zdnd00an1n01x5 FILLER_306_789 ();
 b15zdnd11an1n08x5 FILLER_306_811 ();
 b15zdnd11an1n04x5 FILLER_306_819 ();
 b15zdnd00an1n02x5 FILLER_306_823 ();
 b15zdnd11an1n64x5 FILLER_306_856 ();
 b15zdnd11an1n32x5 FILLER_306_920 ();
 b15zdnd11an1n16x5 FILLER_306_952 ();
 b15zdnd11an1n64x5 FILLER_306_983 ();
 b15zdnd11an1n64x5 FILLER_306_1047 ();
 b15zdnd11an1n04x5 FILLER_306_1111 ();
 b15zdnd00an1n02x5 FILLER_306_1115 ();
 b15zdnd11an1n32x5 FILLER_306_1135 ();
 b15zdnd00an1n01x5 FILLER_306_1167 ();
 b15zdnd11an1n04x5 FILLER_306_1194 ();
 b15zdnd11an1n04x5 FILLER_306_1203 ();
 b15zdnd11an1n16x5 FILLER_306_1212 ();
 b15zdnd11an1n08x5 FILLER_306_1228 ();
 b15zdnd00an1n02x5 FILLER_306_1236 ();
 b15zdnd11an1n16x5 FILLER_306_1249 ();
 b15zdnd00an1n02x5 FILLER_306_1265 ();
 b15zdnd11an1n16x5 FILLER_306_1277 ();
 b15zdnd11an1n08x5 FILLER_306_1293 ();
 b15zdnd11an1n04x5 FILLER_306_1301 ();
 b15zdnd00an1n02x5 FILLER_306_1305 ();
 b15zdnd11an1n64x5 FILLER_306_1323 ();
 b15zdnd11an1n08x5 FILLER_306_1387 ();
 b15zdnd11an1n04x5 FILLER_306_1395 ();
 b15zdnd00an1n02x5 FILLER_306_1399 ();
 b15zdnd00an1n01x5 FILLER_306_1401 ();
 b15zdnd11an1n64x5 FILLER_306_1407 ();
 b15zdnd11an1n16x5 FILLER_306_1478 ();
 b15zdnd11an1n04x5 FILLER_306_1494 ();
 b15zdnd00an1n02x5 FILLER_306_1498 ();
 b15zdnd11an1n64x5 FILLER_306_1509 ();
 b15zdnd11an1n32x5 FILLER_306_1573 ();
 b15zdnd00an1n02x5 FILLER_306_1605 ();
 b15zdnd00an1n01x5 FILLER_306_1607 ();
 b15zdnd11an1n04x5 FILLER_306_1619 ();
 b15zdnd11an1n64x5 FILLER_306_1630 ();
 b15zdnd11an1n64x5 FILLER_306_1694 ();
 b15zdnd11an1n64x5 FILLER_306_1758 ();
 b15zdnd11an1n64x5 FILLER_306_1822 ();
 b15zdnd11an1n32x5 FILLER_306_1886 ();
 b15zdnd11an1n08x5 FILLER_306_1918 ();
 b15zdnd00an1n02x5 FILLER_306_1926 ();
 b15zdnd00an1n01x5 FILLER_306_1928 ();
 b15zdnd11an1n16x5 FILLER_306_1948 ();
 b15zdnd11an1n64x5 FILLER_306_1969 ();
 b15zdnd11an1n16x5 FILLER_306_2033 ();
 b15zdnd11an1n08x5 FILLER_306_2049 ();
 b15zdnd11an1n04x5 FILLER_306_2057 ();
 b15zdnd11an1n64x5 FILLER_306_2067 ();
 b15zdnd11an1n16x5 FILLER_306_2131 ();
 b15zdnd11an1n04x5 FILLER_306_2147 ();
 b15zdnd00an1n02x5 FILLER_306_2151 ();
 b15zdnd00an1n01x5 FILLER_306_2153 ();
 b15zdnd00an1n02x5 FILLER_306_2162 ();
 b15zdnd00an1n01x5 FILLER_306_2164 ();
 b15zdnd11an1n16x5 FILLER_306_2171 ();
 b15zdnd00an1n01x5 FILLER_306_2187 ();
 b15zdnd11an1n04x5 FILLER_306_2194 ();
 b15zdnd11an1n32x5 FILLER_306_2218 ();
 b15zdnd11an1n16x5 FILLER_306_2250 ();
 b15zdnd11an1n08x5 FILLER_306_2266 ();
 b15zdnd00an1n02x5 FILLER_306_2274 ();
 b15zdnd11an1n64x5 FILLER_307_0 ();
 b15zdnd11an1n64x5 FILLER_307_64 ();
 b15zdnd11an1n64x5 FILLER_307_128 ();
 b15zdnd11an1n32x5 FILLER_307_192 ();
 b15zdnd11an1n04x5 FILLER_307_224 ();
 b15zdnd11an1n64x5 FILLER_307_233 ();
 b15zdnd11an1n64x5 FILLER_307_297 ();
 b15zdnd11an1n32x5 FILLER_307_361 ();
 b15zdnd11an1n16x5 FILLER_307_399 ();
 b15zdnd11an1n04x5 FILLER_307_428 ();
 b15zdnd11an1n04x5 FILLER_307_444 ();
 b15zdnd11an1n32x5 FILLER_307_464 ();
 b15zdnd11an1n04x5 FILLER_307_496 ();
 b15zdnd00an1n02x5 FILLER_307_500 ();
 b15zdnd11an1n64x5 FILLER_307_515 ();
 b15zdnd11an1n32x5 FILLER_307_579 ();
 b15zdnd11an1n16x5 FILLER_307_611 ();
 b15zdnd00an1n02x5 FILLER_307_627 ();
 b15zdnd11an1n32x5 FILLER_307_661 ();
 b15zdnd11an1n04x5 FILLER_307_713 ();
 b15zdnd11an1n16x5 FILLER_307_748 ();
 b15zdnd11an1n04x5 FILLER_307_764 ();
 b15zdnd00an1n01x5 FILLER_307_768 ();
 b15zdnd11an1n04x5 FILLER_307_790 ();
 b15zdnd00an1n02x5 FILLER_307_794 ();
 b15zdnd11an1n08x5 FILLER_307_827 ();
 b15zdnd11an1n04x5 FILLER_307_835 ();
 b15zdnd00an1n02x5 FILLER_307_839 ();
 b15zdnd00an1n01x5 FILLER_307_841 ();
 b15zdnd11an1n64x5 FILLER_307_854 ();
 b15zdnd11an1n08x5 FILLER_307_918 ();
 b15zdnd11an1n04x5 FILLER_307_926 ();
 b15zdnd00an1n02x5 FILLER_307_930 ();
 b15zdnd11an1n64x5 FILLER_307_944 ();
 b15zdnd11an1n64x5 FILLER_307_1008 ();
 b15zdnd11an1n04x5 FILLER_307_1072 ();
 b15zdnd00an1n02x5 FILLER_307_1076 ();
 b15zdnd11an1n32x5 FILLER_307_1109 ();
 b15zdnd11an1n16x5 FILLER_307_1141 ();
 b15zdnd11an1n08x5 FILLER_307_1157 ();
 b15zdnd00an1n02x5 FILLER_307_1165 ();
 b15zdnd00an1n01x5 FILLER_307_1167 ();
 b15zdnd11an1n32x5 FILLER_307_1175 ();
 b15zdnd00an1n02x5 FILLER_307_1207 ();
 b15zdnd11an1n16x5 FILLER_307_1214 ();
 b15zdnd00an1n02x5 FILLER_307_1230 ();
 b15zdnd11an1n32x5 FILLER_307_1241 ();
 b15zdnd11an1n16x5 FILLER_307_1273 ();
 b15zdnd11an1n04x5 FILLER_307_1289 ();
 b15zdnd00an1n02x5 FILLER_307_1293 ();
 b15zdnd00an1n01x5 FILLER_307_1295 ();
 b15zdnd11an1n64x5 FILLER_307_1328 ();
 b15zdnd11an1n64x5 FILLER_307_1392 ();
 b15zdnd11an1n08x5 FILLER_307_1456 ();
 b15zdnd11an1n04x5 FILLER_307_1469 ();
 b15zdnd11an1n08x5 FILLER_307_1480 ();
 b15zdnd11an1n04x5 FILLER_307_1488 ();
 b15zdnd11an1n04x5 FILLER_307_1498 ();
 b15zdnd11an1n64x5 FILLER_307_1518 ();
 b15zdnd11an1n64x5 FILLER_307_1582 ();
 b15zdnd11an1n08x5 FILLER_307_1646 ();
 b15zdnd11an1n04x5 FILLER_307_1654 ();
 b15zdnd00an1n01x5 FILLER_307_1658 ();
 b15zdnd11an1n16x5 FILLER_307_1665 ();
 b15zdnd11an1n04x5 FILLER_307_1681 ();
 b15zdnd00an1n02x5 FILLER_307_1685 ();
 b15zdnd00an1n01x5 FILLER_307_1687 ();
 b15zdnd11an1n04x5 FILLER_307_1695 ();
 b15zdnd11an1n04x5 FILLER_307_1703 ();
 b15zdnd11an1n04x5 FILLER_307_1719 ();
 b15zdnd00an1n01x5 FILLER_307_1723 ();
 b15zdnd11an1n04x5 FILLER_307_1736 ();
 b15zdnd00an1n02x5 FILLER_307_1740 ();
 b15zdnd00an1n01x5 FILLER_307_1742 ();
 b15zdnd11an1n16x5 FILLER_307_1759 ();
 b15zdnd11an1n08x5 FILLER_307_1775 ();
 b15zdnd11an1n64x5 FILLER_307_1814 ();
 b15zdnd11an1n08x5 FILLER_307_1878 ();
 b15zdnd11an1n04x5 FILLER_307_1886 ();
 b15zdnd00an1n02x5 FILLER_307_1890 ();
 b15zdnd11an1n16x5 FILLER_307_1918 ();
 b15zdnd11an1n08x5 FILLER_307_1934 ();
 b15zdnd11an1n04x5 FILLER_307_1942 ();
 b15zdnd11an1n32x5 FILLER_307_1962 ();
 b15zdnd11an1n08x5 FILLER_307_1994 ();
 b15zdnd00an1n01x5 FILLER_307_2002 ();
 b15zdnd11an1n04x5 FILLER_307_2009 ();
 b15zdnd11an1n16x5 FILLER_307_2021 ();
 b15zdnd11an1n08x5 FILLER_307_2037 ();
 b15zdnd00an1n01x5 FILLER_307_2045 ();
 b15zdnd11an1n04x5 FILLER_307_2055 ();
 b15zdnd11an1n64x5 FILLER_307_2064 ();
 b15zdnd11an1n32x5 FILLER_307_2128 ();
 b15zdnd11an1n04x5 FILLER_307_2169 ();
 b15zdnd11an1n64x5 FILLER_307_2194 ();
 b15zdnd11an1n16x5 FILLER_307_2258 ();
 b15zdnd11an1n08x5 FILLER_307_2274 ();
 b15zdnd00an1n02x5 FILLER_307_2282 ();
 b15zdnd11an1n64x5 FILLER_308_8 ();
 b15zdnd11an1n64x5 FILLER_308_72 ();
 b15zdnd11an1n64x5 FILLER_308_136 ();
 b15zdnd11an1n16x5 FILLER_308_200 ();
 b15zdnd11an1n08x5 FILLER_308_216 ();
 b15zdnd00an1n02x5 FILLER_308_224 ();
 b15zdnd00an1n01x5 FILLER_308_226 ();
 b15zdnd11an1n16x5 FILLER_308_233 ();
 b15zdnd00an1n02x5 FILLER_308_249 ();
 b15zdnd00an1n01x5 FILLER_308_251 ();
 b15zdnd11an1n64x5 FILLER_308_259 ();
 b15zdnd11an1n16x5 FILLER_308_323 ();
 b15zdnd11an1n08x5 FILLER_308_339 ();
 b15zdnd11an1n04x5 FILLER_308_347 ();
 b15zdnd00an1n02x5 FILLER_308_351 ();
 b15zdnd11an1n16x5 FILLER_308_368 ();
 b15zdnd11an1n08x5 FILLER_308_384 ();
 b15zdnd00an1n02x5 FILLER_308_392 ();
 b15zdnd11an1n16x5 FILLER_308_403 ();
 b15zdnd00an1n01x5 FILLER_308_419 ();
 b15zdnd11an1n32x5 FILLER_308_436 ();
 b15zdnd11an1n04x5 FILLER_308_484 ();
 b15zdnd11an1n64x5 FILLER_308_519 ();
 b15zdnd11an1n64x5 FILLER_308_583 ();
 b15zdnd11an1n64x5 FILLER_308_647 ();
 b15zdnd11an1n04x5 FILLER_308_711 ();
 b15zdnd00an1n02x5 FILLER_308_715 ();
 b15zdnd00an1n01x5 FILLER_308_717 ();
 b15zdnd11an1n64x5 FILLER_308_726 ();
 b15zdnd11an1n64x5 FILLER_308_790 ();
 b15zdnd11an1n32x5 FILLER_308_854 ();
 b15zdnd00an1n02x5 FILLER_308_886 ();
 b15zdnd11an1n16x5 FILLER_308_911 ();
 b15zdnd00an1n02x5 FILLER_308_927 ();
 b15zdnd11an1n64x5 FILLER_308_954 ();
 b15zdnd11an1n32x5 FILLER_308_1018 ();
 b15zdnd11an1n16x5 FILLER_308_1050 ();
 b15zdnd11an1n08x5 FILLER_308_1066 ();
 b15zdnd11an1n04x5 FILLER_308_1074 ();
 b15zdnd00an1n02x5 FILLER_308_1078 ();
 b15zdnd00an1n01x5 FILLER_308_1080 ();
 b15zdnd11an1n32x5 FILLER_308_1085 ();
 b15zdnd11an1n16x5 FILLER_308_1117 ();
 b15zdnd11an1n08x5 FILLER_308_1133 ();
 b15zdnd11an1n04x5 FILLER_308_1141 ();
 b15zdnd00an1n02x5 FILLER_308_1145 ();
 b15zdnd11an1n64x5 FILLER_308_1156 ();
 b15zdnd11an1n04x5 FILLER_308_1220 ();
 b15zdnd00an1n02x5 FILLER_308_1224 ();
 b15zdnd00an1n01x5 FILLER_308_1226 ();
 b15zdnd11an1n04x5 FILLER_308_1233 ();
 b15zdnd11an1n64x5 FILLER_308_1247 ();
 b15zdnd11an1n32x5 FILLER_308_1311 ();
 b15zdnd11an1n08x5 FILLER_308_1343 ();
 b15zdnd11an1n04x5 FILLER_308_1351 ();
 b15zdnd00an1n02x5 FILLER_308_1355 ();
 b15zdnd00an1n01x5 FILLER_308_1357 ();
 b15zdnd11an1n04x5 FILLER_308_1369 ();
 b15zdnd00an1n02x5 FILLER_308_1373 ();
 b15zdnd00an1n01x5 FILLER_308_1375 ();
 b15zdnd11an1n32x5 FILLER_308_1387 ();
 b15zdnd11an1n08x5 FILLER_308_1419 ();
 b15zdnd11an1n04x5 FILLER_308_1427 ();
 b15zdnd00an1n01x5 FILLER_308_1431 ();
 b15zdnd11an1n32x5 FILLER_308_1450 ();
 b15zdnd11an1n04x5 FILLER_308_1482 ();
 b15zdnd00an1n02x5 FILLER_308_1486 ();
 b15zdnd00an1n01x5 FILLER_308_1488 ();
 b15zdnd11an1n32x5 FILLER_308_1499 ();
 b15zdnd11an1n16x5 FILLER_308_1531 ();
 b15zdnd11an1n08x5 FILLER_308_1547 ();
 b15zdnd11an1n04x5 FILLER_308_1555 ();
 b15zdnd00an1n02x5 FILLER_308_1559 ();
 b15zdnd11an1n64x5 FILLER_308_1587 ();
 b15zdnd11an1n08x5 FILLER_308_1651 ();
 b15zdnd11an1n32x5 FILLER_308_1665 ();
 b15zdnd11an1n08x5 FILLER_308_1697 ();
 b15zdnd00an1n02x5 FILLER_308_1705 ();
 b15zdnd11an1n32x5 FILLER_308_1715 ();
 b15zdnd11an1n16x5 FILLER_308_1747 ();
 b15zdnd11an1n04x5 FILLER_308_1763 ();
 b15zdnd00an1n01x5 FILLER_308_1767 ();
 b15zdnd11an1n04x5 FILLER_308_1780 ();
 b15zdnd11an1n32x5 FILLER_308_1788 ();
 b15zdnd11an1n16x5 FILLER_308_1820 ();
 b15zdnd11an1n08x5 FILLER_308_1836 ();
 b15zdnd11an1n04x5 FILLER_308_1844 ();
 b15zdnd00an1n01x5 FILLER_308_1848 ();
 b15zdnd11an1n04x5 FILLER_308_1869 ();
 b15zdnd00an1n02x5 FILLER_308_1873 ();
 b15zdnd11an1n32x5 FILLER_308_1901 ();
 b15zdnd00an1n02x5 FILLER_308_1933 ();
 b15zdnd11an1n32x5 FILLER_308_1961 ();
 b15zdnd11an1n04x5 FILLER_308_1993 ();
 b15zdnd11an1n04x5 FILLER_308_2008 ();
 b15zdnd11an1n08x5 FILLER_308_2028 ();
 b15zdnd11an1n04x5 FILLER_308_2036 ();
 b15zdnd00an1n02x5 FILLER_308_2040 ();
 b15zdnd11an1n16x5 FILLER_308_2054 ();
 b15zdnd00an1n02x5 FILLER_308_2070 ();
 b15zdnd00an1n01x5 FILLER_308_2072 ();
 b15zdnd11an1n32x5 FILLER_308_2078 ();
 b15zdnd11an1n16x5 FILLER_308_2110 ();
 b15zdnd11an1n08x5 FILLER_308_2126 ();
 b15zdnd00an1n02x5 FILLER_308_2134 ();
 b15zdnd00an1n01x5 FILLER_308_2136 ();
 b15zdnd11an1n08x5 FILLER_308_2144 ();
 b15zdnd00an1n02x5 FILLER_308_2152 ();
 b15zdnd11an1n04x5 FILLER_308_2162 ();
 b15zdnd00an1n02x5 FILLER_308_2166 ();
 b15zdnd11an1n16x5 FILLER_308_2173 ();
 b15zdnd11an1n08x5 FILLER_308_2189 ();
 b15zdnd11an1n04x5 FILLER_308_2197 ();
 b15zdnd00an1n01x5 FILLER_308_2201 ();
 b15zdnd11an1n64x5 FILLER_308_2207 ();
 b15zdnd11an1n04x5 FILLER_308_2271 ();
 b15zdnd00an1n01x5 FILLER_308_2275 ();
 b15zdnd11an1n64x5 FILLER_309_0 ();
 b15zdnd11an1n64x5 FILLER_309_64 ();
 b15zdnd11an1n64x5 FILLER_309_128 ();
 b15zdnd11an1n64x5 FILLER_309_192 ();
 b15zdnd11an1n16x5 FILLER_309_256 ();
 b15zdnd11an1n04x5 FILLER_309_272 ();
 b15zdnd00an1n02x5 FILLER_309_276 ();
 b15zdnd11an1n04x5 FILLER_309_292 ();
 b15zdnd11an1n04x5 FILLER_309_309 ();
 b15zdnd11an1n08x5 FILLER_309_345 ();
 b15zdnd11an1n04x5 FILLER_309_353 ();
 b15zdnd11an1n64x5 FILLER_309_369 ();
 b15zdnd11an1n64x5 FILLER_309_433 ();
 b15zdnd11an1n64x5 FILLER_309_497 ();
 b15zdnd11an1n64x5 FILLER_309_561 ();
 b15zdnd11an1n64x5 FILLER_309_625 ();
 b15zdnd11an1n64x5 FILLER_309_689 ();
 b15zdnd11an1n64x5 FILLER_309_753 ();
 b15zdnd11an1n08x5 FILLER_309_817 ();
 b15zdnd11an1n04x5 FILLER_309_825 ();
 b15zdnd00an1n01x5 FILLER_309_829 ();
 b15zdnd11an1n04x5 FILLER_309_840 ();
 b15zdnd11an1n32x5 FILLER_309_853 ();
 b15zdnd11an1n16x5 FILLER_309_885 ();
 b15zdnd11an1n08x5 FILLER_309_901 ();
 b15zdnd11an1n04x5 FILLER_309_914 ();
 b15zdnd11an1n32x5 FILLER_309_922 ();
 b15zdnd00an1n02x5 FILLER_309_954 ();
 b15zdnd00an1n01x5 FILLER_309_956 ();
 b15zdnd11an1n04x5 FILLER_309_978 ();
 b15zdnd11an1n16x5 FILLER_309_993 ();
 b15zdnd00an1n02x5 FILLER_309_1009 ();
 b15zdnd00an1n01x5 FILLER_309_1011 ();
 b15zdnd11an1n04x5 FILLER_309_1037 ();
 b15zdnd11an1n04x5 FILLER_309_1046 ();
 b15zdnd11an1n04x5 FILLER_309_1054 ();
 b15zdnd00an1n01x5 FILLER_309_1058 ();
 b15zdnd11an1n08x5 FILLER_309_1063 ();
 b15zdnd11an1n04x5 FILLER_309_1071 ();
 b15zdnd11an1n04x5 FILLER_309_1080 ();
 b15zdnd11an1n16x5 FILLER_309_1099 ();
 b15zdnd11an1n08x5 FILLER_309_1115 ();
 b15zdnd00an1n01x5 FILLER_309_1123 ();
 b15zdnd11an1n64x5 FILLER_309_1138 ();
 b15zdnd11an1n64x5 FILLER_309_1202 ();
 b15zdnd11an1n64x5 FILLER_309_1266 ();
 b15zdnd11an1n32x5 FILLER_309_1330 ();
 b15zdnd00an1n01x5 FILLER_309_1362 ();
 b15zdnd11an1n32x5 FILLER_309_1383 ();
 b15zdnd00an1n01x5 FILLER_309_1415 ();
 b15zdnd11an1n04x5 FILLER_309_1442 ();
 b15zdnd11an1n32x5 FILLER_309_1463 ();
 b15zdnd11an1n16x5 FILLER_309_1495 ();
 b15zdnd11an1n08x5 FILLER_309_1511 ();
 b15zdnd00an1n02x5 FILLER_309_1519 ();
 b15zdnd00an1n01x5 FILLER_309_1521 ();
 b15zdnd11an1n08x5 FILLER_309_1531 ();
 b15zdnd00an1n02x5 FILLER_309_1539 ();
 b15zdnd00an1n01x5 FILLER_309_1541 ();
 b15zdnd11an1n16x5 FILLER_309_1558 ();
 b15zdnd11an1n04x5 FILLER_309_1574 ();
 b15zdnd11an1n32x5 FILLER_309_1584 ();
 b15zdnd11an1n16x5 FILLER_309_1616 ();
 b15zdnd11an1n08x5 FILLER_309_1632 ();
 b15zdnd11an1n04x5 FILLER_309_1640 ();
 b15zdnd00an1n01x5 FILLER_309_1644 ();
 b15zdnd11an1n04x5 FILLER_309_1649 ();
 b15zdnd00an1n02x5 FILLER_309_1653 ();
 b15zdnd00an1n01x5 FILLER_309_1655 ();
 b15zdnd11an1n64x5 FILLER_309_1661 ();
 b15zdnd11an1n32x5 FILLER_309_1725 ();
 b15zdnd11an1n08x5 FILLER_309_1757 ();
 b15zdnd11an1n04x5 FILLER_309_1765 ();
 b15zdnd00an1n02x5 FILLER_309_1769 ();
 b15zdnd11an1n08x5 FILLER_309_1776 ();
 b15zdnd00an1n01x5 FILLER_309_1784 ();
 b15zdnd11an1n16x5 FILLER_309_1789 ();
 b15zdnd11an1n04x5 FILLER_309_1814 ();
 b15zdnd00an1n01x5 FILLER_309_1818 ();
 b15zdnd11an1n04x5 FILLER_309_1828 ();
 b15zdnd00an1n02x5 FILLER_309_1832 ();
 b15zdnd00an1n01x5 FILLER_309_1834 ();
 b15zdnd11an1n32x5 FILLER_309_1855 ();
 b15zdnd11an1n16x5 FILLER_309_1887 ();
 b15zdnd11an1n08x5 FILLER_309_1903 ();
 b15zdnd11an1n04x5 FILLER_309_1911 ();
 b15zdnd11an1n16x5 FILLER_309_1935 ();
 b15zdnd11an1n04x5 FILLER_309_1951 ();
 b15zdnd00an1n02x5 FILLER_309_1955 ();
 b15zdnd11an1n04x5 FILLER_309_1964 ();
 b15zdnd11an1n08x5 FILLER_309_1984 ();
 b15zdnd00an1n01x5 FILLER_309_1992 ();
 b15zdnd11an1n16x5 FILLER_309_2019 ();
 b15zdnd00an1n01x5 FILLER_309_2035 ();
 b15zdnd11an1n16x5 FILLER_309_2046 ();
 b15zdnd11an1n08x5 FILLER_309_2062 ();
 b15zdnd00an1n02x5 FILLER_309_2070 ();
 b15zdnd11an1n16x5 FILLER_309_2077 ();
 b15zdnd11an1n04x5 FILLER_309_2093 ();
 b15zdnd00an1n01x5 FILLER_309_2097 ();
 b15zdnd11an1n04x5 FILLER_309_2104 ();
 b15zdnd11an1n04x5 FILLER_309_2120 ();
 b15zdnd11an1n16x5 FILLER_309_2138 ();
 b15zdnd11an1n04x5 FILLER_309_2154 ();
 b15zdnd11an1n64x5 FILLER_309_2168 ();
 b15zdnd11an1n32x5 FILLER_309_2232 ();
 b15zdnd11an1n16x5 FILLER_309_2264 ();
 b15zdnd11an1n04x5 FILLER_309_2280 ();
 b15zdnd11an1n64x5 FILLER_310_8 ();
 b15zdnd11an1n64x5 FILLER_310_72 ();
 b15zdnd11an1n64x5 FILLER_310_136 ();
 b15zdnd11an1n64x5 FILLER_310_200 ();
 b15zdnd11an1n08x5 FILLER_310_264 ();
 b15zdnd11an1n04x5 FILLER_310_288 ();
 b15zdnd11an1n32x5 FILLER_310_312 ();
 b15zdnd11an1n16x5 FILLER_310_359 ();
 b15zdnd11an1n08x5 FILLER_310_375 ();
 b15zdnd11an1n16x5 FILLER_310_398 ();
 b15zdnd11an1n08x5 FILLER_310_414 ();
 b15zdnd11an1n04x5 FILLER_310_448 ();
 b15zdnd11an1n64x5 FILLER_310_468 ();
 b15zdnd00an1n01x5 FILLER_310_532 ();
 b15zdnd11an1n04x5 FILLER_310_564 ();
 b15zdnd11an1n16x5 FILLER_310_573 ();
 b15zdnd00an1n01x5 FILLER_310_589 ();
 b15zdnd11an1n16x5 FILLER_310_610 ();
 b15zdnd11an1n08x5 FILLER_310_626 ();
 b15zdnd11an1n64x5 FILLER_310_654 ();
 b15zdnd11an1n64x5 FILLER_310_726 ();
 b15zdnd11an1n32x5 FILLER_310_790 ();
 b15zdnd11an1n16x5 FILLER_310_822 ();
 b15zdnd11an1n64x5 FILLER_310_847 ();
 b15zdnd11an1n64x5 FILLER_310_911 ();
 b15zdnd11an1n04x5 FILLER_310_975 ();
 b15zdnd00an1n02x5 FILLER_310_979 ();
 b15zdnd00an1n01x5 FILLER_310_981 ();
 b15zdnd11an1n32x5 FILLER_310_1002 ();
 b15zdnd00an1n01x5 FILLER_310_1034 ();
 b15zdnd11an1n08x5 FILLER_310_1051 ();
 b15zdnd11an1n04x5 FILLER_310_1059 ();
 b15zdnd00an1n02x5 FILLER_310_1063 ();
 b15zdnd11an1n16x5 FILLER_310_1069 ();
 b15zdnd00an1n02x5 FILLER_310_1085 ();
 b15zdnd00an1n01x5 FILLER_310_1087 ();
 b15zdnd11an1n32x5 FILLER_310_1092 ();
 b15zdnd11an1n16x5 FILLER_310_1124 ();
 b15zdnd11an1n08x5 FILLER_310_1140 ();
 b15zdnd00an1n02x5 FILLER_310_1148 ();
 b15zdnd00an1n01x5 FILLER_310_1150 ();
 b15zdnd11an1n64x5 FILLER_310_1171 ();
 b15zdnd11an1n16x5 FILLER_310_1235 ();
 b15zdnd11an1n08x5 FILLER_310_1251 ();
 b15zdnd11an1n04x5 FILLER_310_1259 ();
 b15zdnd00an1n01x5 FILLER_310_1263 ();
 b15zdnd11an1n64x5 FILLER_310_1273 ();
 b15zdnd11an1n16x5 FILLER_310_1337 ();
 b15zdnd11an1n08x5 FILLER_310_1353 ();
 b15zdnd00an1n01x5 FILLER_310_1361 ();
 b15zdnd11an1n32x5 FILLER_310_1367 ();
 b15zdnd11an1n04x5 FILLER_310_1399 ();
 b15zdnd00an1n02x5 FILLER_310_1403 ();
 b15zdnd00an1n01x5 FILLER_310_1405 ();
 b15zdnd11an1n16x5 FILLER_310_1410 ();
 b15zdnd11an1n08x5 FILLER_310_1426 ();
 b15zdnd11an1n04x5 FILLER_310_1434 ();
 b15zdnd00an1n02x5 FILLER_310_1438 ();
 b15zdnd00an1n01x5 FILLER_310_1440 ();
 b15zdnd11an1n04x5 FILLER_310_1467 ();
 b15zdnd11an1n32x5 FILLER_310_1475 ();
 b15zdnd00an1n02x5 FILLER_310_1507 ();
 b15zdnd11an1n04x5 FILLER_310_1540 ();
 b15zdnd00an1n01x5 FILLER_310_1544 ();
 b15zdnd11an1n04x5 FILLER_310_1571 ();
 b15zdnd11an1n64x5 FILLER_310_1580 ();
 b15zdnd00an1n02x5 FILLER_310_1644 ();
 b15zdnd11an1n04x5 FILLER_310_1652 ();
 b15zdnd00an1n01x5 FILLER_310_1656 ();
 b15zdnd11an1n16x5 FILLER_310_1664 ();
 b15zdnd11an1n04x5 FILLER_310_1680 ();
 b15zdnd11an1n32x5 FILLER_310_1694 ();
 b15zdnd11an1n08x5 FILLER_310_1726 ();
 b15zdnd11an1n64x5 FILLER_310_1765 ();
 b15zdnd11an1n64x5 FILLER_310_1829 ();
 b15zdnd11an1n64x5 FILLER_310_1893 ();
 b15zdnd11an1n16x5 FILLER_310_1957 ();
 b15zdnd11an1n04x5 FILLER_310_1973 ();
 b15zdnd11an1n64x5 FILLER_310_1983 ();
 b15zdnd11an1n08x5 FILLER_310_2047 ();
 b15zdnd11an1n04x5 FILLER_310_2055 ();
 b15zdnd00an1n01x5 FILLER_310_2059 ();
 b15zdnd11an1n16x5 FILLER_310_2071 ();
 b15zdnd11an1n08x5 FILLER_310_2087 ();
 b15zdnd11an1n04x5 FILLER_310_2095 ();
 b15zdnd11an1n08x5 FILLER_310_2106 ();
 b15zdnd00an1n01x5 FILLER_310_2114 ();
 b15zdnd11an1n04x5 FILLER_310_2124 ();
 b15zdnd00an1n01x5 FILLER_310_2128 ();
 b15zdnd11an1n16x5 FILLER_310_2137 ();
 b15zdnd00an1n01x5 FILLER_310_2153 ();
 b15zdnd11an1n64x5 FILLER_310_2162 ();
 b15zdnd11an1n32x5 FILLER_310_2226 ();
 b15zdnd11an1n16x5 FILLER_310_2258 ();
 b15zdnd00an1n02x5 FILLER_310_2274 ();
 b15zdnd11an1n64x5 FILLER_311_0 ();
 b15zdnd11an1n64x5 FILLER_311_64 ();
 b15zdnd11an1n64x5 FILLER_311_128 ();
 b15zdnd11an1n32x5 FILLER_311_192 ();
 b15zdnd00an1n02x5 FILLER_311_224 ();
 b15zdnd11an1n04x5 FILLER_311_257 ();
 b15zdnd11an1n16x5 FILLER_311_277 ();
 b15zdnd11an1n04x5 FILLER_311_293 ();
 b15zdnd00an1n02x5 FILLER_311_297 ();
 b15zdnd11an1n32x5 FILLER_311_305 ();
 b15zdnd00an1n02x5 FILLER_311_337 ();
 b15zdnd00an1n01x5 FILLER_311_339 ();
 b15zdnd11an1n08x5 FILLER_311_347 ();
 b15zdnd00an1n01x5 FILLER_311_355 ();
 b15zdnd11an1n16x5 FILLER_311_363 ();
 b15zdnd11an1n08x5 FILLER_311_379 ();
 b15zdnd00an1n02x5 FILLER_311_387 ();
 b15zdnd00an1n01x5 FILLER_311_389 ();
 b15zdnd11an1n04x5 FILLER_311_396 ();
 b15zdnd11an1n04x5 FILLER_311_405 ();
 b15zdnd00an1n01x5 FILLER_311_409 ();
 b15zdnd11an1n16x5 FILLER_311_415 ();
 b15zdnd00an1n01x5 FILLER_311_431 ();
 b15zdnd11an1n32x5 FILLER_311_436 ();
 b15zdnd00an1n02x5 FILLER_311_468 ();
 b15zdnd11an1n64x5 FILLER_311_480 ();
 b15zdnd11an1n16x5 FILLER_311_544 ();
 b15zdnd11an1n04x5 FILLER_311_560 ();
 b15zdnd00an1n02x5 FILLER_311_564 ();
 b15zdnd00an1n01x5 FILLER_311_566 ();
 b15zdnd11an1n04x5 FILLER_311_581 ();
 b15zdnd11an1n64x5 FILLER_311_611 ();
 b15zdnd11an1n16x5 FILLER_311_675 ();
 b15zdnd11an1n08x5 FILLER_311_691 ();
 b15zdnd11an1n04x5 FILLER_311_699 ();
 b15zdnd11an1n32x5 FILLER_311_723 ();
 b15zdnd00an1n02x5 FILLER_311_755 ();
 b15zdnd11an1n64x5 FILLER_311_769 ();
 b15zdnd11an1n64x5 FILLER_311_833 ();
 b15zdnd11an1n64x5 FILLER_311_897 ();
 b15zdnd11an1n64x5 FILLER_311_961 ();
 b15zdnd11an1n08x5 FILLER_311_1025 ();
 b15zdnd11an1n04x5 FILLER_311_1033 ();
 b15zdnd11an1n64x5 FILLER_311_1046 ();
 b15zdnd11an1n32x5 FILLER_311_1110 ();
 b15zdnd11an1n08x5 FILLER_311_1142 ();
 b15zdnd11an1n32x5 FILLER_311_1155 ();
 b15zdnd11an1n04x5 FILLER_311_1187 ();
 b15zdnd00an1n01x5 FILLER_311_1191 ();
 b15zdnd11an1n64x5 FILLER_311_1202 ();
 b15zdnd11an1n32x5 FILLER_311_1266 ();
 b15zdnd11an1n32x5 FILLER_311_1318 ();
 b15zdnd11an1n04x5 FILLER_311_1350 ();
 b15zdnd00an1n02x5 FILLER_311_1354 ();
 b15zdnd00an1n01x5 FILLER_311_1356 ();
 b15zdnd11an1n32x5 FILLER_311_1369 ();
 b15zdnd11an1n04x5 FILLER_311_1401 ();
 b15zdnd11an1n32x5 FILLER_311_1414 ();
 b15zdnd11an1n08x5 FILLER_311_1446 ();
 b15zdnd11an1n04x5 FILLER_311_1454 ();
 b15zdnd00an1n01x5 FILLER_311_1458 ();
 b15zdnd11an1n04x5 FILLER_311_1468 ();
 b15zdnd11an1n04x5 FILLER_311_1490 ();
 b15zdnd11an1n16x5 FILLER_311_1501 ();
 b15zdnd11an1n08x5 FILLER_311_1517 ();
 b15zdnd00an1n01x5 FILLER_311_1525 ();
 b15zdnd11an1n04x5 FILLER_311_1544 ();
 b15zdnd00an1n02x5 FILLER_311_1548 ();
 b15zdnd11an1n04x5 FILLER_311_1570 ();
 b15zdnd00an1n01x5 FILLER_311_1574 ();
 b15zdnd11an1n08x5 FILLER_311_1580 ();
 b15zdnd00an1n02x5 FILLER_311_1588 ();
 b15zdnd11an1n04x5 FILLER_311_1608 ();
 b15zdnd11an1n16x5 FILLER_311_1617 ();
 b15zdnd11an1n08x5 FILLER_311_1633 ();
 b15zdnd11an1n04x5 FILLER_311_1641 ();
 b15zdnd00an1n02x5 FILLER_311_1645 ();
 b15zdnd00an1n01x5 FILLER_311_1647 ();
 b15zdnd11an1n16x5 FILLER_311_1655 ();
 b15zdnd11an1n04x5 FILLER_311_1671 ();
 b15zdnd11an1n16x5 FILLER_311_1682 ();
 b15zdnd11an1n08x5 FILLER_311_1698 ();
 b15zdnd00an1n02x5 FILLER_311_1706 ();
 b15zdnd00an1n01x5 FILLER_311_1708 ();
 b15zdnd11an1n04x5 FILLER_311_1715 ();
 b15zdnd00an1n02x5 FILLER_311_1719 ();
 b15zdnd00an1n01x5 FILLER_311_1721 ();
 b15zdnd11an1n04x5 FILLER_311_1738 ();
 b15zdnd11an1n32x5 FILLER_311_1755 ();
 b15zdnd11an1n16x5 FILLER_311_1787 ();
 b15zdnd11an1n04x5 FILLER_311_1803 ();
 b15zdnd00an1n02x5 FILLER_311_1807 ();
 b15zdnd11an1n32x5 FILLER_311_1829 ();
 b15zdnd11an1n08x5 FILLER_311_1861 ();
 b15zdnd00an1n01x5 FILLER_311_1869 ();
 b15zdnd11an1n64x5 FILLER_311_1890 ();
 b15zdnd11an1n04x5 FILLER_311_1954 ();
 b15zdnd00an1n02x5 FILLER_311_1958 ();
 b15zdnd00an1n01x5 FILLER_311_1960 ();
 b15zdnd11an1n64x5 FILLER_311_1981 ();
 b15zdnd11an1n64x5 FILLER_311_2045 ();
 b15zdnd11an1n64x5 FILLER_311_2109 ();
 b15zdnd11an1n64x5 FILLER_311_2173 ();
 b15zdnd11an1n32x5 FILLER_311_2237 ();
 b15zdnd11an1n08x5 FILLER_311_2269 ();
 b15zdnd11an1n04x5 FILLER_311_2277 ();
 b15zdnd00an1n02x5 FILLER_311_2281 ();
 b15zdnd00an1n01x5 FILLER_311_2283 ();
 b15zdnd11an1n64x5 FILLER_312_8 ();
 b15zdnd11an1n64x5 FILLER_312_72 ();
 b15zdnd11an1n64x5 FILLER_312_136 ();
 b15zdnd11an1n16x5 FILLER_312_200 ();
 b15zdnd00an1n02x5 FILLER_312_216 ();
 b15zdnd11an1n04x5 FILLER_312_225 ();
 b15zdnd11an1n08x5 FILLER_312_245 ();
 b15zdnd11an1n04x5 FILLER_312_253 ();
 b15zdnd00an1n01x5 FILLER_312_257 ();
 b15zdnd11an1n16x5 FILLER_312_276 ();
 b15zdnd11an1n08x5 FILLER_312_292 ();
 b15zdnd00an1n02x5 FILLER_312_300 ();
 b15zdnd00an1n01x5 FILLER_312_302 ();
 b15zdnd11an1n08x5 FILLER_312_310 ();
 b15zdnd11an1n04x5 FILLER_312_318 ();
 b15zdnd11an1n32x5 FILLER_312_327 ();
 b15zdnd11an1n16x5 FILLER_312_359 ();
 b15zdnd11an1n16x5 FILLER_312_385 ();
 b15zdnd11an1n08x5 FILLER_312_401 ();
 b15zdnd11an1n04x5 FILLER_312_409 ();
 b15zdnd11an1n04x5 FILLER_312_418 ();
 b15zdnd00an1n02x5 FILLER_312_422 ();
 b15zdnd00an1n01x5 FILLER_312_424 ();
 b15zdnd11an1n16x5 FILLER_312_437 ();
 b15zdnd11an1n08x5 FILLER_312_453 ();
 b15zdnd11an1n04x5 FILLER_312_461 ();
 b15zdnd00an1n01x5 FILLER_312_465 ();
 b15zdnd11an1n64x5 FILLER_312_478 ();
 b15zdnd11an1n16x5 FILLER_312_542 ();
 b15zdnd00an1n02x5 FILLER_312_558 ();
 b15zdnd11an1n04x5 FILLER_312_570 ();
 b15zdnd11an1n16x5 FILLER_312_600 ();
 b15zdnd11an1n08x5 FILLER_312_616 ();
 b15zdnd11an1n08x5 FILLER_312_650 ();
 b15zdnd00an1n02x5 FILLER_312_658 ();
 b15zdnd11an1n32x5 FILLER_312_680 ();
 b15zdnd11an1n04x5 FILLER_312_712 ();
 b15zdnd00an1n02x5 FILLER_312_716 ();
 b15zdnd11an1n16x5 FILLER_312_726 ();
 b15zdnd00an1n02x5 FILLER_312_742 ();
 b15zdnd11an1n04x5 FILLER_312_753 ();
 b15zdnd11an1n16x5 FILLER_312_769 ();
 b15zdnd11an1n04x5 FILLER_312_785 ();
 b15zdnd00an1n01x5 FILLER_312_789 ();
 b15zdnd11an1n64x5 FILLER_312_805 ();
 b15zdnd11an1n32x5 FILLER_312_869 ();
 b15zdnd11an1n16x5 FILLER_312_901 ();
 b15zdnd11an1n04x5 FILLER_312_917 ();
 b15zdnd00an1n01x5 FILLER_312_921 ();
 b15zdnd11an1n04x5 FILLER_312_937 ();
 b15zdnd00an1n02x5 FILLER_312_941 ();
 b15zdnd11an1n04x5 FILLER_312_946 ();
 b15zdnd11an1n64x5 FILLER_312_970 ();
 b15zdnd11an1n64x5 FILLER_312_1034 ();
 b15zdnd11an1n32x5 FILLER_312_1098 ();
 b15zdnd11an1n16x5 FILLER_312_1130 ();
 b15zdnd11an1n08x5 FILLER_312_1146 ();
 b15zdnd11an1n04x5 FILLER_312_1154 ();
 b15zdnd11an1n32x5 FILLER_312_1162 ();
 b15zdnd11an1n08x5 FILLER_312_1194 ();
 b15zdnd11an1n04x5 FILLER_312_1202 ();
 b15zdnd11an1n32x5 FILLER_312_1215 ();
 b15zdnd11an1n16x5 FILLER_312_1247 ();
 b15zdnd00an1n02x5 FILLER_312_1263 ();
 b15zdnd11an1n08x5 FILLER_312_1285 ();
 b15zdnd11an1n04x5 FILLER_312_1293 ();
 b15zdnd11an1n32x5 FILLER_312_1302 ();
 b15zdnd11an1n08x5 FILLER_312_1334 ();
 b15zdnd00an1n02x5 FILLER_312_1342 ();
 b15zdnd11an1n04x5 FILLER_312_1364 ();
 b15zdnd11an1n64x5 FILLER_312_1372 ();
 b15zdnd11an1n32x5 FILLER_312_1436 ();
 b15zdnd00an1n02x5 FILLER_312_1468 ();
 b15zdnd00an1n01x5 FILLER_312_1470 ();
 b15zdnd11an1n08x5 FILLER_312_1475 ();
 b15zdnd00an1n01x5 FILLER_312_1483 ();
 b15zdnd11an1n08x5 FILLER_312_1496 ();
 b15zdnd11an1n04x5 FILLER_312_1504 ();
 b15zdnd00an1n01x5 FILLER_312_1508 ();
 b15zdnd11an1n64x5 FILLER_312_1521 ();
 b15zdnd11an1n16x5 FILLER_312_1585 ();
 b15zdnd11an1n08x5 FILLER_312_1601 ();
 b15zdnd11an1n04x5 FILLER_312_1614 ();
 b15zdnd11an1n16x5 FILLER_312_1630 ();
 b15zdnd11an1n04x5 FILLER_312_1646 ();
 b15zdnd00an1n02x5 FILLER_312_1650 ();
 b15zdnd11an1n16x5 FILLER_312_1658 ();
 b15zdnd11an1n08x5 FILLER_312_1674 ();
 b15zdnd11an1n04x5 FILLER_312_1682 ();
 b15zdnd00an1n02x5 FILLER_312_1686 ();
 b15zdnd11an1n08x5 FILLER_312_1693 ();
 b15zdnd11an1n04x5 FILLER_312_1701 ();
 b15zdnd00an1n02x5 FILLER_312_1705 ();
 b15zdnd11an1n08x5 FILLER_312_1711 ();
 b15zdnd00an1n01x5 FILLER_312_1719 ();
 b15zdnd11an1n64x5 FILLER_312_1752 ();
 b15zdnd11an1n64x5 FILLER_312_1816 ();
 b15zdnd11an1n64x5 FILLER_312_1880 ();
 b15zdnd11an1n64x5 FILLER_312_1944 ();
 b15zdnd11an1n64x5 FILLER_312_2008 ();
 b15zdnd11an1n64x5 FILLER_312_2072 ();
 b15zdnd11an1n16x5 FILLER_312_2136 ();
 b15zdnd00an1n02x5 FILLER_312_2152 ();
 b15zdnd11an1n64x5 FILLER_312_2162 ();
 b15zdnd11an1n16x5 FILLER_312_2226 ();
 b15zdnd11an1n08x5 FILLER_312_2242 ();
 b15zdnd11an1n04x5 FILLER_312_2250 ();
 b15zdnd00an1n02x5 FILLER_312_2274 ();
 b15zdnd11an1n64x5 FILLER_313_0 ();
 b15zdnd11an1n64x5 FILLER_313_64 ();
 b15zdnd11an1n64x5 FILLER_313_128 ();
 b15zdnd11an1n32x5 FILLER_313_192 ();
 b15zdnd11an1n04x5 FILLER_313_224 ();
 b15zdnd11an1n64x5 FILLER_313_235 ();
 b15zdnd11an1n04x5 FILLER_313_299 ();
 b15zdnd00an1n02x5 FILLER_313_303 ();
 b15zdnd00an1n01x5 FILLER_313_305 ();
 b15zdnd11an1n64x5 FILLER_313_315 ();
 b15zdnd11an1n32x5 FILLER_313_379 ();
 b15zdnd11an1n04x5 FILLER_313_411 ();
 b15zdnd11an1n08x5 FILLER_313_424 ();
 b15zdnd11an1n08x5 FILLER_313_437 ();
 b15zdnd11an1n04x5 FILLER_313_445 ();
 b15zdnd00an1n01x5 FILLER_313_449 ();
 b15zdnd11an1n16x5 FILLER_313_476 ();
 b15zdnd00an1n02x5 FILLER_313_492 ();
 b15zdnd00an1n01x5 FILLER_313_494 ();
 b15zdnd11an1n08x5 FILLER_313_502 ();
 b15zdnd00an1n01x5 FILLER_313_510 ();
 b15zdnd11an1n04x5 FILLER_313_524 ();
 b15zdnd11an1n04x5 FILLER_313_535 ();
 b15zdnd00an1n01x5 FILLER_313_539 ();
 b15zdnd11an1n04x5 FILLER_313_554 ();
 b15zdnd11an1n04x5 FILLER_313_584 ();
 b15zdnd11an1n04x5 FILLER_313_603 ();
 b15zdnd11an1n64x5 FILLER_313_638 ();
 b15zdnd11an1n32x5 FILLER_313_702 ();
 b15zdnd11an1n04x5 FILLER_313_734 ();
 b15zdnd00an1n02x5 FILLER_313_738 ();
 b15zdnd00an1n01x5 FILLER_313_740 ();
 b15zdnd11an1n04x5 FILLER_313_750 ();
 b15zdnd11an1n16x5 FILLER_313_763 ();
 b15zdnd11an1n08x5 FILLER_313_779 ();
 b15zdnd11an1n04x5 FILLER_313_787 ();
 b15zdnd00an1n02x5 FILLER_313_791 ();
 b15zdnd00an1n01x5 FILLER_313_793 ();
 b15zdnd11an1n16x5 FILLER_313_812 ();
 b15zdnd11an1n04x5 FILLER_313_828 ();
 b15zdnd11an1n16x5 FILLER_313_839 ();
 b15zdnd11an1n08x5 FILLER_313_855 ();
 b15zdnd11an1n04x5 FILLER_313_863 ();
 b15zdnd00an1n02x5 FILLER_313_867 ();
 b15zdnd11an1n04x5 FILLER_313_892 ();
 b15zdnd11an1n16x5 FILLER_313_901 ();
 b15zdnd11an1n04x5 FILLER_313_917 ();
 b15zdnd00an1n02x5 FILLER_313_921 ();
 b15zdnd11an1n64x5 FILLER_313_954 ();
 b15zdnd11an1n32x5 FILLER_313_1018 ();
 b15zdnd11an1n16x5 FILLER_313_1050 ();
 b15zdnd11an1n08x5 FILLER_313_1066 ();
 b15zdnd11an1n04x5 FILLER_313_1074 ();
 b15zdnd11an1n64x5 FILLER_313_1087 ();
 b15zdnd11an1n16x5 FILLER_313_1151 ();
 b15zdnd11an1n08x5 FILLER_313_1167 ();
 b15zdnd00an1n02x5 FILLER_313_1175 ();
 b15zdnd11an1n64x5 FILLER_313_1198 ();
 b15zdnd11an1n64x5 FILLER_313_1262 ();
 b15zdnd11an1n64x5 FILLER_313_1326 ();
 b15zdnd11an1n64x5 FILLER_313_1390 ();
 b15zdnd11an1n04x5 FILLER_313_1454 ();
 b15zdnd00an1n01x5 FILLER_313_1458 ();
 b15zdnd11an1n64x5 FILLER_313_1485 ();
 b15zdnd11an1n64x5 FILLER_313_1549 ();
 b15zdnd11an1n64x5 FILLER_313_1613 ();
 b15zdnd11an1n64x5 FILLER_313_1677 ();
 b15zdnd11an1n08x5 FILLER_313_1741 ();
 b15zdnd11an1n04x5 FILLER_313_1749 ();
 b15zdnd00an1n02x5 FILLER_313_1753 ();
 b15zdnd00an1n01x5 FILLER_313_1755 ();
 b15zdnd11an1n04x5 FILLER_313_1766 ();
 b15zdnd11an1n32x5 FILLER_313_1786 ();
 b15zdnd00an1n01x5 FILLER_313_1818 ();
 b15zdnd11an1n04x5 FILLER_313_1831 ();
 b15zdnd00an1n02x5 FILLER_313_1835 ();
 b15zdnd11an1n64x5 FILLER_313_1857 ();
 b15zdnd11an1n08x5 FILLER_313_1921 ();
 b15zdnd11an1n04x5 FILLER_313_1929 ();
 b15zdnd00an1n02x5 FILLER_313_1933 ();
 b15zdnd11an1n04x5 FILLER_313_1955 ();
 b15zdnd11an1n64x5 FILLER_313_1985 ();
 b15zdnd11an1n64x5 FILLER_313_2049 ();
 b15zdnd11an1n32x5 FILLER_313_2113 ();
 b15zdnd11an1n08x5 FILLER_313_2145 ();
 b15zdnd00an1n01x5 FILLER_313_2153 ();
 b15zdnd11an1n08x5 FILLER_313_2174 ();
 b15zdnd11an1n04x5 FILLER_313_2182 ();
 b15zdnd11an1n16x5 FILLER_313_2206 ();
 b15zdnd11an1n08x5 FILLER_313_2222 ();
 b15zdnd00an1n02x5 FILLER_313_2230 ();
 b15zdnd00an1n01x5 FILLER_313_2232 ();
 b15zdnd11an1n04x5 FILLER_313_2253 ();
 b15zdnd11an1n16x5 FILLER_313_2265 ();
 b15zdnd00an1n02x5 FILLER_313_2281 ();
 b15zdnd00an1n01x5 FILLER_313_2283 ();
 b15zdnd11an1n64x5 FILLER_314_8 ();
 b15zdnd11an1n64x5 FILLER_314_72 ();
 b15zdnd11an1n64x5 FILLER_314_136 ();
 b15zdnd11an1n32x5 FILLER_314_200 ();
 b15zdnd11an1n04x5 FILLER_314_232 ();
 b15zdnd00an1n01x5 FILLER_314_236 ();
 b15zdnd11an1n32x5 FILLER_314_245 ();
 b15zdnd00an1n02x5 FILLER_314_277 ();
 b15zdnd11an1n04x5 FILLER_314_285 ();
 b15zdnd11an1n32x5 FILLER_314_296 ();
 b15zdnd11an1n16x5 FILLER_314_328 ();
 b15zdnd11an1n08x5 FILLER_314_344 ();
 b15zdnd11an1n16x5 FILLER_314_357 ();
 b15zdnd11an1n04x5 FILLER_314_373 ();
 b15zdnd11an1n32x5 FILLER_314_386 ();
 b15zdnd00an1n02x5 FILLER_314_418 ();
 b15zdnd00an1n01x5 FILLER_314_420 ();
 b15zdnd11an1n08x5 FILLER_314_433 ();
 b15zdnd11an1n32x5 FILLER_314_445 ();
 b15zdnd11an1n16x5 FILLER_314_477 ();
 b15zdnd00an1n02x5 FILLER_314_493 ();
 b15zdnd00an1n01x5 FILLER_314_495 ();
 b15zdnd11an1n08x5 FILLER_314_501 ();
 b15zdnd11an1n04x5 FILLER_314_509 ();
 b15zdnd11an1n32x5 FILLER_314_519 ();
 b15zdnd11an1n08x5 FILLER_314_551 ();
 b15zdnd00an1n02x5 FILLER_314_559 ();
 b15zdnd00an1n01x5 FILLER_314_561 ();
 b15zdnd11an1n16x5 FILLER_314_571 ();
 b15zdnd11an1n08x5 FILLER_314_587 ();
 b15zdnd00an1n01x5 FILLER_314_595 ();
 b15zdnd11an1n64x5 FILLER_314_628 ();
 b15zdnd11an1n16x5 FILLER_314_692 ();
 b15zdnd11an1n08x5 FILLER_314_708 ();
 b15zdnd00an1n02x5 FILLER_314_716 ();
 b15zdnd11an1n64x5 FILLER_314_726 ();
 b15zdnd11an1n08x5 FILLER_314_790 ();
 b15zdnd11an1n04x5 FILLER_314_798 ();
 b15zdnd11an1n04x5 FILLER_314_833 ();
 b15zdnd11an1n32x5 FILLER_314_852 ();
 b15zdnd11an1n04x5 FILLER_314_884 ();
 b15zdnd00an1n02x5 FILLER_314_888 ();
 b15zdnd11an1n32x5 FILLER_314_910 ();
 b15zdnd00an1n02x5 FILLER_314_942 ();
 b15zdnd11an1n64x5 FILLER_314_949 ();
 b15zdnd11an1n64x5 FILLER_314_1013 ();
 b15zdnd11an1n32x5 FILLER_314_1077 ();
 b15zdnd11an1n08x5 FILLER_314_1109 ();
 b15zdnd11an1n04x5 FILLER_314_1117 ();
 b15zdnd11an1n64x5 FILLER_314_1130 ();
 b15zdnd11an1n08x5 FILLER_314_1194 ();
 b15zdnd11an1n04x5 FILLER_314_1202 ();
 b15zdnd00an1n02x5 FILLER_314_1206 ();
 b15zdnd11an1n04x5 FILLER_314_1213 ();
 b15zdnd11an1n04x5 FILLER_314_1237 ();
 b15zdnd11an1n04x5 FILLER_314_1263 ();
 b15zdnd11an1n16x5 FILLER_314_1282 ();
 b15zdnd00an1n01x5 FILLER_314_1298 ();
 b15zdnd11an1n32x5 FILLER_314_1303 ();
 b15zdnd11an1n32x5 FILLER_314_1346 ();
 b15zdnd11an1n16x5 FILLER_314_1378 ();
 b15zdnd11an1n04x5 FILLER_314_1394 ();
 b15zdnd11an1n32x5 FILLER_314_1418 ();
 b15zdnd11an1n08x5 FILLER_314_1450 ();
 b15zdnd11an1n04x5 FILLER_314_1458 ();
 b15zdnd11an1n32x5 FILLER_314_1482 ();
 b15zdnd11an1n08x5 FILLER_314_1514 ();
 b15zdnd00an1n01x5 FILLER_314_1522 ();
 b15zdnd11an1n16x5 FILLER_314_1532 ();
 b15zdnd11an1n04x5 FILLER_314_1548 ();
 b15zdnd00an1n02x5 FILLER_314_1552 ();
 b15zdnd00an1n01x5 FILLER_314_1554 ();
 b15zdnd11an1n04x5 FILLER_314_1563 ();
 b15zdnd00an1n01x5 FILLER_314_1567 ();
 b15zdnd11an1n16x5 FILLER_314_1580 ();
 b15zdnd11an1n08x5 FILLER_314_1608 ();
 b15zdnd00an1n02x5 FILLER_314_1616 ();
 b15zdnd11an1n32x5 FILLER_314_1625 ();
 b15zdnd11an1n16x5 FILLER_314_1657 ();
 b15zdnd00an1n02x5 FILLER_314_1673 ();
 b15zdnd00an1n01x5 FILLER_314_1675 ();
 b15zdnd11an1n16x5 FILLER_314_1681 ();
 b15zdnd11an1n08x5 FILLER_314_1697 ();
 b15zdnd00an1n02x5 FILLER_314_1705 ();
 b15zdnd11an1n32x5 FILLER_314_1712 ();
 b15zdnd11an1n16x5 FILLER_314_1744 ();
 b15zdnd11an1n04x5 FILLER_314_1760 ();
 b15zdnd00an1n01x5 FILLER_314_1764 ();
 b15zdnd11an1n16x5 FILLER_314_1783 ();
 b15zdnd11an1n04x5 FILLER_314_1799 ();
 b15zdnd11an1n04x5 FILLER_314_1812 ();
 b15zdnd00an1n02x5 FILLER_314_1816 ();
 b15zdnd11an1n64x5 FILLER_314_1840 ();
 b15zdnd11an1n64x5 FILLER_314_1904 ();
 b15zdnd11an1n64x5 FILLER_314_1968 ();
 b15zdnd11an1n64x5 FILLER_314_2032 ();
 b15zdnd11an1n32x5 FILLER_314_2096 ();
 b15zdnd11an1n16x5 FILLER_314_2128 ();
 b15zdnd11an1n08x5 FILLER_314_2144 ();
 b15zdnd00an1n02x5 FILLER_314_2152 ();
 b15zdnd11an1n04x5 FILLER_314_2162 ();
 b15zdnd00an1n02x5 FILLER_314_2166 ();
 b15zdnd11an1n32x5 FILLER_314_2194 ();
 b15zdnd00an1n01x5 FILLER_314_2226 ();
 b15zdnd11an1n04x5 FILLER_314_2232 ();
 b15zdnd11an1n16x5 FILLER_314_2241 ();
 b15zdnd11an1n08x5 FILLER_314_2261 ();
 b15zdnd11an1n04x5 FILLER_314_2269 ();
 b15zdnd00an1n02x5 FILLER_314_2273 ();
 b15zdnd00an1n01x5 FILLER_314_2275 ();
 b15zdnd11an1n64x5 FILLER_315_0 ();
 b15zdnd11an1n64x5 FILLER_315_64 ();
 b15zdnd11an1n64x5 FILLER_315_128 ();
 b15zdnd11an1n32x5 FILLER_315_192 ();
 b15zdnd11an1n04x5 FILLER_315_224 ();
 b15zdnd00an1n01x5 FILLER_315_228 ();
 b15zdnd11an1n16x5 FILLER_315_234 ();
 b15zdnd11an1n04x5 FILLER_315_250 ();
 b15zdnd11an1n08x5 FILLER_315_266 ();
 b15zdnd11an1n04x5 FILLER_315_274 ();
 b15zdnd00an1n02x5 FILLER_315_278 ();
 b15zdnd00an1n01x5 FILLER_315_280 ();
 b15zdnd11an1n08x5 FILLER_315_287 ();
 b15zdnd11an1n04x5 FILLER_315_295 ();
 b15zdnd00an1n02x5 FILLER_315_299 ();
 b15zdnd11an1n32x5 FILLER_315_305 ();
 b15zdnd11an1n08x5 FILLER_315_337 ();
 b15zdnd11an1n04x5 FILLER_315_345 ();
 b15zdnd00an1n02x5 FILLER_315_349 ();
 b15zdnd00an1n01x5 FILLER_315_351 ();
 b15zdnd11an1n08x5 FILLER_315_358 ();
 b15zdnd00an1n02x5 FILLER_315_366 ();
 b15zdnd00an1n01x5 FILLER_315_368 ();
 b15zdnd11an1n04x5 FILLER_315_383 ();
 b15zdnd00an1n01x5 FILLER_315_387 ();
 b15zdnd11an1n08x5 FILLER_315_393 ();
 b15zdnd11an1n04x5 FILLER_315_401 ();
 b15zdnd00an1n01x5 FILLER_315_405 ();
 b15zdnd11an1n64x5 FILLER_315_411 ();
 b15zdnd11an1n16x5 FILLER_315_475 ();
 b15zdnd00an1n02x5 FILLER_315_491 ();
 b15zdnd00an1n01x5 FILLER_315_493 ();
 b15zdnd11an1n16x5 FILLER_315_501 ();
 b15zdnd11an1n04x5 FILLER_315_517 ();
 b15zdnd11an1n32x5 FILLER_315_547 ();
 b15zdnd11an1n08x5 FILLER_315_579 ();
 b15zdnd00an1n02x5 FILLER_315_587 ();
 b15zdnd00an1n01x5 FILLER_315_589 ();
 b15zdnd11an1n04x5 FILLER_315_622 ();
 b15zdnd11an1n64x5 FILLER_315_652 ();
 b15zdnd11an1n16x5 FILLER_315_716 ();
 b15zdnd11an1n08x5 FILLER_315_732 ();
 b15zdnd00an1n02x5 FILLER_315_740 ();
 b15zdnd11an1n04x5 FILLER_315_767 ();
 b15zdnd11an1n32x5 FILLER_315_792 ();
 b15zdnd11an1n08x5 FILLER_315_824 ();
 b15zdnd00an1n02x5 FILLER_315_832 ();
 b15zdnd11an1n32x5 FILLER_315_842 ();
 b15zdnd11an1n16x5 FILLER_315_874 ();
 b15zdnd11an1n04x5 FILLER_315_890 ();
 b15zdnd11an1n32x5 FILLER_315_900 ();
 b15zdnd11an1n08x5 FILLER_315_932 ();
 b15zdnd11an1n04x5 FILLER_315_940 ();
 b15zdnd00an1n01x5 FILLER_315_944 ();
 b15zdnd11an1n08x5 FILLER_315_949 ();
 b15zdnd11an1n04x5 FILLER_315_957 ();
 b15zdnd00an1n02x5 FILLER_315_961 ();
 b15zdnd11an1n04x5 FILLER_315_974 ();
 b15zdnd11an1n16x5 FILLER_315_987 ();
 b15zdnd11an1n04x5 FILLER_315_1003 ();
 b15zdnd11an1n16x5 FILLER_315_1027 ();
 b15zdnd00an1n02x5 FILLER_315_1043 ();
 b15zdnd11an1n08x5 FILLER_315_1065 ();
 b15zdnd11an1n04x5 FILLER_315_1073 ();
 b15zdnd00an1n02x5 FILLER_315_1077 ();
 b15zdnd11an1n16x5 FILLER_315_1099 ();
 b15zdnd11an1n04x5 FILLER_315_1115 ();
 b15zdnd00an1n02x5 FILLER_315_1119 ();
 b15zdnd00an1n01x5 FILLER_315_1121 ();
 b15zdnd11an1n64x5 FILLER_315_1127 ();
 b15zdnd11an1n32x5 FILLER_315_1191 ();
 b15zdnd11an1n08x5 FILLER_315_1223 ();
 b15zdnd11an1n04x5 FILLER_315_1231 ();
 b15zdnd00an1n02x5 FILLER_315_1235 ();
 b15zdnd11an1n64x5 FILLER_315_1263 ();
 b15zdnd11an1n64x5 FILLER_315_1327 ();
 b15zdnd11an1n16x5 FILLER_315_1391 ();
 b15zdnd00an1n01x5 FILLER_315_1407 ();
 b15zdnd11an1n16x5 FILLER_315_1413 ();
 b15zdnd00an1n02x5 FILLER_315_1429 ();
 b15zdnd11an1n64x5 FILLER_315_1435 ();
 b15zdnd11an1n64x5 FILLER_315_1499 ();
 b15zdnd11an1n08x5 FILLER_315_1572 ();
 b15zdnd11an1n16x5 FILLER_315_1589 ();
 b15zdnd11an1n08x5 FILLER_315_1605 ();
 b15zdnd00an1n01x5 FILLER_315_1613 ();
 b15zdnd11an1n16x5 FILLER_315_1626 ();
 b15zdnd11an1n08x5 FILLER_315_1642 ();
 b15zdnd00an1n02x5 FILLER_315_1650 ();
 b15zdnd00an1n01x5 FILLER_315_1652 ();
 b15zdnd11an1n04x5 FILLER_315_1662 ();
 b15zdnd11an1n16x5 FILLER_315_1678 ();
 b15zdnd11an1n08x5 FILLER_315_1694 ();
 b15zdnd11an1n04x5 FILLER_315_1702 ();
 b15zdnd11an1n08x5 FILLER_315_1715 ();
 b15zdnd00an1n02x5 FILLER_315_1723 ();
 b15zdnd00an1n01x5 FILLER_315_1725 ();
 b15zdnd11an1n64x5 FILLER_315_1744 ();
 b15zdnd11an1n64x5 FILLER_315_1808 ();
 b15zdnd11an1n32x5 FILLER_315_1872 ();
 b15zdnd11an1n04x5 FILLER_315_1904 ();
 b15zdnd11an1n64x5 FILLER_315_1920 ();
 b15zdnd11an1n16x5 FILLER_315_1984 ();
 b15zdnd00an1n02x5 FILLER_315_2000 ();
 b15zdnd00an1n01x5 FILLER_315_2002 ();
 b15zdnd11an1n16x5 FILLER_315_2009 ();
 b15zdnd11an1n08x5 FILLER_315_2025 ();
 b15zdnd00an1n02x5 FILLER_315_2033 ();
 b15zdnd00an1n01x5 FILLER_315_2035 ();
 b15zdnd11an1n04x5 FILLER_315_2051 ();
 b15zdnd11an1n64x5 FILLER_315_2066 ();
 b15zdnd11an1n16x5 FILLER_315_2130 ();
 b15zdnd11an1n08x5 FILLER_315_2146 ();
 b15zdnd11an1n04x5 FILLER_315_2154 ();
 b15zdnd00an1n02x5 FILLER_315_2158 ();
 b15zdnd11an1n64x5 FILLER_315_2169 ();
 b15zdnd11an1n32x5 FILLER_315_2233 ();
 b15zdnd11an1n16x5 FILLER_315_2265 ();
 b15zdnd00an1n02x5 FILLER_315_2281 ();
 b15zdnd00an1n01x5 FILLER_315_2283 ();
 b15zdnd11an1n64x5 FILLER_316_8 ();
 b15zdnd11an1n64x5 FILLER_316_72 ();
 b15zdnd11an1n64x5 FILLER_316_136 ();
 b15zdnd11an1n32x5 FILLER_316_200 ();
 b15zdnd00an1n01x5 FILLER_316_232 ();
 b15zdnd11an1n32x5 FILLER_316_241 ();
 b15zdnd11an1n16x5 FILLER_316_273 ();
 b15zdnd11an1n08x5 FILLER_316_289 ();
 b15zdnd11an1n04x5 FILLER_316_297 ();
 b15zdnd00an1n02x5 FILLER_316_301 ();
 b15zdnd11an1n16x5 FILLER_316_309 ();
 b15zdnd11an1n04x5 FILLER_316_325 ();
 b15zdnd00an1n01x5 FILLER_316_329 ();
 b15zdnd11an1n04x5 FILLER_316_346 ();
 b15zdnd11an1n16x5 FILLER_316_357 ();
 b15zdnd00an1n02x5 FILLER_316_373 ();
 b15zdnd00an1n01x5 FILLER_316_375 ();
 b15zdnd11an1n64x5 FILLER_316_397 ();
 b15zdnd11an1n16x5 FILLER_316_461 ();
 b15zdnd11an1n64x5 FILLER_316_484 ();
 b15zdnd11an1n16x5 FILLER_316_548 ();
 b15zdnd11an1n08x5 FILLER_316_564 ();
 b15zdnd00an1n02x5 FILLER_316_572 ();
 b15zdnd00an1n01x5 FILLER_316_574 ();
 b15zdnd11an1n16x5 FILLER_316_607 ();
 b15zdnd00an1n01x5 FILLER_316_623 ();
 b15zdnd11an1n04x5 FILLER_316_650 ();
 b15zdnd11an1n16x5 FILLER_316_674 ();
 b15zdnd00an1n02x5 FILLER_316_690 ();
 b15zdnd00an1n01x5 FILLER_316_692 ();
 b15zdnd00an1n02x5 FILLER_316_716 ();
 b15zdnd11an1n32x5 FILLER_316_726 ();
 b15zdnd11an1n04x5 FILLER_316_758 ();
 b15zdnd11an1n64x5 FILLER_316_784 ();
 b15zdnd11an1n16x5 FILLER_316_848 ();
 b15zdnd00an1n02x5 FILLER_316_864 ();
 b15zdnd00an1n01x5 FILLER_316_866 ();
 b15zdnd11an1n64x5 FILLER_316_893 ();
 b15zdnd11an1n64x5 FILLER_316_957 ();
 b15zdnd11an1n16x5 FILLER_316_1021 ();
 b15zdnd11an1n08x5 FILLER_316_1037 ();
 b15zdnd00an1n02x5 FILLER_316_1045 ();
 b15zdnd00an1n01x5 FILLER_316_1047 ();
 b15zdnd11an1n64x5 FILLER_316_1059 ();
 b15zdnd00an1n02x5 FILLER_316_1123 ();
 b15zdnd11an1n08x5 FILLER_316_1145 ();
 b15zdnd00an1n02x5 FILLER_316_1153 ();
 b15zdnd00an1n01x5 FILLER_316_1155 ();
 b15zdnd11an1n08x5 FILLER_316_1161 ();
 b15zdnd11an1n04x5 FILLER_316_1169 ();
 b15zdnd00an1n02x5 FILLER_316_1173 ();
 b15zdnd11an1n64x5 FILLER_316_1181 ();
 b15zdnd11an1n64x5 FILLER_316_1245 ();
 b15zdnd00an1n02x5 FILLER_316_1309 ();
 b15zdnd11an1n32x5 FILLER_316_1319 ();
 b15zdnd11an1n16x5 FILLER_316_1351 ();
 b15zdnd00an1n02x5 FILLER_316_1367 ();
 b15zdnd00an1n01x5 FILLER_316_1369 ();
 b15zdnd11an1n64x5 FILLER_316_1390 ();
 b15zdnd11an1n64x5 FILLER_316_1454 ();
 b15zdnd11an1n32x5 FILLER_316_1518 ();
 b15zdnd11an1n08x5 FILLER_316_1550 ();
 b15zdnd00an1n01x5 FILLER_316_1558 ();
 b15zdnd11an1n16x5 FILLER_316_1570 ();
 b15zdnd00an1n01x5 FILLER_316_1586 ();
 b15zdnd11an1n04x5 FILLER_316_1618 ();
 b15zdnd11an1n04x5 FILLER_316_1627 ();
 b15zdnd11an1n16x5 FILLER_316_1635 ();
 b15zdnd11an1n04x5 FILLER_316_1651 ();
 b15zdnd00an1n01x5 FILLER_316_1655 ();
 b15zdnd11an1n08x5 FILLER_316_1663 ();
 b15zdnd11an1n08x5 FILLER_316_1681 ();
 b15zdnd11an1n04x5 FILLER_316_1689 ();
 b15zdnd11an1n04x5 FILLER_316_1705 ();
 b15zdnd11an1n16x5 FILLER_316_1713 ();
 b15zdnd00an1n01x5 FILLER_316_1729 ();
 b15zdnd11an1n64x5 FILLER_316_1756 ();
 b15zdnd11an1n64x5 FILLER_316_1820 ();
 b15zdnd11an1n32x5 FILLER_316_1884 ();
 b15zdnd11an1n16x5 FILLER_316_1916 ();
 b15zdnd00an1n02x5 FILLER_316_1932 ();
 b15zdnd00an1n01x5 FILLER_316_1934 ();
 b15zdnd11an1n32x5 FILLER_316_1940 ();
 b15zdnd11an1n04x5 FILLER_316_1972 ();
 b15zdnd00an1n02x5 FILLER_316_1976 ();
 b15zdnd11an1n16x5 FILLER_316_1992 ();
 b15zdnd11an1n08x5 FILLER_316_2008 ();
 b15zdnd11an1n04x5 FILLER_316_2016 ();
 b15zdnd00an1n02x5 FILLER_316_2020 ();
 b15zdnd11an1n32x5 FILLER_316_2053 ();
 b15zdnd11an1n04x5 FILLER_316_2085 ();
 b15zdnd00an1n02x5 FILLER_316_2089 ();
 b15zdnd00an1n01x5 FILLER_316_2091 ();
 b15zdnd11an1n32x5 FILLER_316_2099 ();
 b15zdnd11an1n16x5 FILLER_316_2131 ();
 b15zdnd11an1n04x5 FILLER_316_2147 ();
 b15zdnd00an1n02x5 FILLER_316_2151 ();
 b15zdnd00an1n01x5 FILLER_316_2153 ();
 b15zdnd00an1n02x5 FILLER_316_2162 ();
 b15zdnd11an1n64x5 FILLER_316_2185 ();
 b15zdnd11an1n16x5 FILLER_316_2249 ();
 b15zdnd11an1n08x5 FILLER_316_2265 ();
 b15zdnd00an1n02x5 FILLER_316_2273 ();
 b15zdnd00an1n01x5 FILLER_316_2275 ();
 b15zdnd11an1n64x5 FILLER_317_0 ();
 b15zdnd11an1n64x5 FILLER_317_64 ();
 b15zdnd11an1n64x5 FILLER_317_128 ();
 b15zdnd11an1n64x5 FILLER_317_192 ();
 b15zdnd11an1n64x5 FILLER_317_256 ();
 b15zdnd11an1n64x5 FILLER_317_320 ();
 b15zdnd11an1n04x5 FILLER_317_384 ();
 b15zdnd00an1n02x5 FILLER_317_388 ();
 b15zdnd00an1n01x5 FILLER_317_390 ();
 b15zdnd11an1n64x5 FILLER_317_397 ();
 b15zdnd11an1n16x5 FILLER_317_461 ();
 b15zdnd11an1n08x5 FILLER_317_477 ();
 b15zdnd11an1n64x5 FILLER_317_497 ();
 b15zdnd11an1n32x5 FILLER_317_561 ();
 b15zdnd11an1n08x5 FILLER_317_593 ();
 b15zdnd11an1n64x5 FILLER_317_617 ();
 b15zdnd11an1n16x5 FILLER_317_681 ();
 b15zdnd11an1n08x5 FILLER_317_697 ();
 b15zdnd00an1n02x5 FILLER_317_705 ();
 b15zdnd00an1n01x5 FILLER_317_707 ();
 b15zdnd11an1n32x5 FILLER_317_717 ();
 b15zdnd11an1n16x5 FILLER_317_749 ();
 b15zdnd11an1n04x5 FILLER_317_765 ();
 b15zdnd00an1n02x5 FILLER_317_769 ();
 b15zdnd00an1n01x5 FILLER_317_771 ();
 b15zdnd11an1n32x5 FILLER_317_797 ();
 b15zdnd11an1n16x5 FILLER_317_829 ();
 b15zdnd11an1n08x5 FILLER_317_845 ();
 b15zdnd00an1n02x5 FILLER_317_853 ();
 b15zdnd11an1n04x5 FILLER_317_864 ();
 b15zdnd11an1n16x5 FILLER_317_891 ();
 b15zdnd11an1n08x5 FILLER_317_907 ();
 b15zdnd00an1n02x5 FILLER_317_915 ();
 b15zdnd00an1n01x5 FILLER_317_917 ();
 b15zdnd11an1n16x5 FILLER_317_927 ();
 b15zdnd11an1n08x5 FILLER_317_943 ();
 b15zdnd00an1n01x5 FILLER_317_951 ();
 b15zdnd11an1n16x5 FILLER_317_961 ();
 b15zdnd00an1n02x5 FILLER_317_977 ();
 b15zdnd11an1n64x5 FILLER_317_999 ();
 b15zdnd11an1n64x5 FILLER_317_1063 ();
 b15zdnd00an1n02x5 FILLER_317_1127 ();
 b15zdnd11an1n08x5 FILLER_317_1133 ();
 b15zdnd11an1n04x5 FILLER_317_1141 ();
 b15zdnd00an1n02x5 FILLER_317_1145 ();
 b15zdnd00an1n01x5 FILLER_317_1147 ();
 b15zdnd11an1n04x5 FILLER_317_1152 ();
 b15zdnd00an1n02x5 FILLER_317_1156 ();
 b15zdnd11an1n08x5 FILLER_317_1178 ();
 b15zdnd11an1n04x5 FILLER_317_1186 ();
 b15zdnd00an1n01x5 FILLER_317_1190 ();
 b15zdnd11an1n08x5 FILLER_317_1199 ();
 b15zdnd00an1n01x5 FILLER_317_1207 ();
 b15zdnd11an1n64x5 FILLER_317_1212 ();
 b15zdnd11an1n16x5 FILLER_317_1276 ();
 b15zdnd00an1n01x5 FILLER_317_1292 ();
 b15zdnd11an1n16x5 FILLER_317_1313 ();
 b15zdnd11an1n08x5 FILLER_317_1329 ();
 b15zdnd00an1n02x5 FILLER_317_1337 ();
 b15zdnd11an1n08x5 FILLER_317_1348 ();
 b15zdnd00an1n02x5 FILLER_317_1356 ();
 b15zdnd00an1n01x5 FILLER_317_1358 ();
 b15zdnd11an1n04x5 FILLER_317_1368 ();
 b15zdnd11an1n64x5 FILLER_317_1377 ();
 b15zdnd11an1n64x5 FILLER_317_1441 ();
 b15zdnd11an1n04x5 FILLER_317_1505 ();
 b15zdnd00an1n02x5 FILLER_317_1509 ();
 b15zdnd00an1n01x5 FILLER_317_1511 ();
 b15zdnd11an1n64x5 FILLER_317_1523 ();
 b15zdnd11an1n64x5 FILLER_317_1587 ();
 b15zdnd11an1n04x5 FILLER_317_1651 ();
 b15zdnd00an1n02x5 FILLER_317_1655 ();
 b15zdnd00an1n01x5 FILLER_317_1657 ();
 b15zdnd11an1n04x5 FILLER_317_1664 ();
 b15zdnd00an1n02x5 FILLER_317_1668 ();
 b15zdnd00an1n01x5 FILLER_317_1670 ();
 b15zdnd11an1n64x5 FILLER_317_1689 ();
 b15zdnd11an1n64x5 FILLER_317_1753 ();
 b15zdnd11an1n32x5 FILLER_317_1817 ();
 b15zdnd11an1n16x5 FILLER_317_1849 ();
 b15zdnd11an1n04x5 FILLER_317_1865 ();
 b15zdnd11an1n16x5 FILLER_317_1875 ();
 b15zdnd11an1n04x5 FILLER_317_1897 ();
 b15zdnd11an1n08x5 FILLER_317_1922 ();
 b15zdnd00an1n02x5 FILLER_317_1930 ();
 b15zdnd11an1n08x5 FILLER_317_1948 ();
 b15zdnd11an1n04x5 FILLER_317_1956 ();
 b15zdnd00an1n01x5 FILLER_317_1960 ();
 b15zdnd11an1n08x5 FILLER_317_1965 ();
 b15zdnd11an1n04x5 FILLER_317_1973 ();
 b15zdnd11an1n04x5 FILLER_317_1981 ();
 b15zdnd11an1n08x5 FILLER_317_1994 ();
 b15zdnd11an1n04x5 FILLER_317_2002 ();
 b15zdnd11an1n16x5 FILLER_317_2013 ();
 b15zdnd11an1n08x5 FILLER_317_2029 ();
 b15zdnd11an1n04x5 FILLER_317_2037 ();
 b15zdnd00an1n01x5 FILLER_317_2041 ();
 b15zdnd11an1n08x5 FILLER_317_2046 ();
 b15zdnd11an1n04x5 FILLER_317_2054 ();
 b15zdnd00an1n02x5 FILLER_317_2058 ();
 b15zdnd11an1n32x5 FILLER_317_2064 ();
 b15zdnd00an1n02x5 FILLER_317_2096 ();
 b15zdnd11an1n16x5 FILLER_317_2113 ();
 b15zdnd11an1n08x5 FILLER_317_2129 ();
 b15zdnd11an1n64x5 FILLER_317_2163 ();
 b15zdnd11an1n04x5 FILLER_317_2227 ();
 b15zdnd00an1n01x5 FILLER_317_2231 ();
 b15zdnd11an1n32x5 FILLER_317_2238 ();
 b15zdnd11an1n08x5 FILLER_317_2270 ();
 b15zdnd11an1n04x5 FILLER_317_2278 ();
 b15zdnd00an1n02x5 FILLER_317_2282 ();
 b15zdnd11an1n64x5 FILLER_318_8 ();
 b15zdnd11an1n64x5 FILLER_318_72 ();
 b15zdnd11an1n64x5 FILLER_318_136 ();
 b15zdnd11an1n32x5 FILLER_318_200 ();
 b15zdnd11an1n08x5 FILLER_318_232 ();
 b15zdnd00an1n01x5 FILLER_318_240 ();
 b15zdnd11an1n04x5 FILLER_318_245 ();
 b15zdnd11an1n64x5 FILLER_318_256 ();
 b15zdnd11an1n64x5 FILLER_318_320 ();
 b15zdnd11an1n16x5 FILLER_318_384 ();
 b15zdnd11an1n08x5 FILLER_318_400 ();
 b15zdnd00an1n02x5 FILLER_318_408 ();
 b15zdnd11an1n04x5 FILLER_318_415 ();
 b15zdnd11an1n16x5 FILLER_318_427 ();
 b15zdnd11an1n08x5 FILLER_318_443 ();
 b15zdnd00an1n02x5 FILLER_318_451 ();
 b15zdnd11an1n32x5 FILLER_318_458 ();
 b15zdnd11an1n16x5 FILLER_318_490 ();
 b15zdnd11an1n04x5 FILLER_318_511 ();
 b15zdnd11an1n32x5 FILLER_318_520 ();
 b15zdnd11an1n04x5 FILLER_318_552 ();
 b15zdnd00an1n02x5 FILLER_318_556 ();
 b15zdnd11an1n04x5 FILLER_318_567 ();
 b15zdnd11an1n08x5 FILLER_318_577 ();
 b15zdnd11an1n04x5 FILLER_318_585 ();
 b15zdnd11an1n08x5 FILLER_318_594 ();
 b15zdnd00an1n02x5 FILLER_318_602 ();
 b15zdnd00an1n01x5 FILLER_318_604 ();
 b15zdnd11an1n64x5 FILLER_318_636 ();
 b15zdnd11an1n08x5 FILLER_318_700 ();
 b15zdnd00an1n01x5 FILLER_318_708 ();
 b15zdnd11an1n04x5 FILLER_318_713 ();
 b15zdnd00an1n01x5 FILLER_318_717 ();
 b15zdnd11an1n32x5 FILLER_318_726 ();
 b15zdnd11an1n16x5 FILLER_318_758 ();
 b15zdnd11an1n08x5 FILLER_318_774 ();
 b15zdnd11an1n64x5 FILLER_318_786 ();
 b15zdnd11an1n32x5 FILLER_318_850 ();
 b15zdnd11an1n16x5 FILLER_318_882 ();
 b15zdnd00an1n01x5 FILLER_318_898 ();
 b15zdnd11an1n16x5 FILLER_318_903 ();
 b15zdnd00an1n01x5 FILLER_318_919 ();
 b15zdnd11an1n64x5 FILLER_318_940 ();
 b15zdnd11an1n64x5 FILLER_318_1004 ();
 b15zdnd11an1n08x5 FILLER_318_1068 ();
 b15zdnd11an1n04x5 FILLER_318_1076 ();
 b15zdnd00an1n01x5 FILLER_318_1080 ();
 b15zdnd11an1n64x5 FILLER_318_1090 ();
 b15zdnd11an1n64x5 FILLER_318_1154 ();
 b15zdnd11an1n16x5 FILLER_318_1218 ();
 b15zdnd11an1n08x5 FILLER_318_1234 ();
 b15zdnd00an1n01x5 FILLER_318_1242 ();
 b15zdnd11an1n16x5 FILLER_318_1252 ();
 b15zdnd11an1n08x5 FILLER_318_1274 ();
 b15zdnd11an1n04x5 FILLER_318_1286 ();
 b15zdnd11an1n64x5 FILLER_318_1295 ();
 b15zdnd11an1n32x5 FILLER_318_1359 ();
 b15zdnd11an1n16x5 FILLER_318_1391 ();
 b15zdnd11an1n08x5 FILLER_318_1407 ();
 b15zdnd11an1n04x5 FILLER_318_1415 ();
 b15zdnd00an1n01x5 FILLER_318_1419 ();
 b15zdnd11an1n64x5 FILLER_318_1429 ();
 b15zdnd11an1n16x5 FILLER_318_1493 ();
 b15zdnd11an1n04x5 FILLER_318_1529 ();
 b15zdnd11an1n32x5 FILLER_318_1559 ();
 b15zdnd11an1n16x5 FILLER_318_1591 ();
 b15zdnd00an1n02x5 FILLER_318_1607 ();
 b15zdnd11an1n32x5 FILLER_318_1623 ();
 b15zdnd11an1n08x5 FILLER_318_1655 ();
 b15zdnd11an1n64x5 FILLER_318_1675 ();
 b15zdnd11an1n64x5 FILLER_318_1739 ();
 b15zdnd11an1n08x5 FILLER_318_1803 ();
 b15zdnd11an1n32x5 FILLER_318_1831 ();
 b15zdnd11an1n16x5 FILLER_318_1863 ();
 b15zdnd11an1n04x5 FILLER_318_1889 ();
 b15zdnd11an1n08x5 FILLER_318_1901 ();
 b15zdnd00an1n02x5 FILLER_318_1909 ();
 b15zdnd00an1n01x5 FILLER_318_1911 ();
 b15zdnd11an1n16x5 FILLER_318_1925 ();
 b15zdnd11an1n04x5 FILLER_318_1953 ();
 b15zdnd00an1n01x5 FILLER_318_1957 ();
 b15zdnd11an1n04x5 FILLER_318_1979 ();
 b15zdnd11an1n32x5 FILLER_318_1993 ();
 b15zdnd11an1n08x5 FILLER_318_2025 ();
 b15zdnd11an1n04x5 FILLER_318_2033 ();
 b15zdnd00an1n01x5 FILLER_318_2037 ();
 b15zdnd11an1n16x5 FILLER_318_2045 ();
 b15zdnd11an1n04x5 FILLER_318_2085 ();
 b15zdnd11an1n16x5 FILLER_318_2100 ();
 b15zdnd11an1n04x5 FILLER_318_2116 ();
 b15zdnd00an1n02x5 FILLER_318_2152 ();
 b15zdnd11an1n16x5 FILLER_318_2162 ();
 b15zdnd11an1n04x5 FILLER_318_2178 ();
 b15zdnd00an1n02x5 FILLER_318_2182 ();
 b15zdnd11an1n04x5 FILLER_318_2215 ();
 b15zdnd00an1n02x5 FILLER_318_2219 ();
 b15zdnd00an1n01x5 FILLER_318_2221 ();
 b15zdnd11an1n04x5 FILLER_318_2242 ();
 b15zdnd11an1n04x5 FILLER_318_2251 ();
 b15zdnd11an1n08x5 FILLER_318_2262 ();
 b15zdnd11an1n04x5 FILLER_318_2270 ();
 b15zdnd00an1n02x5 FILLER_318_2274 ();
 b15zdnd11an1n64x5 FILLER_319_0 ();
 b15zdnd11an1n64x5 FILLER_319_64 ();
 b15zdnd11an1n64x5 FILLER_319_128 ();
 b15zdnd11an1n32x5 FILLER_319_192 ();
 b15zdnd11an1n08x5 FILLER_319_224 ();
 b15zdnd00an1n01x5 FILLER_319_232 ();
 b15zdnd11an1n16x5 FILLER_319_237 ();
 b15zdnd11an1n08x5 FILLER_319_253 ();
 b15zdnd11an1n32x5 FILLER_319_265 ();
 b15zdnd11an1n08x5 FILLER_319_297 ();
 b15zdnd00an1n02x5 FILLER_319_305 ();
 b15zdnd00an1n01x5 FILLER_319_307 ();
 b15zdnd11an1n16x5 FILLER_319_324 ();
 b15zdnd00an1n02x5 FILLER_319_340 ();
 b15zdnd00an1n01x5 FILLER_319_342 ();
 b15zdnd11an1n08x5 FILLER_319_360 ();
 b15zdnd11an1n04x5 FILLER_319_368 ();
 b15zdnd11an1n16x5 FILLER_319_377 ();
 b15zdnd00an1n02x5 FILLER_319_393 ();
 b15zdnd00an1n01x5 FILLER_319_395 ();
 b15zdnd11an1n08x5 FILLER_319_422 ();
 b15zdnd11an1n04x5 FILLER_319_430 ();
 b15zdnd11an1n08x5 FILLER_319_441 ();
 b15zdnd00an1n02x5 FILLER_319_449 ();
 b15zdnd00an1n01x5 FILLER_319_451 ();
 b15zdnd11an1n16x5 FILLER_319_457 ();
 b15zdnd11an1n04x5 FILLER_319_473 ();
 b15zdnd11an1n16x5 FILLER_319_481 ();
 b15zdnd11an1n08x5 FILLER_319_497 ();
 b15zdnd00an1n02x5 FILLER_319_505 ();
 b15zdnd00an1n01x5 FILLER_319_507 ();
 b15zdnd11an1n04x5 FILLER_319_521 ();
 b15zdnd11an1n04x5 FILLER_319_546 ();
 b15zdnd11an1n64x5 FILLER_319_570 ();
 b15zdnd11an1n16x5 FILLER_319_634 ();
 b15zdnd11an1n08x5 FILLER_319_650 ();
 b15zdnd00an1n02x5 FILLER_319_658 ();
 b15zdnd00an1n01x5 FILLER_319_660 ();
 b15zdnd11an1n08x5 FILLER_319_687 ();
 b15zdnd11an1n04x5 FILLER_319_695 ();
 b15zdnd11an1n32x5 FILLER_319_724 ();
 b15zdnd11an1n16x5 FILLER_319_756 ();
 b15zdnd11an1n08x5 FILLER_319_772 ();
 b15zdnd00an1n02x5 FILLER_319_780 ();
 b15zdnd11an1n16x5 FILLER_319_797 ();
 b15zdnd00an1n02x5 FILLER_319_813 ();
 b15zdnd11an1n32x5 FILLER_319_835 ();
 b15zdnd11an1n08x5 FILLER_319_867 ();
 b15zdnd11an1n04x5 FILLER_319_875 ();
 b15zdnd00an1n02x5 FILLER_319_879 ();
 b15zdnd11an1n32x5 FILLER_319_885 ();
 b15zdnd00an1n02x5 FILLER_319_917 ();
 b15zdnd11an1n64x5 FILLER_319_928 ();
 b15zdnd11an1n32x5 FILLER_319_992 ();
 b15zdnd00an1n01x5 FILLER_319_1024 ();
 b15zdnd11an1n32x5 FILLER_319_1034 ();
 b15zdnd11an1n08x5 FILLER_319_1066 ();
 b15zdnd11an1n04x5 FILLER_319_1074 ();
 b15zdnd00an1n01x5 FILLER_319_1078 ();
 b15zdnd11an1n64x5 FILLER_319_1084 ();
 b15zdnd11an1n64x5 FILLER_319_1148 ();
 b15zdnd11an1n64x5 FILLER_319_1212 ();
 b15zdnd11an1n32x5 FILLER_319_1276 ();
 b15zdnd11an1n16x5 FILLER_319_1308 ();
 b15zdnd11an1n08x5 FILLER_319_1324 ();
 b15zdnd11an1n04x5 FILLER_319_1332 ();
 b15zdnd00an1n01x5 FILLER_319_1336 ();
 b15zdnd11an1n64x5 FILLER_319_1342 ();
 b15zdnd11an1n32x5 FILLER_319_1406 ();
 b15zdnd11an1n08x5 FILLER_319_1458 ();
 b15zdnd11an1n04x5 FILLER_319_1466 ();
 b15zdnd00an1n01x5 FILLER_319_1470 ();
 b15zdnd11an1n04x5 FILLER_319_1476 ();
 b15zdnd11an1n64x5 FILLER_319_1493 ();
 b15zdnd11an1n64x5 FILLER_319_1557 ();
 b15zdnd11an1n64x5 FILLER_319_1621 ();
 b15zdnd11an1n64x5 FILLER_319_1685 ();
 b15zdnd11an1n08x5 FILLER_319_1749 ();
 b15zdnd11an1n04x5 FILLER_319_1757 ();
 b15zdnd00an1n02x5 FILLER_319_1761 ();
 b15zdnd00an1n01x5 FILLER_319_1763 ();
 b15zdnd11an1n64x5 FILLER_319_1784 ();
 b15zdnd11an1n04x5 FILLER_319_1848 ();
 b15zdnd00an1n02x5 FILLER_319_1852 ();
 b15zdnd11an1n32x5 FILLER_319_1873 ();
 b15zdnd11an1n08x5 FILLER_319_1905 ();
 b15zdnd00an1n02x5 FILLER_319_1913 ();
 b15zdnd11an1n64x5 FILLER_319_1922 ();
 b15zdnd11an1n16x5 FILLER_319_1986 ();
 b15zdnd11an1n08x5 FILLER_319_2002 ();
 b15zdnd11an1n04x5 FILLER_319_2019 ();
 b15zdnd11an1n04x5 FILLER_319_2035 ();
 b15zdnd11an1n32x5 FILLER_319_2046 ();
 b15zdnd00an1n02x5 FILLER_319_2078 ();
 b15zdnd00an1n01x5 FILLER_319_2080 ();
 b15zdnd11an1n32x5 FILLER_319_2098 ();
 b15zdnd11an1n04x5 FILLER_319_2130 ();
 b15zdnd00an1n01x5 FILLER_319_2134 ();
 b15zdnd11an1n16x5 FILLER_319_2145 ();
 b15zdnd00an1n02x5 FILLER_319_2161 ();
 b15zdnd00an1n01x5 FILLER_319_2163 ();
 b15zdnd11an1n32x5 FILLER_319_2190 ();
 b15zdnd11an1n04x5 FILLER_319_2222 ();
 b15zdnd00an1n01x5 FILLER_319_2226 ();
 b15zdnd11an1n16x5 FILLER_319_2232 ();
 b15zdnd11an1n08x5 FILLER_319_2248 ();
 b15zdnd11an1n04x5 FILLER_319_2256 ();
 b15zdnd00an1n01x5 FILLER_319_2260 ();
 b15zdnd00an1n02x5 FILLER_319_2281 ();
 b15zdnd00an1n01x5 FILLER_319_2283 ();
 b15zdnd11an1n64x5 FILLER_320_8 ();
 b15zdnd11an1n64x5 FILLER_320_72 ();
 b15zdnd11an1n64x5 FILLER_320_136 ();
 b15zdnd11an1n16x5 FILLER_320_200 ();
 b15zdnd11an1n04x5 FILLER_320_216 ();
 b15zdnd00an1n01x5 FILLER_320_220 ();
 b15zdnd11an1n16x5 FILLER_320_233 ();
 b15zdnd11an1n04x5 FILLER_320_249 ();
 b15zdnd00an1n02x5 FILLER_320_253 ();
 b15zdnd00an1n01x5 FILLER_320_255 ();
 b15zdnd11an1n08x5 FILLER_320_266 ();
 b15zdnd11an1n04x5 FILLER_320_274 ();
 b15zdnd00an1n02x5 FILLER_320_278 ();
 b15zdnd00an1n01x5 FILLER_320_280 ();
 b15zdnd11an1n16x5 FILLER_320_288 ();
 b15zdnd11an1n04x5 FILLER_320_304 ();
 b15zdnd00an1n02x5 FILLER_320_308 ();
 b15zdnd00an1n01x5 FILLER_320_310 ();
 b15zdnd11an1n16x5 FILLER_320_324 ();
 b15zdnd11an1n04x5 FILLER_320_340 ();
 b15zdnd00an1n01x5 FILLER_320_344 ();
 b15zdnd11an1n04x5 FILLER_320_350 ();
 b15zdnd11an1n32x5 FILLER_320_364 ();
 b15zdnd11an1n16x5 FILLER_320_408 ();
 b15zdnd11an1n08x5 FILLER_320_424 ();
 b15zdnd00an1n01x5 FILLER_320_432 ();
 b15zdnd11an1n64x5 FILLER_320_442 ();
 b15zdnd00an1n02x5 FILLER_320_506 ();
 b15zdnd00an1n01x5 FILLER_320_508 ();
 b15zdnd11an1n04x5 FILLER_320_515 ();
 b15zdnd11an1n08x5 FILLER_320_532 ();
 b15zdnd11an1n04x5 FILLER_320_540 ();
 b15zdnd00an1n02x5 FILLER_320_544 ();
 b15zdnd00an1n01x5 FILLER_320_546 ();
 b15zdnd11an1n16x5 FILLER_320_561 ();
 b15zdnd11an1n04x5 FILLER_320_577 ();
 b15zdnd00an1n02x5 FILLER_320_581 ();
 b15zdnd11an1n04x5 FILLER_320_604 ();
 b15zdnd11an1n04x5 FILLER_320_634 ();
 b15zdnd11an1n32x5 FILLER_320_658 ();
 b15zdnd11an1n08x5 FILLER_320_690 ();
 b15zdnd11an1n04x5 FILLER_320_698 ();
 b15zdnd00an1n02x5 FILLER_320_702 ();
 b15zdnd00an1n01x5 FILLER_320_704 ();
 b15zdnd00an1n02x5 FILLER_320_715 ();
 b15zdnd00an1n01x5 FILLER_320_717 ();
 b15zdnd11an1n32x5 FILLER_320_726 ();
 b15zdnd11an1n16x5 FILLER_320_758 ();
 b15zdnd11an1n08x5 FILLER_320_774 ();
 b15zdnd00an1n02x5 FILLER_320_782 ();
 b15zdnd11an1n08x5 FILLER_320_815 ();
 b15zdnd11an1n04x5 FILLER_320_823 ();
 b15zdnd00an1n02x5 FILLER_320_827 ();
 b15zdnd11an1n04x5 FILLER_320_834 ();
 b15zdnd11an1n32x5 FILLER_320_843 ();
 b15zdnd11an1n16x5 FILLER_320_875 ();
 b15zdnd11an1n04x5 FILLER_320_891 ();
 b15zdnd11an1n16x5 FILLER_320_935 ();
 b15zdnd11an1n08x5 FILLER_320_951 ();
 b15zdnd00an1n02x5 FILLER_320_959 ();
 b15zdnd11an1n32x5 FILLER_320_973 ();
 b15zdnd11an1n16x5 FILLER_320_1005 ();
 b15zdnd11an1n04x5 FILLER_320_1021 ();
 b15zdnd00an1n01x5 FILLER_320_1025 ();
 b15zdnd11an1n04x5 FILLER_320_1046 ();
 b15zdnd11an1n08x5 FILLER_320_1070 ();
 b15zdnd00an1n02x5 FILLER_320_1078 ();
 b15zdnd11an1n64x5 FILLER_320_1100 ();
 b15zdnd11an1n16x5 FILLER_320_1164 ();
 b15zdnd11an1n08x5 FILLER_320_1180 ();
 b15zdnd11an1n04x5 FILLER_320_1188 ();
 b15zdnd00an1n01x5 FILLER_320_1192 ();
 b15zdnd11an1n04x5 FILLER_320_1199 ();
 b15zdnd00an1n01x5 FILLER_320_1203 ();
 b15zdnd11an1n32x5 FILLER_320_1211 ();
 b15zdnd11an1n08x5 FILLER_320_1243 ();
 b15zdnd11an1n04x5 FILLER_320_1251 ();
 b15zdnd00an1n01x5 FILLER_320_1255 ();
 b15zdnd11an1n04x5 FILLER_320_1261 ();
 b15zdnd00an1n02x5 FILLER_320_1265 ();
 b15zdnd11an1n32x5 FILLER_320_1287 ();
 b15zdnd11an1n08x5 FILLER_320_1319 ();
 b15zdnd00an1n02x5 FILLER_320_1327 ();
 b15zdnd00an1n01x5 FILLER_320_1329 ();
 b15zdnd11an1n16x5 FILLER_320_1350 ();
 b15zdnd11an1n08x5 FILLER_320_1366 ();
 b15zdnd00an1n02x5 FILLER_320_1374 ();
 b15zdnd11an1n64x5 FILLER_320_1380 ();
 b15zdnd11an1n32x5 FILLER_320_1444 ();
 b15zdnd11an1n08x5 FILLER_320_1476 ();
 b15zdnd00an1n02x5 FILLER_320_1484 ();
 b15zdnd11an1n04x5 FILLER_320_1495 ();
 b15zdnd11an1n64x5 FILLER_320_1503 ();
 b15zdnd11an1n64x5 FILLER_320_1567 ();
 b15zdnd11an1n64x5 FILLER_320_1631 ();
 b15zdnd11an1n32x5 FILLER_320_1695 ();
 b15zdnd11an1n08x5 FILLER_320_1727 ();
 b15zdnd11an1n32x5 FILLER_320_1745 ();
 b15zdnd11an1n64x5 FILLER_320_1797 ();
 b15zdnd11an1n32x5 FILLER_320_1861 ();
 b15zdnd11an1n08x5 FILLER_320_1893 ();
 b15zdnd11an1n04x5 FILLER_320_1901 ();
 b15zdnd00an1n02x5 FILLER_320_1905 ();
 b15zdnd11an1n32x5 FILLER_320_1916 ();
 b15zdnd11an1n16x5 FILLER_320_1948 ();
 b15zdnd11an1n08x5 FILLER_320_1964 ();
 b15zdnd11an1n04x5 FILLER_320_1972 ();
 b15zdnd00an1n02x5 FILLER_320_1976 ();
 b15zdnd00an1n01x5 FILLER_320_1978 ();
 b15zdnd11an1n04x5 FILLER_320_1989 ();
 b15zdnd11an1n08x5 FILLER_320_1999 ();
 b15zdnd11an1n04x5 FILLER_320_2007 ();
 b15zdnd00an1n02x5 FILLER_320_2011 ();
 b15zdnd00an1n01x5 FILLER_320_2013 ();
 b15zdnd11an1n64x5 FILLER_320_2019 ();
 b15zdnd11an1n32x5 FILLER_320_2083 ();
 b15zdnd11an1n16x5 FILLER_320_2115 ();
 b15zdnd11an1n04x5 FILLER_320_2131 ();
 b15zdnd11an1n08x5 FILLER_320_2145 ();
 b15zdnd00an1n01x5 FILLER_320_2153 ();
 b15zdnd00an1n02x5 FILLER_320_2162 ();
 b15zdnd00an1n01x5 FILLER_320_2164 ();
 b15zdnd11an1n64x5 FILLER_320_2188 ();
 b15zdnd11an1n16x5 FILLER_320_2252 ();
 b15zdnd11an1n08x5 FILLER_320_2268 ();
 b15zdnd11an1n64x5 FILLER_321_0 ();
 b15zdnd11an1n64x5 FILLER_321_64 ();
 b15zdnd11an1n64x5 FILLER_321_128 ();
 b15zdnd11an1n16x5 FILLER_321_192 ();
 b15zdnd00an1n02x5 FILLER_321_208 ();
 b15zdnd00an1n01x5 FILLER_321_210 ();
 b15zdnd11an1n04x5 FILLER_321_231 ();
 b15zdnd11an1n04x5 FILLER_321_266 ();
 b15zdnd11an1n08x5 FILLER_321_276 ();
 b15zdnd11an1n04x5 FILLER_321_296 ();
 b15zdnd00an1n02x5 FILLER_321_300 ();
 b15zdnd00an1n01x5 FILLER_321_302 ();
 b15zdnd11an1n04x5 FILLER_321_309 ();
 b15zdnd11an1n32x5 FILLER_321_320 ();
 b15zdnd11an1n16x5 FILLER_321_352 ();
 b15zdnd11an1n08x5 FILLER_321_368 ();
 b15zdnd00an1n02x5 FILLER_321_376 ();
 b15zdnd11an1n16x5 FILLER_321_382 ();
 b15zdnd11an1n08x5 FILLER_321_398 ();
 b15zdnd11an1n04x5 FILLER_321_406 ();
 b15zdnd11an1n64x5 FILLER_321_415 ();
 b15zdnd11an1n16x5 FILLER_321_479 ();
 b15zdnd11an1n04x5 FILLER_321_495 ();
 b15zdnd00an1n02x5 FILLER_321_499 ();
 b15zdnd00an1n01x5 FILLER_321_501 ();
 b15zdnd11an1n64x5 FILLER_321_509 ();
 b15zdnd11an1n64x5 FILLER_321_573 ();
 b15zdnd11an1n64x5 FILLER_321_637 ();
 b15zdnd11an1n64x5 FILLER_321_701 ();
 b15zdnd11an1n32x5 FILLER_321_765 ();
 b15zdnd11an1n16x5 FILLER_321_797 ();
 b15zdnd11an1n08x5 FILLER_321_813 ();
 b15zdnd00an1n02x5 FILLER_321_821 ();
 b15zdnd11an1n64x5 FILLER_321_829 ();
 b15zdnd11an1n32x5 FILLER_321_893 ();
 b15zdnd11an1n16x5 FILLER_321_925 ();
 b15zdnd11an1n08x5 FILLER_321_941 ();
 b15zdnd11an1n04x5 FILLER_321_949 ();
 b15zdnd11an1n16x5 FILLER_321_973 ();
 b15zdnd11an1n04x5 FILLER_321_989 ();
 b15zdnd00an1n02x5 FILLER_321_993 ();
 b15zdnd11an1n64x5 FILLER_321_998 ();
 b15zdnd11an1n16x5 FILLER_321_1062 ();
 b15zdnd00an1n01x5 FILLER_321_1078 ();
 b15zdnd11an1n32x5 FILLER_321_1083 ();
 b15zdnd11an1n04x5 FILLER_321_1115 ();
 b15zdnd11an1n32x5 FILLER_321_1139 ();
 b15zdnd11an1n16x5 FILLER_321_1171 ();
 b15zdnd11an1n04x5 FILLER_321_1187 ();
 b15zdnd00an1n01x5 FILLER_321_1191 ();
 b15zdnd11an1n08x5 FILLER_321_1212 ();
 b15zdnd11an1n04x5 FILLER_321_1220 ();
 b15zdnd00an1n02x5 FILLER_321_1224 ();
 b15zdnd11an1n32x5 FILLER_321_1235 ();
 b15zdnd11an1n16x5 FILLER_321_1267 ();
 b15zdnd00an1n02x5 FILLER_321_1283 ();
 b15zdnd11an1n64x5 FILLER_321_1311 ();
 b15zdnd11an1n32x5 FILLER_321_1375 ();
 b15zdnd11an1n04x5 FILLER_321_1407 ();
 b15zdnd11an1n04x5 FILLER_321_1418 ();
 b15zdnd11an1n32x5 FILLER_321_1429 ();
 b15zdnd11an1n16x5 FILLER_321_1461 ();
 b15zdnd00an1n02x5 FILLER_321_1477 ();
 b15zdnd00an1n01x5 FILLER_321_1479 ();
 b15zdnd11an1n64x5 FILLER_321_1496 ();
 b15zdnd11an1n16x5 FILLER_321_1560 ();
 b15zdnd00an1n02x5 FILLER_321_1576 ();
 b15zdnd11an1n32x5 FILLER_321_1610 ();
 b15zdnd00an1n02x5 FILLER_321_1642 ();
 b15zdnd00an1n01x5 FILLER_321_1644 ();
 b15zdnd11an1n64x5 FILLER_321_1665 ();
 b15zdnd11an1n64x5 FILLER_321_1729 ();
 b15zdnd11an1n32x5 FILLER_321_1793 ();
 b15zdnd11an1n16x5 FILLER_321_1825 ();
 b15zdnd11an1n08x5 FILLER_321_1841 ();
 b15zdnd11an1n08x5 FILLER_321_1854 ();
 b15zdnd00an1n02x5 FILLER_321_1862 ();
 b15zdnd00an1n01x5 FILLER_321_1864 ();
 b15zdnd11an1n08x5 FILLER_321_1877 ();
 b15zdnd11an1n04x5 FILLER_321_1885 ();
 b15zdnd11an1n64x5 FILLER_321_1896 ();
 b15zdnd11an1n64x5 FILLER_321_1960 ();
 b15zdnd11an1n16x5 FILLER_321_2029 ();
 b15zdnd11an1n08x5 FILLER_321_2045 ();
 b15zdnd11an1n04x5 FILLER_321_2053 ();
 b15zdnd00an1n02x5 FILLER_321_2057 ();
 b15zdnd11an1n16x5 FILLER_321_2064 ();
 b15zdnd11an1n08x5 FILLER_321_2080 ();
 b15zdnd00an1n02x5 FILLER_321_2088 ();
 b15zdnd00an1n01x5 FILLER_321_2090 ();
 b15zdnd11an1n04x5 FILLER_321_2100 ();
 b15zdnd11an1n64x5 FILLER_321_2109 ();
 b15zdnd11an1n64x5 FILLER_321_2173 ();
 b15zdnd11an1n32x5 FILLER_321_2237 ();
 b15zdnd11an1n08x5 FILLER_321_2269 ();
 b15zdnd00an1n01x5 FILLER_321_2277 ();
 b15zdnd00an1n02x5 FILLER_321_2282 ();
 b15zdnd11an1n64x5 FILLER_322_8 ();
 b15zdnd11an1n64x5 FILLER_322_72 ();
 b15zdnd11an1n64x5 FILLER_322_136 ();
 b15zdnd11an1n32x5 FILLER_322_200 ();
 b15zdnd11an1n08x5 FILLER_322_232 ();
 b15zdnd00an1n02x5 FILLER_322_240 ();
 b15zdnd00an1n01x5 FILLER_322_242 ();
 b15zdnd11an1n04x5 FILLER_322_251 ();
 b15zdnd00an1n02x5 FILLER_322_255 ();
 b15zdnd00an1n01x5 FILLER_322_257 ();
 b15zdnd11an1n64x5 FILLER_322_268 ();
 b15zdnd11an1n08x5 FILLER_322_332 ();
 b15zdnd11an1n16x5 FILLER_322_357 ();
 b15zdnd00an1n02x5 FILLER_322_373 ();
 b15zdnd11an1n32x5 FILLER_322_384 ();
 b15zdnd11an1n16x5 FILLER_322_416 ();
 b15zdnd11an1n04x5 FILLER_322_432 ();
 b15zdnd00an1n01x5 FILLER_322_436 ();
 b15zdnd11an1n04x5 FILLER_322_441 ();
 b15zdnd11an1n32x5 FILLER_322_452 ();
 b15zdnd11an1n04x5 FILLER_322_484 ();
 b15zdnd00an1n02x5 FILLER_322_488 ();
 b15zdnd11an1n16x5 FILLER_322_521 ();
 b15zdnd11an1n08x5 FILLER_322_537 ();
 b15zdnd11an1n04x5 FILLER_322_545 ();
 b15zdnd00an1n02x5 FILLER_322_549 ();
 b15zdnd00an1n01x5 FILLER_322_551 ();
 b15zdnd11an1n16x5 FILLER_322_564 ();
 b15zdnd11an1n08x5 FILLER_322_580 ();
 b15zdnd00an1n01x5 FILLER_322_588 ();
 b15zdnd11an1n64x5 FILLER_322_594 ();
 b15zdnd11an1n32x5 FILLER_322_658 ();
 b15zdnd11an1n16x5 FILLER_322_690 ();
 b15zdnd11an1n08x5 FILLER_322_706 ();
 b15zdnd11an1n04x5 FILLER_322_714 ();
 b15zdnd11an1n16x5 FILLER_322_726 ();
 b15zdnd11an1n08x5 FILLER_322_742 ();
 b15zdnd00an1n01x5 FILLER_322_750 ();
 b15zdnd11an1n64x5 FILLER_322_771 ();
 b15zdnd11an1n64x5 FILLER_322_835 ();
 b15zdnd11an1n64x5 FILLER_322_899 ();
 b15zdnd11an1n16x5 FILLER_322_963 ();
 b15zdnd11an1n04x5 FILLER_322_979 ();
 b15zdnd00an1n02x5 FILLER_322_983 ();
 b15zdnd00an1n01x5 FILLER_322_985 ();
 b15zdnd11an1n64x5 FILLER_322_1006 ();
 b15zdnd11an1n32x5 FILLER_322_1070 ();
 b15zdnd11an1n16x5 FILLER_322_1102 ();
 b15zdnd11an1n08x5 FILLER_322_1118 ();
 b15zdnd11an1n04x5 FILLER_322_1126 ();
 b15zdnd00an1n02x5 FILLER_322_1130 ();
 b15zdnd00an1n01x5 FILLER_322_1132 ();
 b15zdnd11an1n16x5 FILLER_322_1138 ();
 b15zdnd00an1n02x5 FILLER_322_1154 ();
 b15zdnd11an1n16x5 FILLER_322_1165 ();
 b15zdnd11an1n08x5 FILLER_322_1181 ();
 b15zdnd11an1n04x5 FILLER_322_1189 ();
 b15zdnd00an1n02x5 FILLER_322_1193 ();
 b15zdnd11an1n32x5 FILLER_322_1200 ();
 b15zdnd11an1n16x5 FILLER_322_1232 ();
 b15zdnd11an1n08x5 FILLER_322_1248 ();
 b15zdnd11an1n04x5 FILLER_322_1256 ();
 b15zdnd00an1n02x5 FILLER_322_1260 ();
 b15zdnd11an1n32x5 FILLER_322_1266 ();
 b15zdnd11an1n04x5 FILLER_322_1298 ();
 b15zdnd11an1n04x5 FILLER_322_1322 ();
 b15zdnd11an1n04x5 FILLER_322_1334 ();
 b15zdnd00an1n02x5 FILLER_322_1338 ();
 b15zdnd00an1n01x5 FILLER_322_1340 ();
 b15zdnd11an1n32x5 FILLER_322_1345 ();
 b15zdnd11an1n16x5 FILLER_322_1377 ();
 b15zdnd11an1n08x5 FILLER_322_1393 ();
 b15zdnd11an1n04x5 FILLER_322_1401 ();
 b15zdnd00an1n02x5 FILLER_322_1405 ();
 b15zdnd11an1n04x5 FILLER_322_1416 ();
 b15zdnd11an1n04x5 FILLER_322_1429 ();
 b15zdnd11an1n64x5 FILLER_322_1441 ();
 b15zdnd11an1n16x5 FILLER_322_1505 ();
 b15zdnd11an1n08x5 FILLER_322_1521 ();
 b15zdnd11an1n04x5 FILLER_322_1529 ();
 b15zdnd11an1n64x5 FILLER_322_1542 ();
 b15zdnd11an1n32x5 FILLER_322_1606 ();
 b15zdnd11an1n16x5 FILLER_322_1638 ();
 b15zdnd00an1n02x5 FILLER_322_1654 ();
 b15zdnd11an1n32x5 FILLER_322_1666 ();
 b15zdnd11an1n16x5 FILLER_322_1698 ();
 b15zdnd00an1n02x5 FILLER_322_1714 ();
 b15zdnd11an1n04x5 FILLER_322_1732 ();
 b15zdnd11an1n04x5 FILLER_322_1753 ();
 b15zdnd00an1n01x5 FILLER_322_1757 ();
 b15zdnd11an1n32x5 FILLER_322_1778 ();
 b15zdnd11an1n16x5 FILLER_322_1810 ();
 b15zdnd11an1n04x5 FILLER_322_1826 ();
 b15zdnd11an1n04x5 FILLER_322_1856 ();
 b15zdnd11an1n04x5 FILLER_322_1879 ();
 b15zdnd00an1n02x5 FILLER_322_1883 ();
 b15zdnd00an1n01x5 FILLER_322_1885 ();
 b15zdnd11an1n32x5 FILLER_322_1895 ();
 b15zdnd00an1n01x5 FILLER_322_1927 ();
 b15zdnd11an1n16x5 FILLER_322_1932 ();
 b15zdnd11an1n04x5 FILLER_322_1948 ();
 b15zdnd11an1n04x5 FILLER_322_1957 ();
 b15zdnd11an1n04x5 FILLER_322_1981 ();
 b15zdnd11an1n32x5 FILLER_322_1992 ();
 b15zdnd11an1n16x5 FILLER_322_2024 ();
 b15zdnd11an1n08x5 FILLER_322_2040 ();
 b15zdnd11an1n04x5 FILLER_322_2048 ();
 b15zdnd00an1n01x5 FILLER_322_2052 ();
 b15zdnd11an1n04x5 FILLER_322_2060 ();
 b15zdnd11an1n04x5 FILLER_322_2090 ();
 b15zdnd11an1n04x5 FILLER_322_2103 ();
 b15zdnd00an1n02x5 FILLER_322_2107 ();
 b15zdnd11an1n32x5 FILLER_322_2114 ();
 b15zdnd11an1n08x5 FILLER_322_2146 ();
 b15zdnd11an1n16x5 FILLER_322_2162 ();
 b15zdnd11an1n08x5 FILLER_322_2178 ();
 b15zdnd00an1n02x5 FILLER_322_2186 ();
 b15zdnd00an1n01x5 FILLER_322_2188 ();
 b15zdnd11an1n04x5 FILLER_322_2221 ();
 b15zdnd11an1n04x5 FILLER_322_2231 ();
 b15zdnd00an1n01x5 FILLER_322_2235 ();
 b15zdnd11an1n04x5 FILLER_322_2240 ();
 b15zdnd11an1n16x5 FILLER_322_2249 ();
 b15zdnd11an1n08x5 FILLER_322_2265 ();
 b15zdnd00an1n02x5 FILLER_322_2273 ();
 b15zdnd00an1n01x5 FILLER_322_2275 ();
 b15zdnd11an1n64x5 FILLER_323_0 ();
 b15zdnd11an1n64x5 FILLER_323_64 ();
 b15zdnd11an1n64x5 FILLER_323_128 ();
 b15zdnd11an1n64x5 FILLER_323_192 ();
 b15zdnd11an1n64x5 FILLER_323_256 ();
 b15zdnd11an1n08x5 FILLER_323_320 ();
 b15zdnd00an1n01x5 FILLER_323_328 ();
 b15zdnd11an1n04x5 FILLER_323_334 ();
 b15zdnd11an1n16x5 FILLER_323_351 ();
 b15zdnd11an1n08x5 FILLER_323_367 ();
 b15zdnd00an1n02x5 FILLER_323_375 ();
 b15zdnd11an1n08x5 FILLER_323_387 ();
 b15zdnd11an1n04x5 FILLER_323_395 ();
 b15zdnd00an1n01x5 FILLER_323_399 ();
 b15zdnd11an1n16x5 FILLER_323_409 ();
 b15zdnd11an1n32x5 FILLER_323_431 ();
 b15zdnd11an1n08x5 FILLER_323_463 ();
 b15zdnd00an1n02x5 FILLER_323_471 ();
 b15zdnd00an1n01x5 FILLER_323_473 ();
 b15zdnd11an1n04x5 FILLER_323_483 ();
 b15zdnd11an1n04x5 FILLER_323_492 ();
 b15zdnd11an1n32x5 FILLER_323_508 ();
 b15zdnd11an1n08x5 FILLER_323_540 ();
 b15zdnd11an1n04x5 FILLER_323_548 ();
 b15zdnd00an1n02x5 FILLER_323_552 ();
 b15zdnd00an1n01x5 FILLER_323_554 ();
 b15zdnd11an1n16x5 FILLER_323_560 ();
 b15zdnd11an1n08x5 FILLER_323_576 ();
 b15zdnd00an1n02x5 FILLER_323_584 ();
 b15zdnd00an1n01x5 FILLER_323_586 ();
 b15zdnd11an1n64x5 FILLER_323_595 ();
 b15zdnd11an1n32x5 FILLER_323_659 ();
 b15zdnd11an1n16x5 FILLER_323_691 ();
 b15zdnd11an1n08x5 FILLER_323_707 ();
 b15zdnd11an1n04x5 FILLER_323_715 ();
 b15zdnd11an1n16x5 FILLER_323_722 ();
 b15zdnd11an1n08x5 FILLER_323_738 ();
 b15zdnd11an1n04x5 FILLER_323_746 ();
 b15zdnd11an1n04x5 FILLER_323_755 ();
 b15zdnd11an1n32x5 FILLER_323_762 ();
 b15zdnd00an1n02x5 FILLER_323_794 ();
 b15zdnd00an1n01x5 FILLER_323_796 ();
 b15zdnd11an1n32x5 FILLER_323_800 ();
 b15zdnd11an1n08x5 FILLER_323_832 ();
 b15zdnd00an1n01x5 FILLER_323_840 ();
 b15zdnd11an1n16x5 FILLER_323_847 ();
 b15zdnd11an1n08x5 FILLER_323_863 ();
 b15zdnd00an1n01x5 FILLER_323_871 ();
 b15zdnd11an1n64x5 FILLER_323_881 ();
 b15zdnd11an1n32x5 FILLER_323_945 ();
 b15zdnd11an1n08x5 FILLER_323_977 ();
 b15zdnd11an1n04x5 FILLER_323_985 ();
 b15zdnd11an1n04x5 FILLER_323_994 ();
 b15zdnd00an1n02x5 FILLER_323_998 ();
 b15zdnd00an1n01x5 FILLER_323_1000 ();
 b15zdnd11an1n64x5 FILLER_323_1005 ();
 b15zdnd11an1n64x5 FILLER_323_1069 ();
 b15zdnd11an1n08x5 FILLER_323_1139 ();
 b15zdnd11an1n04x5 FILLER_323_1147 ();
 b15zdnd00an1n02x5 FILLER_323_1151 ();
 b15zdnd11an1n32x5 FILLER_323_1164 ();
 b15zdnd00an1n02x5 FILLER_323_1196 ();
 b15zdnd00an1n01x5 FILLER_323_1198 ();
 b15zdnd11an1n32x5 FILLER_323_1203 ();
 b15zdnd11an1n04x5 FILLER_323_1235 ();
 b15zdnd00an1n02x5 FILLER_323_1239 ();
 b15zdnd11an1n32x5 FILLER_323_1261 ();
 b15zdnd11an1n08x5 FILLER_323_1293 ();
 b15zdnd00an1n01x5 FILLER_323_1301 ();
 b15zdnd11an1n64x5 FILLER_323_1307 ();
 b15zdnd11an1n32x5 FILLER_323_1371 ();
 b15zdnd11an1n16x5 FILLER_323_1403 ();
 b15zdnd11an1n08x5 FILLER_323_1419 ();
 b15zdnd11an1n04x5 FILLER_323_1427 ();
 b15zdnd00an1n02x5 FILLER_323_1431 ();
 b15zdnd11an1n08x5 FILLER_323_1439 ();
 b15zdnd11an1n04x5 FILLER_323_1451 ();
 b15zdnd11an1n32x5 FILLER_323_1466 ();
 b15zdnd11an1n16x5 FILLER_323_1498 ();
 b15zdnd00an1n01x5 FILLER_323_1514 ();
 b15zdnd11an1n04x5 FILLER_323_1520 ();
 b15zdnd11an1n16x5 FILLER_323_1528 ();
 b15zdnd00an1n02x5 FILLER_323_1544 ();
 b15zdnd11an1n04x5 FILLER_323_1551 ();
 b15zdnd11an1n04x5 FILLER_323_1561 ();
 b15zdnd11an1n32x5 FILLER_323_1571 ();
 b15zdnd11an1n04x5 FILLER_323_1603 ();
 b15zdnd11an1n08x5 FILLER_323_1614 ();
 b15zdnd11an1n04x5 FILLER_323_1622 ();
 b15zdnd00an1n02x5 FILLER_323_1626 ();
 b15zdnd00an1n01x5 FILLER_323_1628 ();
 b15zdnd11an1n16x5 FILLER_323_1634 ();
 b15zdnd11an1n04x5 FILLER_323_1650 ();
 b15zdnd00an1n02x5 FILLER_323_1654 ();
 b15zdnd11an1n04x5 FILLER_323_1672 ();
 b15zdnd11an1n04x5 FILLER_323_1708 ();
 b15zdnd11an1n64x5 FILLER_323_1733 ();
 b15zdnd11an1n08x5 FILLER_323_1797 ();
 b15zdnd11an1n04x5 FILLER_323_1805 ();
 b15zdnd00an1n01x5 FILLER_323_1809 ();
 b15zdnd11an1n16x5 FILLER_323_1841 ();
 b15zdnd11an1n04x5 FILLER_323_1863 ();
 b15zdnd11an1n08x5 FILLER_323_1872 ();
 b15zdnd00an1n02x5 FILLER_323_1880 ();
 b15zdnd11an1n08x5 FILLER_323_1887 ();
 b15zdnd00an1n01x5 FILLER_323_1895 ();
 b15zdnd11an1n08x5 FILLER_323_1908 ();
 b15zdnd00an1n02x5 FILLER_323_1916 ();
 b15zdnd00an1n01x5 FILLER_323_1918 ();
 b15zdnd11an1n16x5 FILLER_323_1932 ();
 b15zdnd11an1n04x5 FILLER_323_1948 ();
 b15zdnd00an1n02x5 FILLER_323_1952 ();
 b15zdnd00an1n01x5 FILLER_323_1954 ();
 b15zdnd11an1n32x5 FILLER_323_1962 ();
 b15zdnd11an1n16x5 FILLER_323_1994 ();
 b15zdnd11an1n08x5 FILLER_323_2010 ();
 b15zdnd11an1n04x5 FILLER_323_2018 ();
 b15zdnd00an1n01x5 FILLER_323_2022 ();
 b15zdnd11an1n08x5 FILLER_323_2039 ();
 b15zdnd11an1n04x5 FILLER_323_2047 ();
 b15zdnd00an1n02x5 FILLER_323_2051 ();
 b15zdnd00an1n01x5 FILLER_323_2053 ();
 b15zdnd11an1n16x5 FILLER_323_2059 ();
 b15zdnd11an1n08x5 FILLER_323_2075 ();
 b15zdnd11an1n04x5 FILLER_323_2083 ();
 b15zdnd00an1n02x5 FILLER_323_2087 ();
 b15zdnd11an1n16x5 FILLER_323_2094 ();
 b15zdnd11an1n08x5 FILLER_323_2110 ();
 b15zdnd11an1n04x5 FILLER_323_2118 ();
 b15zdnd11an1n16x5 FILLER_323_2132 ();
 b15zdnd11an1n08x5 FILLER_323_2148 ();
 b15zdnd11an1n04x5 FILLER_323_2156 ();
 b15zdnd00an1n02x5 FILLER_323_2160 ();
 b15zdnd00an1n01x5 FILLER_323_2162 ();
 b15zdnd11an1n32x5 FILLER_323_2195 ();
 b15zdnd11an1n04x5 FILLER_323_2232 ();
 b15zdnd11an1n04x5 FILLER_323_2241 ();
 b15zdnd11an1n08x5 FILLER_323_2251 ();
 b15zdnd11an1n04x5 FILLER_323_2259 ();
 b15zdnd11an1n16x5 FILLER_323_2267 ();
 b15zdnd00an1n01x5 FILLER_323_2283 ();
 b15zdnd11an1n64x5 FILLER_324_8 ();
 b15zdnd11an1n64x5 FILLER_324_72 ();
 b15zdnd11an1n64x5 FILLER_324_136 ();
 b15zdnd11an1n08x5 FILLER_324_200 ();
 b15zdnd00an1n01x5 FILLER_324_208 ();
 b15zdnd11an1n16x5 FILLER_324_228 ();
 b15zdnd11an1n04x5 FILLER_324_244 ();
 b15zdnd00an1n02x5 FILLER_324_248 ();
 b15zdnd11an1n32x5 FILLER_324_268 ();
 b15zdnd11an1n32x5 FILLER_324_309 ();
 b15zdnd11an1n08x5 FILLER_324_341 ();
 b15zdnd00an1n02x5 FILLER_324_349 ();
 b15zdnd00an1n01x5 FILLER_324_351 ();
 b15zdnd11an1n08x5 FILLER_324_368 ();
 b15zdnd11an1n04x5 FILLER_324_376 ();
 b15zdnd11an1n08x5 FILLER_324_386 ();
 b15zdnd11an1n04x5 FILLER_324_394 ();
 b15zdnd00an1n02x5 FILLER_324_398 ();
 b15zdnd11an1n16x5 FILLER_324_406 ();
 b15zdnd00an1n02x5 FILLER_324_422 ();
 b15zdnd11an1n64x5 FILLER_324_435 ();
 b15zdnd11an1n08x5 FILLER_324_499 ();
 b15zdnd11an1n04x5 FILLER_324_507 ();
 b15zdnd00an1n02x5 FILLER_324_511 ();
 b15zdnd11an1n16x5 FILLER_324_519 ();
 b15zdnd11an1n04x5 FILLER_324_535 ();
 b15zdnd00an1n02x5 FILLER_324_539 ();
 b15zdnd00an1n01x5 FILLER_324_541 ();
 b15zdnd11an1n04x5 FILLER_324_549 ();
 b15zdnd11an1n16x5 FILLER_324_573 ();
 b15zdnd11an1n08x5 FILLER_324_589 ();
 b15zdnd11an1n08x5 FILLER_324_609 ();
 b15zdnd00an1n02x5 FILLER_324_617 ();
 b15zdnd00an1n01x5 FILLER_324_619 ();
 b15zdnd11an1n16x5 FILLER_324_636 ();
 b15zdnd00an1n02x5 FILLER_324_652 ();
 b15zdnd11an1n08x5 FILLER_324_680 ();
 b15zdnd11an1n08x5 FILLER_324_708 ();
 b15zdnd00an1n02x5 FILLER_324_716 ();
 b15zdnd11an1n32x5 FILLER_324_726 ();
 b15zdnd11an1n16x5 FILLER_324_758 ();
 b15zdnd11an1n04x5 FILLER_324_774 ();
 b15zdnd00an1n01x5 FILLER_324_778 ();
 b15zdnd11an1n04x5 FILLER_324_799 ();
 b15zdnd11an1n32x5 FILLER_324_808 ();
 b15zdnd11an1n16x5 FILLER_324_860 ();
 b15zdnd00an1n01x5 FILLER_324_876 ();
 b15zdnd11an1n08x5 FILLER_324_895 ();
 b15zdnd11an1n04x5 FILLER_324_903 ();
 b15zdnd11an1n64x5 FILLER_324_910 ();
 b15zdnd11an1n64x5 FILLER_324_974 ();
 b15zdnd11an1n64x5 FILLER_324_1038 ();
 b15zdnd11an1n32x5 FILLER_324_1102 ();
 b15zdnd11an1n16x5 FILLER_324_1134 ();
 b15zdnd11an1n04x5 FILLER_324_1150 ();
 b15zdnd00an1n01x5 FILLER_324_1154 ();
 b15zdnd11an1n64x5 FILLER_324_1175 ();
 b15zdnd11an1n32x5 FILLER_324_1239 ();
 b15zdnd11an1n16x5 FILLER_324_1271 ();
 b15zdnd11an1n04x5 FILLER_324_1287 ();
 b15zdnd00an1n02x5 FILLER_324_1291 ();
 b15zdnd00an1n01x5 FILLER_324_1293 ();
 b15zdnd11an1n64x5 FILLER_324_1298 ();
 b15zdnd11an1n32x5 FILLER_324_1362 ();
 b15zdnd11an1n04x5 FILLER_324_1426 ();
 b15zdnd11an1n08x5 FILLER_324_1444 ();
 b15zdnd00an1n02x5 FILLER_324_1452 ();
 b15zdnd00an1n01x5 FILLER_324_1454 ();
 b15zdnd11an1n32x5 FILLER_324_1461 ();
 b15zdnd11an1n08x5 FILLER_324_1493 ();
 b15zdnd11an1n04x5 FILLER_324_1501 ();
 b15zdnd00an1n01x5 FILLER_324_1505 ();
 b15zdnd11an1n04x5 FILLER_324_1510 ();
 b15zdnd00an1n02x5 FILLER_324_1514 ();
 b15zdnd00an1n01x5 FILLER_324_1516 ();
 b15zdnd11an1n16x5 FILLER_324_1529 ();
 b15zdnd11an1n08x5 FILLER_324_1545 ();
 b15zdnd00an1n02x5 FILLER_324_1553 ();
 b15zdnd11an1n32x5 FILLER_324_1562 ();
 b15zdnd11an1n08x5 FILLER_324_1594 ();
 b15zdnd11an1n04x5 FILLER_324_1602 ();
 b15zdnd00an1n01x5 FILLER_324_1606 ();
 b15zdnd11an1n04x5 FILLER_324_1615 ();
 b15zdnd11an1n04x5 FILLER_324_1625 ();
 b15zdnd11an1n32x5 FILLER_324_1635 ();
 b15zdnd11an1n08x5 FILLER_324_1667 ();
 b15zdnd11an1n04x5 FILLER_324_1675 ();
 b15zdnd00an1n01x5 FILLER_324_1679 ();
 b15zdnd11an1n16x5 FILLER_324_1698 ();
 b15zdnd00an1n02x5 FILLER_324_1714 ();
 b15zdnd11an1n64x5 FILLER_324_1742 ();
 b15zdnd11an1n16x5 FILLER_324_1837 ();
 b15zdnd00an1n01x5 FILLER_324_1853 ();
 b15zdnd11an1n16x5 FILLER_324_1862 ();
 b15zdnd11an1n08x5 FILLER_324_1878 ();
 b15zdnd11an1n04x5 FILLER_324_1886 ();
 b15zdnd11an1n04x5 FILLER_324_1910 ();
 b15zdnd11an1n08x5 FILLER_324_1940 ();
 b15zdnd11an1n04x5 FILLER_324_1948 ();
 b15zdnd11an1n32x5 FILLER_324_1971 ();
 b15zdnd11an1n16x5 FILLER_324_2003 ();
 b15zdnd11an1n04x5 FILLER_324_2019 ();
 b15zdnd00an1n02x5 FILLER_324_2023 ();
 b15zdnd11an1n32x5 FILLER_324_2038 ();
 b15zdnd11an1n16x5 FILLER_324_2070 ();
 b15zdnd00an1n02x5 FILLER_324_2086 ();
 b15zdnd11an1n32x5 FILLER_324_2107 ();
 b15zdnd11an1n08x5 FILLER_324_2139 ();
 b15zdnd11an1n04x5 FILLER_324_2147 ();
 b15zdnd00an1n02x5 FILLER_324_2151 ();
 b15zdnd00an1n01x5 FILLER_324_2153 ();
 b15zdnd11an1n04x5 FILLER_324_2162 ();
 b15zdnd11an1n32x5 FILLER_324_2184 ();
 b15zdnd11an1n16x5 FILLER_324_2216 ();
 b15zdnd11an1n08x5 FILLER_324_2232 ();
 b15zdnd11an1n04x5 FILLER_324_2240 ();
 b15zdnd00an1n01x5 FILLER_324_2244 ();
 b15zdnd11an1n16x5 FILLER_324_2252 ();
 b15zdnd11an1n08x5 FILLER_324_2268 ();
 b15zdnd11an1n64x5 FILLER_325_0 ();
 b15zdnd11an1n64x5 FILLER_325_64 ();
 b15zdnd11an1n64x5 FILLER_325_128 ();
 b15zdnd11an1n16x5 FILLER_325_192 ();
 b15zdnd11an1n08x5 FILLER_325_208 ();
 b15zdnd11an1n04x5 FILLER_325_216 ();
 b15zdnd00an1n01x5 FILLER_325_220 ();
 b15zdnd11an1n32x5 FILLER_325_237 ();
 b15zdnd11an1n08x5 FILLER_325_269 ();
 b15zdnd11an1n04x5 FILLER_325_277 ();
 b15zdnd00an1n02x5 FILLER_325_281 ();
 b15zdnd00an1n01x5 FILLER_325_283 ();
 b15zdnd11an1n64x5 FILLER_325_305 ();
 b15zdnd00an1n02x5 FILLER_325_369 ();
 b15zdnd00an1n01x5 FILLER_325_371 ();
 b15zdnd11an1n16x5 FILLER_325_376 ();
 b15zdnd11an1n08x5 FILLER_325_392 ();
 b15zdnd11an1n64x5 FILLER_325_426 ();
 b15zdnd11an1n04x5 FILLER_325_490 ();
 b15zdnd11an1n16x5 FILLER_325_501 ();
 b15zdnd11an1n04x5 FILLER_325_517 ();
 b15zdnd11an1n16x5 FILLER_325_526 ();
 b15zdnd11an1n08x5 FILLER_325_542 ();
 b15zdnd11an1n32x5 FILLER_325_576 ();
 b15zdnd00an1n02x5 FILLER_325_608 ();
 b15zdnd11an1n04x5 FILLER_325_614 ();
 b15zdnd11an1n64x5 FILLER_325_634 ();
 b15zdnd11an1n04x5 FILLER_325_698 ();
 b15zdnd00an1n02x5 FILLER_325_702 ();
 b15zdnd00an1n01x5 FILLER_325_704 ();
 b15zdnd11an1n04x5 FILLER_325_725 ();
 b15zdnd11an1n32x5 FILLER_325_734 ();
 b15zdnd11an1n08x5 FILLER_325_766 ();
 b15zdnd11an1n04x5 FILLER_325_774 ();
 b15zdnd11an1n64x5 FILLER_325_782 ();
 b15zdnd00an1n01x5 FILLER_325_846 ();
 b15zdnd11an1n32x5 FILLER_325_852 ();
 b15zdnd11an1n08x5 FILLER_325_884 ();
 b15zdnd11an1n04x5 FILLER_325_892 ();
 b15zdnd11an1n16x5 FILLER_325_916 ();
 b15zdnd11an1n08x5 FILLER_325_932 ();
 b15zdnd11an1n64x5 FILLER_325_945 ();
 b15zdnd11an1n64x5 FILLER_325_1009 ();
 b15zdnd11an1n08x5 FILLER_325_1073 ();
 b15zdnd11an1n64x5 FILLER_325_1090 ();
 b15zdnd11an1n32x5 FILLER_325_1154 ();
 b15zdnd11an1n16x5 FILLER_325_1186 ();
 b15zdnd11an1n16x5 FILLER_325_1228 ();
 b15zdnd11an1n04x5 FILLER_325_1244 ();
 b15zdnd00an1n02x5 FILLER_325_1248 ();
 b15zdnd00an1n01x5 FILLER_325_1250 ();
 b15zdnd11an1n64x5 FILLER_325_1271 ();
 b15zdnd11an1n32x5 FILLER_325_1335 ();
 b15zdnd11an1n08x5 FILLER_325_1367 ();
 b15zdnd11an1n04x5 FILLER_325_1375 ();
 b15zdnd11an1n08x5 FILLER_325_1387 ();
 b15zdnd11an1n04x5 FILLER_325_1395 ();
 b15zdnd00an1n02x5 FILLER_325_1399 ();
 b15zdnd00an1n01x5 FILLER_325_1401 ();
 b15zdnd11an1n04x5 FILLER_325_1418 ();
 b15zdnd11an1n16x5 FILLER_325_1442 ();
 b15zdnd11an1n08x5 FILLER_325_1458 ();
 b15zdnd11an1n04x5 FILLER_325_1466 ();
 b15zdnd00an1n02x5 FILLER_325_1470 ();
 b15zdnd11an1n04x5 FILLER_325_1477 ();
 b15zdnd11an1n04x5 FILLER_325_1488 ();
 b15zdnd00an1n02x5 FILLER_325_1492 ();
 b15zdnd11an1n32x5 FILLER_325_1499 ();
 b15zdnd11an1n16x5 FILLER_325_1531 ();
 b15zdnd11an1n08x5 FILLER_325_1547 ();
 b15zdnd11an1n16x5 FILLER_325_1561 ();
 b15zdnd11an1n04x5 FILLER_325_1577 ();
 b15zdnd11an1n16x5 FILLER_325_1586 ();
 b15zdnd11an1n04x5 FILLER_325_1602 ();
 b15zdnd00an1n02x5 FILLER_325_1606 ();
 b15zdnd00an1n01x5 FILLER_325_1608 ();
 b15zdnd11an1n08x5 FILLER_325_1614 ();
 b15zdnd11an1n04x5 FILLER_325_1622 ();
 b15zdnd00an1n01x5 FILLER_325_1626 ();
 b15zdnd11an1n64x5 FILLER_325_1643 ();
 b15zdnd11an1n08x5 FILLER_325_1707 ();
 b15zdnd00an1n02x5 FILLER_325_1715 ();
 b15zdnd11an1n32x5 FILLER_325_1748 ();
 b15zdnd00an1n02x5 FILLER_325_1780 ();
 b15zdnd00an1n01x5 FILLER_325_1782 ();
 b15zdnd11an1n04x5 FILLER_325_1809 ();
 b15zdnd11an1n32x5 FILLER_325_1831 ();
 b15zdnd11an1n16x5 FILLER_325_1863 ();
 b15zdnd11an1n04x5 FILLER_325_1879 ();
 b15zdnd00an1n02x5 FILLER_325_1883 ();
 b15zdnd00an1n01x5 FILLER_325_1885 ();
 b15zdnd11an1n04x5 FILLER_325_1898 ();
 b15zdnd11an1n32x5 FILLER_325_1908 ();
 b15zdnd11an1n16x5 FILLER_325_1940 ();
 b15zdnd11an1n04x5 FILLER_325_1956 ();
 b15zdnd00an1n02x5 FILLER_325_1960 ();
 b15zdnd11an1n04x5 FILLER_325_1969 ();
 b15zdnd00an1n02x5 FILLER_325_1973 ();
 b15zdnd11an1n04x5 FILLER_325_1981 ();
 b15zdnd11an1n64x5 FILLER_325_1989 ();
 b15zdnd11an1n04x5 FILLER_325_2053 ();
 b15zdnd11an1n32x5 FILLER_325_2064 ();
 b15zdnd11an1n16x5 FILLER_325_2096 ();
 b15zdnd11an1n08x5 FILLER_325_2112 ();
 b15zdnd11an1n04x5 FILLER_325_2120 ();
 b15zdnd11an1n32x5 FILLER_325_2129 ();
 b15zdnd11an1n16x5 FILLER_325_2161 ();
 b15zdnd11an1n08x5 FILLER_325_2177 ();
 b15zdnd00an1n02x5 FILLER_325_2185 ();
 b15zdnd00an1n01x5 FILLER_325_2187 ();
 b15zdnd11an1n32x5 FILLER_325_2204 ();
 b15zdnd11an1n04x5 FILLER_325_2236 ();
 b15zdnd00an1n02x5 FILLER_325_2240 ();
 b15zdnd00an1n01x5 FILLER_325_2242 ();
 b15zdnd11an1n16x5 FILLER_325_2263 ();
 b15zdnd11an1n04x5 FILLER_325_2279 ();
 b15zdnd00an1n01x5 FILLER_325_2283 ();
 b15zdnd11an1n64x5 FILLER_326_8 ();
 b15zdnd11an1n64x5 FILLER_326_72 ();
 b15zdnd11an1n64x5 FILLER_326_136 ();
 b15zdnd11an1n32x5 FILLER_326_200 ();
 b15zdnd11an1n16x5 FILLER_326_232 ();
 b15zdnd00an1n01x5 FILLER_326_248 ();
 b15zdnd11an1n04x5 FILLER_326_257 ();
 b15zdnd11an1n08x5 FILLER_326_287 ();
 b15zdnd11an1n04x5 FILLER_326_295 ();
 b15zdnd00an1n02x5 FILLER_326_299 ();
 b15zdnd00an1n01x5 FILLER_326_301 ();
 b15zdnd11an1n32x5 FILLER_326_307 ();
 b15zdnd11an1n16x5 FILLER_326_339 ();
 b15zdnd00an1n02x5 FILLER_326_355 ();
 b15zdnd11an1n04x5 FILLER_326_370 ();
 b15zdnd11an1n32x5 FILLER_326_379 ();
 b15zdnd11an1n08x5 FILLER_326_411 ();
 b15zdnd11an1n04x5 FILLER_326_419 ();
 b15zdnd00an1n02x5 FILLER_326_423 ();
 b15zdnd11an1n08x5 FILLER_326_431 ();
 b15zdnd11an1n04x5 FILLER_326_439 ();
 b15zdnd00an1n02x5 FILLER_326_443 ();
 b15zdnd00an1n01x5 FILLER_326_445 ();
 b15zdnd11an1n04x5 FILLER_326_451 ();
 b15zdnd11an1n08x5 FILLER_326_467 ();
 b15zdnd00an1n02x5 FILLER_326_475 ();
 b15zdnd00an1n01x5 FILLER_326_477 ();
 b15zdnd11an1n16x5 FILLER_326_488 ();
 b15zdnd11an1n08x5 FILLER_326_504 ();
 b15zdnd00an1n02x5 FILLER_326_512 ();
 b15zdnd11an1n32x5 FILLER_326_520 ();
 b15zdnd00an1n02x5 FILLER_326_552 ();
 b15zdnd00an1n01x5 FILLER_326_554 ();
 b15zdnd11an1n04x5 FILLER_326_574 ();
 b15zdnd11an1n64x5 FILLER_326_585 ();
 b15zdnd11an1n64x5 FILLER_326_649 ();
 b15zdnd11an1n04x5 FILLER_326_713 ();
 b15zdnd00an1n01x5 FILLER_326_717 ();
 b15zdnd11an1n08x5 FILLER_326_726 ();
 b15zdnd11an1n04x5 FILLER_326_734 ();
 b15zdnd11an1n64x5 FILLER_326_742 ();
 b15zdnd11an1n08x5 FILLER_326_806 ();
 b15zdnd11an1n04x5 FILLER_326_814 ();
 b15zdnd00an1n01x5 FILLER_326_818 ();
 b15zdnd11an1n64x5 FILLER_326_823 ();
 b15zdnd11an1n08x5 FILLER_326_887 ();
 b15zdnd00an1n02x5 FILLER_326_895 ();
 b15zdnd00an1n01x5 FILLER_326_897 ();
 b15zdnd11an1n16x5 FILLER_326_903 ();
 b15zdnd11an1n04x5 FILLER_326_919 ();
 b15zdnd00an1n02x5 FILLER_326_923 ();
 b15zdnd00an1n01x5 FILLER_326_925 ();
 b15zdnd11an1n04x5 FILLER_326_930 ();
 b15zdnd11an1n16x5 FILLER_326_954 ();
 b15zdnd00an1n01x5 FILLER_326_970 ();
 b15zdnd11an1n16x5 FILLER_326_980 ();
 b15zdnd11an1n08x5 FILLER_326_996 ();
 b15zdnd11an1n04x5 FILLER_326_1004 ();
 b15zdnd11an1n32x5 FILLER_326_1019 ();
 b15zdnd11an1n08x5 FILLER_326_1051 ();
 b15zdnd00an1n02x5 FILLER_326_1059 ();
 b15zdnd11an1n08x5 FILLER_326_1070 ();
 b15zdnd00an1n02x5 FILLER_326_1078 ();
 b15zdnd00an1n01x5 FILLER_326_1080 ();
 b15zdnd11an1n64x5 FILLER_326_1101 ();
 b15zdnd11an1n32x5 FILLER_326_1165 ();
 b15zdnd11an1n16x5 FILLER_326_1197 ();
 b15zdnd11an1n08x5 FILLER_326_1213 ();
 b15zdnd00an1n02x5 FILLER_326_1221 ();
 b15zdnd11an1n08x5 FILLER_326_1243 ();
 b15zdnd00an1n02x5 FILLER_326_1251 ();
 b15zdnd11an1n64x5 FILLER_326_1258 ();
 b15zdnd11an1n16x5 FILLER_326_1322 ();
 b15zdnd00an1n02x5 FILLER_326_1338 ();
 b15zdnd11an1n16x5 FILLER_326_1356 ();
 b15zdnd11an1n08x5 FILLER_326_1372 ();
 b15zdnd00an1n01x5 FILLER_326_1380 ();
 b15zdnd11an1n32x5 FILLER_326_1394 ();
 b15zdnd00an1n01x5 FILLER_326_1426 ();
 b15zdnd11an1n64x5 FILLER_326_1453 ();
 b15zdnd11an1n64x5 FILLER_326_1517 ();
 b15zdnd11an1n32x5 FILLER_326_1593 ();
 b15zdnd00an1n02x5 FILLER_326_1625 ();
 b15zdnd00an1n01x5 FILLER_326_1627 ();
 b15zdnd11an1n64x5 FILLER_326_1637 ();
 b15zdnd11an1n64x5 FILLER_326_1701 ();
 b15zdnd11an1n64x5 FILLER_326_1765 ();
 b15zdnd11an1n64x5 FILLER_326_1829 ();
 b15zdnd11an1n08x5 FILLER_326_1893 ();
 b15zdnd00an1n01x5 FILLER_326_1901 ();
 b15zdnd11an1n04x5 FILLER_326_1907 ();
 b15zdnd11an1n32x5 FILLER_326_1924 ();
 b15zdnd00an1n02x5 FILLER_326_1956 ();
 b15zdnd00an1n01x5 FILLER_326_1958 ();
 b15zdnd11an1n08x5 FILLER_326_1965 ();
 b15zdnd11an1n04x5 FILLER_326_1973 ();
 b15zdnd00an1n02x5 FILLER_326_1977 ();
 b15zdnd11an1n16x5 FILLER_326_1983 ();
 b15zdnd11an1n04x5 FILLER_326_1999 ();
 b15zdnd11an1n04x5 FILLER_326_2015 ();
 b15zdnd11an1n16x5 FILLER_326_2024 ();
 b15zdnd11an1n08x5 FILLER_326_2040 ();
 b15zdnd11an1n04x5 FILLER_326_2048 ();
 b15zdnd00an1n01x5 FILLER_326_2052 ();
 b15zdnd11an1n32x5 FILLER_326_2062 ();
 b15zdnd11an1n16x5 FILLER_326_2094 ();
 b15zdnd11an1n04x5 FILLER_326_2110 ();
 b15zdnd00an1n02x5 FILLER_326_2114 ();
 b15zdnd00an1n01x5 FILLER_326_2116 ();
 b15zdnd11an1n16x5 FILLER_326_2128 ();
 b15zdnd11an1n08x5 FILLER_326_2144 ();
 b15zdnd00an1n02x5 FILLER_326_2152 ();
 b15zdnd00an1n02x5 FILLER_326_2162 ();
 b15zdnd11an1n64x5 FILLER_326_2195 ();
 b15zdnd11an1n16x5 FILLER_326_2259 ();
 b15zdnd00an1n01x5 FILLER_326_2275 ();
 b15zdnd11an1n64x5 FILLER_327_0 ();
 b15zdnd11an1n64x5 FILLER_327_64 ();
 b15zdnd11an1n64x5 FILLER_327_128 ();
 b15zdnd11an1n16x5 FILLER_327_192 ();
 b15zdnd11an1n08x5 FILLER_327_208 ();
 b15zdnd11an1n04x5 FILLER_327_236 ();
 b15zdnd00an1n01x5 FILLER_327_240 ();
 b15zdnd11an1n04x5 FILLER_327_250 ();
 b15zdnd00an1n01x5 FILLER_327_254 ();
 b15zdnd11an1n04x5 FILLER_327_261 ();
 b15zdnd00an1n02x5 FILLER_327_265 ();
 b15zdnd00an1n01x5 FILLER_327_267 ();
 b15zdnd11an1n08x5 FILLER_327_292 ();
 b15zdnd00an1n01x5 FILLER_327_300 ();
 b15zdnd11an1n64x5 FILLER_327_313 ();
 b15zdnd11an1n64x5 FILLER_327_377 ();
 b15zdnd11an1n32x5 FILLER_327_441 ();
 b15zdnd11an1n08x5 FILLER_327_473 ();
 b15zdnd11an1n04x5 FILLER_327_481 ();
 b15zdnd11an1n16x5 FILLER_327_490 ();
 b15zdnd11an1n04x5 FILLER_327_506 ();
 b15zdnd11an1n64x5 FILLER_327_514 ();
 b15zdnd00an1n02x5 FILLER_327_578 ();
 b15zdnd00an1n01x5 FILLER_327_580 ();
 b15zdnd11an1n16x5 FILLER_327_586 ();
 b15zdnd11an1n08x5 FILLER_327_602 ();
 b15zdnd00an1n02x5 FILLER_327_610 ();
 b15zdnd11an1n64x5 FILLER_327_624 ();
 b15zdnd11an1n64x5 FILLER_327_688 ();
 b15zdnd11an1n64x5 FILLER_327_752 ();
 b15zdnd11an1n64x5 FILLER_327_816 ();
 b15zdnd11an1n32x5 FILLER_327_880 ();
 b15zdnd11an1n16x5 FILLER_327_912 ();
 b15zdnd11an1n08x5 FILLER_327_928 ();
 b15zdnd00an1n02x5 FILLER_327_936 ();
 b15zdnd11an1n64x5 FILLER_327_944 ();
 b15zdnd11an1n04x5 FILLER_327_1008 ();
 b15zdnd00an1n02x5 FILLER_327_1012 ();
 b15zdnd00an1n01x5 FILLER_327_1014 ();
 b15zdnd11an1n64x5 FILLER_327_1035 ();
 b15zdnd11an1n08x5 FILLER_327_1099 ();
 b15zdnd11an1n04x5 FILLER_327_1107 ();
 b15zdnd00an1n01x5 FILLER_327_1111 ();
 b15zdnd11an1n32x5 FILLER_327_1132 ();
 b15zdnd11an1n16x5 FILLER_327_1164 ();
 b15zdnd11an1n08x5 FILLER_327_1180 ();
 b15zdnd11an1n04x5 FILLER_327_1188 ();
 b15zdnd00an1n02x5 FILLER_327_1192 ();
 b15zdnd11an1n32x5 FILLER_327_1214 ();
 b15zdnd11an1n04x5 FILLER_327_1246 ();
 b15zdnd00an1n01x5 FILLER_327_1250 ();
 b15zdnd11an1n64x5 FILLER_327_1257 ();
 b15zdnd11an1n32x5 FILLER_327_1321 ();
 b15zdnd00an1n02x5 FILLER_327_1353 ();
 b15zdnd00an1n01x5 FILLER_327_1355 ();
 b15zdnd11an1n32x5 FILLER_327_1365 ();
 b15zdnd00an1n02x5 FILLER_327_1397 ();
 b15zdnd11an1n04x5 FILLER_327_1406 ();
 b15zdnd00an1n01x5 FILLER_327_1410 ();
 b15zdnd11an1n04x5 FILLER_327_1416 ();
 b15zdnd11an1n64x5 FILLER_327_1428 ();
 b15zdnd11an1n64x5 FILLER_327_1492 ();
 b15zdnd11an1n32x5 FILLER_327_1556 ();
 b15zdnd11an1n16x5 FILLER_327_1588 ();
 b15zdnd11an1n08x5 FILLER_327_1604 ();
 b15zdnd00an1n01x5 FILLER_327_1612 ();
 b15zdnd11an1n08x5 FILLER_327_1618 ();
 b15zdnd00an1n01x5 FILLER_327_1626 ();
 b15zdnd11an1n64x5 FILLER_327_1633 ();
 b15zdnd11an1n16x5 FILLER_327_1697 ();
 b15zdnd11an1n04x5 FILLER_327_1713 ();
 b15zdnd00an1n02x5 FILLER_327_1717 ();
 b15zdnd11an1n32x5 FILLER_327_1737 ();
 b15zdnd11an1n16x5 FILLER_327_1769 ();
 b15zdnd11an1n08x5 FILLER_327_1785 ();
 b15zdnd00an1n02x5 FILLER_327_1793 ();
 b15zdnd11an1n04x5 FILLER_327_1811 ();
 b15zdnd11an1n08x5 FILLER_327_1841 ();
 b15zdnd00an1n02x5 FILLER_327_1849 ();
 b15zdnd11an1n32x5 FILLER_327_1874 ();
 b15zdnd11an1n08x5 FILLER_327_1906 ();
 b15zdnd11an1n04x5 FILLER_327_1914 ();
 b15zdnd11an1n64x5 FILLER_327_1932 ();
 b15zdnd11an1n08x5 FILLER_327_1996 ();
 b15zdnd00an1n02x5 FILLER_327_2004 ();
 b15zdnd00an1n01x5 FILLER_327_2006 ();
 b15zdnd11an1n04x5 FILLER_327_2020 ();
 b15zdnd00an1n01x5 FILLER_327_2024 ();
 b15zdnd11an1n32x5 FILLER_327_2042 ();
 b15zdnd00an1n02x5 FILLER_327_2074 ();
 b15zdnd00an1n01x5 FILLER_327_2076 ();
 b15zdnd11an1n64x5 FILLER_327_2082 ();
 b15zdnd11an1n08x5 FILLER_327_2146 ();
 b15zdnd11an1n04x5 FILLER_327_2154 ();
 b15zdnd00an1n02x5 FILLER_327_2158 ();
 b15zdnd00an1n01x5 FILLER_327_2160 ();
 b15zdnd11an1n04x5 FILLER_327_2166 ();
 b15zdnd11an1n16x5 FILLER_327_2180 ();
 b15zdnd11an1n04x5 FILLER_327_2196 ();
 b15zdnd00an1n02x5 FILLER_327_2200 ();
 b15zdnd00an1n01x5 FILLER_327_2202 ();
 b15zdnd11an1n64x5 FILLER_327_2219 ();
 b15zdnd00an1n01x5 FILLER_327_2283 ();
 b15zdnd11an1n64x5 FILLER_328_8 ();
 b15zdnd11an1n64x5 FILLER_328_72 ();
 b15zdnd11an1n64x5 FILLER_328_136 ();
 b15zdnd11an1n16x5 FILLER_328_200 ();
 b15zdnd11an1n08x5 FILLER_328_216 ();
 b15zdnd00an1n01x5 FILLER_328_224 ();
 b15zdnd11an1n64x5 FILLER_328_241 ();
 b15zdnd11an1n16x5 FILLER_328_305 ();
 b15zdnd00an1n02x5 FILLER_328_321 ();
 b15zdnd00an1n01x5 FILLER_328_323 ();
 b15zdnd11an1n32x5 FILLER_328_329 ();
 b15zdnd11an1n08x5 FILLER_328_361 ();
 b15zdnd00an1n02x5 FILLER_328_369 ();
 b15zdnd00an1n01x5 FILLER_328_371 ();
 b15zdnd11an1n64x5 FILLER_328_381 ();
 b15zdnd11an1n32x5 FILLER_328_445 ();
 b15zdnd11an1n04x5 FILLER_328_477 ();
 b15zdnd00an1n02x5 FILLER_328_481 ();
 b15zdnd11an1n16x5 FILLER_328_495 ();
 b15zdnd11an1n08x5 FILLER_328_511 ();
 b15zdnd00an1n01x5 FILLER_328_519 ();
 b15zdnd11an1n16x5 FILLER_328_540 ();
 b15zdnd11an1n04x5 FILLER_328_556 ();
 b15zdnd00an1n01x5 FILLER_328_560 ();
 b15zdnd11an1n04x5 FILLER_328_570 ();
 b15zdnd00an1n02x5 FILLER_328_574 ();
 b15zdnd11an1n16x5 FILLER_328_588 ();
 b15zdnd00an1n01x5 FILLER_328_604 ();
 b15zdnd11an1n64x5 FILLER_328_614 ();
 b15zdnd11an1n32x5 FILLER_328_678 ();
 b15zdnd11an1n08x5 FILLER_328_710 ();
 b15zdnd11an1n64x5 FILLER_328_726 ();
 b15zdnd11an1n16x5 FILLER_328_790 ();
 b15zdnd11an1n08x5 FILLER_328_806 ();
 b15zdnd11an1n04x5 FILLER_328_814 ();
 b15zdnd00an1n01x5 FILLER_328_818 ();
 b15zdnd11an1n08x5 FILLER_328_828 ();
 b15zdnd11an1n04x5 FILLER_328_836 ();
 b15zdnd00an1n02x5 FILLER_328_840 ();
 b15zdnd11an1n64x5 FILLER_328_874 ();
 b15zdnd11an1n32x5 FILLER_328_938 ();
 b15zdnd00an1n02x5 FILLER_328_970 ();
 b15zdnd11an1n64x5 FILLER_328_992 ();
 b15zdnd11an1n08x5 FILLER_328_1056 ();
 b15zdnd11an1n04x5 FILLER_328_1064 ();
 b15zdnd11an1n16x5 FILLER_328_1088 ();
 b15zdnd11an1n08x5 FILLER_328_1104 ();
 b15zdnd11an1n04x5 FILLER_328_1115 ();
 b15zdnd11an1n16x5 FILLER_328_1124 ();
 b15zdnd11an1n08x5 FILLER_328_1140 ();
 b15zdnd00an1n02x5 FILLER_328_1148 ();
 b15zdnd11an1n64x5 FILLER_328_1156 ();
 b15zdnd11an1n64x5 FILLER_328_1220 ();
 b15zdnd11an1n64x5 FILLER_328_1284 ();
 b15zdnd11an1n64x5 FILLER_328_1348 ();
 b15zdnd11an1n08x5 FILLER_328_1412 ();
 b15zdnd11an1n04x5 FILLER_328_1420 ();
 b15zdnd00an1n02x5 FILLER_328_1424 ();
 b15zdnd00an1n01x5 FILLER_328_1426 ();
 b15zdnd11an1n04x5 FILLER_328_1433 ();
 b15zdnd11an1n32x5 FILLER_328_1449 ();
 b15zdnd00an1n02x5 FILLER_328_1481 ();
 b15zdnd11an1n16x5 FILLER_328_1504 ();
 b15zdnd11an1n04x5 FILLER_328_1520 ();
 b15zdnd11an1n32x5 FILLER_328_1545 ();
 b15zdnd11an1n16x5 FILLER_328_1577 ();
 b15zdnd00an1n02x5 FILLER_328_1593 ();
 b15zdnd11an1n08x5 FILLER_328_1610 ();
 b15zdnd11an1n04x5 FILLER_328_1618 ();
 b15zdnd11an1n64x5 FILLER_328_1628 ();
 b15zdnd11an1n04x5 FILLER_328_1692 ();
 b15zdnd00an1n02x5 FILLER_328_1696 ();
 b15zdnd00an1n01x5 FILLER_328_1698 ();
 b15zdnd11an1n04x5 FILLER_328_1705 ();
 b15zdnd11an1n64x5 FILLER_328_1713 ();
 b15zdnd11an1n16x5 FILLER_328_1777 ();
 b15zdnd00an1n02x5 FILLER_328_1793 ();
 b15zdnd11an1n16x5 FILLER_328_1821 ();
 b15zdnd11an1n08x5 FILLER_328_1837 ();
 b15zdnd00an1n02x5 FILLER_328_1845 ();
 b15zdnd00an1n01x5 FILLER_328_1847 ();
 b15zdnd11an1n08x5 FILLER_328_1861 ();
 b15zdnd11an1n04x5 FILLER_328_1869 ();
 b15zdnd00an1n02x5 FILLER_328_1873 ();
 b15zdnd00an1n01x5 FILLER_328_1875 ();
 b15zdnd11an1n08x5 FILLER_328_1890 ();
 b15zdnd11an1n32x5 FILLER_328_1902 ();
 b15zdnd00an1n02x5 FILLER_328_1934 ();
 b15zdnd11an1n08x5 FILLER_328_1950 ();
 b15zdnd00an1n02x5 FILLER_328_1958 ();
 b15zdnd11an1n64x5 FILLER_328_1964 ();
 b15zdnd11an1n16x5 FILLER_328_2028 ();
 b15zdnd00an1n02x5 FILLER_328_2044 ();
 b15zdnd11an1n16x5 FILLER_328_2066 ();
 b15zdnd11an1n32x5 FILLER_328_2088 ();
 b15zdnd11an1n04x5 FILLER_328_2120 ();
 b15zdnd11an1n16x5 FILLER_328_2136 ();
 b15zdnd00an1n02x5 FILLER_328_2152 ();
 b15zdnd11an1n32x5 FILLER_328_2162 ();
 b15zdnd11an1n08x5 FILLER_328_2194 ();
 b15zdnd00an1n01x5 FILLER_328_2202 ();
 b15zdnd11an1n32x5 FILLER_328_2223 ();
 b15zdnd11an1n16x5 FILLER_328_2255 ();
 b15zdnd11an1n04x5 FILLER_328_2271 ();
 b15zdnd00an1n01x5 FILLER_328_2275 ();
 b15zdnd11an1n64x5 FILLER_329_0 ();
 b15zdnd11an1n64x5 FILLER_329_64 ();
 b15zdnd11an1n64x5 FILLER_329_128 ();
 b15zdnd11an1n64x5 FILLER_329_192 ();
 b15zdnd11an1n32x5 FILLER_329_256 ();
 b15zdnd11an1n16x5 FILLER_329_288 ();
 b15zdnd11an1n08x5 FILLER_329_304 ();
 b15zdnd11an1n04x5 FILLER_329_312 ();
 b15zdnd00an1n02x5 FILLER_329_316 ();
 b15zdnd00an1n01x5 FILLER_329_318 ();
 b15zdnd11an1n16x5 FILLER_329_334 ();
 b15zdnd11an1n04x5 FILLER_329_350 ();
 b15zdnd00an1n02x5 FILLER_329_354 ();
 b15zdnd00an1n01x5 FILLER_329_356 ();
 b15zdnd11an1n04x5 FILLER_329_378 ();
 b15zdnd11an1n04x5 FILLER_329_392 ();
 b15zdnd11an1n32x5 FILLER_329_406 ();
 b15zdnd11an1n16x5 FILLER_329_438 ();
 b15zdnd11an1n08x5 FILLER_329_454 ();
 b15zdnd00an1n01x5 FILLER_329_462 ();
 b15zdnd11an1n16x5 FILLER_329_483 ();
 b15zdnd11an1n04x5 FILLER_329_499 ();
 b15zdnd00an1n02x5 FILLER_329_503 ();
 b15zdnd00an1n01x5 FILLER_329_505 ();
 b15zdnd11an1n08x5 FILLER_329_510 ();
 b15zdnd00an1n02x5 FILLER_329_518 ();
 b15zdnd00an1n01x5 FILLER_329_520 ();
 b15zdnd11an1n32x5 FILLER_329_534 ();
 b15zdnd11an1n08x5 FILLER_329_566 ();
 b15zdnd00an1n02x5 FILLER_329_574 ();
 b15zdnd00an1n01x5 FILLER_329_576 ();
 b15zdnd11an1n04x5 FILLER_329_581 ();
 b15zdnd11an1n04x5 FILLER_329_605 ();
 b15zdnd11an1n04x5 FILLER_329_623 ();
 b15zdnd11an1n32x5 FILLER_329_636 ();
 b15zdnd00an1n02x5 FILLER_329_668 ();
 b15zdnd11an1n08x5 FILLER_329_682 ();
 b15zdnd00an1n02x5 FILLER_329_690 ();
 b15zdnd11an1n16x5 FILLER_329_710 ();
 b15zdnd11an1n04x5 FILLER_329_726 ();
 b15zdnd00an1n02x5 FILLER_329_730 ();
 b15zdnd11an1n04x5 FILLER_329_744 ();
 b15zdnd11an1n04x5 FILLER_329_755 ();
 b15zdnd00an1n02x5 FILLER_329_759 ();
 b15zdnd11an1n64x5 FILLER_329_767 ();
 b15zdnd11an1n04x5 FILLER_329_831 ();
 b15zdnd11an1n64x5 FILLER_329_844 ();
 b15zdnd11an1n64x5 FILLER_329_908 ();
 b15zdnd11an1n64x5 FILLER_329_972 ();
 b15zdnd11an1n64x5 FILLER_329_1036 ();
 b15zdnd11an1n32x5 FILLER_329_1100 ();
 b15zdnd11an1n16x5 FILLER_329_1152 ();
 b15zdnd11an1n04x5 FILLER_329_1168 ();
 b15zdnd00an1n01x5 FILLER_329_1172 ();
 b15zdnd11an1n16x5 FILLER_329_1193 ();
 b15zdnd11an1n08x5 FILLER_329_1209 ();
 b15zdnd11an1n04x5 FILLER_329_1217 ();
 b15zdnd00an1n02x5 FILLER_329_1221 ();
 b15zdnd11an1n32x5 FILLER_329_1243 ();
 b15zdnd11an1n08x5 FILLER_329_1275 ();
 b15zdnd11an1n04x5 FILLER_329_1283 ();
 b15zdnd00an1n01x5 FILLER_329_1287 ();
 b15zdnd11an1n04x5 FILLER_329_1297 ();
 b15zdnd00an1n02x5 FILLER_329_1301 ();
 b15zdnd00an1n01x5 FILLER_329_1303 ();
 b15zdnd11an1n04x5 FILLER_329_1324 ();
 b15zdnd11an1n04x5 FILLER_329_1335 ();
 b15zdnd11an1n64x5 FILLER_329_1346 ();
 b15zdnd11an1n04x5 FILLER_329_1410 ();
 b15zdnd00an1n02x5 FILLER_329_1414 ();
 b15zdnd11an1n08x5 FILLER_329_1425 ();
 b15zdnd00an1n02x5 FILLER_329_1433 ();
 b15zdnd11an1n08x5 FILLER_329_1447 ();
 b15zdnd11an1n04x5 FILLER_329_1455 ();
 b15zdnd00an1n01x5 FILLER_329_1459 ();
 b15zdnd11an1n32x5 FILLER_329_1464 ();
 b15zdnd11an1n16x5 FILLER_329_1496 ();
 b15zdnd11an1n08x5 FILLER_329_1512 ();
 b15zdnd00an1n01x5 FILLER_329_1520 ();
 b15zdnd11an1n32x5 FILLER_329_1530 ();
 b15zdnd11an1n16x5 FILLER_329_1562 ();
 b15zdnd11an1n04x5 FILLER_329_1578 ();
 b15zdnd11an1n16x5 FILLER_329_1586 ();
 b15zdnd00an1n01x5 FILLER_329_1602 ();
 b15zdnd11an1n16x5 FILLER_329_1629 ();
 b15zdnd11an1n04x5 FILLER_329_1645 ();
 b15zdnd00an1n02x5 FILLER_329_1649 ();
 b15zdnd11an1n04x5 FILLER_329_1656 ();
 b15zdnd00an1n02x5 FILLER_329_1660 ();
 b15zdnd00an1n01x5 FILLER_329_1662 ();
 b15zdnd11an1n04x5 FILLER_329_1667 ();
 b15zdnd11an1n16x5 FILLER_329_1684 ();
 b15zdnd11an1n08x5 FILLER_329_1700 ();
 b15zdnd00an1n01x5 FILLER_329_1708 ();
 b15zdnd11an1n04x5 FILLER_329_1741 ();
 b15zdnd11an1n32x5 FILLER_329_1749 ();
 b15zdnd11an1n16x5 FILLER_329_1781 ();
 b15zdnd11an1n04x5 FILLER_329_1797 ();
 b15zdnd11an1n04x5 FILLER_329_1827 ();
 b15zdnd11an1n16x5 FILLER_329_1847 ();
 b15zdnd11an1n04x5 FILLER_329_1863 ();
 b15zdnd00an1n02x5 FILLER_329_1867 ();
 b15zdnd00an1n01x5 FILLER_329_1869 ();
 b15zdnd11an1n04x5 FILLER_329_1893 ();
 b15zdnd11an1n64x5 FILLER_329_1903 ();
 b15zdnd11an1n32x5 FILLER_329_1967 ();
 b15zdnd11an1n08x5 FILLER_329_1999 ();
 b15zdnd11an1n04x5 FILLER_329_2007 ();
 b15zdnd00an1n02x5 FILLER_329_2011 ();
 b15zdnd11an1n16x5 FILLER_329_2034 ();
 b15zdnd00an1n02x5 FILLER_329_2050 ();
 b15zdnd11an1n08x5 FILLER_329_2061 ();
 b15zdnd11an1n04x5 FILLER_329_2069 ();
 b15zdnd11an1n32x5 FILLER_329_2081 ();
 b15zdnd11an1n08x5 FILLER_329_2113 ();
 b15zdnd00an1n02x5 FILLER_329_2121 ();
 b15zdnd00an1n01x5 FILLER_329_2123 ();
 b15zdnd11an1n16x5 FILLER_329_2134 ();
 b15zdnd11an1n08x5 FILLER_329_2150 ();
 b15zdnd11an1n08x5 FILLER_329_2174 ();
 b15zdnd00an1n02x5 FILLER_329_2182 ();
 b15zdnd00an1n01x5 FILLER_329_2184 ();
 b15zdnd11an1n64x5 FILLER_329_2191 ();
 b15zdnd11an1n16x5 FILLER_329_2255 ();
 b15zdnd11an1n08x5 FILLER_329_2271 ();
 b15zdnd11an1n04x5 FILLER_329_2279 ();
 b15zdnd00an1n01x5 FILLER_329_2283 ();
 b15zdnd11an1n64x5 FILLER_330_8 ();
 b15zdnd11an1n64x5 FILLER_330_72 ();
 b15zdnd11an1n64x5 FILLER_330_136 ();
 b15zdnd11an1n64x5 FILLER_330_200 ();
 b15zdnd11an1n32x5 FILLER_330_264 ();
 b15zdnd11an1n08x5 FILLER_330_296 ();
 b15zdnd11an1n04x5 FILLER_330_316 ();
 b15zdnd11an1n32x5 FILLER_330_324 ();
 b15zdnd11an1n16x5 FILLER_330_356 ();
 b15zdnd11an1n04x5 FILLER_330_372 ();
 b15zdnd11an1n04x5 FILLER_330_382 ();
 b15zdnd11an1n08x5 FILLER_330_391 ();
 b15zdnd11an1n04x5 FILLER_330_399 ();
 b15zdnd11an1n04x5 FILLER_330_415 ();
 b15zdnd11an1n04x5 FILLER_330_425 ();
 b15zdnd11an1n04x5 FILLER_330_434 ();
 b15zdnd11an1n08x5 FILLER_330_442 ();
 b15zdnd00an1n02x5 FILLER_330_450 ();
 b15zdnd11an1n16x5 FILLER_330_466 ();
 b15zdnd11an1n08x5 FILLER_330_482 ();
 b15zdnd00an1n01x5 FILLER_330_490 ();
 b15zdnd11an1n04x5 FILLER_330_503 ();
 b15zdnd11an1n32x5 FILLER_330_513 ();
 b15zdnd11an1n08x5 FILLER_330_545 ();
 b15zdnd11an1n04x5 FILLER_330_553 ();
 b15zdnd00an1n02x5 FILLER_330_557 ();
 b15zdnd00an1n01x5 FILLER_330_559 ();
 b15zdnd11an1n64x5 FILLER_330_580 ();
 b15zdnd11an1n32x5 FILLER_330_644 ();
 b15zdnd11an1n04x5 FILLER_330_676 ();
 b15zdnd11an1n16x5 FILLER_330_701 ();
 b15zdnd00an1n01x5 FILLER_330_717 ();
 b15zdnd11an1n08x5 FILLER_330_726 ();
 b15zdnd00an1n02x5 FILLER_330_734 ();
 b15zdnd11an1n08x5 FILLER_330_750 ();
 b15zdnd00an1n02x5 FILLER_330_758 ();
 b15zdnd11an1n04x5 FILLER_330_778 ();
 b15zdnd11an1n32x5 FILLER_330_790 ();
 b15zdnd11an1n04x5 FILLER_330_822 ();
 b15zdnd00an1n02x5 FILLER_330_826 ();
 b15zdnd00an1n01x5 FILLER_330_828 ();
 b15zdnd11an1n08x5 FILLER_330_836 ();
 b15zdnd00an1n02x5 FILLER_330_844 ();
 b15zdnd00an1n01x5 FILLER_330_846 ();
 b15zdnd11an1n04x5 FILLER_330_857 ();
 b15zdnd00an1n02x5 FILLER_330_861 ();
 b15zdnd11an1n04x5 FILLER_330_879 ();
 b15zdnd00an1n02x5 FILLER_330_883 ();
 b15zdnd00an1n01x5 FILLER_330_885 ();
 b15zdnd11an1n64x5 FILLER_330_891 ();
 b15zdnd11an1n64x5 FILLER_330_955 ();
 b15zdnd11an1n32x5 FILLER_330_1019 ();
 b15zdnd11an1n16x5 FILLER_330_1051 ();
 b15zdnd11an1n08x5 FILLER_330_1067 ();
 b15zdnd00an1n02x5 FILLER_330_1075 ();
 b15zdnd11an1n32x5 FILLER_330_1095 ();
 b15zdnd11an1n08x5 FILLER_330_1127 ();
 b15zdnd11an1n04x5 FILLER_330_1135 ();
 b15zdnd11an1n16x5 FILLER_330_1144 ();
 b15zdnd11an1n08x5 FILLER_330_1160 ();
 b15zdnd00an1n01x5 FILLER_330_1168 ();
 b15zdnd11an1n08x5 FILLER_330_1175 ();
 b15zdnd11an1n04x5 FILLER_330_1183 ();
 b15zdnd00an1n01x5 FILLER_330_1187 ();
 b15zdnd11an1n16x5 FILLER_330_1193 ();
 b15zdnd11an1n08x5 FILLER_330_1209 ();
 b15zdnd11an1n04x5 FILLER_330_1217 ();
 b15zdnd00an1n01x5 FILLER_330_1221 ();
 b15zdnd11an1n08x5 FILLER_330_1227 ();
 b15zdnd11an1n04x5 FILLER_330_1235 ();
 b15zdnd00an1n02x5 FILLER_330_1239 ();
 b15zdnd11an1n64x5 FILLER_330_1245 ();
 b15zdnd11an1n32x5 FILLER_330_1309 ();
 b15zdnd00an1n02x5 FILLER_330_1341 ();
 b15zdnd00an1n01x5 FILLER_330_1343 ();
 b15zdnd11an1n32x5 FILLER_330_1350 ();
 b15zdnd11an1n08x5 FILLER_330_1382 ();
 b15zdnd11an1n04x5 FILLER_330_1390 ();
 b15zdnd00an1n01x5 FILLER_330_1394 ();
 b15zdnd11an1n04x5 FILLER_330_1399 ();
 b15zdnd11an1n08x5 FILLER_330_1410 ();
 b15zdnd11an1n04x5 FILLER_330_1418 ();
 b15zdnd11an1n04x5 FILLER_330_1428 ();
 b15zdnd11an1n08x5 FILLER_330_1437 ();
 b15zdnd11an1n04x5 FILLER_330_1445 ();
 b15zdnd00an1n02x5 FILLER_330_1449 ();
 b15zdnd11an1n04x5 FILLER_330_1477 ();
 b15zdnd11an1n04x5 FILLER_330_1488 ();
 b15zdnd11an1n16x5 FILLER_330_1498 ();
 b15zdnd11an1n04x5 FILLER_330_1514 ();
 b15zdnd11an1n16x5 FILLER_330_1525 ();
 b15zdnd11an1n04x5 FILLER_330_1541 ();
 b15zdnd11an1n16x5 FILLER_330_1551 ();
 b15zdnd11an1n08x5 FILLER_330_1567 ();
 b15zdnd11an1n04x5 FILLER_330_1575 ();
 b15zdnd11an1n08x5 FILLER_330_1585 ();
 b15zdnd11an1n04x5 FILLER_330_1593 ();
 b15zdnd00an1n01x5 FILLER_330_1597 ();
 b15zdnd11an1n04x5 FILLER_330_1629 ();
 b15zdnd11an1n08x5 FILLER_330_1639 ();
 b15zdnd00an1n02x5 FILLER_330_1647 ();
 b15zdnd11an1n32x5 FILLER_330_1665 ();
 b15zdnd11an1n08x5 FILLER_330_1697 ();
 b15zdnd00an1n02x5 FILLER_330_1705 ();
 b15zdnd11an1n16x5 FILLER_330_1718 ();
 b15zdnd11an1n04x5 FILLER_330_1734 ();
 b15zdnd00an1n02x5 FILLER_330_1738 ();
 b15zdnd11an1n04x5 FILLER_330_1745 ();
 b15zdnd00an1n02x5 FILLER_330_1749 ();
 b15zdnd11an1n32x5 FILLER_330_1757 ();
 b15zdnd11an1n08x5 FILLER_330_1789 ();
 b15zdnd11an1n04x5 FILLER_330_1797 ();
 b15zdnd11an1n32x5 FILLER_330_1819 ();
 b15zdnd11an1n16x5 FILLER_330_1851 ();
 b15zdnd11an1n08x5 FILLER_330_1867 ();
 b15zdnd11an1n04x5 FILLER_330_1875 ();
 b15zdnd11an1n04x5 FILLER_330_1885 ();
 b15zdnd00an1n02x5 FILLER_330_1889 ();
 b15zdnd11an1n32x5 FILLER_330_1905 ();
 b15zdnd11an1n16x5 FILLER_330_1937 ();
 b15zdnd11an1n08x5 FILLER_330_1953 ();
 b15zdnd11an1n04x5 FILLER_330_1961 ();
 b15zdnd00an1n02x5 FILLER_330_1965 ();
 b15zdnd00an1n01x5 FILLER_330_1967 ();
 b15zdnd11an1n64x5 FILLER_330_1978 ();
 b15zdnd00an1n02x5 FILLER_330_2042 ();
 b15zdnd11an1n16x5 FILLER_330_2051 ();
 b15zdnd00an1n01x5 FILLER_330_2067 ();
 b15zdnd11an1n04x5 FILLER_330_2074 ();
 b15zdnd11an1n08x5 FILLER_330_2083 ();
 b15zdnd00an1n02x5 FILLER_330_2091 ();
 b15zdnd00an1n01x5 FILLER_330_2093 ();
 b15zdnd11an1n16x5 FILLER_330_2100 ();
 b15zdnd00an1n02x5 FILLER_330_2116 ();
 b15zdnd00an1n01x5 FILLER_330_2118 ();
 b15zdnd11an1n16x5 FILLER_330_2131 ();
 b15zdnd11an1n04x5 FILLER_330_2147 ();
 b15zdnd00an1n02x5 FILLER_330_2151 ();
 b15zdnd00an1n01x5 FILLER_330_2153 ();
 b15zdnd11an1n04x5 FILLER_330_2162 ();
 b15zdnd00an1n02x5 FILLER_330_2166 ();
 b15zdnd11an1n04x5 FILLER_330_2174 ();
 b15zdnd11an1n08x5 FILLER_330_2182 ();
 b15zdnd00an1n02x5 FILLER_330_2190 ();
 b15zdnd11an1n04x5 FILLER_330_2197 ();
 b15zdnd11an1n32x5 FILLER_330_2213 ();
 b15zdnd11an1n16x5 FILLER_330_2245 ();
 b15zdnd11an1n08x5 FILLER_330_2261 ();
 b15zdnd11an1n04x5 FILLER_330_2269 ();
 b15zdnd00an1n02x5 FILLER_330_2273 ();
 b15zdnd00an1n01x5 FILLER_330_2275 ();
 b15zdnd11an1n64x5 FILLER_331_0 ();
 b15zdnd11an1n64x5 FILLER_331_64 ();
 b15zdnd11an1n64x5 FILLER_331_128 ();
 b15zdnd11an1n16x5 FILLER_331_192 ();
 b15zdnd11an1n08x5 FILLER_331_208 ();
 b15zdnd11an1n04x5 FILLER_331_216 ();
 b15zdnd11an1n08x5 FILLER_331_229 ();
 b15zdnd11an1n04x5 FILLER_331_252 ();
 b15zdnd11an1n32x5 FILLER_331_272 ();
 b15zdnd11an1n16x5 FILLER_331_304 ();
 b15zdnd11an1n04x5 FILLER_331_320 ();
 b15zdnd00an1n02x5 FILLER_331_324 ();
 b15zdnd11an1n32x5 FILLER_331_330 ();
 b15zdnd11an1n16x5 FILLER_331_362 ();
 b15zdnd11an1n08x5 FILLER_331_378 ();
 b15zdnd00an1n02x5 FILLER_331_386 ();
 b15zdnd00an1n01x5 FILLER_331_388 ();
 b15zdnd11an1n64x5 FILLER_331_413 ();
 b15zdnd11an1n64x5 FILLER_331_477 ();
 b15zdnd11an1n08x5 FILLER_331_541 ();
 b15zdnd11an1n04x5 FILLER_331_549 ();
 b15zdnd00an1n02x5 FILLER_331_553 ();
 b15zdnd00an1n01x5 FILLER_331_555 ();
 b15zdnd11an1n04x5 FILLER_331_566 ();
 b15zdnd11an1n64x5 FILLER_331_582 ();
 b15zdnd11an1n32x5 FILLER_331_646 ();
 b15zdnd11an1n08x5 FILLER_331_678 ();
 b15zdnd11an1n64x5 FILLER_331_702 ();
 b15zdnd11an1n08x5 FILLER_331_766 ();
 b15zdnd00an1n02x5 FILLER_331_774 ();
 b15zdnd11an1n04x5 FILLER_331_788 ();
 b15zdnd11an1n04x5 FILLER_331_803 ();
 b15zdnd11an1n64x5 FILLER_331_812 ();
 b15zdnd11an1n04x5 FILLER_331_876 ();
 b15zdnd00an1n01x5 FILLER_331_880 ();
 b15zdnd11an1n04x5 FILLER_331_886 ();
 b15zdnd11an1n08x5 FILLER_331_902 ();
 b15zdnd11an1n04x5 FILLER_331_910 ();
 b15zdnd00an1n02x5 FILLER_331_914 ();
 b15zdnd00an1n01x5 FILLER_331_916 ();
 b15zdnd11an1n32x5 FILLER_331_935 ();
 b15zdnd11an1n16x5 FILLER_331_967 ();
 b15zdnd11an1n04x5 FILLER_331_983 ();
 b15zdnd00an1n02x5 FILLER_331_987 ();
 b15zdnd00an1n01x5 FILLER_331_989 ();
 b15zdnd11an1n32x5 FILLER_331_998 ();
 b15zdnd11an1n04x5 FILLER_331_1030 ();
 b15zdnd00an1n02x5 FILLER_331_1034 ();
 b15zdnd00an1n01x5 FILLER_331_1036 ();
 b15zdnd11an1n04x5 FILLER_331_1041 ();
 b15zdnd11an1n04x5 FILLER_331_1063 ();
 b15zdnd11an1n32x5 FILLER_331_1093 ();
 b15zdnd11an1n08x5 FILLER_331_1129 ();
 b15zdnd11an1n04x5 FILLER_331_1137 ();
 b15zdnd00an1n02x5 FILLER_331_1141 ();
 b15zdnd11an1n64x5 FILLER_331_1147 ();
 b15zdnd11an1n16x5 FILLER_331_1211 ();
 b15zdnd00an1n01x5 FILLER_331_1227 ();
 b15zdnd11an1n64x5 FILLER_331_1232 ();
 b15zdnd11an1n32x5 FILLER_331_1296 ();
 b15zdnd11an1n16x5 FILLER_331_1328 ();
 b15zdnd11an1n08x5 FILLER_331_1344 ();
 b15zdnd11an1n04x5 FILLER_331_1352 ();
 b15zdnd00an1n01x5 FILLER_331_1356 ();
 b15zdnd11an1n04x5 FILLER_331_1369 ();
 b15zdnd11an1n08x5 FILLER_331_1389 ();
 b15zdnd11an1n04x5 FILLER_331_1397 ();
 b15zdnd00an1n02x5 FILLER_331_1401 ();
 b15zdnd00an1n01x5 FILLER_331_1403 ();
 b15zdnd11an1n08x5 FILLER_331_1410 ();
 b15zdnd11an1n04x5 FILLER_331_1418 ();
 b15zdnd00an1n02x5 FILLER_331_1422 ();
 b15zdnd00an1n01x5 FILLER_331_1424 ();
 b15zdnd11an1n16x5 FILLER_331_1445 ();
 b15zdnd11an1n04x5 FILLER_331_1461 ();
 b15zdnd00an1n02x5 FILLER_331_1465 ();
 b15zdnd00an1n01x5 FILLER_331_1467 ();
 b15zdnd11an1n08x5 FILLER_331_1482 ();
 b15zdnd00an1n01x5 FILLER_331_1490 ();
 b15zdnd11an1n08x5 FILLER_331_1508 ();
 b15zdnd00an1n01x5 FILLER_331_1516 ();
 b15zdnd11an1n04x5 FILLER_331_1523 ();
 b15zdnd00an1n01x5 FILLER_331_1527 ();
 b15zdnd11an1n16x5 FILLER_331_1532 ();
 b15zdnd11an1n08x5 FILLER_331_1548 ();
 b15zdnd11an1n32x5 FILLER_331_1566 ();
 b15zdnd11an1n16x5 FILLER_331_1598 ();
 b15zdnd11an1n32x5 FILLER_331_1628 ();
 b15zdnd11an1n16x5 FILLER_331_1660 ();
 b15zdnd11an1n08x5 FILLER_331_1676 ();
 b15zdnd11an1n04x5 FILLER_331_1684 ();
 b15zdnd00an1n01x5 FILLER_331_1688 ();
 b15zdnd11an1n04x5 FILLER_331_1693 ();
 b15zdnd00an1n02x5 FILLER_331_1697 ();
 b15zdnd11an1n32x5 FILLER_331_1706 ();
 b15zdnd11an1n04x5 FILLER_331_1738 ();
 b15zdnd00an1n02x5 FILLER_331_1742 ();
 b15zdnd00an1n01x5 FILLER_331_1744 ();
 b15zdnd11an1n08x5 FILLER_331_1749 ();
 b15zdnd00an1n02x5 FILLER_331_1757 ();
 b15zdnd00an1n01x5 FILLER_331_1759 ();
 b15zdnd11an1n16x5 FILLER_331_1786 ();
 b15zdnd11an1n08x5 FILLER_331_1823 ();
 b15zdnd11an1n04x5 FILLER_331_1831 ();
 b15zdnd11an1n16x5 FILLER_331_1851 ();
 b15zdnd11an1n08x5 FILLER_331_1867 ();
 b15zdnd00an1n02x5 FILLER_331_1875 ();
 b15zdnd00an1n01x5 FILLER_331_1877 ();
 b15zdnd11an1n04x5 FILLER_331_1890 ();
 b15zdnd11an1n16x5 FILLER_331_1925 ();
 b15zdnd00an1n02x5 FILLER_331_1941 ();
 b15zdnd00an1n01x5 FILLER_331_1943 ();
 b15zdnd11an1n08x5 FILLER_331_1949 ();
 b15zdnd11an1n04x5 FILLER_331_1957 ();
 b15zdnd00an1n01x5 FILLER_331_1961 ();
 b15zdnd11an1n08x5 FILLER_331_1967 ();
 b15zdnd00an1n02x5 FILLER_331_1975 ();
 b15zdnd00an1n01x5 FILLER_331_1977 ();
 b15zdnd11an1n32x5 FILLER_331_1993 ();
 b15zdnd11an1n16x5 FILLER_331_2025 ();
 b15zdnd00an1n01x5 FILLER_331_2041 ();
 b15zdnd11an1n08x5 FILLER_331_2049 ();
 b15zdnd00an1n02x5 FILLER_331_2057 ();
 b15zdnd00an1n01x5 FILLER_331_2059 ();
 b15zdnd11an1n16x5 FILLER_331_2068 ();
 b15zdnd11an1n08x5 FILLER_331_2084 ();
 b15zdnd00an1n02x5 FILLER_331_2092 ();
 b15zdnd00an1n01x5 FILLER_331_2094 ();
 b15zdnd11an1n04x5 FILLER_331_2104 ();
 b15zdnd11an1n08x5 FILLER_331_2119 ();
 b15zdnd11an1n04x5 FILLER_331_2127 ();
 b15zdnd11an1n16x5 FILLER_331_2136 ();
 b15zdnd11an1n04x5 FILLER_331_2152 ();
 b15zdnd11an1n04x5 FILLER_331_2162 ();
 b15zdnd00an1n02x5 FILLER_331_2166 ();
 b15zdnd11an1n08x5 FILLER_331_2194 ();
 b15zdnd00an1n02x5 FILLER_331_2202 ();
 b15zdnd11an1n04x5 FILLER_331_2209 ();
 b15zdnd00an1n02x5 FILLER_331_2213 ();
 b15zdnd11an1n04x5 FILLER_331_2221 ();
 b15zdnd11an1n32x5 FILLER_331_2231 ();
 b15zdnd11an1n16x5 FILLER_331_2263 ();
 b15zdnd11an1n04x5 FILLER_331_2279 ();
 b15zdnd00an1n01x5 FILLER_331_2283 ();
 b15zdnd11an1n64x5 FILLER_332_8 ();
 b15zdnd11an1n64x5 FILLER_332_72 ();
 b15zdnd11an1n64x5 FILLER_332_136 ();
 b15zdnd11an1n32x5 FILLER_332_200 ();
 b15zdnd11an1n16x5 FILLER_332_232 ();
 b15zdnd11an1n04x5 FILLER_332_248 ();
 b15zdnd11an1n16x5 FILLER_332_256 ();
 b15zdnd11an1n16x5 FILLER_332_278 ();
 b15zdnd11an1n08x5 FILLER_332_294 ();
 b15zdnd11an1n04x5 FILLER_332_302 ();
 b15zdnd00an1n01x5 FILLER_332_306 ();
 b15zdnd11an1n08x5 FILLER_332_311 ();
 b15zdnd11an1n04x5 FILLER_332_319 ();
 b15zdnd00an1n02x5 FILLER_332_323 ();
 b15zdnd00an1n01x5 FILLER_332_325 ();
 b15zdnd11an1n64x5 FILLER_332_335 ();
 b15zdnd11an1n32x5 FILLER_332_399 ();
 b15zdnd11an1n16x5 FILLER_332_431 ();
 b15zdnd11an1n04x5 FILLER_332_447 ();
 b15zdnd00an1n02x5 FILLER_332_451 ();
 b15zdnd00an1n01x5 FILLER_332_453 ();
 b15zdnd11an1n64x5 FILLER_332_460 ();
 b15zdnd11an1n16x5 FILLER_332_524 ();
 b15zdnd11an1n08x5 FILLER_332_540 ();
 b15zdnd11an1n04x5 FILLER_332_548 ();
 b15zdnd00an1n02x5 FILLER_332_552 ();
 b15zdnd11an1n04x5 FILLER_332_568 ();
 b15zdnd11an1n04x5 FILLER_332_578 ();
 b15zdnd11an1n08x5 FILLER_332_602 ();
 b15zdnd11an1n32x5 FILLER_332_616 ();
 b15zdnd11an1n16x5 FILLER_332_648 ();
 b15zdnd11an1n08x5 FILLER_332_664 ();
 b15zdnd00an1n01x5 FILLER_332_672 ();
 b15zdnd11an1n04x5 FILLER_332_677 ();
 b15zdnd11an1n32x5 FILLER_332_686 ();
 b15zdnd11an1n04x5 FILLER_332_726 ();
 b15zdnd00an1n02x5 FILLER_332_730 ();
 b15zdnd00an1n01x5 FILLER_332_732 ();
 b15zdnd11an1n64x5 FILLER_332_743 ();
 b15zdnd11an1n08x5 FILLER_332_807 ();
 b15zdnd11an1n04x5 FILLER_332_815 ();
 b15zdnd00an1n02x5 FILLER_332_819 ();
 b15zdnd11an1n16x5 FILLER_332_833 ();
 b15zdnd11an1n08x5 FILLER_332_849 ();
 b15zdnd00an1n02x5 FILLER_332_857 ();
 b15zdnd00an1n01x5 FILLER_332_859 ();
 b15zdnd11an1n04x5 FILLER_332_866 ();
 b15zdnd00an1n01x5 FILLER_332_870 ();
 b15zdnd11an1n32x5 FILLER_332_877 ();
 b15zdnd11an1n08x5 FILLER_332_909 ();
 b15zdnd11an1n64x5 FILLER_332_949 ();
 b15zdnd11an1n08x5 FILLER_332_1013 ();
 b15zdnd11an1n04x5 FILLER_332_1021 ();
 b15zdnd00an1n02x5 FILLER_332_1025 ();
 b15zdnd00an1n01x5 FILLER_332_1027 ();
 b15zdnd11an1n04x5 FILLER_332_1032 ();
 b15zdnd11an1n32x5 FILLER_332_1043 ();
 b15zdnd11an1n16x5 FILLER_332_1075 ();
 b15zdnd00an1n02x5 FILLER_332_1091 ();
 b15zdnd11an1n64x5 FILLER_332_1116 ();
 b15zdnd11an1n64x5 FILLER_332_1180 ();
 b15zdnd11an1n64x5 FILLER_332_1244 ();
 b15zdnd11an1n16x5 FILLER_332_1308 ();
 b15zdnd00an1n01x5 FILLER_332_1324 ();
 b15zdnd11an1n04x5 FILLER_332_1341 ();
 b15zdnd11an1n08x5 FILLER_332_1371 ();
 b15zdnd11an1n04x5 FILLER_332_1379 ();
 b15zdnd00an1n01x5 FILLER_332_1383 ();
 b15zdnd11an1n32x5 FILLER_332_1398 ();
 b15zdnd11an1n04x5 FILLER_332_1430 ();
 b15zdnd00an1n02x5 FILLER_332_1434 ();
 b15zdnd11an1n08x5 FILLER_332_1444 ();
 b15zdnd11an1n04x5 FILLER_332_1452 ();
 b15zdnd00an1n02x5 FILLER_332_1456 ();
 b15zdnd00an1n01x5 FILLER_332_1458 ();
 b15zdnd11an1n64x5 FILLER_332_1464 ();
 b15zdnd11an1n16x5 FILLER_332_1528 ();
 b15zdnd11an1n08x5 FILLER_332_1550 ();
 b15zdnd00an1n02x5 FILLER_332_1558 ();
 b15zdnd11an1n64x5 FILLER_332_1567 ();
 b15zdnd11an1n32x5 FILLER_332_1631 ();
 b15zdnd11an1n08x5 FILLER_332_1663 ();
 b15zdnd00an1n02x5 FILLER_332_1671 ();
 b15zdnd00an1n01x5 FILLER_332_1673 ();
 b15zdnd11an1n32x5 FILLER_332_1692 ();
 b15zdnd11an1n08x5 FILLER_332_1724 ();
 b15zdnd00an1n02x5 FILLER_332_1732 ();
 b15zdnd11an1n32x5 FILLER_332_1744 ();
 b15zdnd11an1n16x5 FILLER_332_1776 ();
 b15zdnd11an1n04x5 FILLER_332_1792 ();
 b15zdnd00an1n02x5 FILLER_332_1796 ();
 b15zdnd00an1n01x5 FILLER_332_1798 ();
 b15zdnd11an1n32x5 FILLER_332_1825 ();
 b15zdnd11an1n16x5 FILLER_332_1857 ();
 b15zdnd11an1n08x5 FILLER_332_1873 ();
 b15zdnd11an1n04x5 FILLER_332_1881 ();
 b15zdnd00an1n01x5 FILLER_332_1885 ();
 b15zdnd11an1n32x5 FILLER_332_1895 ();
 b15zdnd11an1n08x5 FILLER_332_1927 ();
 b15zdnd11an1n04x5 FILLER_332_1935 ();
 b15zdnd00an1n02x5 FILLER_332_1939 ();
 b15zdnd11an1n08x5 FILLER_332_1947 ();
 b15zdnd11an1n08x5 FILLER_332_1965 ();
 b15zdnd00an1n02x5 FILLER_332_1973 ();
 b15zdnd11an1n04x5 FILLER_332_1979 ();
 b15zdnd11an1n64x5 FILLER_332_1998 ();
 b15zdnd11an1n64x5 FILLER_332_2062 ();
 b15zdnd11an1n16x5 FILLER_332_2126 ();
 b15zdnd11an1n08x5 FILLER_332_2142 ();
 b15zdnd11an1n04x5 FILLER_332_2150 ();
 b15zdnd11an1n04x5 FILLER_332_2162 ();
 b15zdnd00an1n01x5 FILLER_332_2166 ();
 b15zdnd11an1n04x5 FILLER_332_2179 ();
 b15zdnd11an1n04x5 FILLER_332_2215 ();
 b15zdnd11an1n32x5 FILLER_332_2224 ();
 b15zdnd11an1n16x5 FILLER_332_2256 ();
 b15zdnd11an1n04x5 FILLER_332_2272 ();
 b15zdnd11an1n64x5 FILLER_333_0 ();
 b15zdnd11an1n64x5 FILLER_333_64 ();
 b15zdnd11an1n64x5 FILLER_333_128 ();
 b15zdnd11an1n08x5 FILLER_333_192 ();
 b15zdnd11an1n04x5 FILLER_333_200 ();
 b15zdnd00an1n01x5 FILLER_333_204 ();
 b15zdnd11an1n04x5 FILLER_333_221 ();
 b15zdnd11an1n04x5 FILLER_333_234 ();
 b15zdnd11an1n04x5 FILLER_333_253 ();
 b15zdnd00an1n02x5 FILLER_333_257 ();
 b15zdnd00an1n01x5 FILLER_333_259 ();
 b15zdnd11an1n04x5 FILLER_333_269 ();
 b15zdnd11an1n64x5 FILLER_333_279 ();
 b15zdnd11an1n08x5 FILLER_333_343 ();
 b15zdnd11an1n04x5 FILLER_333_351 ();
 b15zdnd00an1n02x5 FILLER_333_355 ();
 b15zdnd11an1n04x5 FILLER_333_367 ();
 b15zdnd11an1n64x5 FILLER_333_377 ();
 b15zdnd00an1n02x5 FILLER_333_441 ();
 b15zdnd00an1n01x5 FILLER_333_443 ();
 b15zdnd11an1n08x5 FILLER_333_456 ();
 b15zdnd00an1n01x5 FILLER_333_464 ();
 b15zdnd11an1n04x5 FILLER_333_478 ();
 b15zdnd11an1n16x5 FILLER_333_494 ();
 b15zdnd11an1n32x5 FILLER_333_517 ();
 b15zdnd11an1n08x5 FILLER_333_549 ();
 b15zdnd00an1n01x5 FILLER_333_557 ();
 b15zdnd11an1n64x5 FILLER_333_563 ();
 b15zdnd11an1n08x5 FILLER_333_627 ();
 b15zdnd11an1n04x5 FILLER_333_635 ();
 b15zdnd00an1n02x5 FILLER_333_639 ();
 b15zdnd11an1n64x5 FILLER_333_664 ();
 b15zdnd11an1n64x5 FILLER_333_728 ();
 b15zdnd11an1n32x5 FILLER_333_792 ();
 b15zdnd11an1n16x5 FILLER_333_824 ();
 b15zdnd11an1n04x5 FILLER_333_840 ();
 b15zdnd11an1n08x5 FILLER_333_860 ();
 b15zdnd00an1n01x5 FILLER_333_868 ();
 b15zdnd11an1n32x5 FILLER_333_878 ();
 b15zdnd11an1n04x5 FILLER_333_910 ();
 b15zdnd00an1n01x5 FILLER_333_914 ();
 b15zdnd11an1n32x5 FILLER_333_923 ();
 b15zdnd11an1n08x5 FILLER_333_955 ();
 b15zdnd00an1n01x5 FILLER_333_963 ();
 b15zdnd11an1n16x5 FILLER_333_981 ();
 b15zdnd11an1n08x5 FILLER_333_997 ();
 b15zdnd11an1n04x5 FILLER_333_1005 ();
 b15zdnd00an1n01x5 FILLER_333_1009 ();
 b15zdnd11an1n16x5 FILLER_333_1014 ();
 b15zdnd11an1n08x5 FILLER_333_1030 ();
 b15zdnd11an1n04x5 FILLER_333_1038 ();
 b15zdnd00an1n02x5 FILLER_333_1042 ();
 b15zdnd11an1n16x5 FILLER_333_1062 ();
 b15zdnd11an1n04x5 FILLER_333_1078 ();
 b15zdnd00an1n02x5 FILLER_333_1082 ();
 b15zdnd11an1n08x5 FILLER_333_1110 ();
 b15zdnd00an1n01x5 FILLER_333_1118 ();
 b15zdnd11an1n08x5 FILLER_333_1150 ();
 b15zdnd00an1n01x5 FILLER_333_1158 ();
 b15zdnd11an1n64x5 FILLER_333_1175 ();
 b15zdnd11an1n16x5 FILLER_333_1239 ();
 b15zdnd11an1n08x5 FILLER_333_1255 ();
 b15zdnd00an1n02x5 FILLER_333_1263 ();
 b15zdnd11an1n08x5 FILLER_333_1291 ();
 b15zdnd00an1n02x5 FILLER_333_1299 ();
 b15zdnd11an1n04x5 FILLER_333_1326 ();
 b15zdnd11an1n64x5 FILLER_333_1334 ();
 b15zdnd11an1n64x5 FILLER_333_1398 ();
 b15zdnd11an1n64x5 FILLER_333_1462 ();
 b15zdnd11an1n64x5 FILLER_333_1526 ();
 b15zdnd11an1n16x5 FILLER_333_1590 ();
 b15zdnd11an1n08x5 FILLER_333_1606 ();
 b15zdnd00an1n01x5 FILLER_333_1614 ();
 b15zdnd11an1n16x5 FILLER_333_1625 ();
 b15zdnd11an1n08x5 FILLER_333_1641 ();
 b15zdnd00an1n02x5 FILLER_333_1649 ();
 b15zdnd00an1n01x5 FILLER_333_1651 ();
 b15zdnd11an1n64x5 FILLER_333_1664 ();
 b15zdnd11an1n64x5 FILLER_333_1728 ();
 b15zdnd11an1n32x5 FILLER_333_1792 ();
 b15zdnd11an1n16x5 FILLER_333_1824 ();
 b15zdnd11an1n04x5 FILLER_333_1852 ();
 b15zdnd00an1n01x5 FILLER_333_1856 ();
 b15zdnd11an1n04x5 FILLER_333_1881 ();
 b15zdnd11an1n32x5 FILLER_333_1895 ();
 b15zdnd11an1n16x5 FILLER_333_1927 ();
 b15zdnd00an1n02x5 FILLER_333_1943 ();
 b15zdnd11an1n04x5 FILLER_333_1950 ();
 b15zdnd11an1n32x5 FILLER_333_1960 ();
 b15zdnd11an1n16x5 FILLER_333_1992 ();
 b15zdnd11an1n04x5 FILLER_333_2008 ();
 b15zdnd00an1n01x5 FILLER_333_2012 ();
 b15zdnd11an1n64x5 FILLER_333_2022 ();
 b15zdnd11an1n64x5 FILLER_333_2086 ();
 b15zdnd11an1n64x5 FILLER_333_2150 ();
 b15zdnd11an1n64x5 FILLER_333_2214 ();
 b15zdnd11an1n04x5 FILLER_333_2278 ();
 b15zdnd00an1n02x5 FILLER_333_2282 ();
 b15zdnd11an1n64x5 FILLER_334_8 ();
 b15zdnd11an1n64x5 FILLER_334_72 ();
 b15zdnd11an1n64x5 FILLER_334_136 ();
 b15zdnd11an1n16x5 FILLER_334_200 ();
 b15zdnd00an1n02x5 FILLER_334_216 ();
 b15zdnd00an1n01x5 FILLER_334_218 ();
 b15zdnd11an1n64x5 FILLER_334_229 ();
 b15zdnd11an1n16x5 FILLER_334_293 ();
 b15zdnd00an1n01x5 FILLER_334_309 ();
 b15zdnd11an1n64x5 FILLER_334_320 ();
 b15zdnd11an1n64x5 FILLER_334_384 ();
 b15zdnd11an1n08x5 FILLER_334_448 ();
 b15zdnd11an1n04x5 FILLER_334_456 ();
 b15zdnd11an1n16x5 FILLER_334_465 ();
 b15zdnd11an1n08x5 FILLER_334_481 ();
 b15zdnd11an1n64x5 FILLER_334_495 ();
 b15zdnd11an1n64x5 FILLER_334_559 ();
 b15zdnd11an1n32x5 FILLER_334_623 ();
 b15zdnd00an1n02x5 FILLER_334_655 ();
 b15zdnd00an1n01x5 FILLER_334_657 ();
 b15zdnd11an1n04x5 FILLER_334_664 ();
 b15zdnd11an1n04x5 FILLER_334_673 ();
 b15zdnd11an1n32x5 FILLER_334_684 ();
 b15zdnd00an1n02x5 FILLER_334_716 ();
 b15zdnd11an1n04x5 FILLER_334_726 ();
 b15zdnd11an1n64x5 FILLER_334_739 ();
 b15zdnd11an1n16x5 FILLER_334_803 ();
 b15zdnd00an1n02x5 FILLER_334_819 ();
 b15zdnd11an1n32x5 FILLER_334_836 ();
 b15zdnd11an1n16x5 FILLER_334_868 ();
 b15zdnd11an1n04x5 FILLER_334_884 ();
 b15zdnd00an1n02x5 FILLER_334_888 ();
 b15zdnd11an1n16x5 FILLER_334_902 ();
 b15zdnd00an1n01x5 FILLER_334_918 ();
 b15zdnd11an1n32x5 FILLER_334_926 ();
 b15zdnd11an1n04x5 FILLER_334_958 ();
 b15zdnd00an1n02x5 FILLER_334_962 ();
 b15zdnd11an1n04x5 FILLER_334_978 ();
 b15zdnd00an1n02x5 FILLER_334_982 ();
 b15zdnd11an1n08x5 FILLER_334_996 ();
 b15zdnd00an1n02x5 FILLER_334_1004 ();
 b15zdnd00an1n01x5 FILLER_334_1006 ();
 b15zdnd11an1n04x5 FILLER_334_1028 ();
 b15zdnd00an1n02x5 FILLER_334_1032 ();
 b15zdnd11an1n08x5 FILLER_334_1043 ();
 b15zdnd11an1n04x5 FILLER_334_1051 ();
 b15zdnd11an1n04x5 FILLER_334_1067 ();
 b15zdnd11an1n32x5 FILLER_334_1076 ();
 b15zdnd11an1n08x5 FILLER_334_1108 ();
 b15zdnd00an1n02x5 FILLER_334_1116 ();
 b15zdnd00an1n01x5 FILLER_334_1118 ();
 b15zdnd11an1n64x5 FILLER_334_1126 ();
 b15zdnd11an1n08x5 FILLER_334_1190 ();
 b15zdnd00an1n01x5 FILLER_334_1198 ();
 b15zdnd11an1n32x5 FILLER_334_1206 ();
 b15zdnd11an1n04x5 FILLER_334_1238 ();
 b15zdnd11an1n08x5 FILLER_334_1262 ();
 b15zdnd00an1n02x5 FILLER_334_1270 ();
 b15zdnd00an1n01x5 FILLER_334_1272 ();
 b15zdnd11an1n64x5 FILLER_334_1286 ();
 b15zdnd11an1n16x5 FILLER_334_1350 ();
 b15zdnd00an1n02x5 FILLER_334_1366 ();
 b15zdnd11an1n16x5 FILLER_334_1384 ();
 b15zdnd11an1n08x5 FILLER_334_1400 ();
 b15zdnd11an1n04x5 FILLER_334_1408 ();
 b15zdnd00an1n02x5 FILLER_334_1412 ();
 b15zdnd11an1n32x5 FILLER_334_1418 ();
 b15zdnd11an1n04x5 FILLER_334_1450 ();
 b15zdnd00an1n02x5 FILLER_334_1454 ();
 b15zdnd00an1n01x5 FILLER_334_1456 ();
 b15zdnd11an1n32x5 FILLER_334_1461 ();
 b15zdnd11an1n16x5 FILLER_334_1493 ();
 b15zdnd11an1n64x5 FILLER_334_1523 ();
 b15zdnd11an1n08x5 FILLER_334_1587 ();
 b15zdnd00an1n02x5 FILLER_334_1595 ();
 b15zdnd00an1n01x5 FILLER_334_1597 ();
 b15zdnd11an1n32x5 FILLER_334_1602 ();
 b15zdnd00an1n02x5 FILLER_334_1634 ();
 b15zdnd00an1n01x5 FILLER_334_1636 ();
 b15zdnd11an1n04x5 FILLER_334_1658 ();
 b15zdnd11an1n16x5 FILLER_334_1668 ();
 b15zdnd11an1n04x5 FILLER_334_1684 ();
 b15zdnd00an1n01x5 FILLER_334_1688 ();
 b15zdnd11an1n08x5 FILLER_334_1693 ();
 b15zdnd11an1n04x5 FILLER_334_1701 ();
 b15zdnd00an1n01x5 FILLER_334_1705 ();
 b15zdnd11an1n08x5 FILLER_334_1714 ();
 b15zdnd11an1n04x5 FILLER_334_1722 ();
 b15zdnd00an1n02x5 FILLER_334_1726 ();
 b15zdnd11an1n32x5 FILLER_334_1744 ();
 b15zdnd11an1n16x5 FILLER_334_1776 ();
 b15zdnd11an1n08x5 FILLER_334_1792 ();
 b15zdnd00an1n02x5 FILLER_334_1800 ();
 b15zdnd11an1n04x5 FILLER_334_1822 ();
 b15zdnd00an1n01x5 FILLER_334_1826 ();
 b15zdnd11an1n04x5 FILLER_334_1837 ();
 b15zdnd11an1n04x5 FILLER_334_1846 ();
 b15zdnd11an1n32x5 FILLER_334_1863 ();
 b15zdnd11an1n08x5 FILLER_334_1895 ();
 b15zdnd00an1n02x5 FILLER_334_1903 ();
 b15zdnd00an1n01x5 FILLER_334_1905 ();
 b15zdnd11an1n32x5 FILLER_334_1912 ();
 b15zdnd00an1n01x5 FILLER_334_1944 ();
 b15zdnd11an1n32x5 FILLER_334_1952 ();
 b15zdnd11an1n16x5 FILLER_334_1984 ();
 b15zdnd11an1n08x5 FILLER_334_2000 ();
 b15zdnd00an1n02x5 FILLER_334_2008 ();
 b15zdnd00an1n01x5 FILLER_334_2010 ();
 b15zdnd11an1n32x5 FILLER_334_2031 ();
 b15zdnd11an1n16x5 FILLER_334_2063 ();
 b15zdnd11an1n08x5 FILLER_334_2079 ();
 b15zdnd00an1n02x5 FILLER_334_2087 ();
 b15zdnd11an1n32x5 FILLER_334_2105 ();
 b15zdnd11an1n16x5 FILLER_334_2137 ();
 b15zdnd00an1n01x5 FILLER_334_2153 ();
 b15zdnd00an1n02x5 FILLER_334_2162 ();
 b15zdnd11an1n64x5 FILLER_334_2190 ();
 b15zdnd11an1n16x5 FILLER_334_2254 ();
 b15zdnd11an1n04x5 FILLER_334_2270 ();
 b15zdnd00an1n02x5 FILLER_334_2274 ();
 b15zdnd11an1n64x5 FILLER_335_0 ();
 b15zdnd11an1n64x5 FILLER_335_64 ();
 b15zdnd11an1n64x5 FILLER_335_128 ();
 b15zdnd11an1n32x5 FILLER_335_192 ();
 b15zdnd11an1n04x5 FILLER_335_224 ();
 b15zdnd11an1n32x5 FILLER_335_244 ();
 b15zdnd11an1n16x5 FILLER_335_276 ();
 b15zdnd11an1n08x5 FILLER_335_292 ();
 b15zdnd11an1n04x5 FILLER_335_300 ();
 b15zdnd00an1n01x5 FILLER_335_304 ();
 b15zdnd11an1n16x5 FILLER_335_315 ();
 b15zdnd11an1n08x5 FILLER_335_331 ();
 b15zdnd00an1n01x5 FILLER_335_339 ();
 b15zdnd11an1n32x5 FILLER_335_345 ();
 b15zdnd11an1n16x5 FILLER_335_377 ();
 b15zdnd11an1n08x5 FILLER_335_393 ();
 b15zdnd11an1n04x5 FILLER_335_401 ();
 b15zdnd00an1n02x5 FILLER_335_405 ();
 b15zdnd00an1n01x5 FILLER_335_407 ();
 b15zdnd11an1n08x5 FILLER_335_420 ();
 b15zdnd11an1n04x5 FILLER_335_428 ();
 b15zdnd00an1n02x5 FILLER_335_432 ();
 b15zdnd00an1n01x5 FILLER_335_434 ();
 b15zdnd11an1n16x5 FILLER_335_445 ();
 b15zdnd11an1n08x5 FILLER_335_461 ();
 b15zdnd11an1n04x5 FILLER_335_469 ();
 b15zdnd00an1n01x5 FILLER_335_473 ();
 b15zdnd11an1n08x5 FILLER_335_482 ();
 b15zdnd11an1n04x5 FILLER_335_490 ();
 b15zdnd11an1n08x5 FILLER_335_498 ();
 b15zdnd00an1n02x5 FILLER_335_506 ();
 b15zdnd11an1n16x5 FILLER_335_515 ();
 b15zdnd11an1n08x5 FILLER_335_531 ();
 b15zdnd11an1n04x5 FILLER_335_539 ();
 b15zdnd00an1n01x5 FILLER_335_543 ();
 b15zdnd11an1n64x5 FILLER_335_555 ();
 b15zdnd11an1n16x5 FILLER_335_619 ();
 b15zdnd11an1n08x5 FILLER_335_635 ();
 b15zdnd11an1n04x5 FILLER_335_643 ();
 b15zdnd00an1n02x5 FILLER_335_647 ();
 b15zdnd00an1n01x5 FILLER_335_649 ();
 b15zdnd11an1n08x5 FILLER_335_662 ();
 b15zdnd11an1n04x5 FILLER_335_670 ();
 b15zdnd11an1n32x5 FILLER_335_679 ();
 b15zdnd11an1n16x5 FILLER_335_711 ();
 b15zdnd11an1n08x5 FILLER_335_727 ();
 b15zdnd00an1n02x5 FILLER_335_735 ();
 b15zdnd11an1n04x5 FILLER_335_749 ();
 b15zdnd11an1n04x5 FILLER_335_758 ();
 b15zdnd11an1n04x5 FILLER_335_769 ();
 b15zdnd11an1n64x5 FILLER_335_778 ();
 b15zdnd11an1n64x5 FILLER_335_842 ();
 b15zdnd11an1n32x5 FILLER_335_906 ();
 b15zdnd11an1n16x5 FILLER_335_938 ();
 b15zdnd11an1n08x5 FILLER_335_954 ();
 b15zdnd11an1n04x5 FILLER_335_962 ();
 b15zdnd00an1n02x5 FILLER_335_966 ();
 b15zdnd11an1n64x5 FILLER_335_984 ();
 b15zdnd11an1n64x5 FILLER_335_1048 ();
 b15zdnd00an1n01x5 FILLER_335_1112 ();
 b15zdnd11an1n32x5 FILLER_335_1125 ();
 b15zdnd11an1n08x5 FILLER_335_1157 ();
 b15zdnd11an1n04x5 FILLER_335_1165 ();
 b15zdnd00an1n02x5 FILLER_335_1169 ();
 b15zdnd11an1n04x5 FILLER_335_1203 ();
 b15zdnd00an1n01x5 FILLER_335_1207 ();
 b15zdnd11an1n08x5 FILLER_335_1226 ();
 b15zdnd11an1n04x5 FILLER_335_1234 ();
 b15zdnd11an1n04x5 FILLER_335_1248 ();
 b15zdnd00an1n02x5 FILLER_335_1252 ();
 b15zdnd11an1n04x5 FILLER_335_1263 ();
 b15zdnd00an1n01x5 FILLER_335_1267 ();
 b15zdnd11an1n08x5 FILLER_335_1272 ();
 b15zdnd00an1n02x5 FILLER_335_1280 ();
 b15zdnd00an1n01x5 FILLER_335_1282 ();
 b15zdnd11an1n64x5 FILLER_335_1289 ();
 b15zdnd11an1n04x5 FILLER_335_1353 ();
 b15zdnd00an1n02x5 FILLER_335_1357 ();
 b15zdnd00an1n01x5 FILLER_335_1359 ();
 b15zdnd11an1n04x5 FILLER_335_1372 ();
 b15zdnd11an1n08x5 FILLER_335_1380 ();
 b15zdnd11an1n04x5 FILLER_335_1388 ();
 b15zdnd00an1n02x5 FILLER_335_1392 ();
 b15zdnd11an1n08x5 FILLER_335_1400 ();
 b15zdnd11an1n04x5 FILLER_335_1413 ();
 b15zdnd11an1n08x5 FILLER_335_1422 ();
 b15zdnd11an1n04x5 FILLER_335_1430 ();
 b15zdnd00an1n01x5 FILLER_335_1434 ();
 b15zdnd11an1n08x5 FILLER_335_1440 ();
 b15zdnd00an1n02x5 FILLER_335_1448 ();
 b15zdnd11an1n04x5 FILLER_335_1463 ();
 b15zdnd11an1n64x5 FILLER_335_1472 ();
 b15zdnd11an1n08x5 FILLER_335_1536 ();
 b15zdnd11an1n32x5 FILLER_335_1549 ();
 b15zdnd11an1n08x5 FILLER_335_1581 ();
 b15zdnd11an1n08x5 FILLER_335_1595 ();
 b15zdnd00an1n02x5 FILLER_335_1603 ();
 b15zdnd11an1n16x5 FILLER_335_1614 ();
 b15zdnd11an1n08x5 FILLER_335_1630 ();
 b15zdnd00an1n02x5 FILLER_335_1638 ();
 b15zdnd11an1n08x5 FILLER_335_1652 ();
 b15zdnd11an1n04x5 FILLER_335_1660 ();
 b15zdnd00an1n02x5 FILLER_335_1664 ();
 b15zdnd00an1n01x5 FILLER_335_1666 ();
 b15zdnd11an1n32x5 FILLER_335_1673 ();
 b15zdnd11an1n16x5 FILLER_335_1711 ();
 b15zdnd00an1n02x5 FILLER_335_1727 ();
 b15zdnd00an1n01x5 FILLER_335_1729 ();
 b15zdnd11an1n64x5 FILLER_335_1762 ();
 b15zdnd11an1n08x5 FILLER_335_1826 ();
 b15zdnd11an1n04x5 FILLER_335_1834 ();
 b15zdnd00an1n01x5 FILLER_335_1838 ();
 b15zdnd11an1n16x5 FILLER_335_1849 ();
 b15zdnd11an1n08x5 FILLER_335_1865 ();
 b15zdnd11an1n04x5 FILLER_335_1873 ();
 b15zdnd00an1n01x5 FILLER_335_1877 ();
 b15zdnd11an1n04x5 FILLER_335_1885 ();
 b15zdnd11an1n32x5 FILLER_335_1909 ();
 b15zdnd00an1n01x5 FILLER_335_1941 ();
 b15zdnd11an1n64x5 FILLER_335_1949 ();
 b15zdnd11an1n08x5 FILLER_335_2013 ();
 b15zdnd00an1n01x5 FILLER_335_2021 ();
 b15zdnd11an1n16x5 FILLER_335_2029 ();
 b15zdnd11an1n04x5 FILLER_335_2045 ();
 b15zdnd00an1n02x5 FILLER_335_2049 ();
 b15zdnd11an1n16x5 FILLER_335_2061 ();
 b15zdnd11an1n04x5 FILLER_335_2077 ();
 b15zdnd00an1n01x5 FILLER_335_2081 ();
 b15zdnd11an1n08x5 FILLER_335_2089 ();
 b15zdnd00an1n02x5 FILLER_335_2097 ();
 b15zdnd11an1n04x5 FILLER_335_2117 ();
 b15zdnd11an1n32x5 FILLER_335_2137 ();
 b15zdnd11an1n08x5 FILLER_335_2169 ();
 b15zdnd11an1n64x5 FILLER_335_2183 ();
 b15zdnd11an1n32x5 FILLER_335_2247 ();
 b15zdnd11an1n04x5 FILLER_335_2279 ();
 b15zdnd00an1n01x5 FILLER_335_2283 ();
 b15zdnd11an1n64x5 FILLER_336_8 ();
 b15zdnd11an1n64x5 FILLER_336_72 ();
 b15zdnd11an1n64x5 FILLER_336_136 ();
 b15zdnd11an1n64x5 FILLER_336_200 ();
 b15zdnd00an1n01x5 FILLER_336_264 ();
 b15zdnd11an1n64x5 FILLER_336_269 ();
 b15zdnd11an1n08x5 FILLER_336_333 ();
 b15zdnd11an1n04x5 FILLER_336_341 ();
 b15zdnd00an1n01x5 FILLER_336_345 ();
 b15zdnd11an1n04x5 FILLER_336_353 ();
 b15zdnd11an1n16x5 FILLER_336_369 ();
 b15zdnd11an1n04x5 FILLER_336_385 ();
 b15zdnd11an1n04x5 FILLER_336_396 ();
 b15zdnd00an1n02x5 FILLER_336_400 ();
 b15zdnd00an1n01x5 FILLER_336_402 ();
 b15zdnd11an1n16x5 FILLER_336_410 ();
 b15zdnd11an1n04x5 FILLER_336_426 ();
 b15zdnd00an1n01x5 FILLER_336_430 ();
 b15zdnd11an1n04x5 FILLER_336_438 ();
 b15zdnd00an1n02x5 FILLER_336_442 ();
 b15zdnd11an1n16x5 FILLER_336_470 ();
 b15zdnd11an1n08x5 FILLER_336_498 ();
 b15zdnd00an1n02x5 FILLER_336_506 ();
 b15zdnd00an1n01x5 FILLER_336_508 ();
 b15zdnd11an1n04x5 FILLER_336_521 ();
 b15zdnd11an1n32x5 FILLER_336_539 ();
 b15zdnd11an1n08x5 FILLER_336_571 ();
 b15zdnd11an1n04x5 FILLER_336_579 ();
 b15zdnd00an1n02x5 FILLER_336_583 ();
 b15zdnd11an1n64x5 FILLER_336_591 ();
 b15zdnd00an1n02x5 FILLER_336_655 ();
 b15zdnd00an1n01x5 FILLER_336_657 ();
 b15zdnd11an1n32x5 FILLER_336_669 ();
 b15zdnd00an1n02x5 FILLER_336_701 ();
 b15zdnd11an1n04x5 FILLER_336_713 ();
 b15zdnd00an1n01x5 FILLER_336_717 ();
 b15zdnd11an1n08x5 FILLER_336_726 ();
 b15zdnd00an1n02x5 FILLER_336_734 ();
 b15zdnd00an1n01x5 FILLER_336_736 ();
 b15zdnd11an1n16x5 FILLER_336_742 ();
 b15zdnd11an1n04x5 FILLER_336_758 ();
 b15zdnd00an1n02x5 FILLER_336_762 ();
 b15zdnd11an1n16x5 FILLER_336_773 ();
 b15zdnd11an1n08x5 FILLER_336_789 ();
 b15zdnd00an1n01x5 FILLER_336_797 ();
 b15zdnd11an1n04x5 FILLER_336_803 ();
 b15zdnd11an1n16x5 FILLER_336_813 ();
 b15zdnd00an1n01x5 FILLER_336_829 ();
 b15zdnd11an1n04x5 FILLER_336_845 ();
 b15zdnd11an1n64x5 FILLER_336_856 ();
 b15zdnd11an1n64x5 FILLER_336_920 ();
 b15zdnd11an1n64x5 FILLER_336_984 ();
 b15zdnd11an1n32x5 FILLER_336_1048 ();
 b15zdnd11an1n16x5 FILLER_336_1080 ();
 b15zdnd11an1n08x5 FILLER_336_1096 ();
 b15zdnd11an1n04x5 FILLER_336_1130 ();
 b15zdnd11an1n04x5 FILLER_336_1160 ();
 b15zdnd11an1n04x5 FILLER_336_1190 ();
 b15zdnd11an1n16x5 FILLER_336_1220 ();
 b15zdnd11an1n04x5 FILLER_336_1236 ();
 b15zdnd00an1n02x5 FILLER_336_1240 ();
 b15zdnd11an1n16x5 FILLER_336_1268 ();
 b15zdnd00an1n01x5 FILLER_336_1284 ();
 b15zdnd11an1n08x5 FILLER_336_1290 ();
 b15zdnd11an1n04x5 FILLER_336_1298 ();
 b15zdnd00an1n02x5 FILLER_336_1302 ();
 b15zdnd00an1n01x5 FILLER_336_1304 ();
 b15zdnd11an1n04x5 FILLER_336_1315 ();
 b15zdnd11an1n16x5 FILLER_336_1327 ();
 b15zdnd11an1n08x5 FILLER_336_1343 ();
 b15zdnd00an1n02x5 FILLER_336_1351 ();
 b15zdnd11an1n04x5 FILLER_336_1359 ();
 b15zdnd11an1n08x5 FILLER_336_1383 ();
 b15zdnd00an1n02x5 FILLER_336_1391 ();
 b15zdnd00an1n01x5 FILLER_336_1393 ();
 b15zdnd11an1n08x5 FILLER_336_1398 ();
 b15zdnd11an1n08x5 FILLER_336_1418 ();
 b15zdnd11an1n04x5 FILLER_336_1426 ();
 b15zdnd00an1n02x5 FILLER_336_1430 ();
 b15zdnd11an1n08x5 FILLER_336_1448 ();
 b15zdnd11an1n04x5 FILLER_336_1456 ();
 b15zdnd00an1n02x5 FILLER_336_1460 ();
 b15zdnd11an1n08x5 FILLER_336_1468 ();
 b15zdnd00an1n02x5 FILLER_336_1476 ();
 b15zdnd11an1n04x5 FILLER_336_1489 ();
 b15zdnd11an1n16x5 FILLER_336_1513 ();
 b15zdnd11an1n04x5 FILLER_336_1529 ();
 b15zdnd00an1n02x5 FILLER_336_1533 ();
 b15zdnd11an1n04x5 FILLER_336_1544 ();
 b15zdnd11an1n04x5 FILLER_336_1560 ();
 b15zdnd00an1n02x5 FILLER_336_1564 ();
 b15zdnd11an1n08x5 FILLER_336_1576 ();
 b15zdnd11an1n04x5 FILLER_336_1584 ();
 b15zdnd11an1n04x5 FILLER_336_1600 ();
 b15zdnd11an1n04x5 FILLER_336_1616 ();
 b15zdnd11an1n16x5 FILLER_336_1626 ();
 b15zdnd11an1n16x5 FILLER_336_1654 ();
 b15zdnd11an1n04x5 FILLER_336_1690 ();
 b15zdnd11an1n16x5 FILLER_336_1706 ();
 b15zdnd11an1n08x5 FILLER_336_1722 ();
 b15zdnd00an1n02x5 FILLER_336_1730 ();
 b15zdnd11an1n64x5 FILLER_336_1736 ();
 b15zdnd11an1n16x5 FILLER_336_1800 ();
 b15zdnd00an1n01x5 FILLER_336_1816 ();
 b15zdnd11an1n32x5 FILLER_336_1826 ();
 b15zdnd11an1n08x5 FILLER_336_1858 ();
 b15zdnd11an1n04x5 FILLER_336_1866 ();
 b15zdnd00an1n02x5 FILLER_336_1870 ();
 b15zdnd00an1n01x5 FILLER_336_1872 ();
 b15zdnd11an1n16x5 FILLER_336_1888 ();
 b15zdnd00an1n02x5 FILLER_336_1904 ();
 b15zdnd11an1n16x5 FILLER_336_1912 ();
 b15zdnd11an1n08x5 FILLER_336_1928 ();
 b15zdnd11an1n04x5 FILLER_336_1936 ();
 b15zdnd00an1n02x5 FILLER_336_1940 ();
 b15zdnd11an1n08x5 FILLER_336_1946 ();
 b15zdnd11an1n04x5 FILLER_336_1954 ();
 b15zdnd00an1n01x5 FILLER_336_1958 ();
 b15zdnd11an1n32x5 FILLER_336_1971 ();
 b15zdnd11an1n16x5 FILLER_336_2003 ();
 b15zdnd11an1n08x5 FILLER_336_2019 ();
 b15zdnd11an1n04x5 FILLER_336_2041 ();
 b15zdnd00an1n01x5 FILLER_336_2045 ();
 b15zdnd11an1n32x5 FILLER_336_2056 ();
 b15zdnd00an1n02x5 FILLER_336_2088 ();
 b15zdnd00an1n01x5 FILLER_336_2090 ();
 b15zdnd11an1n16x5 FILLER_336_2105 ();
 b15zdnd11an1n08x5 FILLER_336_2121 ();
 b15zdnd00an1n02x5 FILLER_336_2129 ();
 b15zdnd00an1n02x5 FILLER_336_2152 ();
 b15zdnd11an1n16x5 FILLER_336_2162 ();
 b15zdnd11an1n04x5 FILLER_336_2178 ();
 b15zdnd00an1n02x5 FILLER_336_2182 ();
 b15zdnd00an1n01x5 FILLER_336_2184 ();
 b15zdnd11an1n16x5 FILLER_336_2190 ();
 b15zdnd00an1n02x5 FILLER_336_2206 ();
 b15zdnd00an1n01x5 FILLER_336_2208 ();
 b15zdnd11an1n04x5 FILLER_336_2215 ();
 b15zdnd11an1n32x5 FILLER_336_2224 ();
 b15zdnd11an1n16x5 FILLER_336_2256 ();
 b15zdnd11an1n04x5 FILLER_336_2272 ();
 b15zdnd11an1n64x5 FILLER_337_0 ();
 b15zdnd11an1n64x5 FILLER_337_64 ();
 b15zdnd11an1n64x5 FILLER_337_128 ();
 b15zdnd11an1n64x5 FILLER_337_192 ();
 b15zdnd11an1n04x5 FILLER_337_256 ();
 b15zdnd00an1n02x5 FILLER_337_260 ();
 b15zdnd00an1n01x5 FILLER_337_262 ();
 b15zdnd11an1n64x5 FILLER_337_269 ();
 b15zdnd11an1n04x5 FILLER_337_333 ();
 b15zdnd00an1n02x5 FILLER_337_337 ();
 b15zdnd00an1n01x5 FILLER_337_339 ();
 b15zdnd11an1n04x5 FILLER_337_346 ();
 b15zdnd00an1n01x5 FILLER_337_350 ();
 b15zdnd11an1n04x5 FILLER_337_355 ();
 b15zdnd11an1n04x5 FILLER_337_364 ();
 b15zdnd11an1n08x5 FILLER_337_379 ();
 b15zdnd11an1n04x5 FILLER_337_387 ();
 b15zdnd00an1n01x5 FILLER_337_391 ();
 b15zdnd11an1n64x5 FILLER_337_413 ();
 b15zdnd11an1n08x5 FILLER_337_477 ();
 b15zdnd11an1n04x5 FILLER_337_485 ();
 b15zdnd11an1n08x5 FILLER_337_509 ();
 b15zdnd11an1n04x5 FILLER_337_517 ();
 b15zdnd00an1n02x5 FILLER_337_521 ();
 b15zdnd11an1n16x5 FILLER_337_537 ();
 b15zdnd11an1n08x5 FILLER_337_553 ();
 b15zdnd11an1n04x5 FILLER_337_561 ();
 b15zdnd11an1n64x5 FILLER_337_573 ();
 b15zdnd11an1n16x5 FILLER_337_637 ();
 b15zdnd11an1n04x5 FILLER_337_653 ();
 b15zdnd11an1n32x5 FILLER_337_664 ();
 b15zdnd11an1n08x5 FILLER_337_696 ();
 b15zdnd00an1n02x5 FILLER_337_704 ();
 b15zdnd00an1n01x5 FILLER_337_706 ();
 b15zdnd11an1n16x5 FILLER_337_728 ();
 b15zdnd11an1n08x5 FILLER_337_744 ();
 b15zdnd11an1n04x5 FILLER_337_752 ();
 b15zdnd00an1n02x5 FILLER_337_756 ();
 b15zdnd00an1n01x5 FILLER_337_758 ();
 b15zdnd11an1n16x5 FILLER_337_777 ();
 b15zdnd11an1n08x5 FILLER_337_793 ();
 b15zdnd11an1n04x5 FILLER_337_801 ();
 b15zdnd00an1n02x5 FILLER_337_805 ();
 b15zdnd00an1n01x5 FILLER_337_807 ();
 b15zdnd11an1n08x5 FILLER_337_834 ();
 b15zdnd11an1n04x5 FILLER_337_842 ();
 b15zdnd00an1n02x5 FILLER_337_846 ();
 b15zdnd00an1n01x5 FILLER_337_848 ();
 b15zdnd11an1n08x5 FILLER_337_854 ();
 b15zdnd00an1n01x5 FILLER_337_862 ();
 b15zdnd11an1n16x5 FILLER_337_894 ();
 b15zdnd11an1n04x5 FILLER_337_910 ();
 b15zdnd00an1n02x5 FILLER_337_914 ();
 b15zdnd00an1n01x5 FILLER_337_916 ();
 b15zdnd11an1n04x5 FILLER_337_922 ();
 b15zdnd11an1n16x5 FILLER_337_933 ();
 b15zdnd00an1n02x5 FILLER_337_949 ();
 b15zdnd00an1n01x5 FILLER_337_951 ();
 b15zdnd11an1n16x5 FILLER_337_959 ();
 b15zdnd11an1n16x5 FILLER_337_1007 ();
 b15zdnd00an1n02x5 FILLER_337_1023 ();
 b15zdnd00an1n01x5 FILLER_337_1025 ();
 b15zdnd11an1n32x5 FILLER_337_1036 ();
 b15zdnd11an1n16x5 FILLER_337_1068 ();
 b15zdnd00an1n01x5 FILLER_337_1084 ();
 b15zdnd11an1n08x5 FILLER_337_1105 ();
 b15zdnd00an1n02x5 FILLER_337_1113 ();
 b15zdnd00an1n01x5 FILLER_337_1115 ();
 b15zdnd11an1n04x5 FILLER_337_1133 ();
 b15zdnd00an1n01x5 FILLER_337_1137 ();
 b15zdnd11an1n04x5 FILLER_337_1145 ();
 b15zdnd11an1n16x5 FILLER_337_1163 ();
 b15zdnd11an1n08x5 FILLER_337_1205 ();
 b15zdnd11an1n04x5 FILLER_337_1213 ();
 b15zdnd11an1n08x5 FILLER_337_1223 ();
 b15zdnd00an1n02x5 FILLER_337_1231 ();
 b15zdnd11an1n08x5 FILLER_337_1259 ();
 b15zdnd11an1n04x5 FILLER_337_1267 ();
 b15zdnd00an1n02x5 FILLER_337_1271 ();
 b15zdnd11an1n04x5 FILLER_337_1277 ();
 b15zdnd00an1n02x5 FILLER_337_1281 ();
 b15zdnd00an1n01x5 FILLER_337_1283 ();
 b15zdnd11an1n64x5 FILLER_337_1291 ();
 b15zdnd11an1n32x5 FILLER_337_1355 ();
 b15zdnd11an1n04x5 FILLER_337_1387 ();
 b15zdnd00an1n02x5 FILLER_337_1391 ();
 b15zdnd00an1n01x5 FILLER_337_1393 ();
 b15zdnd11an1n64x5 FILLER_337_1404 ();
 b15zdnd11an1n32x5 FILLER_337_1468 ();
 b15zdnd00an1n01x5 FILLER_337_1500 ();
 b15zdnd11an1n04x5 FILLER_337_1507 ();
 b15zdnd11an1n08x5 FILLER_337_1523 ();
 b15zdnd11an1n04x5 FILLER_337_1531 ();
 b15zdnd00an1n01x5 FILLER_337_1535 ();
 b15zdnd11an1n64x5 FILLER_337_1541 ();
 b15zdnd11an1n64x5 FILLER_337_1605 ();
 b15zdnd11an1n04x5 FILLER_337_1669 ();
 b15zdnd00an1n02x5 FILLER_337_1673 ();
 b15zdnd11an1n16x5 FILLER_337_1679 ();
 b15zdnd00an1n01x5 FILLER_337_1695 ();
 b15zdnd11an1n64x5 FILLER_337_1701 ();
 b15zdnd11an1n32x5 FILLER_337_1765 ();
 b15zdnd11an1n08x5 FILLER_337_1797 ();
 b15zdnd11an1n04x5 FILLER_337_1805 ();
 b15zdnd11an1n04x5 FILLER_337_1827 ();
 b15zdnd11an1n04x5 FILLER_337_1851 ();
 b15zdnd11an1n16x5 FILLER_337_1861 ();
 b15zdnd11an1n08x5 FILLER_337_1877 ();
 b15zdnd00an1n02x5 FILLER_337_1885 ();
 b15zdnd11an1n04x5 FILLER_337_1892 ();
 b15zdnd11an1n08x5 FILLER_337_1902 ();
 b15zdnd11an1n32x5 FILLER_337_1915 ();
 b15zdnd11an1n04x5 FILLER_337_1947 ();
 b15zdnd00an1n02x5 FILLER_337_1951 ();
 b15zdnd00an1n01x5 FILLER_337_1953 ();
 b15zdnd11an1n16x5 FILLER_337_1966 ();
 b15zdnd11an1n08x5 FILLER_337_1982 ();
 b15zdnd11an1n04x5 FILLER_337_1996 ();
 b15zdnd11an1n32x5 FILLER_337_2006 ();
 b15zdnd11an1n08x5 FILLER_337_2038 ();
 b15zdnd11an1n04x5 FILLER_337_2046 ();
 b15zdnd11an1n04x5 FILLER_337_2064 ();
 b15zdnd00an1n01x5 FILLER_337_2068 ();
 b15zdnd11an1n16x5 FILLER_337_2078 ();
 b15zdnd00an1n02x5 FILLER_337_2094 ();
 b15zdnd00an1n01x5 FILLER_337_2096 ();
 b15zdnd11an1n32x5 FILLER_337_2107 ();
 b15zdnd11an1n04x5 FILLER_337_2139 ();
 b15zdnd00an1n02x5 FILLER_337_2143 ();
 b15zdnd11an1n32x5 FILLER_337_2155 ();
 b15zdnd11an1n16x5 FILLER_337_2187 ();
 b15zdnd00an1n01x5 FILLER_337_2203 ();
 b15zdnd11an1n04x5 FILLER_337_2213 ();
 b15zdnd11an1n32x5 FILLER_337_2223 ();
 b15zdnd11an1n16x5 FILLER_337_2255 ();
 b15zdnd11an1n08x5 FILLER_337_2271 ();
 b15zdnd11an1n04x5 FILLER_337_2279 ();
 b15zdnd00an1n01x5 FILLER_337_2283 ();
 b15zdnd11an1n64x5 FILLER_338_8 ();
 b15zdnd11an1n64x5 FILLER_338_72 ();
 b15zdnd11an1n64x5 FILLER_338_136 ();
 b15zdnd11an1n32x5 FILLER_338_200 ();
 b15zdnd11an1n16x5 FILLER_338_232 ();
 b15zdnd00an1n02x5 FILLER_338_248 ();
 b15zdnd00an1n01x5 FILLER_338_250 ();
 b15zdnd11an1n04x5 FILLER_338_255 ();
 b15zdnd11an1n16x5 FILLER_338_273 ();
 b15zdnd00an1n01x5 FILLER_338_289 ();
 b15zdnd11an1n04x5 FILLER_338_300 ();
 b15zdnd11an1n16x5 FILLER_338_317 ();
 b15zdnd11an1n08x5 FILLER_338_333 ();
 b15zdnd00an1n02x5 FILLER_338_341 ();
 b15zdnd11an1n16x5 FILLER_338_357 ();
 b15zdnd00an1n01x5 FILLER_338_373 ();
 b15zdnd11an1n32x5 FILLER_338_395 ();
 b15zdnd11an1n08x5 FILLER_338_427 ();
 b15zdnd00an1n02x5 FILLER_338_435 ();
 b15zdnd00an1n01x5 FILLER_338_437 ();
 b15zdnd11an1n32x5 FILLER_338_444 ();
 b15zdnd11an1n08x5 FILLER_338_476 ();
 b15zdnd11an1n04x5 FILLER_338_484 ();
 b15zdnd11an1n04x5 FILLER_338_494 ();
 b15zdnd11an1n04x5 FILLER_338_504 ();
 b15zdnd00an1n01x5 FILLER_338_508 ();
 b15zdnd11an1n16x5 FILLER_338_521 ();
 b15zdnd11an1n08x5 FILLER_338_537 ();
 b15zdnd00an1n02x5 FILLER_338_545 ();
 b15zdnd11an1n16x5 FILLER_338_556 ();
 b15zdnd00an1n02x5 FILLER_338_572 ();
 b15zdnd11an1n64x5 FILLER_338_578 ();
 b15zdnd11an1n08x5 FILLER_338_642 ();
 b15zdnd11an1n32x5 FILLER_338_656 ();
 b15zdnd11an1n16x5 FILLER_338_688 ();
 b15zdnd11an1n08x5 FILLER_338_704 ();
 b15zdnd11an1n04x5 FILLER_338_712 ();
 b15zdnd00an1n02x5 FILLER_338_716 ();
 b15zdnd11an1n64x5 FILLER_338_726 ();
 b15zdnd11an1n04x5 FILLER_338_790 ();
 b15zdnd00an1n02x5 FILLER_338_794 ();
 b15zdnd11an1n16x5 FILLER_338_815 ();
 b15zdnd00an1n02x5 FILLER_338_831 ();
 b15zdnd00an1n01x5 FILLER_338_833 ();
 b15zdnd11an1n16x5 FILLER_338_838 ();
 b15zdnd00an1n01x5 FILLER_338_854 ();
 b15zdnd11an1n08x5 FILLER_338_867 ();
 b15zdnd11an1n04x5 FILLER_338_875 ();
 b15zdnd11an1n08x5 FILLER_338_892 ();
 b15zdnd00an1n02x5 FILLER_338_900 ();
 b15zdnd11an1n04x5 FILLER_338_914 ();
 b15zdnd11an1n08x5 FILLER_338_938 ();
 b15zdnd11an1n04x5 FILLER_338_946 ();
 b15zdnd00an1n02x5 FILLER_338_950 ();
 b15zdnd00an1n01x5 FILLER_338_952 ();
 b15zdnd11an1n04x5 FILLER_338_960 ();
 b15zdnd11an1n16x5 FILLER_338_971 ();
 b15zdnd11an1n04x5 FILLER_338_987 ();
 b15zdnd11an1n16x5 FILLER_338_1002 ();
 b15zdnd00an1n01x5 FILLER_338_1018 ();
 b15zdnd11an1n04x5 FILLER_338_1023 ();
 b15zdnd11an1n04x5 FILLER_338_1033 ();
 b15zdnd11an1n16x5 FILLER_338_1043 ();
 b15zdnd11an1n04x5 FILLER_338_1059 ();
 b15zdnd00an1n02x5 FILLER_338_1063 ();
 b15zdnd11an1n04x5 FILLER_338_1069 ();
 b15zdnd11an1n16x5 FILLER_338_1079 ();
 b15zdnd11an1n04x5 FILLER_338_1095 ();
 b15zdnd11an1n04x5 FILLER_338_1103 ();
 b15zdnd11an1n08x5 FILLER_338_1113 ();
 b15zdnd11an1n16x5 FILLER_338_1147 ();
 b15zdnd11an1n04x5 FILLER_338_1163 ();
 b15zdnd11an1n04x5 FILLER_338_1171 ();
 b15zdnd11an1n04x5 FILLER_338_1187 ();
 b15zdnd11an1n08x5 FILLER_338_1214 ();
 b15zdnd11an1n04x5 FILLER_338_1248 ();
 b15zdnd11an1n04x5 FILLER_338_1278 ();
 b15zdnd11an1n64x5 FILLER_338_1292 ();
 b15zdnd11an1n16x5 FILLER_338_1356 ();
 b15zdnd11an1n08x5 FILLER_338_1372 ();
 b15zdnd11an1n04x5 FILLER_338_1380 ();
 b15zdnd00an1n02x5 FILLER_338_1384 ();
 b15zdnd00an1n01x5 FILLER_338_1386 ();
 b15zdnd11an1n64x5 FILLER_338_1394 ();
 b15zdnd11an1n64x5 FILLER_338_1458 ();
 b15zdnd11an1n64x5 FILLER_338_1522 ();
 b15zdnd11an1n32x5 FILLER_338_1586 ();
 b15zdnd11an1n16x5 FILLER_338_1618 ();
 b15zdnd11an1n04x5 FILLER_338_1634 ();
 b15zdnd00an1n01x5 FILLER_338_1638 ();
 b15zdnd11an1n04x5 FILLER_338_1645 ();
 b15zdnd00an1n02x5 FILLER_338_1649 ();
 b15zdnd11an1n32x5 FILLER_338_1656 ();
 b15zdnd11an1n04x5 FILLER_338_1688 ();
 b15zdnd00an1n01x5 FILLER_338_1692 ();
 b15zdnd11an1n64x5 FILLER_338_1725 ();
 b15zdnd11an1n16x5 FILLER_338_1789 ();
 b15zdnd11an1n08x5 FILLER_338_1805 ();
 b15zdnd11an1n04x5 FILLER_338_1813 ();
 b15zdnd11an1n64x5 FILLER_338_1837 ();
 b15zdnd11an1n32x5 FILLER_338_1901 ();
 b15zdnd11an1n08x5 FILLER_338_1933 ();
 b15zdnd11an1n04x5 FILLER_338_1941 ();
 b15zdnd00an1n01x5 FILLER_338_1945 ();
 b15zdnd11an1n16x5 FILLER_338_1970 ();
 b15zdnd11an1n04x5 FILLER_338_1986 ();
 b15zdnd00an1n02x5 FILLER_338_1990 ();
 b15zdnd11an1n08x5 FILLER_338_1998 ();
 b15zdnd00an1n01x5 FILLER_338_2006 ();
 b15zdnd11an1n64x5 FILLER_338_2012 ();
 b15zdnd11an1n64x5 FILLER_338_2076 ();
 b15zdnd11an1n08x5 FILLER_338_2140 ();
 b15zdnd11an1n04x5 FILLER_338_2148 ();
 b15zdnd00an1n02x5 FILLER_338_2152 ();
 b15zdnd11an1n32x5 FILLER_338_2162 ();
 b15zdnd11an1n08x5 FILLER_338_2194 ();
 b15zdnd11an1n04x5 FILLER_338_2207 ();
 b15zdnd00an1n01x5 FILLER_338_2211 ();
 b15zdnd11an1n32x5 FILLER_338_2220 ();
 b15zdnd11an1n16x5 FILLER_338_2252 ();
 b15zdnd11an1n08x5 FILLER_338_2268 ();
 b15zdnd11an1n64x5 FILLER_339_0 ();
 b15zdnd11an1n64x5 FILLER_339_64 ();
 b15zdnd11an1n64x5 FILLER_339_128 ();
 b15zdnd11an1n32x5 FILLER_339_192 ();
 b15zdnd11an1n16x5 FILLER_339_224 ();
 b15zdnd11an1n08x5 FILLER_339_240 ();
 b15zdnd00an1n02x5 FILLER_339_248 ();
 b15zdnd00an1n01x5 FILLER_339_250 ();
 b15zdnd11an1n04x5 FILLER_339_262 ();
 b15zdnd11an1n16x5 FILLER_339_271 ();
 b15zdnd11an1n04x5 FILLER_339_287 ();
 b15zdnd00an1n02x5 FILLER_339_291 ();
 b15zdnd00an1n01x5 FILLER_339_293 ();
 b15zdnd11an1n64x5 FILLER_339_314 ();
 b15zdnd11an1n32x5 FILLER_339_378 ();
 b15zdnd11an1n16x5 FILLER_339_410 ();
 b15zdnd11an1n04x5 FILLER_339_426 ();
 b15zdnd11an1n16x5 FILLER_339_435 ();
 b15zdnd11an1n04x5 FILLER_339_451 ();
 b15zdnd11an1n16x5 FILLER_339_461 ();
 b15zdnd11an1n08x5 FILLER_339_477 ();
 b15zdnd11an1n04x5 FILLER_339_485 ();
 b15zdnd00an1n02x5 FILLER_339_489 ();
 b15zdnd11an1n64x5 FILLER_339_501 ();
 b15zdnd11an1n16x5 FILLER_339_565 ();
 b15zdnd11an1n04x5 FILLER_339_587 ();
 b15zdnd11an1n04x5 FILLER_339_598 ();
 b15zdnd11an1n64x5 FILLER_339_608 ();
 b15zdnd11an1n64x5 FILLER_339_672 ();
 b15zdnd11an1n16x5 FILLER_339_736 ();
 b15zdnd11an1n08x5 FILLER_339_752 ();
 b15zdnd11an1n04x5 FILLER_339_760 ();
 b15zdnd11an1n64x5 FILLER_339_769 ();
 b15zdnd11an1n32x5 FILLER_339_833 ();
 b15zdnd11an1n08x5 FILLER_339_865 ();
 b15zdnd11an1n04x5 FILLER_339_882 ();
 b15zdnd00an1n02x5 FILLER_339_886 ();
 b15zdnd00an1n01x5 FILLER_339_888 ();
 b15zdnd11an1n04x5 FILLER_339_894 ();
 b15zdnd11an1n64x5 FILLER_339_908 ();
 b15zdnd11an1n16x5 FILLER_339_972 ();
 b15zdnd00an1n02x5 FILLER_339_988 ();
 b15zdnd11an1n16x5 FILLER_339_1000 ();
 b15zdnd11an1n04x5 FILLER_339_1016 ();
 b15zdnd00an1n02x5 FILLER_339_1020 ();
 b15zdnd00an1n01x5 FILLER_339_1022 ();
 b15zdnd11an1n04x5 FILLER_339_1030 ();
 b15zdnd11an1n16x5 FILLER_339_1040 ();
 b15zdnd11an1n08x5 FILLER_339_1056 ();
 b15zdnd11an1n04x5 FILLER_339_1064 ();
 b15zdnd11an1n16x5 FILLER_339_1075 ();
 b15zdnd11an1n08x5 FILLER_339_1091 ();
 b15zdnd00an1n02x5 FILLER_339_1099 ();
 b15zdnd00an1n01x5 FILLER_339_1101 ();
 b15zdnd11an1n04x5 FILLER_339_1115 ();
 b15zdnd11an1n08x5 FILLER_339_1126 ();
 b15zdnd11an1n04x5 FILLER_339_1134 ();
 b15zdnd00an1n01x5 FILLER_339_1138 ();
 b15zdnd11an1n04x5 FILLER_339_1165 ();
 b15zdnd11an1n64x5 FILLER_339_1195 ();
 b15zdnd11an1n16x5 FILLER_339_1259 ();
 b15zdnd11an1n04x5 FILLER_339_1275 ();
 b15zdnd00an1n02x5 FILLER_339_1279 ();
 b15zdnd11an1n64x5 FILLER_339_1288 ();
 b15zdnd11an1n04x5 FILLER_339_1352 ();
 b15zdnd00an1n02x5 FILLER_339_1356 ();
 b15zdnd00an1n01x5 FILLER_339_1358 ();
 b15zdnd11an1n16x5 FILLER_339_1366 ();
 b15zdnd11an1n04x5 FILLER_339_1382 ();
 b15zdnd00an1n02x5 FILLER_339_1386 ();
 b15zdnd00an1n01x5 FILLER_339_1388 ();
 b15zdnd11an1n64x5 FILLER_339_1394 ();
 b15zdnd11an1n16x5 FILLER_339_1458 ();
 b15zdnd11an1n04x5 FILLER_339_1474 ();
 b15zdnd00an1n01x5 FILLER_339_1478 ();
 b15zdnd11an1n32x5 FILLER_339_1486 ();
 b15zdnd11an1n16x5 FILLER_339_1518 ();
 b15zdnd11an1n16x5 FILLER_339_1544 ();
 b15zdnd11an1n04x5 FILLER_339_1560 ();
 b15zdnd00an1n01x5 FILLER_339_1564 ();
 b15zdnd11an1n32x5 FILLER_339_1570 ();
 b15zdnd11an1n16x5 FILLER_339_1602 ();
 b15zdnd11an1n08x5 FILLER_339_1618 ();
 b15zdnd11an1n04x5 FILLER_339_1626 ();
 b15zdnd00an1n02x5 FILLER_339_1630 ();
 b15zdnd00an1n01x5 FILLER_339_1632 ();
 b15zdnd11an1n04x5 FILLER_339_1639 ();
 b15zdnd11an1n32x5 FILLER_339_1655 ();
 b15zdnd11an1n16x5 FILLER_339_1696 ();
 b15zdnd00an1n02x5 FILLER_339_1712 ();
 b15zdnd00an1n01x5 FILLER_339_1714 ();
 b15zdnd11an1n64x5 FILLER_339_1725 ();
 b15zdnd11an1n64x5 FILLER_339_1789 ();
 b15zdnd11an1n16x5 FILLER_339_1853 ();
 b15zdnd11an1n04x5 FILLER_339_1869 ();
 b15zdnd11an1n64x5 FILLER_339_1882 ();
 b15zdnd11an1n64x5 FILLER_339_1946 ();
 b15zdnd11an1n32x5 FILLER_339_2010 ();
 b15zdnd11an1n08x5 FILLER_339_2042 ();
 b15zdnd00an1n01x5 FILLER_339_2050 ();
 b15zdnd11an1n04x5 FILLER_339_2056 ();
 b15zdnd11an1n04x5 FILLER_339_2065 ();
 b15zdnd11an1n32x5 FILLER_339_2077 ();
 b15zdnd11an1n16x5 FILLER_339_2109 ();
 b15zdnd11an1n08x5 FILLER_339_2125 ();
 b15zdnd00an1n02x5 FILLER_339_2133 ();
 b15zdnd00an1n01x5 FILLER_339_2135 ();
 b15zdnd11an1n16x5 FILLER_339_2142 ();
 b15zdnd11an1n04x5 FILLER_339_2158 ();
 b15zdnd00an1n02x5 FILLER_339_2162 ();
 b15zdnd11an1n04x5 FILLER_339_2170 ();
 b15zdnd11an1n16x5 FILLER_339_2179 ();
 b15zdnd11an1n08x5 FILLER_339_2195 ();
 b15zdnd11an1n04x5 FILLER_339_2203 ();
 b15zdnd00an1n02x5 FILLER_339_2207 ();
 b15zdnd11an1n32x5 FILLER_339_2225 ();
 b15zdnd11an1n16x5 FILLER_339_2257 ();
 b15zdnd11an1n08x5 FILLER_339_2273 ();
 b15zdnd00an1n02x5 FILLER_339_2281 ();
 b15zdnd00an1n01x5 FILLER_339_2283 ();
 b15zdnd11an1n64x5 FILLER_340_8 ();
 b15zdnd11an1n64x5 FILLER_340_72 ();
 b15zdnd11an1n64x5 FILLER_340_136 ();
 b15zdnd11an1n16x5 FILLER_340_200 ();
 b15zdnd11an1n08x5 FILLER_340_216 ();
 b15zdnd11an1n04x5 FILLER_340_224 ();
 b15zdnd00an1n02x5 FILLER_340_228 ();
 b15zdnd11an1n08x5 FILLER_340_244 ();
 b15zdnd00an1n01x5 FILLER_340_252 ();
 b15zdnd11an1n64x5 FILLER_340_260 ();
 b15zdnd11an1n32x5 FILLER_340_324 ();
 b15zdnd11an1n08x5 FILLER_340_356 ();
 b15zdnd00an1n02x5 FILLER_340_364 ();
 b15zdnd11an1n32x5 FILLER_340_397 ();
 b15zdnd11an1n08x5 FILLER_340_429 ();
 b15zdnd11an1n04x5 FILLER_340_437 ();
 b15zdnd00an1n01x5 FILLER_340_441 ();
 b15zdnd11an1n04x5 FILLER_340_449 ();
 b15zdnd11an1n32x5 FILLER_340_468 ();
 b15zdnd11an1n08x5 FILLER_340_500 ();
 b15zdnd11an1n16x5 FILLER_340_518 ();
 b15zdnd11an1n04x5 FILLER_340_534 ();
 b15zdnd00an1n01x5 FILLER_340_538 ();
 b15zdnd11an1n32x5 FILLER_340_558 ();
 b15zdnd00an1n02x5 FILLER_340_590 ();
 b15zdnd11an1n64x5 FILLER_340_599 ();
 b15zdnd11an1n16x5 FILLER_340_663 ();
 b15zdnd00an1n01x5 FILLER_340_679 ();
 b15zdnd11an1n08x5 FILLER_340_687 ();
 b15zdnd11an1n04x5 FILLER_340_695 ();
 b15zdnd00an1n01x5 FILLER_340_699 ();
 b15zdnd11an1n04x5 FILLER_340_712 ();
 b15zdnd00an1n02x5 FILLER_340_716 ();
 b15zdnd00an1n02x5 FILLER_340_726 ();
 b15zdnd11an1n08x5 FILLER_340_742 ();
 b15zdnd00an1n02x5 FILLER_340_750 ();
 b15zdnd11an1n08x5 FILLER_340_756 ();
 b15zdnd00an1n01x5 FILLER_340_764 ();
 b15zdnd11an1n16x5 FILLER_340_771 ();
 b15zdnd11an1n08x5 FILLER_340_787 ();
 b15zdnd11an1n04x5 FILLER_340_795 ();
 b15zdnd00an1n02x5 FILLER_340_799 ();
 b15zdnd00an1n01x5 FILLER_340_801 ();
 b15zdnd11an1n64x5 FILLER_340_808 ();
 b15zdnd11an1n64x5 FILLER_340_872 ();
 b15zdnd11an1n16x5 FILLER_340_936 ();
 b15zdnd11an1n04x5 FILLER_340_952 ();
 b15zdnd11an1n16x5 FILLER_340_968 ();
 b15zdnd11an1n04x5 FILLER_340_984 ();
 b15zdnd00an1n02x5 FILLER_340_988 ();
 b15zdnd00an1n01x5 FILLER_340_990 ();
 b15zdnd11an1n64x5 FILLER_340_999 ();
 b15zdnd11an1n32x5 FILLER_340_1063 ();
 b15zdnd11an1n08x5 FILLER_340_1095 ();
 b15zdnd00an1n02x5 FILLER_340_1103 ();
 b15zdnd11an1n08x5 FILLER_340_1125 ();
 b15zdnd00an1n01x5 FILLER_340_1133 ();
 b15zdnd11an1n08x5 FILLER_340_1140 ();
 b15zdnd11an1n04x5 FILLER_340_1148 ();
 b15zdnd00an1n01x5 FILLER_340_1152 ();
 b15zdnd11an1n16x5 FILLER_340_1169 ();
 b15zdnd11an1n04x5 FILLER_340_1185 ();
 b15zdnd11an1n32x5 FILLER_340_1197 ();
 b15zdnd11an1n08x5 FILLER_340_1229 ();
 b15zdnd00an1n01x5 FILLER_340_1237 ();
 b15zdnd11an1n64x5 FILLER_340_1264 ();
 b15zdnd11an1n16x5 FILLER_340_1328 ();
 b15zdnd11an1n04x5 FILLER_340_1344 ();
 b15zdnd11an1n32x5 FILLER_340_1363 ();
 b15zdnd11an1n04x5 FILLER_340_1409 ();
 b15zdnd00an1n01x5 FILLER_340_1413 ();
 b15zdnd11an1n04x5 FILLER_340_1424 ();
 b15zdnd11an1n08x5 FILLER_340_1437 ();
 b15zdnd00an1n01x5 FILLER_340_1445 ();
 b15zdnd11an1n08x5 FILLER_340_1460 ();
 b15zdnd11an1n08x5 FILLER_340_1484 ();
 b15zdnd00an1n02x5 FILLER_340_1492 ();
 b15zdnd00an1n01x5 FILLER_340_1494 ();
 b15zdnd11an1n16x5 FILLER_340_1504 ();
 b15zdnd11an1n08x5 FILLER_340_1520 ();
 b15zdnd00an1n02x5 FILLER_340_1528 ();
 b15zdnd11an1n08x5 FILLER_340_1547 ();
 b15zdnd11an1n04x5 FILLER_340_1555 ();
 b15zdnd00an1n02x5 FILLER_340_1559 ();
 b15zdnd11an1n04x5 FILLER_340_1570 ();
 b15zdnd00an1n02x5 FILLER_340_1574 ();
 b15zdnd00an1n01x5 FILLER_340_1576 ();
 b15zdnd11an1n04x5 FILLER_340_1593 ();
 b15zdnd11an1n04x5 FILLER_340_1604 ();
 b15zdnd00an1n02x5 FILLER_340_1608 ();
 b15zdnd00an1n01x5 FILLER_340_1610 ();
 b15zdnd11an1n16x5 FILLER_340_1616 ();
 b15zdnd11an1n64x5 FILLER_340_1636 ();
 b15zdnd00an1n02x5 FILLER_340_1700 ();
 b15zdnd00an1n01x5 FILLER_340_1702 ();
 b15zdnd11an1n08x5 FILLER_340_1713 ();
 b15zdnd11an1n04x5 FILLER_340_1721 ();
 b15zdnd00an1n02x5 FILLER_340_1725 ();
 b15zdnd11an1n64x5 FILLER_340_1735 ();
 b15zdnd11an1n32x5 FILLER_340_1799 ();
 b15zdnd11an1n16x5 FILLER_340_1831 ();
 b15zdnd00an1n02x5 FILLER_340_1847 ();
 b15zdnd11an1n64x5 FILLER_340_1854 ();
 b15zdnd11an1n32x5 FILLER_340_1918 ();
 b15zdnd11an1n08x5 FILLER_340_1950 ();
 b15zdnd11an1n04x5 FILLER_340_1958 ();
 b15zdnd00an1n02x5 FILLER_340_1962 ();
 b15zdnd11an1n32x5 FILLER_340_1977 ();
 b15zdnd11an1n04x5 FILLER_340_2009 ();
 b15zdnd00an1n02x5 FILLER_340_2013 ();
 b15zdnd00an1n01x5 FILLER_340_2015 ();
 b15zdnd11an1n64x5 FILLER_340_2028 ();
 b15zdnd11an1n04x5 FILLER_340_2092 ();
 b15zdnd00an1n02x5 FILLER_340_2096 ();
 b15zdnd00an1n01x5 FILLER_340_2098 ();
 b15zdnd11an1n16x5 FILLER_340_2115 ();
 b15zdnd11an1n04x5 FILLER_340_2131 ();
 b15zdnd11an1n08x5 FILLER_340_2140 ();
 b15zdnd11an1n04x5 FILLER_340_2148 ();
 b15zdnd00an1n02x5 FILLER_340_2152 ();
 b15zdnd11an1n64x5 FILLER_340_2162 ();
 b15zdnd11an1n32x5 FILLER_340_2226 ();
 b15zdnd11an1n16x5 FILLER_340_2258 ();
 b15zdnd00an1n02x5 FILLER_340_2274 ();
 b15zdnd11an1n64x5 FILLER_341_0 ();
 b15zdnd11an1n64x5 FILLER_341_64 ();
 b15zdnd11an1n64x5 FILLER_341_128 ();
 b15zdnd11an1n16x5 FILLER_341_192 ();
 b15zdnd11an1n08x5 FILLER_341_208 ();
 b15zdnd00an1n02x5 FILLER_341_216 ();
 b15zdnd11an1n04x5 FILLER_341_231 ();
 b15zdnd00an1n01x5 FILLER_341_235 ();
 b15zdnd11an1n04x5 FILLER_341_242 ();
 b15zdnd11an1n32x5 FILLER_341_258 ();
 b15zdnd11an1n04x5 FILLER_341_290 ();
 b15zdnd00an1n01x5 FILLER_341_294 ();
 b15zdnd11an1n32x5 FILLER_341_299 ();
 b15zdnd11an1n16x5 FILLER_341_331 ();
 b15zdnd00an1n01x5 FILLER_341_347 ();
 b15zdnd11an1n04x5 FILLER_341_357 ();
 b15zdnd11an1n08x5 FILLER_341_377 ();
 b15zdnd11an1n04x5 FILLER_341_385 ();
 b15zdnd11an1n04x5 FILLER_341_404 ();
 b15zdnd11an1n08x5 FILLER_341_417 ();
 b15zdnd11an1n04x5 FILLER_341_425 ();
 b15zdnd00an1n02x5 FILLER_341_429 ();
 b15zdnd11an1n32x5 FILLER_341_437 ();
 b15zdnd11an1n08x5 FILLER_341_469 ();
 b15zdnd11an1n04x5 FILLER_341_477 ();
 b15zdnd00an1n01x5 FILLER_341_481 ();
 b15zdnd11an1n32x5 FILLER_341_491 ();
 b15zdnd11an1n16x5 FILLER_341_523 ();
 b15zdnd11an1n64x5 FILLER_341_550 ();
 b15zdnd11an1n64x5 FILLER_341_614 ();
 b15zdnd11an1n04x5 FILLER_341_678 ();
 b15zdnd00an1n02x5 FILLER_341_682 ();
 b15zdnd00an1n01x5 FILLER_341_684 ();
 b15zdnd11an1n08x5 FILLER_341_691 ();
 b15zdnd00an1n01x5 FILLER_341_699 ();
 b15zdnd11an1n32x5 FILLER_341_705 ();
 b15zdnd11an1n16x5 FILLER_341_737 ();
 b15zdnd00an1n02x5 FILLER_341_753 ();
 b15zdnd00an1n01x5 FILLER_341_755 ();
 b15zdnd11an1n64x5 FILLER_341_768 ();
 b15zdnd11an1n04x5 FILLER_341_832 ();
 b15zdnd00an1n02x5 FILLER_341_836 ();
 b15zdnd11an1n64x5 FILLER_341_851 ();
 b15zdnd11an1n64x5 FILLER_341_915 ();
 b15zdnd11an1n64x5 FILLER_341_979 ();
 b15zdnd11an1n64x5 FILLER_341_1043 ();
 b15zdnd11an1n16x5 FILLER_341_1107 ();
 b15zdnd11an1n08x5 FILLER_341_1123 ();
 b15zdnd11an1n04x5 FILLER_341_1131 ();
 b15zdnd11an1n64x5 FILLER_341_1142 ();
 b15zdnd11an1n16x5 FILLER_341_1211 ();
 b15zdnd11an1n08x5 FILLER_341_1227 ();
 b15zdnd00an1n02x5 FILLER_341_1235 ();
 b15zdnd11an1n04x5 FILLER_341_1249 ();
 b15zdnd11an1n08x5 FILLER_341_1257 ();
 b15zdnd11an1n04x5 FILLER_341_1265 ();
 b15zdnd11an1n32x5 FILLER_341_1279 ();
 b15zdnd11an1n04x5 FILLER_341_1311 ();
 b15zdnd11an1n04x5 FILLER_341_1333 ();
 b15zdnd11an1n04x5 FILLER_341_1349 ();
 b15zdnd00an1n02x5 FILLER_341_1353 ();
 b15zdnd11an1n32x5 FILLER_341_1360 ();
 b15zdnd11an1n16x5 FILLER_341_1392 ();
 b15zdnd00an1n01x5 FILLER_341_1408 ();
 b15zdnd11an1n16x5 FILLER_341_1418 ();
 b15zdnd00an1n02x5 FILLER_341_1434 ();
 b15zdnd11an1n32x5 FILLER_341_1443 ();
 b15zdnd11an1n08x5 FILLER_341_1475 ();
 b15zdnd00an1n02x5 FILLER_341_1483 ();
 b15zdnd11an1n08x5 FILLER_341_1499 ();
 b15zdnd00an1n01x5 FILLER_341_1507 ();
 b15zdnd11an1n08x5 FILLER_341_1512 ();
 b15zdnd11an1n04x5 FILLER_341_1520 ();
 b15zdnd00an1n01x5 FILLER_341_1524 ();
 b15zdnd11an1n32x5 FILLER_341_1531 ();
 b15zdnd11an1n04x5 FILLER_341_1563 ();
 b15zdnd00an1n01x5 FILLER_341_1567 ();
 b15zdnd11an1n08x5 FILLER_341_1574 ();
 b15zdnd11an1n04x5 FILLER_341_1602 ();
 b15zdnd11an1n04x5 FILLER_341_1616 ();
 b15zdnd11an1n32x5 FILLER_341_1624 ();
 b15zdnd11an1n16x5 FILLER_341_1656 ();
 b15zdnd11an1n04x5 FILLER_341_1672 ();
 b15zdnd00an1n02x5 FILLER_341_1676 ();
 b15zdnd11an1n08x5 FILLER_341_1685 ();
 b15zdnd11an1n04x5 FILLER_341_1693 ();
 b15zdnd00an1n02x5 FILLER_341_1697 ();
 b15zdnd00an1n01x5 FILLER_341_1699 ();
 b15zdnd11an1n04x5 FILLER_341_1704 ();
 b15zdnd11an1n64x5 FILLER_341_1721 ();
 b15zdnd11an1n16x5 FILLER_341_1785 ();
 b15zdnd11an1n08x5 FILLER_341_1801 ();
 b15zdnd11an1n04x5 FILLER_341_1809 ();
 b15zdnd11an1n16x5 FILLER_341_1818 ();
 b15zdnd00an1n02x5 FILLER_341_1834 ();
 b15zdnd00an1n01x5 FILLER_341_1836 ();
 b15zdnd11an1n04x5 FILLER_341_1842 ();
 b15zdnd00an1n02x5 FILLER_341_1846 ();
 b15zdnd11an1n16x5 FILLER_341_1858 ();
 b15zdnd11an1n08x5 FILLER_341_1874 ();
 b15zdnd11an1n04x5 FILLER_341_1902 ();
 b15zdnd11an1n04x5 FILLER_341_1911 ();
 b15zdnd11an1n04x5 FILLER_341_1919 ();
 b15zdnd11an1n08x5 FILLER_341_1927 ();
 b15zdnd11an1n16x5 FILLER_341_1940 ();
 b15zdnd11an1n08x5 FILLER_341_1956 ();
 b15zdnd11an1n04x5 FILLER_341_1964 ();
 b15zdnd00an1n02x5 FILLER_341_1968 ();
 b15zdnd00an1n01x5 FILLER_341_1970 ();
 b15zdnd11an1n16x5 FILLER_341_1993 ();
 b15zdnd11an1n04x5 FILLER_341_2009 ();
 b15zdnd00an1n01x5 FILLER_341_2013 ();
 b15zdnd11an1n16x5 FILLER_341_2029 ();
 b15zdnd00an1n02x5 FILLER_341_2045 ();
 b15zdnd00an1n01x5 FILLER_341_2047 ();
 b15zdnd11an1n64x5 FILLER_341_2052 ();
 b15zdnd11an1n64x5 FILLER_341_2116 ();
 b15zdnd11an1n64x5 FILLER_341_2180 ();
 b15zdnd11an1n32x5 FILLER_341_2244 ();
 b15zdnd11an1n08x5 FILLER_341_2276 ();
 b15zdnd11an1n64x5 FILLER_342_8 ();
 b15zdnd11an1n64x5 FILLER_342_72 ();
 b15zdnd11an1n64x5 FILLER_342_136 ();
 b15zdnd11an1n32x5 FILLER_342_200 ();
 b15zdnd11an1n16x5 FILLER_342_232 ();
 b15zdnd11an1n04x5 FILLER_342_248 ();
 b15zdnd00an1n01x5 FILLER_342_252 ();
 b15zdnd11an1n16x5 FILLER_342_257 ();
 b15zdnd00an1n02x5 FILLER_342_273 ();
 b15zdnd00an1n01x5 FILLER_342_275 ();
 b15zdnd11an1n04x5 FILLER_342_288 ();
 b15zdnd00an1n02x5 FILLER_342_292 ();
 b15zdnd00an1n01x5 FILLER_342_294 ();
 b15zdnd11an1n08x5 FILLER_342_305 ();
 b15zdnd11an1n04x5 FILLER_342_313 ();
 b15zdnd11an1n04x5 FILLER_342_326 ();
 b15zdnd11an1n16x5 FILLER_342_334 ();
 b15zdnd00an1n02x5 FILLER_342_350 ();
 b15zdnd00an1n01x5 FILLER_342_352 ();
 b15zdnd11an1n32x5 FILLER_342_360 ();
 b15zdnd11an1n16x5 FILLER_342_392 ();
 b15zdnd11an1n04x5 FILLER_342_408 ();
 b15zdnd00an1n02x5 FILLER_342_412 ();
 b15zdnd00an1n01x5 FILLER_342_414 ();
 b15zdnd11an1n32x5 FILLER_342_422 ();
 b15zdnd00an1n02x5 FILLER_342_454 ();
 b15zdnd11an1n32x5 FILLER_342_462 ();
 b15zdnd11an1n16x5 FILLER_342_494 ();
 b15zdnd11an1n16x5 FILLER_342_515 ();
 b15zdnd11an1n08x5 FILLER_342_531 ();
 b15zdnd11an1n64x5 FILLER_342_547 ();
 b15zdnd11an1n32x5 FILLER_342_611 ();
 b15zdnd11an1n16x5 FILLER_342_643 ();
 b15zdnd00an1n02x5 FILLER_342_659 ();
 b15zdnd00an1n01x5 FILLER_342_661 ();
 b15zdnd11an1n08x5 FILLER_342_667 ();
 b15zdnd11an1n04x5 FILLER_342_675 ();
 b15zdnd00an1n02x5 FILLER_342_679 ();
 b15zdnd11an1n08x5 FILLER_342_688 ();
 b15zdnd11an1n04x5 FILLER_342_696 ();
 b15zdnd00an1n02x5 FILLER_342_700 ();
 b15zdnd11an1n04x5 FILLER_342_714 ();
 b15zdnd11an1n32x5 FILLER_342_726 ();
 b15zdnd11an1n16x5 FILLER_342_758 ();
 b15zdnd00an1n02x5 FILLER_342_774 ();
 b15zdnd11an1n32x5 FILLER_342_787 ();
 b15zdnd11an1n04x5 FILLER_342_819 ();
 b15zdnd11an1n08x5 FILLER_342_829 ();
 b15zdnd11an1n08x5 FILLER_342_847 ();
 b15zdnd00an1n02x5 FILLER_342_855 ();
 b15zdnd00an1n01x5 FILLER_342_857 ();
 b15zdnd11an1n32x5 FILLER_342_865 ();
 b15zdnd00an1n02x5 FILLER_342_897 ();
 b15zdnd00an1n01x5 FILLER_342_899 ();
 b15zdnd11an1n04x5 FILLER_342_914 ();
 b15zdnd00an1n01x5 FILLER_342_918 ();
 b15zdnd11an1n08x5 FILLER_342_924 ();
 b15zdnd11an1n04x5 FILLER_342_932 ();
 b15zdnd00an1n02x5 FILLER_342_936 ();
 b15zdnd00an1n01x5 FILLER_342_938 ();
 b15zdnd11an1n04x5 FILLER_342_951 ();
 b15zdnd00an1n02x5 FILLER_342_955 ();
 b15zdnd00an1n01x5 FILLER_342_957 ();
 b15zdnd11an1n64x5 FILLER_342_970 ();
 b15zdnd11an1n32x5 FILLER_342_1034 ();
 b15zdnd11an1n04x5 FILLER_342_1066 ();
 b15zdnd11an1n32x5 FILLER_342_1077 ();
 b15zdnd11an1n16x5 FILLER_342_1109 ();
 b15zdnd00an1n02x5 FILLER_342_1125 ();
 b15zdnd00an1n01x5 FILLER_342_1127 ();
 b15zdnd11an1n32x5 FILLER_342_1138 ();
 b15zdnd11an1n16x5 FILLER_342_1170 ();
 b15zdnd11an1n08x5 FILLER_342_1186 ();
 b15zdnd11an1n04x5 FILLER_342_1194 ();
 b15zdnd00an1n02x5 FILLER_342_1198 ();
 b15zdnd11an1n32x5 FILLER_342_1210 ();
 b15zdnd11an1n08x5 FILLER_342_1242 ();
 b15zdnd11an1n04x5 FILLER_342_1250 ();
 b15zdnd11an1n04x5 FILLER_342_1270 ();
 b15zdnd11an1n32x5 FILLER_342_1278 ();
 b15zdnd11an1n16x5 FILLER_342_1310 ();
 b15zdnd11an1n08x5 FILLER_342_1326 ();
 b15zdnd11an1n04x5 FILLER_342_1334 ();
 b15zdnd00an1n02x5 FILLER_342_1338 ();
 b15zdnd11an1n08x5 FILLER_342_1354 ();
 b15zdnd00an1n01x5 FILLER_342_1362 ();
 b15zdnd11an1n04x5 FILLER_342_1379 ();
 b15zdnd11an1n16x5 FILLER_342_1389 ();
 b15zdnd11an1n04x5 FILLER_342_1405 ();
 b15zdnd00an1n01x5 FILLER_342_1409 ();
 b15zdnd11an1n08x5 FILLER_342_1417 ();
 b15zdnd00an1n01x5 FILLER_342_1425 ();
 b15zdnd11an1n08x5 FILLER_342_1431 ();
 b15zdnd11an1n04x5 FILLER_342_1439 ();
 b15zdnd00an1n01x5 FILLER_342_1443 ();
 b15zdnd11an1n32x5 FILLER_342_1448 ();
 b15zdnd00an1n01x5 FILLER_342_1480 ();
 b15zdnd11an1n32x5 FILLER_342_1491 ();
 b15zdnd11an1n04x5 FILLER_342_1523 ();
 b15zdnd11an1n04x5 FILLER_342_1539 ();
 b15zdnd11an1n08x5 FILLER_342_1549 ();
 b15zdnd00an1n02x5 FILLER_342_1557 ();
 b15zdnd11an1n04x5 FILLER_342_1564 ();
 b15zdnd11an1n32x5 FILLER_342_1577 ();
 b15zdnd11an1n16x5 FILLER_342_1609 ();
 b15zdnd11an1n32x5 FILLER_342_1645 ();
 b15zdnd11an1n04x5 FILLER_342_1690 ();
 b15zdnd11an1n32x5 FILLER_342_1704 ();
 b15zdnd00an1n01x5 FILLER_342_1736 ();
 b15zdnd11an1n64x5 FILLER_342_1742 ();
 b15zdnd11an1n04x5 FILLER_342_1806 ();
 b15zdnd11an1n04x5 FILLER_342_1821 ();
 b15zdnd11an1n04x5 FILLER_342_1834 ();
 b15zdnd11an1n08x5 FILLER_342_1844 ();
 b15zdnd00an1n02x5 FILLER_342_1852 ();
 b15zdnd11an1n08x5 FILLER_342_1861 ();
 b15zdnd11an1n04x5 FILLER_342_1869 ();
 b15zdnd00an1n02x5 FILLER_342_1873 ();
 b15zdnd11an1n32x5 FILLER_342_1882 ();
 b15zdnd11an1n08x5 FILLER_342_1914 ();
 b15zdnd00an1n02x5 FILLER_342_1922 ();
 b15zdnd11an1n08x5 FILLER_342_1938 ();
 b15zdnd00an1n02x5 FILLER_342_1946 ();
 b15zdnd00an1n01x5 FILLER_342_1948 ();
 b15zdnd11an1n64x5 FILLER_342_1956 ();
 b15zdnd11an1n04x5 FILLER_342_2020 ();
 b15zdnd11an1n16x5 FILLER_342_2032 ();
 b15zdnd11an1n08x5 FILLER_342_2048 ();
 b15zdnd11an1n04x5 FILLER_342_2056 ();
 b15zdnd00an1n02x5 FILLER_342_2060 ();
 b15zdnd11an1n08x5 FILLER_342_2067 ();
 b15zdnd11an1n04x5 FILLER_342_2075 ();
 b15zdnd11an1n04x5 FILLER_342_2086 ();
 b15zdnd00an1n02x5 FILLER_342_2090 ();
 b15zdnd00an1n01x5 FILLER_342_2092 ();
 b15zdnd11an1n16x5 FILLER_342_2099 ();
 b15zdnd11an1n08x5 FILLER_342_2115 ();
 b15zdnd00an1n01x5 FILLER_342_2123 ();
 b15zdnd11an1n16x5 FILLER_342_2129 ();
 b15zdnd11an1n08x5 FILLER_342_2145 ();
 b15zdnd00an1n01x5 FILLER_342_2153 ();
 b15zdnd00an1n02x5 FILLER_342_2162 ();
 b15zdnd11an1n08x5 FILLER_342_2169 ();
 b15zdnd11an1n08x5 FILLER_342_2197 ();
 b15zdnd00an1n02x5 FILLER_342_2205 ();
 b15zdnd11an1n32x5 FILLER_342_2219 ();
 b15zdnd11an1n16x5 FILLER_342_2251 ();
 b15zdnd11an1n08x5 FILLER_342_2267 ();
 b15zdnd00an1n01x5 FILLER_342_2275 ();
 b15zdnd11an1n64x5 FILLER_343_0 ();
 b15zdnd11an1n64x5 FILLER_343_64 ();
 b15zdnd11an1n64x5 FILLER_343_128 ();
 b15zdnd11an1n32x5 FILLER_343_192 ();
 b15zdnd11an1n16x5 FILLER_343_224 ();
 b15zdnd00an1n02x5 FILLER_343_240 ();
 b15zdnd11an1n08x5 FILLER_343_256 ();
 b15zdnd11an1n04x5 FILLER_343_264 ();
 b15zdnd00an1n01x5 FILLER_343_268 ();
 b15zdnd11an1n32x5 FILLER_343_274 ();
 b15zdnd11an1n08x5 FILLER_343_306 ();
 b15zdnd11an1n04x5 FILLER_343_314 ();
 b15zdnd00an1n02x5 FILLER_343_318 ();
 b15zdnd11an1n64x5 FILLER_343_338 ();
 b15zdnd11an1n64x5 FILLER_343_402 ();
 b15zdnd11an1n32x5 FILLER_343_466 ();
 b15zdnd00an1n02x5 FILLER_343_498 ();
 b15zdnd00an1n01x5 FILLER_343_500 ();
 b15zdnd11an1n32x5 FILLER_343_508 ();
 b15zdnd11an1n08x5 FILLER_343_540 ();
 b15zdnd11an1n04x5 FILLER_343_548 ();
 b15zdnd11an1n16x5 FILLER_343_556 ();
 b15zdnd11an1n08x5 FILLER_343_572 ();
 b15zdnd11an1n04x5 FILLER_343_580 ();
 b15zdnd00an1n02x5 FILLER_343_584 ();
 b15zdnd11an1n64x5 FILLER_343_595 ();
 b15zdnd11an1n04x5 FILLER_343_659 ();
 b15zdnd11an1n04x5 FILLER_343_672 ();
 b15zdnd00an1n02x5 FILLER_343_676 ();
 b15zdnd00an1n01x5 FILLER_343_678 ();
 b15zdnd11an1n16x5 FILLER_343_685 ();
 b15zdnd11an1n04x5 FILLER_343_701 ();
 b15zdnd00an1n02x5 FILLER_343_705 ();
 b15zdnd11an1n04x5 FILLER_343_711 ();
 b15zdnd11an1n08x5 FILLER_343_721 ();
 b15zdnd00an1n02x5 FILLER_343_729 ();
 b15zdnd00an1n01x5 FILLER_343_731 ();
 b15zdnd11an1n64x5 FILLER_343_739 ();
 b15zdnd11an1n16x5 FILLER_343_803 ();
 b15zdnd00an1n01x5 FILLER_343_819 ();
 b15zdnd11an1n16x5 FILLER_343_826 ();
 b15zdnd11an1n08x5 FILLER_343_842 ();
 b15zdnd11an1n04x5 FILLER_343_850 ();
 b15zdnd00an1n01x5 FILLER_343_854 ();
 b15zdnd11an1n04x5 FILLER_343_859 ();
 b15zdnd11an1n16x5 FILLER_343_875 ();
 b15zdnd00an1n02x5 FILLER_343_891 ();
 b15zdnd11an1n08x5 FILLER_343_903 ();
 b15zdnd11an1n04x5 FILLER_343_911 ();
 b15zdnd00an1n02x5 FILLER_343_915 ();
 b15zdnd11an1n08x5 FILLER_343_928 ();
 b15zdnd00an1n02x5 FILLER_343_936 ();
 b15zdnd11an1n04x5 FILLER_343_958 ();
 b15zdnd11an1n04x5 FILLER_343_978 ();
 b15zdnd11an1n64x5 FILLER_343_988 ();
 b15zdnd11an1n04x5 FILLER_343_1052 ();
 b15zdnd00an1n02x5 FILLER_343_1056 ();
 b15zdnd00an1n01x5 FILLER_343_1058 ();
 b15zdnd11an1n16x5 FILLER_343_1066 ();
 b15zdnd11an1n04x5 FILLER_343_1095 ();
 b15zdnd11an1n32x5 FILLER_343_1103 ();
 b15zdnd11an1n08x5 FILLER_343_1135 ();
 b15zdnd11an1n04x5 FILLER_343_1143 ();
 b15zdnd00an1n02x5 FILLER_343_1147 ();
 b15zdnd11an1n16x5 FILLER_343_1163 ();
 b15zdnd11an1n04x5 FILLER_343_1179 ();
 b15zdnd00an1n02x5 FILLER_343_1183 ();
 b15zdnd00an1n01x5 FILLER_343_1185 ();
 b15zdnd11an1n04x5 FILLER_343_1200 ();
 b15zdnd11an1n32x5 FILLER_343_1216 ();
 b15zdnd11an1n16x5 FILLER_343_1248 ();
 b15zdnd11an1n04x5 FILLER_343_1264 ();
 b15zdnd11an1n16x5 FILLER_343_1272 ();
 b15zdnd11an1n08x5 FILLER_343_1288 ();
 b15zdnd11an1n04x5 FILLER_343_1296 ();
 b15zdnd00an1n02x5 FILLER_343_1300 ();
 b15zdnd11an1n32x5 FILLER_343_1322 ();
 b15zdnd11an1n04x5 FILLER_343_1354 ();
 b15zdnd00an1n02x5 FILLER_343_1358 ();
 b15zdnd00an1n01x5 FILLER_343_1360 ();
 b15zdnd11an1n64x5 FILLER_343_1388 ();
 b15zdnd11an1n64x5 FILLER_343_1452 ();
 b15zdnd11an1n64x5 FILLER_343_1516 ();
 b15zdnd11an1n64x5 FILLER_343_1580 ();
 b15zdnd11an1n16x5 FILLER_343_1644 ();
 b15zdnd00an1n02x5 FILLER_343_1660 ();
 b15zdnd00an1n01x5 FILLER_343_1662 ();
 b15zdnd11an1n32x5 FILLER_343_1669 ();
 b15zdnd11an1n16x5 FILLER_343_1701 ();
 b15zdnd00an1n01x5 FILLER_343_1717 ();
 b15zdnd11an1n08x5 FILLER_343_1723 ();
 b15zdnd11an1n04x5 FILLER_343_1731 ();
 b15zdnd00an1n02x5 FILLER_343_1735 ();
 b15zdnd11an1n64x5 FILLER_343_1749 ();
 b15zdnd00an1n02x5 FILLER_343_1813 ();
 b15zdnd11an1n08x5 FILLER_343_1827 ();
 b15zdnd11an1n04x5 FILLER_343_1835 ();
 b15zdnd00an1n01x5 FILLER_343_1839 ();
 b15zdnd11an1n64x5 FILLER_343_1847 ();
 b15zdnd11an1n32x5 FILLER_343_1911 ();
 b15zdnd11an1n08x5 FILLER_343_1943 ();
 b15zdnd11an1n32x5 FILLER_343_1957 ();
 b15zdnd11an1n16x5 FILLER_343_1989 ();
 b15zdnd00an1n02x5 FILLER_343_2005 ();
 b15zdnd00an1n01x5 FILLER_343_2007 ();
 b15zdnd11an1n08x5 FILLER_343_2015 ();
 b15zdnd00an1n02x5 FILLER_343_2023 ();
 b15zdnd00an1n01x5 FILLER_343_2025 ();
 b15zdnd11an1n04x5 FILLER_343_2041 ();
 b15zdnd11an1n04x5 FILLER_343_2071 ();
 b15zdnd11an1n16x5 FILLER_343_2083 ();
 b15zdnd11an1n04x5 FILLER_343_2099 ();
 b15zdnd00an1n02x5 FILLER_343_2103 ();
 b15zdnd11an1n08x5 FILLER_343_2110 ();
 b15zdnd11an1n04x5 FILLER_343_2118 ();
 b15zdnd00an1n02x5 FILLER_343_2122 ();
 b15zdnd11an1n16x5 FILLER_343_2133 ();
 b15zdnd00an1n02x5 FILLER_343_2149 ();
 b15zdnd00an1n01x5 FILLER_343_2151 ();
 b15zdnd11an1n08x5 FILLER_343_2156 ();
 b15zdnd11an1n16x5 FILLER_343_2172 ();
 b15zdnd11an1n08x5 FILLER_343_2188 ();
 b15zdnd11an1n04x5 FILLER_343_2196 ();
 b15zdnd00an1n01x5 FILLER_343_2200 ();
 b15zdnd11an1n64x5 FILLER_343_2213 ();
 b15zdnd11an1n04x5 FILLER_343_2277 ();
 b15zdnd00an1n02x5 FILLER_343_2281 ();
 b15zdnd00an1n01x5 FILLER_343_2283 ();
 b15zdnd11an1n64x5 FILLER_344_8 ();
 b15zdnd11an1n64x5 FILLER_344_72 ();
 b15zdnd11an1n64x5 FILLER_344_136 ();
 b15zdnd11an1n08x5 FILLER_344_200 ();
 b15zdnd11an1n04x5 FILLER_344_208 ();
 b15zdnd11an1n04x5 FILLER_344_225 ();
 b15zdnd11an1n08x5 FILLER_344_245 ();
 b15zdnd11an1n04x5 FILLER_344_253 ();
 b15zdnd00an1n02x5 FILLER_344_257 ();
 b15zdnd11an1n32x5 FILLER_344_271 ();
 b15zdnd11an1n04x5 FILLER_344_303 ();
 b15zdnd00an1n01x5 FILLER_344_307 ();
 b15zdnd11an1n08x5 FILLER_344_313 ();
 b15zdnd00an1n02x5 FILLER_344_321 ();
 b15zdnd00an1n01x5 FILLER_344_323 ();
 b15zdnd11an1n32x5 FILLER_344_336 ();
 b15zdnd11an1n16x5 FILLER_344_368 ();
 b15zdnd11an1n08x5 FILLER_344_384 ();
 b15zdnd00an1n02x5 FILLER_344_392 ();
 b15zdnd11an1n04x5 FILLER_344_405 ();
 b15zdnd11an1n64x5 FILLER_344_414 ();
 b15zdnd11an1n16x5 FILLER_344_478 ();
 b15zdnd00an1n02x5 FILLER_344_494 ();
 b15zdnd11an1n04x5 FILLER_344_504 ();
 b15zdnd11an1n16x5 FILLER_344_514 ();
 b15zdnd11an1n08x5 FILLER_344_530 ();
 b15zdnd11an1n04x5 FILLER_344_538 ();
 b15zdnd00an1n02x5 FILLER_344_542 ();
 b15zdnd11an1n08x5 FILLER_344_570 ();
 b15zdnd11an1n04x5 FILLER_344_578 ();
 b15zdnd11an1n04x5 FILLER_344_587 ();
 b15zdnd00an1n02x5 FILLER_344_591 ();
 b15zdnd11an1n64x5 FILLER_344_598 ();
 b15zdnd00an1n01x5 FILLER_344_662 ();
 b15zdnd11an1n32x5 FILLER_344_667 ();
 b15zdnd00an1n02x5 FILLER_344_699 ();
 b15zdnd00an1n01x5 FILLER_344_701 ();
 b15zdnd11an1n08x5 FILLER_344_708 ();
 b15zdnd00an1n02x5 FILLER_344_716 ();
 b15zdnd11an1n64x5 FILLER_344_726 ();
 b15zdnd11an1n04x5 FILLER_344_790 ();
 b15zdnd11an1n16x5 FILLER_344_808 ();
 b15zdnd11an1n04x5 FILLER_344_824 ();
 b15zdnd11an1n16x5 FILLER_344_834 ();
 b15zdnd11an1n08x5 FILLER_344_850 ();
 b15zdnd00an1n02x5 FILLER_344_858 ();
 b15zdnd00an1n01x5 FILLER_344_860 ();
 b15zdnd11an1n32x5 FILLER_344_866 ();
 b15zdnd11an1n08x5 FILLER_344_898 ();
 b15zdnd11an1n04x5 FILLER_344_906 ();
 b15zdnd00an1n01x5 FILLER_344_910 ();
 b15zdnd11an1n16x5 FILLER_344_915 ();
 b15zdnd11an1n08x5 FILLER_344_931 ();
 b15zdnd11an1n04x5 FILLER_344_939 ();
 b15zdnd00an1n02x5 FILLER_344_943 ();
 b15zdnd00an1n01x5 FILLER_344_945 ();
 b15zdnd11an1n04x5 FILLER_344_954 ();
 b15zdnd11an1n16x5 FILLER_344_984 ();
 b15zdnd11an1n08x5 FILLER_344_1000 ();
 b15zdnd00an1n01x5 FILLER_344_1008 ();
 b15zdnd11an1n08x5 FILLER_344_1013 ();
 b15zdnd00an1n01x5 FILLER_344_1021 ();
 b15zdnd11an1n04x5 FILLER_344_1042 ();
 b15zdnd11an1n08x5 FILLER_344_1055 ();
 b15zdnd11an1n04x5 FILLER_344_1063 ();
 b15zdnd00an1n01x5 FILLER_344_1067 ();
 b15zdnd11an1n16x5 FILLER_344_1074 ();
 b15zdnd11an1n08x5 FILLER_344_1090 ();
 b15zdnd11an1n32x5 FILLER_344_1105 ();
 b15zdnd11an1n04x5 FILLER_344_1137 ();
 b15zdnd00an1n02x5 FILLER_344_1141 ();
 b15zdnd00an1n01x5 FILLER_344_1143 ();
 b15zdnd11an1n04x5 FILLER_344_1149 ();
 b15zdnd11an1n04x5 FILLER_344_1172 ();
 b15zdnd00an1n02x5 FILLER_344_1176 ();
 b15zdnd11an1n64x5 FILLER_344_1204 ();
 b15zdnd11an1n32x5 FILLER_344_1268 ();
 b15zdnd11an1n16x5 FILLER_344_1300 ();
 b15zdnd00an1n02x5 FILLER_344_1316 ();
 b15zdnd00an1n01x5 FILLER_344_1318 ();
 b15zdnd11an1n08x5 FILLER_344_1324 ();
 b15zdnd00an1n02x5 FILLER_344_1332 ();
 b15zdnd11an1n64x5 FILLER_344_1344 ();
 b15zdnd11an1n64x5 FILLER_344_1408 ();
 b15zdnd11an1n32x5 FILLER_344_1472 ();
 b15zdnd11an1n16x5 FILLER_344_1504 ();
 b15zdnd11an1n04x5 FILLER_344_1520 ();
 b15zdnd11an1n04x5 FILLER_344_1531 ();
 b15zdnd00an1n02x5 FILLER_344_1535 ();
 b15zdnd00an1n01x5 FILLER_344_1537 ();
 b15zdnd11an1n32x5 FILLER_344_1549 ();
 b15zdnd11an1n16x5 FILLER_344_1581 ();
 b15zdnd00an1n02x5 FILLER_344_1597 ();
 b15zdnd00an1n01x5 FILLER_344_1599 ();
 b15zdnd11an1n16x5 FILLER_344_1606 ();
 b15zdnd11an1n08x5 FILLER_344_1622 ();
 b15zdnd11an1n04x5 FILLER_344_1630 ();
 b15zdnd00an1n01x5 FILLER_344_1634 ();
 b15zdnd11an1n32x5 FILLER_344_1639 ();
 b15zdnd11an1n16x5 FILLER_344_1671 ();
 b15zdnd11an1n04x5 FILLER_344_1687 ();
 b15zdnd00an1n02x5 FILLER_344_1691 ();
 b15zdnd11an1n04x5 FILLER_344_1701 ();
 b15zdnd11an1n04x5 FILLER_344_1717 ();
 b15zdnd11an1n04x5 FILLER_344_1739 ();
 b15zdnd11an1n64x5 FILLER_344_1757 ();
 b15zdnd11an1n64x5 FILLER_344_1821 ();
 b15zdnd11an1n16x5 FILLER_344_1885 ();
 b15zdnd11an1n08x5 FILLER_344_1901 ();
 b15zdnd00an1n02x5 FILLER_344_1909 ();
 b15zdnd00an1n01x5 FILLER_344_1911 ();
 b15zdnd11an1n04x5 FILLER_344_1918 ();
 b15zdnd00an1n02x5 FILLER_344_1922 ();
 b15zdnd11an1n64x5 FILLER_344_1929 ();
 b15zdnd11an1n64x5 FILLER_344_1993 ();
 b15zdnd11an1n64x5 FILLER_344_2064 ();
 b15zdnd11an1n16x5 FILLER_344_2128 ();
 b15zdnd11an1n08x5 FILLER_344_2144 ();
 b15zdnd00an1n02x5 FILLER_344_2152 ();
 b15zdnd11an1n32x5 FILLER_344_2162 ();
 b15zdnd11an1n04x5 FILLER_344_2194 ();
 b15zdnd00an1n02x5 FILLER_344_2198 ();
 b15zdnd00an1n01x5 FILLER_344_2200 ();
 b15zdnd11an1n04x5 FILLER_344_2207 ();
 b15zdnd11an1n32x5 FILLER_344_2217 ();
 b15zdnd11an1n16x5 FILLER_344_2249 ();
 b15zdnd11an1n08x5 FILLER_344_2265 ();
 b15zdnd00an1n02x5 FILLER_344_2273 ();
 b15zdnd00an1n01x5 FILLER_344_2275 ();
 b15zdnd11an1n64x5 FILLER_345_0 ();
 b15zdnd11an1n64x5 FILLER_345_64 ();
 b15zdnd11an1n64x5 FILLER_345_128 ();
 b15zdnd11an1n32x5 FILLER_345_192 ();
 b15zdnd00an1n02x5 FILLER_345_224 ();
 b15zdnd11an1n08x5 FILLER_345_236 ();
 b15zdnd00an1n01x5 FILLER_345_244 ();
 b15zdnd11an1n04x5 FILLER_345_252 ();
 b15zdnd11an1n32x5 FILLER_345_268 ();
 b15zdnd11an1n08x5 FILLER_345_300 ();
 b15zdnd11an1n64x5 FILLER_345_313 ();
 b15zdnd11an1n16x5 FILLER_345_377 ();
 b15zdnd11an1n04x5 FILLER_345_405 ();
 b15zdnd11an1n08x5 FILLER_345_419 ();
 b15zdnd00an1n01x5 FILLER_345_427 ();
 b15zdnd11an1n04x5 FILLER_345_454 ();
 b15zdnd11an1n16x5 FILLER_345_467 ();
 b15zdnd11an1n16x5 FILLER_345_489 ();
 b15zdnd11an1n04x5 FILLER_345_505 ();
 b15zdnd00an1n02x5 FILLER_345_509 ();
 b15zdnd11an1n64x5 FILLER_345_520 ();
 b15zdnd11an1n64x5 FILLER_345_584 ();
 b15zdnd11an1n32x5 FILLER_345_648 ();
 b15zdnd11an1n04x5 FILLER_345_680 ();
 b15zdnd00an1n02x5 FILLER_345_684 ();
 b15zdnd11an1n32x5 FILLER_345_696 ();
 b15zdnd11an1n08x5 FILLER_345_728 ();
 b15zdnd11an1n32x5 FILLER_345_742 ();
 b15zdnd11an1n16x5 FILLER_345_774 ();
 b15zdnd11an1n04x5 FILLER_345_790 ();
 b15zdnd00an1n01x5 FILLER_345_794 ();
 b15zdnd11an1n08x5 FILLER_345_810 ();
 b15zdnd00an1n01x5 FILLER_345_818 ();
 b15zdnd11an1n04x5 FILLER_345_836 ();
 b15zdnd11an1n32x5 FILLER_345_862 ();
 b15zdnd11an1n04x5 FILLER_345_894 ();
 b15zdnd00an1n02x5 FILLER_345_898 ();
 b15zdnd00an1n01x5 FILLER_345_900 ();
 b15zdnd11an1n04x5 FILLER_345_905 ();
 b15zdnd11an1n32x5 FILLER_345_922 ();
 b15zdnd00an1n01x5 FILLER_345_954 ();
 b15zdnd11an1n04x5 FILLER_345_963 ();
 b15zdnd11an1n04x5 FILLER_345_979 ();
 b15zdnd11an1n08x5 FILLER_345_990 ();
 b15zdnd11an1n04x5 FILLER_345_998 ();
 b15zdnd00an1n01x5 FILLER_345_1002 ();
 b15zdnd11an1n32x5 FILLER_345_1009 ();
 b15zdnd11an1n08x5 FILLER_345_1041 ();
 b15zdnd11an1n04x5 FILLER_345_1049 ();
 b15zdnd00an1n02x5 FILLER_345_1053 ();
 b15zdnd00an1n01x5 FILLER_345_1055 ();
 b15zdnd11an1n04x5 FILLER_345_1067 ();
 b15zdnd11an1n16x5 FILLER_345_1076 ();
 b15zdnd11an1n08x5 FILLER_345_1092 ();
 b15zdnd11an1n16x5 FILLER_345_1105 ();
 b15zdnd11an1n08x5 FILLER_345_1121 ();
 b15zdnd11an1n04x5 FILLER_345_1129 ();
 b15zdnd00an1n01x5 FILLER_345_1133 ();
 b15zdnd11an1n04x5 FILLER_345_1142 ();
 b15zdnd11an1n04x5 FILLER_345_1151 ();
 b15zdnd11an1n64x5 FILLER_345_1181 ();
 b15zdnd11an1n16x5 FILLER_345_1245 ();
 b15zdnd00an1n02x5 FILLER_345_1261 ();
 b15zdnd11an1n16x5 FILLER_345_1279 ();
 b15zdnd00an1n02x5 FILLER_345_1295 ();
 b15zdnd00an1n01x5 FILLER_345_1297 ();
 b15zdnd11an1n32x5 FILLER_345_1314 ();
 b15zdnd11an1n16x5 FILLER_345_1346 ();
 b15zdnd00an1n01x5 FILLER_345_1362 ();
 b15zdnd11an1n16x5 FILLER_345_1372 ();
 b15zdnd11an1n04x5 FILLER_345_1388 ();
 b15zdnd11an1n16x5 FILLER_345_1401 ();
 b15zdnd11an1n08x5 FILLER_345_1417 ();
 b15zdnd11an1n04x5 FILLER_345_1425 ();
 b15zdnd00an1n01x5 FILLER_345_1429 ();
 b15zdnd11an1n32x5 FILLER_345_1436 ();
 b15zdnd11an1n08x5 FILLER_345_1468 ();
 b15zdnd11an1n04x5 FILLER_345_1476 ();
 b15zdnd11an1n04x5 FILLER_345_1486 ();
 b15zdnd11an1n04x5 FILLER_345_1494 ();
 b15zdnd00an1n01x5 FILLER_345_1498 ();
 b15zdnd11an1n64x5 FILLER_345_1505 ();
 b15zdnd11an1n16x5 FILLER_345_1569 ();
 b15zdnd11an1n08x5 FILLER_345_1585 ();
 b15zdnd11an1n04x5 FILLER_345_1593 ();
 b15zdnd00an1n02x5 FILLER_345_1597 ();
 b15zdnd11an1n32x5 FILLER_345_1604 ();
 b15zdnd11an1n64x5 FILLER_345_1642 ();
 b15zdnd11an1n16x5 FILLER_345_1706 ();
 b15zdnd00an1n02x5 FILLER_345_1722 ();
 b15zdnd00an1n01x5 FILLER_345_1724 ();
 b15zdnd11an1n64x5 FILLER_345_1734 ();
 b15zdnd11an1n04x5 FILLER_345_1798 ();
 b15zdnd11an1n08x5 FILLER_345_1807 ();
 b15zdnd11an1n16x5 FILLER_345_1833 ();
 b15zdnd00an1n02x5 FILLER_345_1849 ();
 b15zdnd00an1n01x5 FILLER_345_1851 ();
 b15zdnd11an1n32x5 FILLER_345_1857 ();
 b15zdnd11an1n04x5 FILLER_345_1889 ();
 b15zdnd11an1n64x5 FILLER_345_1908 ();
 b15zdnd11an1n04x5 FILLER_345_1972 ();
 b15zdnd00an1n02x5 FILLER_345_1976 ();
 b15zdnd11an1n16x5 FILLER_345_1985 ();
 b15zdnd11an1n08x5 FILLER_345_2001 ();
 b15zdnd11an1n04x5 FILLER_345_2009 ();
 b15zdnd00an1n01x5 FILLER_345_2013 ();
 b15zdnd11an1n64x5 FILLER_345_2018 ();
 b15zdnd11an1n32x5 FILLER_345_2082 ();
 b15zdnd11an1n16x5 FILLER_345_2114 ();
 b15zdnd11an1n08x5 FILLER_345_2130 ();
 b15zdnd11an1n04x5 FILLER_345_2138 ();
 b15zdnd11an1n32x5 FILLER_345_2150 ();
 b15zdnd11an1n08x5 FILLER_345_2182 ();
 b15zdnd11an1n04x5 FILLER_345_2190 ();
 b15zdnd11an1n04x5 FILLER_345_2199 ();
 b15zdnd11an1n04x5 FILLER_345_2208 ();
 b15zdnd11an1n64x5 FILLER_345_2218 ();
 b15zdnd00an1n02x5 FILLER_345_2282 ();
 b15zdnd11an1n64x5 FILLER_346_8 ();
 b15zdnd11an1n64x5 FILLER_346_72 ();
 b15zdnd11an1n64x5 FILLER_346_136 ();
 b15zdnd11an1n32x5 FILLER_346_200 ();
 b15zdnd11an1n08x5 FILLER_346_232 ();
 b15zdnd11an1n04x5 FILLER_346_240 ();
 b15zdnd00an1n02x5 FILLER_346_244 ();
 b15zdnd00an1n01x5 FILLER_346_246 ();
 b15zdnd11an1n16x5 FILLER_346_270 ();
 b15zdnd11an1n32x5 FILLER_346_298 ();
 b15zdnd11an1n16x5 FILLER_346_330 ();
 b15zdnd11an1n04x5 FILLER_346_346 ();
 b15zdnd11an1n08x5 FILLER_346_359 ();
 b15zdnd11an1n04x5 FILLER_346_367 ();
 b15zdnd00an1n01x5 FILLER_346_371 ();
 b15zdnd11an1n64x5 FILLER_346_376 ();
 b15zdnd11an1n16x5 FILLER_346_440 ();
 b15zdnd11an1n08x5 FILLER_346_456 ();
 b15zdnd11an1n16x5 FILLER_346_480 ();
 b15zdnd11an1n08x5 FILLER_346_496 ();
 b15zdnd00an1n02x5 FILLER_346_504 ();
 b15zdnd11an1n04x5 FILLER_346_527 ();
 b15zdnd11an1n08x5 FILLER_346_537 ();
 b15zdnd11an1n04x5 FILLER_346_550 ();
 b15zdnd11an1n64x5 FILLER_346_558 ();
 b15zdnd11an1n32x5 FILLER_346_622 ();
 b15zdnd11an1n16x5 FILLER_346_654 ();
 b15zdnd11an1n08x5 FILLER_346_670 ();
 b15zdnd11an1n04x5 FILLER_346_678 ();
 b15zdnd00an1n01x5 FILLER_346_682 ();
 b15zdnd11an1n08x5 FILLER_346_689 ();
 b15zdnd00an1n02x5 FILLER_346_697 ();
 b15zdnd11an1n04x5 FILLER_346_711 ();
 b15zdnd00an1n02x5 FILLER_346_715 ();
 b15zdnd00an1n01x5 FILLER_346_717 ();
 b15zdnd11an1n32x5 FILLER_346_726 ();
 b15zdnd11an1n04x5 FILLER_346_758 ();
 b15zdnd00an1n02x5 FILLER_346_762 ();
 b15zdnd11an1n64x5 FILLER_346_772 ();
 b15zdnd11an1n64x5 FILLER_346_836 ();
 b15zdnd11an1n16x5 FILLER_346_900 ();
 b15zdnd11an1n08x5 FILLER_346_916 ();
 b15zdnd11an1n04x5 FILLER_346_924 ();
 b15zdnd00an1n02x5 FILLER_346_928 ();
 b15zdnd00an1n01x5 FILLER_346_930 ();
 b15zdnd11an1n08x5 FILLER_346_938 ();
 b15zdnd11an1n04x5 FILLER_346_946 ();
 b15zdnd00an1n01x5 FILLER_346_950 ();
 b15zdnd11an1n04x5 FILLER_346_960 ();
 b15zdnd11an1n32x5 FILLER_346_969 ();
 b15zdnd11an1n04x5 FILLER_346_1001 ();
 b15zdnd00an1n02x5 FILLER_346_1005 ();
 b15zdnd00an1n01x5 FILLER_346_1007 ();
 b15zdnd11an1n64x5 FILLER_346_1024 ();
 b15zdnd11an1n16x5 FILLER_346_1088 ();
 b15zdnd00an1n02x5 FILLER_346_1104 ();
 b15zdnd00an1n01x5 FILLER_346_1106 ();
 b15zdnd11an1n16x5 FILLER_346_1118 ();
 b15zdnd11an1n04x5 FILLER_346_1141 ();
 b15zdnd11an1n16x5 FILLER_346_1150 ();
 b15zdnd11an1n04x5 FILLER_346_1166 ();
 b15zdnd00an1n01x5 FILLER_346_1170 ();
 b15zdnd11an1n64x5 FILLER_346_1181 ();
 b15zdnd11an1n04x5 FILLER_346_1245 ();
 b15zdnd00an1n01x5 FILLER_346_1249 ();
 b15zdnd11an1n64x5 FILLER_346_1270 ();
 b15zdnd11an1n08x5 FILLER_346_1334 ();
 b15zdnd11an1n04x5 FILLER_346_1342 ();
 b15zdnd11an1n04x5 FILLER_346_1356 ();
 b15zdnd11an1n16x5 FILLER_346_1380 ();
 b15zdnd00an1n01x5 FILLER_346_1396 ();
 b15zdnd11an1n16x5 FILLER_346_1409 ();
 b15zdnd00an1n01x5 FILLER_346_1425 ();
 b15zdnd11an1n32x5 FILLER_346_1438 ();
 b15zdnd11an1n04x5 FILLER_346_1470 ();
 b15zdnd00an1n02x5 FILLER_346_1474 ();
 b15zdnd00an1n01x5 FILLER_346_1476 ();
 b15zdnd11an1n64x5 FILLER_346_1483 ();
 b15zdnd11an1n16x5 FILLER_346_1547 ();
 b15zdnd00an1n02x5 FILLER_346_1563 ();
 b15zdnd11an1n16x5 FILLER_346_1570 ();
 b15zdnd11an1n08x5 FILLER_346_1586 ();
 b15zdnd00an1n02x5 FILLER_346_1594 ();
 b15zdnd00an1n01x5 FILLER_346_1596 ();
 b15zdnd11an1n16x5 FILLER_346_1611 ();
 b15zdnd00an1n02x5 FILLER_346_1627 ();
 b15zdnd11an1n04x5 FILLER_346_1641 ();
 b15zdnd11an1n08x5 FILLER_346_1650 ();
 b15zdnd11an1n04x5 FILLER_346_1658 ();
 b15zdnd00an1n02x5 FILLER_346_1662 ();
 b15zdnd00an1n01x5 FILLER_346_1664 ();
 b15zdnd11an1n64x5 FILLER_346_1669 ();
 b15zdnd11an1n32x5 FILLER_346_1747 ();
 b15zdnd11an1n16x5 FILLER_346_1779 ();
 b15zdnd11an1n08x5 FILLER_346_1795 ();
 b15zdnd11an1n04x5 FILLER_346_1803 ();
 b15zdnd00an1n01x5 FILLER_346_1807 ();
 b15zdnd11an1n16x5 FILLER_346_1817 ();
 b15zdnd11an1n08x5 FILLER_346_1833 ();
 b15zdnd11an1n04x5 FILLER_346_1841 ();
 b15zdnd00an1n02x5 FILLER_346_1845 ();
 b15zdnd11an1n16x5 FILLER_346_1854 ();
 b15zdnd11an1n04x5 FILLER_346_1870 ();
 b15zdnd00an1n02x5 FILLER_346_1874 ();
 b15zdnd00an1n01x5 FILLER_346_1876 ();
 b15zdnd11an1n32x5 FILLER_346_1883 ();
 b15zdnd11an1n08x5 FILLER_346_1915 ();
 b15zdnd00an1n01x5 FILLER_346_1923 ();
 b15zdnd11an1n16x5 FILLER_346_1935 ();
 b15zdnd11an1n04x5 FILLER_346_1957 ();
 b15zdnd11an1n08x5 FILLER_346_1966 ();
 b15zdnd00an1n02x5 FILLER_346_1974 ();
 b15zdnd11an1n16x5 FILLER_346_1984 ();
 b15zdnd11an1n04x5 FILLER_346_2000 ();
 b15zdnd00an1n01x5 FILLER_346_2004 ();
 b15zdnd11an1n32x5 FILLER_346_2012 ();
 b15zdnd11an1n04x5 FILLER_346_2044 ();
 b15zdnd00an1n02x5 FILLER_346_2048 ();
 b15zdnd00an1n01x5 FILLER_346_2050 ();
 b15zdnd11an1n16x5 FILLER_346_2057 ();
 b15zdnd00an1n02x5 FILLER_346_2073 ();
 b15zdnd11an1n32x5 FILLER_346_2100 ();
 b15zdnd11an1n16x5 FILLER_346_2132 ();
 b15zdnd11an1n04x5 FILLER_346_2148 ();
 b15zdnd00an1n02x5 FILLER_346_2152 ();
 b15zdnd11an1n32x5 FILLER_346_2162 ();
 b15zdnd00an1n02x5 FILLER_346_2194 ();
 b15zdnd11an1n64x5 FILLER_346_2208 ();
 b15zdnd11an1n04x5 FILLER_346_2272 ();
 b15zdnd11an1n64x5 FILLER_347_0 ();
 b15zdnd11an1n64x5 FILLER_347_64 ();
 b15zdnd11an1n64x5 FILLER_347_128 ();
 b15zdnd11an1n64x5 FILLER_347_192 ();
 b15zdnd11an1n32x5 FILLER_347_256 ();
 b15zdnd11an1n04x5 FILLER_347_288 ();
 b15zdnd11an1n04x5 FILLER_347_308 ();
 b15zdnd11an1n16x5 FILLER_347_317 ();
 b15zdnd11an1n04x5 FILLER_347_333 ();
 b15zdnd00an1n01x5 FILLER_347_337 ();
 b15zdnd11an1n04x5 FILLER_347_347 ();
 b15zdnd11an1n04x5 FILLER_347_372 ();
 b15zdnd11an1n04x5 FILLER_347_386 ();
 b15zdnd11an1n64x5 FILLER_347_397 ();
 b15zdnd11an1n64x5 FILLER_347_461 ();
 b15zdnd11an1n16x5 FILLER_347_525 ();
 b15zdnd11an1n04x5 FILLER_347_541 ();
 b15zdnd00an1n02x5 FILLER_347_545 ();
 b15zdnd00an1n01x5 FILLER_347_547 ();
 b15zdnd11an1n16x5 FILLER_347_558 ();
 b15zdnd11an1n04x5 FILLER_347_574 ();
 b15zdnd11an1n64x5 FILLER_347_584 ();
 b15zdnd11an1n04x5 FILLER_347_648 ();
 b15zdnd00an1n02x5 FILLER_347_652 ();
 b15zdnd11an1n32x5 FILLER_347_659 ();
 b15zdnd11an1n04x5 FILLER_347_691 ();
 b15zdnd00an1n02x5 FILLER_347_695 ();
 b15zdnd00an1n01x5 FILLER_347_697 ();
 b15zdnd11an1n32x5 FILLER_347_712 ();
 b15zdnd11an1n08x5 FILLER_347_744 ();
 b15zdnd11an1n04x5 FILLER_347_752 ();
 b15zdnd11an1n04x5 FILLER_347_767 ();
 b15zdnd00an1n01x5 FILLER_347_771 ();
 b15zdnd11an1n64x5 FILLER_347_777 ();
 b15zdnd11an1n64x5 FILLER_347_841 ();
 b15zdnd11an1n08x5 FILLER_347_905 ();
 b15zdnd11an1n04x5 FILLER_347_913 ();
 b15zdnd11an1n04x5 FILLER_347_932 ();
 b15zdnd11an1n08x5 FILLER_347_941 ();
 b15zdnd11an1n04x5 FILLER_347_949 ();
 b15zdnd00an1n02x5 FILLER_347_953 ();
 b15zdnd11an1n64x5 FILLER_347_959 ();
 b15zdnd11an1n64x5 FILLER_347_1023 ();
 b15zdnd11an1n32x5 FILLER_347_1087 ();
 b15zdnd11an1n16x5 FILLER_347_1119 ();
 b15zdnd00an1n01x5 FILLER_347_1135 ();
 b15zdnd11an1n64x5 FILLER_347_1143 ();
 b15zdnd11an1n32x5 FILLER_347_1207 ();
 b15zdnd11an1n08x5 FILLER_347_1239 ();
 b15zdnd11an1n04x5 FILLER_347_1247 ();
 b15zdnd00an1n02x5 FILLER_347_1251 ();
 b15zdnd00an1n01x5 FILLER_347_1253 ();
 b15zdnd11an1n04x5 FILLER_347_1258 ();
 b15zdnd11an1n16x5 FILLER_347_1268 ();
 b15zdnd00an1n02x5 FILLER_347_1284 ();
 b15zdnd11an1n32x5 FILLER_347_1295 ();
 b15zdnd11an1n16x5 FILLER_347_1327 ();
 b15zdnd11an1n04x5 FILLER_347_1354 ();
 b15zdnd11an1n08x5 FILLER_347_1364 ();
 b15zdnd11an1n04x5 FILLER_347_1372 ();
 b15zdnd11an1n08x5 FILLER_347_1382 ();
 b15zdnd00an1n02x5 FILLER_347_1390 ();
 b15zdnd11an1n08x5 FILLER_347_1418 ();
 b15zdnd00an1n02x5 FILLER_347_1426 ();
 b15zdnd00an1n01x5 FILLER_347_1428 ();
 b15zdnd11an1n32x5 FILLER_347_1441 ();
 b15zdnd00an1n02x5 FILLER_347_1473 ();
 b15zdnd00an1n01x5 FILLER_347_1475 ();
 b15zdnd11an1n64x5 FILLER_347_1482 ();
 b15zdnd00an1n01x5 FILLER_347_1546 ();
 b15zdnd11an1n04x5 FILLER_347_1552 ();
 b15zdnd11an1n04x5 FILLER_347_1563 ();
 b15zdnd11an1n16x5 FILLER_347_1581 ();
 b15zdnd11an1n04x5 FILLER_347_1597 ();
 b15zdnd11an1n04x5 FILLER_347_1620 ();
 b15zdnd11an1n16x5 FILLER_347_1639 ();
 b15zdnd11an1n08x5 FILLER_347_1655 ();
 b15zdnd00an1n02x5 FILLER_347_1663 ();
 b15zdnd11an1n04x5 FILLER_347_1677 ();
 b15zdnd11an1n32x5 FILLER_347_1685 ();
 b15zdnd11an1n16x5 FILLER_347_1717 ();
 b15zdnd00an1n02x5 FILLER_347_1733 ();
 b15zdnd00an1n01x5 FILLER_347_1735 ();
 b15zdnd11an1n64x5 FILLER_347_1752 ();
 b15zdnd00an1n02x5 FILLER_347_1816 ();
 b15zdnd00an1n01x5 FILLER_347_1818 ();
 b15zdnd11an1n16x5 FILLER_347_1824 ();
 b15zdnd11an1n04x5 FILLER_347_1840 ();
 b15zdnd00an1n02x5 FILLER_347_1844 ();
 b15zdnd00an1n01x5 FILLER_347_1846 ();
 b15zdnd11an1n32x5 FILLER_347_1853 ();
 b15zdnd11an1n16x5 FILLER_347_1885 ();
 b15zdnd00an1n01x5 FILLER_347_1901 ();
 b15zdnd11an1n64x5 FILLER_347_1907 ();
 b15zdnd11an1n32x5 FILLER_347_1971 ();
 b15zdnd00an1n01x5 FILLER_347_2003 ();
 b15zdnd11an1n16x5 FILLER_347_2017 ();
 b15zdnd11an1n04x5 FILLER_347_2033 ();
 b15zdnd11an1n04x5 FILLER_347_2049 ();
 b15zdnd11an1n04x5 FILLER_347_2071 ();
 b15zdnd11an1n04x5 FILLER_347_2088 ();
 b15zdnd11an1n04x5 FILLER_347_2102 ();
 b15zdnd11an1n64x5 FILLER_347_2110 ();
 b15zdnd00an1n01x5 FILLER_347_2174 ();
 b15zdnd11an1n16x5 FILLER_347_2180 ();
 b15zdnd11an1n08x5 FILLER_347_2196 ();
 b15zdnd00an1n02x5 FILLER_347_2204 ();
 b15zdnd11an1n64x5 FILLER_347_2212 ();
 b15zdnd11an1n08x5 FILLER_347_2276 ();
 b15zdnd11an1n64x5 FILLER_348_8 ();
 b15zdnd11an1n64x5 FILLER_348_72 ();
 b15zdnd11an1n64x5 FILLER_348_136 ();
 b15zdnd11an1n16x5 FILLER_348_200 ();
 b15zdnd11an1n08x5 FILLER_348_216 ();
 b15zdnd11an1n08x5 FILLER_348_228 ();
 b15zdnd11an1n08x5 FILLER_348_240 ();
 b15zdnd11an1n16x5 FILLER_348_260 ();
 b15zdnd11an1n08x5 FILLER_348_276 ();
 b15zdnd11an1n64x5 FILLER_348_304 ();
 b15zdnd11an1n64x5 FILLER_348_368 ();
 b15zdnd11an1n16x5 FILLER_348_432 ();
 b15zdnd11an1n04x5 FILLER_348_448 ();
 b15zdnd00an1n02x5 FILLER_348_452 ();
 b15zdnd00an1n01x5 FILLER_348_454 ();
 b15zdnd11an1n04x5 FILLER_348_471 ();
 b15zdnd11an1n08x5 FILLER_348_481 ();
 b15zdnd11an1n04x5 FILLER_348_489 ();
 b15zdnd00an1n02x5 FILLER_348_493 ();
 b15zdnd11an1n16x5 FILLER_348_502 ();
 b15zdnd11an1n08x5 FILLER_348_518 ();
 b15zdnd11an1n04x5 FILLER_348_526 ();
 b15zdnd00an1n01x5 FILLER_348_530 ();
 b15zdnd11an1n32x5 FILLER_348_540 ();
 b15zdnd11an1n04x5 FILLER_348_581 ();
 b15zdnd00an1n01x5 FILLER_348_585 ();
 b15zdnd11an1n32x5 FILLER_348_592 ();
 b15zdnd11an1n16x5 FILLER_348_624 ();
 b15zdnd11an1n08x5 FILLER_348_640 ();
 b15zdnd11an1n04x5 FILLER_348_648 ();
 b15zdnd00an1n02x5 FILLER_348_652 ();
 b15zdnd00an1n01x5 FILLER_348_654 ();
 b15zdnd11an1n32x5 FILLER_348_665 ();
 b15zdnd11an1n08x5 FILLER_348_697 ();
 b15zdnd11an1n04x5 FILLER_348_705 ();
 b15zdnd00an1n02x5 FILLER_348_709 ();
 b15zdnd00an1n01x5 FILLER_348_711 ();
 b15zdnd00an1n02x5 FILLER_348_716 ();
 b15zdnd11an1n32x5 FILLER_348_726 ();
 b15zdnd11an1n04x5 FILLER_348_758 ();
 b15zdnd00an1n02x5 FILLER_348_762 ();
 b15zdnd00an1n01x5 FILLER_348_764 ();
 b15zdnd11an1n04x5 FILLER_348_771 ();
 b15zdnd11an1n04x5 FILLER_348_787 ();
 b15zdnd00an1n01x5 FILLER_348_791 ();
 b15zdnd11an1n08x5 FILLER_348_796 ();
 b15zdnd11an1n64x5 FILLER_348_809 ();
 b15zdnd11an1n32x5 FILLER_348_873 ();
 b15zdnd11an1n16x5 FILLER_348_905 ();
 b15zdnd11an1n04x5 FILLER_348_921 ();
 b15zdnd00an1n02x5 FILLER_348_925 ();
 b15zdnd11an1n64x5 FILLER_348_943 ();
 b15zdnd11an1n64x5 FILLER_348_1007 ();
 b15zdnd11an1n64x5 FILLER_348_1071 ();
 b15zdnd11an1n32x5 FILLER_348_1135 ();
 b15zdnd11an1n08x5 FILLER_348_1167 ();
 b15zdnd11an1n04x5 FILLER_348_1175 ();
 b15zdnd00an1n02x5 FILLER_348_1179 ();
 b15zdnd00an1n01x5 FILLER_348_1181 ();
 b15zdnd11an1n64x5 FILLER_348_1189 ();
 b15zdnd11an1n16x5 FILLER_348_1253 ();
 b15zdnd00an1n01x5 FILLER_348_1269 ();
 b15zdnd11an1n32x5 FILLER_348_1275 ();
 b15zdnd11an1n08x5 FILLER_348_1307 ();
 b15zdnd00an1n02x5 FILLER_348_1315 ();
 b15zdnd00an1n01x5 FILLER_348_1317 ();
 b15zdnd11an1n32x5 FILLER_348_1327 ();
 b15zdnd11an1n16x5 FILLER_348_1365 ();
 b15zdnd11an1n04x5 FILLER_348_1381 ();
 b15zdnd00an1n01x5 FILLER_348_1385 ();
 b15zdnd11an1n32x5 FILLER_348_1396 ();
 b15zdnd00an1n02x5 FILLER_348_1428 ();
 b15zdnd11an1n32x5 FILLER_348_1442 ();
 b15zdnd11an1n16x5 FILLER_348_1474 ();
 b15zdnd11an1n04x5 FILLER_348_1490 ();
 b15zdnd00an1n02x5 FILLER_348_1494 ();
 b15zdnd11an1n32x5 FILLER_348_1502 ();
 b15zdnd11an1n04x5 FILLER_348_1534 ();
 b15zdnd00an1n02x5 FILLER_348_1538 ();
 b15zdnd11an1n08x5 FILLER_348_1554 ();
 b15zdnd00an1n02x5 FILLER_348_1562 ();
 b15zdnd11an1n16x5 FILLER_348_1568 ();
 b15zdnd11an1n08x5 FILLER_348_1584 ();
 b15zdnd11an1n04x5 FILLER_348_1592 ();
 b15zdnd00an1n02x5 FILLER_348_1596 ();
 b15zdnd00an1n01x5 FILLER_348_1598 ();
 b15zdnd11an1n32x5 FILLER_348_1619 ();
 b15zdnd11an1n16x5 FILLER_348_1651 ();
 b15zdnd11an1n08x5 FILLER_348_1667 ();
 b15zdnd11an1n04x5 FILLER_348_1675 ();
 b15zdnd11an1n16x5 FILLER_348_1695 ();
 b15zdnd11an1n64x5 FILLER_348_1721 ();
 b15zdnd11an1n32x5 FILLER_348_1785 ();
 b15zdnd11an1n16x5 FILLER_348_1817 ();
 b15zdnd11an1n08x5 FILLER_348_1833 ();
 b15zdnd00an1n02x5 FILLER_348_1841 ();
 b15zdnd00an1n01x5 FILLER_348_1843 ();
 b15zdnd11an1n04x5 FILLER_348_1853 ();
 b15zdnd00an1n02x5 FILLER_348_1857 ();
 b15zdnd11an1n16x5 FILLER_348_1885 ();
 b15zdnd11an1n32x5 FILLER_348_1908 ();
 b15zdnd11an1n04x5 FILLER_348_1945 ();
 b15zdnd00an1n02x5 FILLER_348_1949 ();
 b15zdnd00an1n01x5 FILLER_348_1951 ();
 b15zdnd11an1n16x5 FILLER_348_1961 ();
 b15zdnd00an1n02x5 FILLER_348_1977 ();
 b15zdnd11an1n32x5 FILLER_348_1999 ();
 b15zdnd11an1n08x5 FILLER_348_2031 ();
 b15zdnd11an1n04x5 FILLER_348_2039 ();
 b15zdnd00an1n02x5 FILLER_348_2043 ();
 b15zdnd00an1n01x5 FILLER_348_2045 ();
 b15zdnd11an1n04x5 FILLER_348_2052 ();
 b15zdnd00an1n02x5 FILLER_348_2056 ();
 b15zdnd11an1n08x5 FILLER_348_2063 ();
 b15zdnd00an1n02x5 FILLER_348_2071 ();
 b15zdnd00an1n01x5 FILLER_348_2073 ();
 b15zdnd11an1n16x5 FILLER_348_2080 ();
 b15zdnd00an1n02x5 FILLER_348_2096 ();
 b15zdnd00an1n01x5 FILLER_348_2098 ();
 b15zdnd11an1n16x5 FILLER_348_2105 ();
 b15zdnd11an1n04x5 FILLER_348_2121 ();
 b15zdnd00an1n01x5 FILLER_348_2125 ();
 b15zdnd11an1n04x5 FILLER_348_2133 ();
 b15zdnd00an1n02x5 FILLER_348_2152 ();
 b15zdnd11an1n04x5 FILLER_348_2162 ();
 b15zdnd00an1n01x5 FILLER_348_2166 ();
 b15zdnd11an1n16x5 FILLER_348_2171 ();
 b15zdnd11an1n04x5 FILLER_348_2187 ();
 b15zdnd00an1n02x5 FILLER_348_2191 ();
 b15zdnd11an1n16x5 FILLER_348_2200 ();
 b15zdnd00an1n01x5 FILLER_348_2216 ();
 b15zdnd11an1n32x5 FILLER_348_2226 ();
 b15zdnd11an1n16x5 FILLER_348_2258 ();
 b15zdnd00an1n02x5 FILLER_348_2274 ();
 b15zdnd11an1n64x5 FILLER_349_0 ();
 b15zdnd11an1n64x5 FILLER_349_64 ();
 b15zdnd11an1n64x5 FILLER_349_128 ();
 b15zdnd11an1n16x5 FILLER_349_192 ();
 b15zdnd11an1n08x5 FILLER_349_208 ();
 b15zdnd11an1n04x5 FILLER_349_216 ();
 b15zdnd00an1n01x5 FILLER_349_220 ();
 b15zdnd11an1n32x5 FILLER_349_228 ();
 b15zdnd11an1n04x5 FILLER_349_260 ();
 b15zdnd00an1n01x5 FILLER_349_264 ();
 b15zdnd11an1n32x5 FILLER_349_270 ();
 b15zdnd00an1n02x5 FILLER_349_302 ();
 b15zdnd11an1n16x5 FILLER_349_309 ();
 b15zdnd11an1n04x5 FILLER_349_325 ();
 b15zdnd00an1n01x5 FILLER_349_329 ();
 b15zdnd11an1n32x5 FILLER_349_337 ();
 b15zdnd11an1n08x5 FILLER_349_369 ();
 b15zdnd00an1n02x5 FILLER_349_377 ();
 b15zdnd00an1n01x5 FILLER_349_379 ();
 b15zdnd11an1n04x5 FILLER_349_386 ();
 b15zdnd11an1n08x5 FILLER_349_402 ();
 b15zdnd11an1n04x5 FILLER_349_410 ();
 b15zdnd00an1n02x5 FILLER_349_414 ();
 b15zdnd11an1n32x5 FILLER_349_420 ();
 b15zdnd00an1n02x5 FILLER_349_452 ();
 b15zdnd00an1n01x5 FILLER_349_454 ();
 b15zdnd11an1n04x5 FILLER_349_460 ();
 b15zdnd11an1n16x5 FILLER_349_468 ();
 b15zdnd11an1n04x5 FILLER_349_490 ();
 b15zdnd11an1n08x5 FILLER_349_499 ();
 b15zdnd11an1n04x5 FILLER_349_507 ();
 b15zdnd00an1n01x5 FILLER_349_511 ();
 b15zdnd11an1n32x5 FILLER_349_516 ();
 b15zdnd11an1n16x5 FILLER_349_548 ();
 b15zdnd11an1n04x5 FILLER_349_564 ();
 b15zdnd00an1n02x5 FILLER_349_568 ();
 b15zdnd00an1n01x5 FILLER_349_570 ();
 b15zdnd11an1n04x5 FILLER_349_580 ();
 b15zdnd11an1n32x5 FILLER_349_594 ();
 b15zdnd11an1n16x5 FILLER_349_626 ();
 b15zdnd11an1n08x5 FILLER_349_642 ();
 b15zdnd11an1n04x5 FILLER_349_650 ();
 b15zdnd00an1n02x5 FILLER_349_654 ();
 b15zdnd00an1n01x5 FILLER_349_656 ();
 b15zdnd11an1n04x5 FILLER_349_670 ();
 b15zdnd11an1n04x5 FILLER_349_683 ();
 b15zdnd11an1n08x5 FILLER_349_693 ();
 b15zdnd11an1n04x5 FILLER_349_701 ();
 b15zdnd11an1n16x5 FILLER_349_720 ();
 b15zdnd11an1n08x5 FILLER_349_736 ();
 b15zdnd11an1n04x5 FILLER_349_744 ();
 b15zdnd11an1n32x5 FILLER_349_756 ();
 b15zdnd11an1n16x5 FILLER_349_788 ();
 b15zdnd00an1n01x5 FILLER_349_804 ();
 b15zdnd11an1n08x5 FILLER_349_810 ();
 b15zdnd11an1n04x5 FILLER_349_818 ();
 b15zdnd00an1n02x5 FILLER_349_822 ();
 b15zdnd00an1n01x5 FILLER_349_824 ();
 b15zdnd11an1n04x5 FILLER_349_835 ();
 b15zdnd11an1n16x5 FILLER_349_844 ();
 b15zdnd11an1n08x5 FILLER_349_860 ();
 b15zdnd11an1n04x5 FILLER_349_868 ();
 b15zdnd00an1n01x5 FILLER_349_872 ();
 b15zdnd11an1n08x5 FILLER_349_882 ();
 b15zdnd11an1n64x5 FILLER_349_894 ();
 b15zdnd11an1n64x5 FILLER_349_958 ();
 b15zdnd11an1n08x5 FILLER_349_1022 ();
 b15zdnd00an1n02x5 FILLER_349_1030 ();
 b15zdnd00an1n01x5 FILLER_349_1032 ();
 b15zdnd11an1n64x5 FILLER_349_1037 ();
 b15zdnd11an1n08x5 FILLER_349_1101 ();
 b15zdnd11an1n16x5 FILLER_349_1113 ();
 b15zdnd11an1n08x5 FILLER_349_1129 ();
 b15zdnd00an1n01x5 FILLER_349_1137 ();
 b15zdnd11an1n16x5 FILLER_349_1146 ();
 b15zdnd00an1n01x5 FILLER_349_1162 ();
 b15zdnd11an1n08x5 FILLER_349_1170 ();
 b15zdnd00an1n01x5 FILLER_349_1178 ();
 b15zdnd11an1n04x5 FILLER_349_1185 ();
 b15zdnd11an1n64x5 FILLER_349_1194 ();
 b15zdnd00an1n02x5 FILLER_349_1258 ();
 b15zdnd00an1n01x5 FILLER_349_1260 ();
 b15zdnd11an1n32x5 FILLER_349_1271 ();
 b15zdnd11an1n08x5 FILLER_349_1303 ();
 b15zdnd11an1n04x5 FILLER_349_1311 ();
 b15zdnd11an1n64x5 FILLER_349_1322 ();
 b15zdnd11an1n64x5 FILLER_349_1386 ();
 b15zdnd11an1n16x5 FILLER_349_1450 ();
 b15zdnd00an1n02x5 FILLER_349_1466 ();
 b15zdnd11an1n08x5 FILLER_349_1489 ();
 b15zdnd00an1n02x5 FILLER_349_1497 ();
 b15zdnd11an1n08x5 FILLER_349_1511 ();
 b15zdnd11an1n04x5 FILLER_349_1519 ();
 b15zdnd00an1n02x5 FILLER_349_1523 ();
 b15zdnd11an1n16x5 FILLER_349_1534 ();
 b15zdnd11an1n16x5 FILLER_349_1556 ();
 b15zdnd00an1n02x5 FILLER_349_1572 ();
 b15zdnd00an1n01x5 FILLER_349_1574 ();
 b15zdnd11an1n16x5 FILLER_349_1584 ();
 b15zdnd11an1n08x5 FILLER_349_1600 ();
 b15zdnd11an1n04x5 FILLER_349_1608 ();
 b15zdnd00an1n02x5 FILLER_349_1612 ();
 b15zdnd00an1n01x5 FILLER_349_1614 ();
 b15zdnd11an1n32x5 FILLER_349_1625 ();
 b15zdnd11an1n04x5 FILLER_349_1657 ();
 b15zdnd00an1n02x5 FILLER_349_1661 ();
 b15zdnd11an1n16x5 FILLER_349_1679 ();
 b15zdnd11an1n04x5 FILLER_349_1719 ();
 b15zdnd11an1n64x5 FILLER_349_1733 ();
 b15zdnd11an1n32x5 FILLER_349_1797 ();
 b15zdnd11an1n04x5 FILLER_349_1829 ();
 b15zdnd00an1n02x5 FILLER_349_1833 ();
 b15zdnd11an1n32x5 FILLER_349_1845 ();
 b15zdnd11an1n16x5 FILLER_349_1877 ();
 b15zdnd11an1n04x5 FILLER_349_1907 ();
 b15zdnd11an1n16x5 FILLER_349_1918 ();
 b15zdnd00an1n02x5 FILLER_349_1934 ();
 b15zdnd00an1n01x5 FILLER_349_1936 ();
 b15zdnd11an1n08x5 FILLER_349_1945 ();
 b15zdnd11an1n04x5 FILLER_349_1953 ();
 b15zdnd00an1n02x5 FILLER_349_1957 ();
 b15zdnd00an1n01x5 FILLER_349_1959 ();
 b15zdnd11an1n04x5 FILLER_349_1966 ();
 b15zdnd00an1n02x5 FILLER_349_1970 ();
 b15zdnd11an1n04x5 FILLER_349_1983 ();
 b15zdnd11an1n16x5 FILLER_349_1994 ();
 b15zdnd11an1n04x5 FILLER_349_2010 ();
 b15zdnd00an1n02x5 FILLER_349_2014 ();
 b15zdnd00an1n01x5 FILLER_349_2016 ();
 b15zdnd11an1n64x5 FILLER_349_2022 ();
 b15zdnd11an1n32x5 FILLER_349_2086 ();
 b15zdnd11an1n08x5 FILLER_349_2118 ();
 b15zdnd00an1n02x5 FILLER_349_2126 ();
 b15zdnd11an1n32x5 FILLER_349_2134 ();
 b15zdnd11an1n04x5 FILLER_349_2166 ();
 b15zdnd00an1n02x5 FILLER_349_2170 ();
 b15zdnd11an1n08x5 FILLER_349_2178 ();
 b15zdnd11an1n04x5 FILLER_349_2186 ();
 b15zdnd00an1n02x5 FILLER_349_2190 ();
 b15zdnd11an1n04x5 FILLER_349_2197 ();
 b15zdnd00an1n01x5 FILLER_349_2201 ();
 b15zdnd11an1n64x5 FILLER_349_2207 ();
 b15zdnd11an1n08x5 FILLER_349_2271 ();
 b15zdnd11an1n04x5 FILLER_349_2279 ();
 b15zdnd00an1n01x5 FILLER_349_2283 ();
 b15zdnd11an1n64x5 FILLER_350_8 ();
 b15zdnd11an1n64x5 FILLER_350_72 ();
 b15zdnd11an1n64x5 FILLER_350_136 ();
 b15zdnd11an1n16x5 FILLER_350_200 ();
 b15zdnd00an1n01x5 FILLER_350_216 ();
 b15zdnd11an1n64x5 FILLER_350_224 ();
 b15zdnd11an1n16x5 FILLER_350_288 ();
 b15zdnd00an1n02x5 FILLER_350_304 ();
 b15zdnd11an1n08x5 FILLER_350_316 ();
 b15zdnd11an1n04x5 FILLER_350_324 ();
 b15zdnd11an1n32x5 FILLER_350_332 ();
 b15zdnd11an1n16x5 FILLER_350_364 ();
 b15zdnd11an1n08x5 FILLER_350_380 ();
 b15zdnd00an1n02x5 FILLER_350_388 ();
 b15zdnd11an1n04x5 FILLER_350_411 ();
 b15zdnd11an1n04x5 FILLER_350_421 ();
 b15zdnd11an1n64x5 FILLER_350_446 ();
 b15zdnd11an1n16x5 FILLER_350_510 ();
 b15zdnd11an1n08x5 FILLER_350_526 ();
 b15zdnd11an1n04x5 FILLER_350_534 ();
 b15zdnd00an1n02x5 FILLER_350_538 ();
 b15zdnd00an1n01x5 FILLER_350_540 ();
 b15zdnd11an1n64x5 FILLER_350_558 ();
 b15zdnd11an1n16x5 FILLER_350_622 ();
 b15zdnd11an1n08x5 FILLER_350_638 ();
 b15zdnd11an1n04x5 FILLER_350_646 ();
 b15zdnd11an1n16x5 FILLER_350_667 ();
 b15zdnd11an1n08x5 FILLER_350_683 ();
 b15zdnd11an1n04x5 FILLER_350_691 ();
 b15zdnd00an1n02x5 FILLER_350_695 ();
 b15zdnd00an1n01x5 FILLER_350_697 ();
 b15zdnd11an1n08x5 FILLER_350_709 ();
 b15zdnd00an1n01x5 FILLER_350_717 ();
 b15zdnd11an1n32x5 FILLER_350_726 ();
 b15zdnd11an1n32x5 FILLER_350_766 ();
 b15zdnd11an1n16x5 FILLER_350_798 ();
 b15zdnd11an1n08x5 FILLER_350_814 ();
 b15zdnd11an1n04x5 FILLER_350_822 ();
 b15zdnd11an1n08x5 FILLER_350_832 ();
 b15zdnd00an1n01x5 FILLER_350_840 ();
 b15zdnd11an1n16x5 FILLER_350_847 ();
 b15zdnd11an1n08x5 FILLER_350_863 ();
 b15zdnd00an1n02x5 FILLER_350_871 ();
 b15zdnd11an1n04x5 FILLER_350_878 ();
 b15zdnd11an1n32x5 FILLER_350_891 ();
 b15zdnd11an1n16x5 FILLER_350_923 ();
 b15zdnd11an1n04x5 FILLER_350_939 ();
 b15zdnd00an1n02x5 FILLER_350_943 ();
 b15zdnd11an1n16x5 FILLER_350_957 ();
 b15zdnd11an1n04x5 FILLER_350_973 ();
 b15zdnd11an1n16x5 FILLER_350_983 ();
 b15zdnd00an1n02x5 FILLER_350_999 ();
 b15zdnd00an1n01x5 FILLER_350_1001 ();
 b15zdnd11an1n08x5 FILLER_350_1014 ();
 b15zdnd11an1n04x5 FILLER_350_1029 ();
 b15zdnd11an1n04x5 FILLER_350_1039 ();
 b15zdnd00an1n02x5 FILLER_350_1043 ();
 b15zdnd11an1n04x5 FILLER_350_1054 ();
 b15zdnd11an1n04x5 FILLER_350_1070 ();
 b15zdnd11an1n64x5 FILLER_350_1082 ();
 b15zdnd11an1n16x5 FILLER_350_1146 ();
 b15zdnd11an1n08x5 FILLER_350_1162 ();
 b15zdnd11an1n64x5 FILLER_350_1191 ();
 b15zdnd11an1n16x5 FILLER_350_1255 ();
 b15zdnd11an1n08x5 FILLER_350_1271 ();
 b15zdnd11an1n04x5 FILLER_350_1279 ();
 b15zdnd00an1n01x5 FILLER_350_1283 ();
 b15zdnd11an1n08x5 FILLER_350_1303 ();
 b15zdnd11an1n04x5 FILLER_350_1311 ();
 b15zdnd00an1n02x5 FILLER_350_1315 ();
 b15zdnd00an1n01x5 FILLER_350_1317 ();
 b15zdnd11an1n32x5 FILLER_350_1331 ();
 b15zdnd11an1n08x5 FILLER_350_1363 ();
 b15zdnd11an1n04x5 FILLER_350_1371 ();
 b15zdnd00an1n02x5 FILLER_350_1375 ();
 b15zdnd11an1n04x5 FILLER_350_1388 ();
 b15zdnd11an1n64x5 FILLER_350_1396 ();
 b15zdnd11an1n16x5 FILLER_350_1460 ();
 b15zdnd11an1n08x5 FILLER_350_1488 ();
 b15zdnd11an1n04x5 FILLER_350_1496 ();
 b15zdnd00an1n02x5 FILLER_350_1500 ();
 b15zdnd11an1n08x5 FILLER_350_1509 ();
 b15zdnd11an1n04x5 FILLER_350_1517 ();
 b15zdnd00an1n02x5 FILLER_350_1521 ();
 b15zdnd00an1n01x5 FILLER_350_1523 ();
 b15zdnd11an1n64x5 FILLER_350_1536 ();
 b15zdnd11an1n04x5 FILLER_350_1600 ();
 b15zdnd00an1n01x5 FILLER_350_1604 ();
 b15zdnd11an1n16x5 FILLER_350_1625 ();
 b15zdnd11an1n08x5 FILLER_350_1641 ();
 b15zdnd11an1n04x5 FILLER_350_1649 ();
 b15zdnd00an1n02x5 FILLER_350_1653 ();
 b15zdnd00an1n01x5 FILLER_350_1655 ();
 b15zdnd11an1n16x5 FILLER_350_1677 ();
 b15zdnd11an1n04x5 FILLER_350_1693 ();
 b15zdnd00an1n02x5 FILLER_350_1697 ();
 b15zdnd11an1n64x5 FILLER_350_1712 ();
 b15zdnd11an1n64x5 FILLER_350_1776 ();
 b15zdnd11an1n04x5 FILLER_350_1840 ();
 b15zdnd00an1n01x5 FILLER_350_1844 ();
 b15zdnd11an1n16x5 FILLER_350_1859 ();
 b15zdnd11an1n32x5 FILLER_350_1882 ();
 b15zdnd11an1n08x5 FILLER_350_1919 ();
 b15zdnd00an1n01x5 FILLER_350_1927 ();
 b15zdnd11an1n08x5 FILLER_350_1940 ();
 b15zdnd00an1n01x5 FILLER_350_1948 ();
 b15zdnd11an1n64x5 FILLER_350_1969 ();
 b15zdnd11an1n64x5 FILLER_350_2033 ();
 b15zdnd11an1n32x5 FILLER_350_2097 ();
 b15zdnd11an1n08x5 FILLER_350_2129 ();
 b15zdnd00an1n01x5 FILLER_350_2137 ();
 b15zdnd00an1n02x5 FILLER_350_2152 ();
 b15zdnd11an1n32x5 FILLER_350_2162 ();
 b15zdnd11an1n08x5 FILLER_350_2194 ();
 b15zdnd00an1n02x5 FILLER_350_2202 ();
 b15zdnd00an1n01x5 FILLER_350_2204 ();
 b15zdnd11an1n32x5 FILLER_350_2218 ();
 b15zdnd11an1n16x5 FILLER_350_2250 ();
 b15zdnd11an1n08x5 FILLER_350_2266 ();
 b15zdnd00an1n02x5 FILLER_350_2274 ();
 b15zdnd11an1n64x5 FILLER_351_0 ();
 b15zdnd11an1n64x5 FILLER_351_64 ();
 b15zdnd11an1n64x5 FILLER_351_128 ();
 b15zdnd11an1n16x5 FILLER_351_192 ();
 b15zdnd11an1n08x5 FILLER_351_208 ();
 b15zdnd11an1n04x5 FILLER_351_216 ();
 b15zdnd00an1n02x5 FILLER_351_220 ();
 b15zdnd11an1n08x5 FILLER_351_229 ();
 b15zdnd11an1n04x5 FILLER_351_237 ();
 b15zdnd00an1n02x5 FILLER_351_241 ();
 b15zdnd11an1n16x5 FILLER_351_252 ();
 b15zdnd11an1n08x5 FILLER_351_268 ();
 b15zdnd11an1n04x5 FILLER_351_276 ();
 b15zdnd11an1n04x5 FILLER_351_284 ();
 b15zdnd11an1n16x5 FILLER_351_294 ();
 b15zdnd11an1n08x5 FILLER_351_310 ();
 b15zdnd00an1n02x5 FILLER_351_318 ();
 b15zdnd11an1n32x5 FILLER_351_328 ();
 b15zdnd00an1n02x5 FILLER_351_360 ();
 b15zdnd11an1n64x5 FILLER_351_382 ();
 b15zdnd11an1n04x5 FILLER_351_446 ();
 b15zdnd11an1n16x5 FILLER_351_456 ();
 b15zdnd11an1n16x5 FILLER_351_478 ();
 b15zdnd00an1n01x5 FILLER_351_494 ();
 b15zdnd11an1n04x5 FILLER_351_502 ();
 b15zdnd11an1n32x5 FILLER_351_519 ();
 b15zdnd11an1n08x5 FILLER_351_551 ();
 b15zdnd11an1n64x5 FILLER_351_570 ();
 b15zdnd11an1n16x5 FILLER_351_634 ();
 b15zdnd11an1n08x5 FILLER_351_650 ();
 b15zdnd11an1n04x5 FILLER_351_658 ();
 b15zdnd11an1n16x5 FILLER_351_674 ();
 b15zdnd11an1n08x5 FILLER_351_690 ();
 b15zdnd00an1n02x5 FILLER_351_698 ();
 b15zdnd11an1n32x5 FILLER_351_704 ();
 b15zdnd11an1n16x5 FILLER_351_736 ();
 b15zdnd11an1n08x5 FILLER_351_752 ();
 b15zdnd11an1n16x5 FILLER_351_771 ();
 b15zdnd11an1n08x5 FILLER_351_787 ();
 b15zdnd11an1n04x5 FILLER_351_795 ();
 b15zdnd00an1n01x5 FILLER_351_799 ();
 b15zdnd11an1n08x5 FILLER_351_810 ();
 b15zdnd00an1n02x5 FILLER_351_818 ();
 b15zdnd00an1n01x5 FILLER_351_820 ();
 b15zdnd11an1n64x5 FILLER_351_832 ();
 b15zdnd11an1n16x5 FILLER_351_896 ();
 b15zdnd11an1n32x5 FILLER_351_926 ();
 b15zdnd11an1n16x5 FILLER_351_958 ();
 b15zdnd00an1n02x5 FILLER_351_974 ();
 b15zdnd11an1n16x5 FILLER_351_982 ();
 b15zdnd00an1n02x5 FILLER_351_998 ();
 b15zdnd11an1n08x5 FILLER_351_1021 ();
 b15zdnd11an1n32x5 FILLER_351_1033 ();
 b15zdnd11an1n08x5 FILLER_351_1065 ();
 b15zdnd11an1n16x5 FILLER_351_1078 ();
 b15zdnd00an1n02x5 FILLER_351_1094 ();
 b15zdnd11an1n04x5 FILLER_351_1101 ();
 b15zdnd00an1n01x5 FILLER_351_1105 ();
 b15zdnd11an1n64x5 FILLER_351_1111 ();
 b15zdnd11an1n08x5 FILLER_351_1175 ();
 b15zdnd11an1n04x5 FILLER_351_1183 ();
 b15zdnd00an1n02x5 FILLER_351_1187 ();
 b15zdnd00an1n01x5 FILLER_351_1189 ();
 b15zdnd11an1n32x5 FILLER_351_1199 ();
 b15zdnd11an1n16x5 FILLER_351_1231 ();
 b15zdnd11an1n08x5 FILLER_351_1247 ();
 b15zdnd11an1n04x5 FILLER_351_1255 ();
 b15zdnd11an1n32x5 FILLER_351_1276 ();
 b15zdnd11an1n08x5 FILLER_351_1308 ();
 b15zdnd11an1n04x5 FILLER_351_1316 ();
 b15zdnd11an1n64x5 FILLER_351_1325 ();
 b15zdnd11an1n32x5 FILLER_351_1389 ();
 b15zdnd11an1n08x5 FILLER_351_1421 ();
 b15zdnd11an1n04x5 FILLER_351_1429 ();
 b15zdnd00an1n02x5 FILLER_351_1433 ();
 b15zdnd11an1n16x5 FILLER_351_1445 ();
 b15zdnd11an1n04x5 FILLER_351_1461 ();
 b15zdnd00an1n02x5 FILLER_351_1465 ();
 b15zdnd11an1n16x5 FILLER_351_1474 ();
 b15zdnd11an1n04x5 FILLER_351_1490 ();
 b15zdnd00an1n02x5 FILLER_351_1494 ();
 b15zdnd11an1n16x5 FILLER_351_1501 ();
 b15zdnd11an1n04x5 FILLER_351_1517 ();
 b15zdnd00an1n02x5 FILLER_351_1521 ();
 b15zdnd00an1n01x5 FILLER_351_1523 ();
 b15zdnd11an1n16x5 FILLER_351_1530 ();
 b15zdnd11an1n04x5 FILLER_351_1546 ();
 b15zdnd11an1n32x5 FILLER_351_1556 ();
 b15zdnd11an1n16x5 FILLER_351_1588 ();
 b15zdnd11an1n04x5 FILLER_351_1604 ();
 b15zdnd00an1n02x5 FILLER_351_1608 ();
 b15zdnd11an1n32x5 FILLER_351_1614 ();
 b15zdnd11an1n04x5 FILLER_351_1646 ();
 b15zdnd00an1n02x5 FILLER_351_1650 ();
 b15zdnd00an1n01x5 FILLER_351_1652 ();
 b15zdnd11an1n32x5 FILLER_351_1658 ();
 b15zdnd11an1n16x5 FILLER_351_1690 ();
 b15zdnd11an1n04x5 FILLER_351_1706 ();
 b15zdnd00an1n02x5 FILLER_351_1710 ();
 b15zdnd11an1n04x5 FILLER_351_1725 ();
 b15zdnd11an1n64x5 FILLER_351_1735 ();
 b15zdnd11an1n04x5 FILLER_351_1799 ();
 b15zdnd00an1n02x5 FILLER_351_1803 ();
 b15zdnd11an1n16x5 FILLER_351_1817 ();
 b15zdnd11an1n08x5 FILLER_351_1833 ();
 b15zdnd00an1n02x5 FILLER_351_1841 ();
 b15zdnd11an1n08x5 FILLER_351_1852 ();
 b15zdnd00an1n02x5 FILLER_351_1860 ();
 b15zdnd00an1n01x5 FILLER_351_1862 ();
 b15zdnd11an1n04x5 FILLER_351_1875 ();
 b15zdnd11an1n32x5 FILLER_351_1884 ();
 b15zdnd11an1n08x5 FILLER_351_1916 ();
 b15zdnd11an1n04x5 FILLER_351_1924 ();
 b15zdnd00an1n02x5 FILLER_351_1928 ();
 b15zdnd00an1n01x5 FILLER_351_1930 ();
 b15zdnd11an1n64x5 FILLER_351_1935 ();
 b15zdnd11an1n64x5 FILLER_351_1999 ();
 b15zdnd11an1n64x5 FILLER_351_2063 ();
 b15zdnd00an1n01x5 FILLER_351_2127 ();
 b15zdnd11an1n08x5 FILLER_351_2141 ();
 b15zdnd00an1n01x5 FILLER_351_2149 ();
 b15zdnd11an1n04x5 FILLER_351_2159 ();
 b15zdnd11an1n32x5 FILLER_351_2167 ();
 b15zdnd11an1n08x5 FILLER_351_2199 ();
 b15zdnd00an1n01x5 FILLER_351_2207 ();
 b15zdnd11an1n64x5 FILLER_351_2214 ();
 b15zdnd11an1n04x5 FILLER_351_2278 ();
 b15zdnd00an1n02x5 FILLER_351_2282 ();
 b15zdnd11an1n64x5 FILLER_352_8 ();
 b15zdnd11an1n64x5 FILLER_352_72 ();
 b15zdnd11an1n64x5 FILLER_352_136 ();
 b15zdnd11an1n16x5 FILLER_352_200 ();
 b15zdnd11an1n08x5 FILLER_352_216 ();
 b15zdnd11an1n04x5 FILLER_352_224 ();
 b15zdnd00an1n02x5 FILLER_352_228 ();
 b15zdnd00an1n01x5 FILLER_352_230 ();
 b15zdnd11an1n16x5 FILLER_352_244 ();
 b15zdnd11an1n04x5 FILLER_352_260 ();
 b15zdnd00an1n01x5 FILLER_352_264 ();
 b15zdnd11an1n08x5 FILLER_352_283 ();
 b15zdnd00an1n02x5 FILLER_352_291 ();
 b15zdnd00an1n01x5 FILLER_352_293 ();
 b15zdnd11an1n32x5 FILLER_352_300 ();
 b15zdnd11an1n16x5 FILLER_352_332 ();
 b15zdnd11an1n08x5 FILLER_352_348 ();
 b15zdnd11an1n04x5 FILLER_352_356 ();
 b15zdnd00an1n02x5 FILLER_352_360 ();
 b15zdnd00an1n01x5 FILLER_352_362 ();
 b15zdnd11an1n04x5 FILLER_352_375 ();
 b15zdnd00an1n01x5 FILLER_352_379 ();
 b15zdnd11an1n32x5 FILLER_352_395 ();
 b15zdnd11an1n16x5 FILLER_352_427 ();
 b15zdnd11an1n08x5 FILLER_352_443 ();
 b15zdnd11an1n32x5 FILLER_352_463 ();
 b15zdnd11an1n16x5 FILLER_352_495 ();
 b15zdnd00an1n02x5 FILLER_352_511 ();
 b15zdnd11an1n32x5 FILLER_352_517 ();
 b15zdnd11an1n04x5 FILLER_352_549 ();
 b15zdnd00an1n01x5 FILLER_352_553 ();
 b15zdnd11an1n64x5 FILLER_352_563 ();
 b15zdnd11an1n32x5 FILLER_352_627 ();
 b15zdnd00an1n02x5 FILLER_352_659 ();
 b15zdnd00an1n01x5 FILLER_352_661 ();
 b15zdnd11an1n32x5 FILLER_352_666 ();
 b15zdnd11an1n16x5 FILLER_352_698 ();
 b15zdnd11an1n04x5 FILLER_352_714 ();
 b15zdnd11an1n08x5 FILLER_352_726 ();
 b15zdnd00an1n02x5 FILLER_352_734 ();
 b15zdnd11an1n16x5 FILLER_352_741 ();
 b15zdnd11an1n08x5 FILLER_352_757 ();
 b15zdnd00an1n02x5 FILLER_352_765 ();
 b15zdnd00an1n01x5 FILLER_352_767 ();
 b15zdnd11an1n64x5 FILLER_352_784 ();
 b15zdnd11an1n32x5 FILLER_352_848 ();
 b15zdnd11an1n16x5 FILLER_352_880 ();
 b15zdnd11an1n08x5 FILLER_352_896 ();
 b15zdnd00an1n01x5 FILLER_352_904 ();
 b15zdnd11an1n16x5 FILLER_352_918 ();
 b15zdnd11an1n04x5 FILLER_352_934 ();
 b15zdnd11an1n16x5 FILLER_352_949 ();
 b15zdnd11an1n08x5 FILLER_352_965 ();
 b15zdnd00an1n02x5 FILLER_352_973 ();
 b15zdnd11an1n32x5 FILLER_352_984 ();
 b15zdnd11an1n16x5 FILLER_352_1016 ();
 b15zdnd11an1n04x5 FILLER_352_1032 ();
 b15zdnd00an1n02x5 FILLER_352_1036 ();
 b15zdnd11an1n32x5 FILLER_352_1042 ();
 b15zdnd11an1n04x5 FILLER_352_1074 ();
 b15zdnd11an1n08x5 FILLER_352_1083 ();
 b15zdnd11an1n04x5 FILLER_352_1091 ();
 b15zdnd00an1n02x5 FILLER_352_1095 ();
 b15zdnd00an1n01x5 FILLER_352_1097 ();
 b15zdnd11an1n16x5 FILLER_352_1103 ();
 b15zdnd00an1n02x5 FILLER_352_1119 ();
 b15zdnd11an1n64x5 FILLER_352_1129 ();
 b15zdnd11an1n64x5 FILLER_352_1193 ();
 b15zdnd11an1n64x5 FILLER_352_1257 ();
 b15zdnd11an1n32x5 FILLER_352_1321 ();
 b15zdnd11an1n16x5 FILLER_352_1353 ();
 b15zdnd00an1n02x5 FILLER_352_1369 ();
 b15zdnd11an1n16x5 FILLER_352_1385 ();
 b15zdnd11an1n04x5 FILLER_352_1401 ();
 b15zdnd00an1n01x5 FILLER_352_1405 ();
 b15zdnd11an1n08x5 FILLER_352_1416 ();
 b15zdnd00an1n01x5 FILLER_352_1424 ();
 b15zdnd11an1n08x5 FILLER_352_1444 ();
 b15zdnd00an1n02x5 FILLER_352_1452 ();
 b15zdnd11an1n08x5 FILLER_352_1475 ();
 b15zdnd11an1n04x5 FILLER_352_1483 ();
 b15zdnd00an1n02x5 FILLER_352_1487 ();
 b15zdnd00an1n01x5 FILLER_352_1489 ();
 b15zdnd11an1n32x5 FILLER_352_1504 ();
 b15zdnd11an1n08x5 FILLER_352_1536 ();
 b15zdnd11an1n04x5 FILLER_352_1544 ();
 b15zdnd00an1n02x5 FILLER_352_1548 ();
 b15zdnd11an1n32x5 FILLER_352_1554 ();
 b15zdnd11an1n04x5 FILLER_352_1586 ();
 b15zdnd11an1n08x5 FILLER_352_1594 ();
 b15zdnd00an1n02x5 FILLER_352_1602 ();
 b15zdnd00an1n01x5 FILLER_352_1604 ();
 b15zdnd11an1n32x5 FILLER_352_1617 ();
 b15zdnd11an1n04x5 FILLER_352_1649 ();
 b15zdnd00an1n01x5 FILLER_352_1653 ();
 b15zdnd11an1n16x5 FILLER_352_1660 ();
 b15zdnd00an1n02x5 FILLER_352_1676 ();
 b15zdnd00an1n01x5 FILLER_352_1678 ();
 b15zdnd11an1n16x5 FILLER_352_1684 ();
 b15zdnd11an1n08x5 FILLER_352_1700 ();
 b15zdnd11an1n04x5 FILLER_352_1708 ();
 b15zdnd00an1n01x5 FILLER_352_1712 ();
 b15zdnd11an1n64x5 FILLER_352_1716 ();
 b15zdnd11an1n16x5 FILLER_352_1780 ();
 b15zdnd11an1n04x5 FILLER_352_1796 ();
 b15zdnd00an1n02x5 FILLER_352_1800 ();
 b15zdnd11an1n16x5 FILLER_352_1807 ();
 b15zdnd00an1n02x5 FILLER_352_1823 ();
 b15zdnd11an1n04x5 FILLER_352_1840 ();
 b15zdnd00an1n02x5 FILLER_352_1844 ();
 b15zdnd00an1n01x5 FILLER_352_1846 ();
 b15zdnd11an1n16x5 FILLER_352_1853 ();
 b15zdnd11an1n04x5 FILLER_352_1869 ();
 b15zdnd00an1n02x5 FILLER_352_1873 ();
 b15zdnd00an1n01x5 FILLER_352_1875 ();
 b15zdnd11an1n32x5 FILLER_352_1881 ();
 b15zdnd11an1n08x5 FILLER_352_1913 ();
 b15zdnd11an1n04x5 FILLER_352_1921 ();
 b15zdnd00an1n01x5 FILLER_352_1925 ();
 b15zdnd11an1n64x5 FILLER_352_1931 ();
 b15zdnd11an1n16x5 FILLER_352_1995 ();
 b15zdnd11an1n08x5 FILLER_352_2011 ();
 b15zdnd11an1n04x5 FILLER_352_2019 ();
 b15zdnd11an1n32x5 FILLER_352_2030 ();
 b15zdnd11an1n16x5 FILLER_352_2062 ();
 b15zdnd11an1n08x5 FILLER_352_2078 ();
 b15zdnd11an1n16x5 FILLER_352_2092 ();
 b15zdnd11an1n08x5 FILLER_352_2113 ();
 b15zdnd11an1n04x5 FILLER_352_2121 ();
 b15zdnd11an1n04x5 FILLER_352_2132 ();
 b15zdnd11an1n04x5 FILLER_352_2148 ();
 b15zdnd00an1n02x5 FILLER_352_2152 ();
 b15zdnd11an1n16x5 FILLER_352_2162 ();
 b15zdnd11an1n08x5 FILLER_352_2178 ();
 b15zdnd11an1n04x5 FILLER_352_2186 ();
 b15zdnd00an1n02x5 FILLER_352_2190 ();
 b15zdnd11an1n64x5 FILLER_352_2198 ();
 b15zdnd11an1n08x5 FILLER_352_2262 ();
 b15zdnd11an1n04x5 FILLER_352_2270 ();
 b15zdnd00an1n02x5 FILLER_352_2274 ();
 b15zdnd11an1n64x5 FILLER_353_0 ();
 b15zdnd11an1n64x5 FILLER_353_64 ();
 b15zdnd11an1n64x5 FILLER_353_128 ();
 b15zdnd11an1n64x5 FILLER_353_192 ();
 b15zdnd11an1n08x5 FILLER_353_256 ();
 b15zdnd11an1n04x5 FILLER_353_264 ();
 b15zdnd00an1n02x5 FILLER_353_268 ();
 b15zdnd11an1n08x5 FILLER_353_284 ();
 b15zdnd00an1n02x5 FILLER_353_292 ();
 b15zdnd11an1n16x5 FILLER_353_303 ();
 b15zdnd11an1n08x5 FILLER_353_319 ();
 b15zdnd11an1n16x5 FILLER_353_334 ();
 b15zdnd11an1n08x5 FILLER_353_350 ();
 b15zdnd11an1n04x5 FILLER_353_358 ();
 b15zdnd11an1n64x5 FILLER_353_366 ();
 b15zdnd00an1n01x5 FILLER_353_430 ();
 b15zdnd11an1n64x5 FILLER_353_439 ();
 b15zdnd11an1n64x5 FILLER_353_503 ();
 b15zdnd11an1n16x5 FILLER_353_567 ();
 b15zdnd00an1n02x5 FILLER_353_583 ();
 b15zdnd11an1n64x5 FILLER_353_591 ();
 b15zdnd11an1n32x5 FILLER_353_655 ();
 b15zdnd11an1n08x5 FILLER_353_687 ();
 b15zdnd11an1n04x5 FILLER_353_695 ();
 b15zdnd00an1n02x5 FILLER_353_699 ();
 b15zdnd11an1n32x5 FILLER_353_706 ();
 b15zdnd11an1n16x5 FILLER_353_738 ();
 b15zdnd11an1n08x5 FILLER_353_754 ();
 b15zdnd11an1n04x5 FILLER_353_774 ();
 b15zdnd00an1n02x5 FILLER_353_778 ();
 b15zdnd00an1n01x5 FILLER_353_780 ();
 b15zdnd11an1n64x5 FILLER_353_792 ();
 b15zdnd11an1n04x5 FILLER_353_856 ();
 b15zdnd11an1n32x5 FILLER_353_864 ();
 b15zdnd11an1n08x5 FILLER_353_896 ();
 b15zdnd11an1n04x5 FILLER_353_904 ();
 b15zdnd00an1n02x5 FILLER_353_908 ();
 b15zdnd00an1n01x5 FILLER_353_910 ();
 b15zdnd11an1n08x5 FILLER_353_932 ();
 b15zdnd11an1n04x5 FILLER_353_940 ();
 b15zdnd00an1n01x5 FILLER_353_944 ();
 b15zdnd11an1n08x5 FILLER_353_957 ();
 b15zdnd11an1n04x5 FILLER_353_965 ();
 b15zdnd00an1n02x5 FILLER_353_969 ();
 b15zdnd00an1n01x5 FILLER_353_971 ();
 b15zdnd11an1n08x5 FILLER_353_992 ();
 b15zdnd00an1n02x5 FILLER_353_1000 ();
 b15zdnd11an1n32x5 FILLER_353_1014 ();
 b15zdnd11an1n16x5 FILLER_353_1046 ();
 b15zdnd11an1n08x5 FILLER_353_1062 ();
 b15zdnd00an1n02x5 FILLER_353_1070 ();
 b15zdnd00an1n01x5 FILLER_353_1072 ();
 b15zdnd11an1n04x5 FILLER_353_1079 ();
 b15zdnd11an1n08x5 FILLER_353_1096 ();
 b15zdnd11an1n32x5 FILLER_353_1111 ();
 b15zdnd11an1n04x5 FILLER_353_1143 ();
 b15zdnd00an1n02x5 FILLER_353_1147 ();
 b15zdnd11an1n64x5 FILLER_353_1161 ();
 b15zdnd11an1n32x5 FILLER_353_1225 ();
 b15zdnd00an1n02x5 FILLER_353_1257 ();
 b15zdnd00an1n01x5 FILLER_353_1259 ();
 b15zdnd11an1n16x5 FILLER_353_1265 ();
 b15zdnd00an1n01x5 FILLER_353_1281 ();
 b15zdnd11an1n16x5 FILLER_353_1294 ();
 b15zdnd11an1n04x5 FILLER_353_1310 ();
 b15zdnd00an1n02x5 FILLER_353_1314 ();
 b15zdnd00an1n01x5 FILLER_353_1316 ();
 b15zdnd11an1n32x5 FILLER_353_1322 ();
 b15zdnd11an1n04x5 FILLER_353_1354 ();
 b15zdnd00an1n01x5 FILLER_353_1358 ();
 b15zdnd11an1n04x5 FILLER_353_1367 ();
 b15zdnd11an1n32x5 FILLER_353_1377 ();
 b15zdnd11an1n64x5 FILLER_353_1420 ();
 b15zdnd11an1n64x5 FILLER_353_1484 ();
 b15zdnd11an1n08x5 FILLER_353_1548 ();
 b15zdnd11an1n04x5 FILLER_353_1556 ();
 b15zdnd11an1n04x5 FILLER_353_1572 ();
 b15zdnd11an1n32x5 FILLER_353_1581 ();
 b15zdnd11an1n16x5 FILLER_353_1613 ();
 b15zdnd11an1n08x5 FILLER_353_1629 ();
 b15zdnd11an1n32x5 FILLER_353_1641 ();
 b15zdnd00an1n02x5 FILLER_353_1673 ();
 b15zdnd00an1n01x5 FILLER_353_1675 ();
 b15zdnd11an1n64x5 FILLER_353_1688 ();
 b15zdnd11an1n64x5 FILLER_353_1752 ();
 b15zdnd11an1n64x5 FILLER_353_1816 ();
 b15zdnd11an1n32x5 FILLER_353_1880 ();
 b15zdnd11an1n16x5 FILLER_353_1912 ();
 b15zdnd00an1n02x5 FILLER_353_1928 ();
 b15zdnd00an1n01x5 FILLER_353_1930 ();
 b15zdnd11an1n16x5 FILLER_353_1938 ();
 b15zdnd00an1n02x5 FILLER_353_1954 ();
 b15zdnd11an1n32x5 FILLER_353_1972 ();
 b15zdnd11an1n08x5 FILLER_353_2004 ();
 b15zdnd00an1n01x5 FILLER_353_2012 ();
 b15zdnd11an1n04x5 FILLER_353_2018 ();
 b15zdnd11an1n16x5 FILLER_353_2028 ();
 b15zdnd00an1n02x5 FILLER_353_2044 ();
 b15zdnd00an1n01x5 FILLER_353_2046 ();
 b15zdnd11an1n16x5 FILLER_353_2052 ();
 b15zdnd11an1n08x5 FILLER_353_2068 ();
 b15zdnd00an1n01x5 FILLER_353_2076 ();
 b15zdnd11an1n04x5 FILLER_353_2082 ();
 b15zdnd11an1n08x5 FILLER_353_2093 ();
 b15zdnd00an1n02x5 FILLER_353_2101 ();
 b15zdnd00an1n01x5 FILLER_353_2103 ();
 b15zdnd11an1n64x5 FILLER_353_2117 ();
 b15zdnd11an1n64x5 FILLER_353_2181 ();
 b15zdnd11an1n32x5 FILLER_353_2245 ();
 b15zdnd11an1n04x5 FILLER_353_2277 ();
 b15zdnd00an1n02x5 FILLER_353_2281 ();
 b15zdnd00an1n01x5 FILLER_353_2283 ();
 b15zdnd11an1n64x5 FILLER_354_8 ();
 b15zdnd11an1n64x5 FILLER_354_72 ();
 b15zdnd11an1n64x5 FILLER_354_136 ();
 b15zdnd11an1n32x5 FILLER_354_200 ();
 b15zdnd00an1n02x5 FILLER_354_232 ();
 b15zdnd00an1n01x5 FILLER_354_234 ();
 b15zdnd11an1n16x5 FILLER_354_245 ();
 b15zdnd11an1n08x5 FILLER_354_261 ();
 b15zdnd00an1n02x5 FILLER_354_269 ();
 b15zdnd11an1n16x5 FILLER_354_278 ();
 b15zdnd00an1n01x5 FILLER_354_294 ();
 b15zdnd11an1n16x5 FILLER_354_299 ();
 b15zdnd11an1n08x5 FILLER_354_315 ();
 b15zdnd11an1n04x5 FILLER_354_323 ();
 b15zdnd11an1n32x5 FILLER_354_336 ();
 b15zdnd11an1n16x5 FILLER_354_368 ();
 b15zdnd11an1n08x5 FILLER_354_384 ();
 b15zdnd11an1n04x5 FILLER_354_392 ();
 b15zdnd00an1n02x5 FILLER_354_396 ();
 b15zdnd00an1n01x5 FILLER_354_398 ();
 b15zdnd11an1n04x5 FILLER_354_406 ();
 b15zdnd11an1n32x5 FILLER_354_414 ();
 b15zdnd11an1n16x5 FILLER_354_446 ();
 b15zdnd11an1n04x5 FILLER_354_462 ();
 b15zdnd00an1n01x5 FILLER_354_466 ();
 b15zdnd11an1n16x5 FILLER_354_476 ();
 b15zdnd11an1n08x5 FILLER_354_497 ();
 b15zdnd00an1n02x5 FILLER_354_505 ();
 b15zdnd11an1n08x5 FILLER_354_513 ();
 b15zdnd11an1n64x5 FILLER_354_526 ();
 b15zdnd11an1n32x5 FILLER_354_590 ();
 b15zdnd11an1n16x5 FILLER_354_622 ();
 b15zdnd11an1n04x5 FILLER_354_638 ();
 b15zdnd00an1n02x5 FILLER_354_642 ();
 b15zdnd11an1n08x5 FILLER_354_656 ();
 b15zdnd00an1n01x5 FILLER_354_664 ();
 b15zdnd11an1n16x5 FILLER_354_671 ();
 b15zdnd11an1n08x5 FILLER_354_687 ();
 b15zdnd11an1n04x5 FILLER_354_695 ();
 b15zdnd11an1n08x5 FILLER_354_704 ();
 b15zdnd11an1n04x5 FILLER_354_712 ();
 b15zdnd00an1n02x5 FILLER_354_716 ();
 b15zdnd11an1n08x5 FILLER_354_726 ();
 b15zdnd00an1n02x5 FILLER_354_734 ();
 b15zdnd11an1n32x5 FILLER_354_742 ();
 b15zdnd11an1n16x5 FILLER_354_774 ();
 b15zdnd11an1n08x5 FILLER_354_790 ();
 b15zdnd11an1n04x5 FILLER_354_798 ();
 b15zdnd00an1n02x5 FILLER_354_802 ();
 b15zdnd00an1n01x5 FILLER_354_804 ();
 b15zdnd11an1n32x5 FILLER_354_825 ();
 b15zdnd11an1n04x5 FILLER_354_866 ();
 b15zdnd11an1n32x5 FILLER_354_883 ();
 b15zdnd11an1n04x5 FILLER_354_915 ();
 b15zdnd11an1n64x5 FILLER_354_928 ();
 b15zdnd11an1n16x5 FILLER_354_992 ();
 b15zdnd11an1n08x5 FILLER_354_1008 ();
 b15zdnd11an1n04x5 FILLER_354_1016 ();
 b15zdnd11an1n04x5 FILLER_354_1025 ();
 b15zdnd11an1n64x5 FILLER_354_1035 ();
 b15zdnd11an1n32x5 FILLER_354_1099 ();
 b15zdnd00an1n02x5 FILLER_354_1131 ();
 b15zdnd11an1n16x5 FILLER_354_1143 ();
 b15zdnd11an1n08x5 FILLER_354_1159 ();
 b15zdnd11an1n04x5 FILLER_354_1173 ();
 b15zdnd11an1n64x5 FILLER_354_1181 ();
 b15zdnd11an1n08x5 FILLER_354_1245 ();
 b15zdnd11an1n04x5 FILLER_354_1253 ();
 b15zdnd00an1n02x5 FILLER_354_1257 ();
 b15zdnd00an1n01x5 FILLER_354_1259 ();
 b15zdnd11an1n04x5 FILLER_354_1270 ();
 b15zdnd00an1n02x5 FILLER_354_1274 ();
 b15zdnd00an1n01x5 FILLER_354_1276 ();
 b15zdnd11an1n04x5 FILLER_354_1283 ();
 b15zdnd11an1n08x5 FILLER_354_1291 ();
 b15zdnd11an1n08x5 FILLER_354_1304 ();
 b15zdnd00an1n02x5 FILLER_354_1312 ();
 b15zdnd11an1n08x5 FILLER_354_1326 ();
 b15zdnd11an1n04x5 FILLER_354_1334 ();
 b15zdnd00an1n02x5 FILLER_354_1338 ();
 b15zdnd00an1n01x5 FILLER_354_1340 ();
 b15zdnd11an1n16x5 FILLER_354_1347 ();
 b15zdnd11an1n04x5 FILLER_354_1363 ();
 b15zdnd00an1n02x5 FILLER_354_1367 ();
 b15zdnd11an1n04x5 FILLER_354_1374 ();
 b15zdnd11an1n32x5 FILLER_354_1384 ();
 b15zdnd11an1n16x5 FILLER_354_1416 ();
 b15zdnd00an1n02x5 FILLER_354_1432 ();
 b15zdnd11an1n16x5 FILLER_354_1444 ();
 b15zdnd11an1n04x5 FILLER_354_1460 ();
 b15zdnd00an1n01x5 FILLER_354_1464 ();
 b15zdnd11an1n32x5 FILLER_354_1475 ();
 b15zdnd11an1n04x5 FILLER_354_1507 ();
 b15zdnd11an1n32x5 FILLER_354_1523 ();
 b15zdnd11an1n16x5 FILLER_354_1555 ();
 b15zdnd11an1n04x5 FILLER_354_1571 ();
 b15zdnd11an1n16x5 FILLER_354_1584 ();
 b15zdnd11an1n04x5 FILLER_354_1600 ();
 b15zdnd00an1n02x5 FILLER_354_1604 ();
 b15zdnd11an1n04x5 FILLER_354_1616 ();
 b15zdnd11an1n32x5 FILLER_354_1625 ();
 b15zdnd11an1n16x5 FILLER_354_1657 ();
 b15zdnd11an1n08x5 FILLER_354_1673 ();
 b15zdnd11an1n16x5 FILLER_354_1693 ();
 b15zdnd00an1n02x5 FILLER_354_1709 ();
 b15zdnd00an1n01x5 FILLER_354_1711 ();
 b15zdnd11an1n16x5 FILLER_354_1722 ();
 b15zdnd11an1n04x5 FILLER_354_1738 ();
 b15zdnd00an1n01x5 FILLER_354_1742 ();
 b15zdnd11an1n08x5 FILLER_354_1748 ();
 b15zdnd00an1n02x5 FILLER_354_1756 ();
 b15zdnd11an1n32x5 FILLER_354_1762 ();
 b15zdnd11an1n16x5 FILLER_354_1794 ();
 b15zdnd11an1n04x5 FILLER_354_1810 ();
 b15zdnd00an1n02x5 FILLER_354_1814 ();
 b15zdnd11an1n04x5 FILLER_354_1836 ();
 b15zdnd11an1n04x5 FILLER_354_1848 ();
 b15zdnd00an1n02x5 FILLER_354_1852 ();
 b15zdnd11an1n16x5 FILLER_354_1860 ();
 b15zdnd11an1n08x5 FILLER_354_1876 ();
 b15zdnd11an1n04x5 FILLER_354_1884 ();
 b15zdnd00an1n02x5 FILLER_354_1888 ();
 b15zdnd00an1n01x5 FILLER_354_1890 ();
 b15zdnd11an1n04x5 FILLER_354_1900 ();
 b15zdnd00an1n02x5 FILLER_354_1904 ();
 b15zdnd00an1n01x5 FILLER_354_1906 ();
 b15zdnd11an1n32x5 FILLER_354_1919 ();
 b15zdnd11an1n16x5 FILLER_354_1951 ();
 b15zdnd11an1n04x5 FILLER_354_1967 ();
 b15zdnd00an1n01x5 FILLER_354_1971 ();
 b15zdnd11an1n08x5 FILLER_354_1984 ();
 b15zdnd11an1n04x5 FILLER_354_1992 ();
 b15zdnd00an1n02x5 FILLER_354_1996 ();
 b15zdnd11an1n04x5 FILLER_354_2010 ();
 b15zdnd00an1n01x5 FILLER_354_2014 ();
 b15zdnd11an1n08x5 FILLER_354_2036 ();
 b15zdnd00an1n01x5 FILLER_354_2044 ();
 b15zdnd11an1n04x5 FILLER_354_2055 ();
 b15zdnd11an1n08x5 FILLER_354_2065 ();
 b15zdnd11an1n04x5 FILLER_354_2073 ();
 b15zdnd00an1n02x5 FILLER_354_2077 ();
 b15zdnd00an1n01x5 FILLER_354_2079 ();
 b15zdnd11an1n16x5 FILLER_354_2092 ();
 b15zdnd11an1n16x5 FILLER_354_2128 ();
 b15zdnd11an1n08x5 FILLER_354_2144 ();
 b15zdnd00an1n02x5 FILLER_354_2152 ();
 b15zdnd11an1n16x5 FILLER_354_2162 ();
 b15zdnd11an1n08x5 FILLER_354_2178 ();
 b15zdnd00an1n02x5 FILLER_354_2186 ();
 b15zdnd00an1n01x5 FILLER_354_2188 ();
 b15zdnd11an1n04x5 FILLER_354_2195 ();
 b15zdnd11an1n64x5 FILLER_354_2203 ();
 b15zdnd11an1n08x5 FILLER_354_2267 ();
 b15zdnd00an1n01x5 FILLER_354_2275 ();
 b15zdnd11an1n64x5 FILLER_355_0 ();
 b15zdnd11an1n64x5 FILLER_355_64 ();
 b15zdnd11an1n64x5 FILLER_355_128 ();
 b15zdnd11an1n64x5 FILLER_355_192 ();
 b15zdnd11an1n04x5 FILLER_355_256 ();
 b15zdnd00an1n01x5 FILLER_355_260 ();
 b15zdnd11an1n16x5 FILLER_355_273 ();
 b15zdnd11an1n08x5 FILLER_355_289 ();
 b15zdnd11an1n04x5 FILLER_355_297 ();
 b15zdnd11an1n16x5 FILLER_355_315 ();
 b15zdnd11an1n08x5 FILLER_355_331 ();
 b15zdnd00an1n01x5 FILLER_355_339 ();
 b15zdnd11an1n08x5 FILLER_355_361 ();
 b15zdnd11an1n04x5 FILLER_355_369 ();
 b15zdnd00an1n02x5 FILLER_355_373 ();
 b15zdnd00an1n01x5 FILLER_355_375 ();
 b15zdnd11an1n08x5 FILLER_355_381 ();
 b15zdnd11an1n04x5 FILLER_355_389 ();
 b15zdnd00an1n02x5 FILLER_355_393 ();
 b15zdnd00an1n01x5 FILLER_355_395 ();
 b15zdnd11an1n16x5 FILLER_355_405 ();
 b15zdnd11an1n04x5 FILLER_355_421 ();
 b15zdnd11an1n64x5 FILLER_355_440 ();
 b15zdnd11an1n16x5 FILLER_355_504 ();
 b15zdnd00an1n01x5 FILLER_355_520 ();
 b15zdnd11an1n16x5 FILLER_355_531 ();
 b15zdnd11an1n08x5 FILLER_355_547 ();
 b15zdnd11an1n04x5 FILLER_355_560 ();
 b15zdnd11an1n32x5 FILLER_355_588 ();
 b15zdnd11an1n16x5 FILLER_355_620 ();
 b15zdnd11an1n08x5 FILLER_355_636 ();
 b15zdnd00an1n01x5 FILLER_355_644 ();
 b15zdnd11an1n08x5 FILLER_355_650 ();
 b15zdnd00an1n01x5 FILLER_355_658 ();
 b15zdnd11an1n16x5 FILLER_355_671 ();
 b15zdnd00an1n02x5 FILLER_355_687 ();
 b15zdnd00an1n01x5 FILLER_355_689 ();
 b15zdnd11an1n16x5 FILLER_355_708 ();
 b15zdnd11an1n04x5 FILLER_355_724 ();
 b15zdnd11an1n04x5 FILLER_355_734 ();
 b15zdnd11an1n64x5 FILLER_355_745 ();
 b15zdnd11an1n32x5 FILLER_355_809 ();
 b15zdnd11an1n16x5 FILLER_355_841 ();
 b15zdnd11an1n08x5 FILLER_355_857 ();
 b15zdnd00an1n02x5 FILLER_355_865 ();
 b15zdnd11an1n04x5 FILLER_355_881 ();
 b15zdnd11an1n64x5 FILLER_355_890 ();
 b15zdnd11an1n08x5 FILLER_355_954 ();
 b15zdnd00an1n02x5 FILLER_355_962 ();
 b15zdnd00an1n01x5 FILLER_355_964 ();
 b15zdnd11an1n64x5 FILLER_355_975 ();
 b15zdnd11an1n16x5 FILLER_355_1039 ();
 b15zdnd11an1n04x5 FILLER_355_1055 ();
 b15zdnd00an1n02x5 FILLER_355_1059 ();
 b15zdnd11an1n08x5 FILLER_355_1071 ();
 b15zdnd11an1n04x5 FILLER_355_1079 ();
 b15zdnd00an1n02x5 FILLER_355_1083 ();
 b15zdnd00an1n01x5 FILLER_355_1085 ();
 b15zdnd11an1n32x5 FILLER_355_1092 ();
 b15zdnd11an1n08x5 FILLER_355_1124 ();
 b15zdnd11an1n32x5 FILLER_355_1138 ();
 b15zdnd00an1n01x5 FILLER_355_1170 ();
 b15zdnd11an1n04x5 FILLER_355_1185 ();
 b15zdnd00an1n02x5 FILLER_355_1189 ();
 b15zdnd00an1n01x5 FILLER_355_1191 ();
 b15zdnd11an1n32x5 FILLER_355_1204 ();
 b15zdnd11an1n16x5 FILLER_355_1236 ();
 b15zdnd00an1n02x5 FILLER_355_1252 ();
 b15zdnd11an1n64x5 FILLER_355_1265 ();
 b15zdnd11an1n08x5 FILLER_355_1329 ();
 b15zdnd11an1n04x5 FILLER_355_1343 ();
 b15zdnd11an1n04x5 FILLER_355_1365 ();
 b15zdnd11an1n32x5 FILLER_355_1381 ();
 b15zdnd11an1n64x5 FILLER_355_1418 ();
 b15zdnd11an1n32x5 FILLER_355_1482 ();
 b15zdnd11an1n04x5 FILLER_355_1514 ();
 b15zdnd00an1n02x5 FILLER_355_1518 ();
 b15zdnd11an1n16x5 FILLER_355_1527 ();
 b15zdnd11an1n04x5 FILLER_355_1543 ();
 b15zdnd11an1n32x5 FILLER_355_1552 ();
 b15zdnd00an1n01x5 FILLER_355_1584 ();
 b15zdnd11an1n16x5 FILLER_355_1590 ();
 b15zdnd11an1n08x5 FILLER_355_1606 ();
 b15zdnd11an1n04x5 FILLER_355_1614 ();
 b15zdnd00an1n02x5 FILLER_355_1618 ();
 b15zdnd00an1n01x5 FILLER_355_1620 ();
 b15zdnd11an1n32x5 FILLER_355_1627 ();
 b15zdnd11an1n16x5 FILLER_355_1659 ();
 b15zdnd11an1n04x5 FILLER_355_1675 ();
 b15zdnd00an1n02x5 FILLER_355_1679 ();
 b15zdnd00an1n01x5 FILLER_355_1681 ();
 b15zdnd11an1n04x5 FILLER_355_1698 ();
 b15zdnd11an1n08x5 FILLER_355_1716 ();
 b15zdnd00an1n01x5 FILLER_355_1724 ();
 b15zdnd11an1n16x5 FILLER_355_1732 ();
 b15zdnd00an1n02x5 FILLER_355_1748 ();
 b15zdnd00an1n01x5 FILLER_355_1750 ();
 b15zdnd11an1n04x5 FILLER_355_1755 ();
 b15zdnd11an1n64x5 FILLER_355_1767 ();
 b15zdnd11an1n04x5 FILLER_355_1831 ();
 b15zdnd00an1n01x5 FILLER_355_1835 ();
 b15zdnd11an1n32x5 FILLER_355_1841 ();
 b15zdnd11an1n16x5 FILLER_355_1873 ();
 b15zdnd11an1n08x5 FILLER_355_1889 ();
 b15zdnd00an1n02x5 FILLER_355_1897 ();
 b15zdnd11an1n04x5 FILLER_355_1903 ();
 b15zdnd00an1n02x5 FILLER_355_1907 ();
 b15zdnd00an1n01x5 FILLER_355_1909 ();
 b15zdnd11an1n16x5 FILLER_355_1915 ();
 b15zdnd11an1n04x5 FILLER_355_1931 ();
 b15zdnd00an1n01x5 FILLER_355_1935 ();
 b15zdnd11an1n16x5 FILLER_355_1944 ();
 b15zdnd11an1n08x5 FILLER_355_1960 ();
 b15zdnd00an1n02x5 FILLER_355_1968 ();
 b15zdnd11an1n16x5 FILLER_355_1975 ();
 b15zdnd11an1n08x5 FILLER_355_1991 ();
 b15zdnd11an1n04x5 FILLER_355_1999 ();
 b15zdnd00an1n02x5 FILLER_355_2003 ();
 b15zdnd00an1n01x5 FILLER_355_2005 ();
 b15zdnd11an1n64x5 FILLER_355_2013 ();
 b15zdnd11an1n64x5 FILLER_355_2077 ();
 b15zdnd11an1n32x5 FILLER_355_2141 ();
 b15zdnd00an1n02x5 FILLER_355_2173 ();
 b15zdnd11an1n08x5 FILLER_355_2182 ();
 b15zdnd11an1n08x5 FILLER_355_2202 ();
 b15zdnd00an1n01x5 FILLER_355_2210 ();
 b15zdnd11an1n32x5 FILLER_355_2229 ();
 b15zdnd11an1n16x5 FILLER_355_2261 ();
 b15zdnd11an1n04x5 FILLER_355_2277 ();
 b15zdnd00an1n02x5 FILLER_355_2281 ();
 b15zdnd00an1n01x5 FILLER_355_2283 ();
 b15zdnd11an1n64x5 FILLER_356_8 ();
 b15zdnd11an1n64x5 FILLER_356_72 ();
 b15zdnd11an1n64x5 FILLER_356_136 ();
 b15zdnd11an1n16x5 FILLER_356_200 ();
 b15zdnd11an1n08x5 FILLER_356_216 ();
 b15zdnd11an1n04x5 FILLER_356_231 ();
 b15zdnd11an1n08x5 FILLER_356_242 ();
 b15zdnd11an1n04x5 FILLER_356_250 ();
 b15zdnd00an1n01x5 FILLER_356_254 ();
 b15zdnd11an1n04x5 FILLER_356_271 ();
 b15zdnd00an1n02x5 FILLER_356_275 ();
 b15zdnd00an1n01x5 FILLER_356_277 ();
 b15zdnd11an1n16x5 FILLER_356_301 ();
 b15zdnd11an1n04x5 FILLER_356_317 ();
 b15zdnd00an1n01x5 FILLER_356_321 ();
 b15zdnd11an1n32x5 FILLER_356_331 ();
 b15zdnd11an1n04x5 FILLER_356_363 ();
 b15zdnd11an1n32x5 FILLER_356_379 ();
 b15zdnd11an1n16x5 FILLER_356_411 ();
 b15zdnd11an1n04x5 FILLER_356_427 ();
 b15zdnd00an1n02x5 FILLER_356_431 ();
 b15zdnd00an1n01x5 FILLER_356_433 ();
 b15zdnd11an1n16x5 FILLER_356_439 ();
 b15zdnd11an1n04x5 FILLER_356_455 ();
 b15zdnd00an1n01x5 FILLER_356_459 ();
 b15zdnd11an1n04x5 FILLER_356_466 ();
 b15zdnd11an1n16x5 FILLER_356_482 ();
 b15zdnd00an1n02x5 FILLER_356_498 ();
 b15zdnd11an1n04x5 FILLER_356_510 ();
 b15zdnd00an1n02x5 FILLER_356_514 ();
 b15zdnd00an1n01x5 FILLER_356_516 ();
 b15zdnd11an1n16x5 FILLER_356_523 ();
 b15zdnd11an1n08x5 FILLER_356_539 ();
 b15zdnd00an1n02x5 FILLER_356_547 ();
 b15zdnd11an1n04x5 FILLER_356_559 ();
 b15zdnd00an1n01x5 FILLER_356_563 ();
 b15zdnd11an1n64x5 FILLER_356_569 ();
 b15zdnd11an1n08x5 FILLER_356_633 ();
 b15zdnd11an1n04x5 FILLER_356_641 ();
 b15zdnd11an1n32x5 FILLER_356_650 ();
 b15zdnd11an1n16x5 FILLER_356_682 ();
 b15zdnd00an1n02x5 FILLER_356_698 ();
 b15zdnd00an1n01x5 FILLER_356_700 ();
 b15zdnd11an1n08x5 FILLER_356_707 ();
 b15zdnd00an1n02x5 FILLER_356_715 ();
 b15zdnd00an1n01x5 FILLER_356_717 ();
 b15zdnd11an1n04x5 FILLER_356_726 ();
 b15zdnd00an1n01x5 FILLER_356_730 ();
 b15zdnd11an1n32x5 FILLER_356_735 ();
 b15zdnd11an1n16x5 FILLER_356_767 ();
 b15zdnd11an1n04x5 FILLER_356_783 ();
 b15zdnd00an1n02x5 FILLER_356_787 ();
 b15zdnd00an1n01x5 FILLER_356_789 ();
 b15zdnd11an1n16x5 FILLER_356_800 ();
 b15zdnd11an1n08x5 FILLER_356_816 ();
 b15zdnd00an1n02x5 FILLER_356_824 ();
 b15zdnd00an1n01x5 FILLER_356_826 ();
 b15zdnd11an1n04x5 FILLER_356_841 ();
 b15zdnd11an1n08x5 FILLER_356_871 ();
 b15zdnd00an1n01x5 FILLER_356_879 ();
 b15zdnd11an1n32x5 FILLER_356_888 ();
 b15zdnd11an1n08x5 FILLER_356_920 ();
 b15zdnd00an1n02x5 FILLER_356_928 ();
 b15zdnd11an1n04x5 FILLER_356_944 ();
 b15zdnd00an1n01x5 FILLER_356_948 ();
 b15zdnd11an1n32x5 FILLER_356_960 ();
 b15zdnd11an1n16x5 FILLER_356_992 ();
 b15zdnd11an1n32x5 FILLER_356_1014 ();
 b15zdnd11an1n08x5 FILLER_356_1046 ();
 b15zdnd11an1n04x5 FILLER_356_1054 ();
 b15zdnd00an1n01x5 FILLER_356_1058 ();
 b15zdnd11an1n64x5 FILLER_356_1065 ();
 b15zdnd11an1n32x5 FILLER_356_1129 ();
 b15zdnd11an1n16x5 FILLER_356_1161 ();
 b15zdnd00an1n01x5 FILLER_356_1177 ();
 b15zdnd11an1n04x5 FILLER_356_1183 ();
 b15zdnd00an1n02x5 FILLER_356_1187 ();
 b15zdnd00an1n01x5 FILLER_356_1189 ();
 b15zdnd11an1n32x5 FILLER_356_1199 ();
 b15zdnd11an1n16x5 FILLER_356_1231 ();
 b15zdnd11an1n08x5 FILLER_356_1247 ();
 b15zdnd00an1n02x5 FILLER_356_1255 ();
 b15zdnd00an1n01x5 FILLER_356_1257 ();
 b15zdnd11an1n64x5 FILLER_356_1269 ();
 b15zdnd11an1n32x5 FILLER_356_1333 ();
 b15zdnd00an1n02x5 FILLER_356_1365 ();
 b15zdnd11an1n04x5 FILLER_356_1375 ();
 b15zdnd00an1n02x5 FILLER_356_1379 ();
 b15zdnd11an1n64x5 FILLER_356_1387 ();
 b15zdnd11an1n16x5 FILLER_356_1451 ();
 b15zdnd11an1n08x5 FILLER_356_1467 ();
 b15zdnd11an1n64x5 FILLER_356_1482 ();
 b15zdnd11an1n64x5 FILLER_356_1553 ();
 b15zdnd11an1n16x5 FILLER_356_1617 ();
 b15zdnd11an1n16x5 FILLER_356_1637 ();
 b15zdnd11an1n08x5 FILLER_356_1653 ();
 b15zdnd11an1n04x5 FILLER_356_1661 ();
 b15zdnd11an1n64x5 FILLER_356_1678 ();
 b15zdnd11an1n08x5 FILLER_356_1742 ();
 b15zdnd00an1n02x5 FILLER_356_1750 ();
 b15zdnd00an1n01x5 FILLER_356_1752 ();
 b15zdnd11an1n64x5 FILLER_356_1766 ();
 b15zdnd11an1n16x5 FILLER_356_1830 ();
 b15zdnd11an1n08x5 FILLER_356_1846 ();
 b15zdnd00an1n02x5 FILLER_356_1854 ();
 b15zdnd11an1n32x5 FILLER_356_1862 ();
 b15zdnd00an1n02x5 FILLER_356_1894 ();
 b15zdnd11an1n32x5 FILLER_356_1900 ();
 b15zdnd11an1n16x5 FILLER_356_1932 ();
 b15zdnd11an1n04x5 FILLER_356_1948 ();
 b15zdnd00an1n02x5 FILLER_356_1952 ();
 b15zdnd11an1n64x5 FILLER_356_1960 ();
 b15zdnd11an1n64x5 FILLER_356_2024 ();
 b15zdnd11an1n04x5 FILLER_356_2088 ();
 b15zdnd11an1n32x5 FILLER_356_2099 ();
 b15zdnd11an1n16x5 FILLER_356_2131 ();
 b15zdnd11an1n04x5 FILLER_356_2147 ();
 b15zdnd00an1n02x5 FILLER_356_2151 ();
 b15zdnd00an1n01x5 FILLER_356_2153 ();
 b15zdnd11an1n04x5 FILLER_356_2162 ();
 b15zdnd00an1n02x5 FILLER_356_2166 ();
 b15zdnd00an1n01x5 FILLER_356_2168 ();
 b15zdnd11an1n08x5 FILLER_356_2178 ();
 b15zdnd00an1n02x5 FILLER_356_2186 ();
 b15zdnd00an1n01x5 FILLER_356_2188 ();
 b15zdnd11an1n16x5 FILLER_356_2196 ();
 b15zdnd11an1n32x5 FILLER_356_2228 ();
 b15zdnd11an1n16x5 FILLER_356_2260 ();
 b15zdnd11an1n64x5 FILLER_357_0 ();
 b15zdnd11an1n64x5 FILLER_357_64 ();
 b15zdnd11an1n64x5 FILLER_357_128 ();
 b15zdnd11an1n16x5 FILLER_357_192 ();
 b15zdnd11an1n08x5 FILLER_357_208 ();
 b15zdnd00an1n01x5 FILLER_357_216 ();
 b15zdnd11an1n32x5 FILLER_357_230 ();
 b15zdnd11an1n16x5 FILLER_357_262 ();
 b15zdnd11an1n08x5 FILLER_357_278 ();
 b15zdnd11an1n04x5 FILLER_357_286 ();
 b15zdnd11an1n64x5 FILLER_357_300 ();
 b15zdnd11an1n64x5 FILLER_357_364 ();
 b15zdnd11an1n32x5 FILLER_357_428 ();
 b15zdnd11an1n16x5 FILLER_357_460 ();
 b15zdnd00an1n01x5 FILLER_357_476 ();
 b15zdnd11an1n64x5 FILLER_357_491 ();
 b15zdnd11an1n64x5 FILLER_357_555 ();
 b15zdnd11an1n32x5 FILLER_357_619 ();
 b15zdnd00an1n02x5 FILLER_357_651 ();
 b15zdnd00an1n01x5 FILLER_357_653 ();
 b15zdnd11an1n04x5 FILLER_357_657 ();
 b15zdnd11an1n32x5 FILLER_357_666 ();
 b15zdnd00an1n01x5 FILLER_357_698 ();
 b15zdnd11an1n64x5 FILLER_357_713 ();
 b15zdnd11an1n16x5 FILLER_357_777 ();
 b15zdnd11an1n08x5 FILLER_357_793 ();
 b15zdnd11an1n04x5 FILLER_357_801 ();
 b15zdnd00an1n01x5 FILLER_357_805 ();
 b15zdnd11an1n08x5 FILLER_357_816 ();
 b15zdnd00an1n02x5 FILLER_357_824 ();
 b15zdnd00an1n01x5 FILLER_357_826 ();
 b15zdnd11an1n32x5 FILLER_357_848 ();
 b15zdnd11an1n08x5 FILLER_357_880 ();
 b15zdnd00an1n02x5 FILLER_357_888 ();
 b15zdnd00an1n01x5 FILLER_357_890 ();
 b15zdnd11an1n08x5 FILLER_357_896 ();
 b15zdnd11an1n04x5 FILLER_357_904 ();
 b15zdnd11an1n16x5 FILLER_357_920 ();
 b15zdnd11an1n08x5 FILLER_357_936 ();
 b15zdnd11an1n04x5 FILLER_357_944 ();
 b15zdnd00an1n02x5 FILLER_357_948 ();
 b15zdnd00an1n01x5 FILLER_357_950 ();
 b15zdnd11an1n16x5 FILLER_357_955 ();
 b15zdnd11an1n04x5 FILLER_357_971 ();
 b15zdnd00an1n02x5 FILLER_357_975 ();
 b15zdnd11an1n04x5 FILLER_357_985 ();
 b15zdnd11an1n04x5 FILLER_357_1001 ();
 b15zdnd11an1n04x5 FILLER_357_1020 ();
 b15zdnd11an1n04x5 FILLER_357_1028 ();
 b15zdnd00an1n02x5 FILLER_357_1032 ();
 b15zdnd00an1n01x5 FILLER_357_1034 ();
 b15zdnd11an1n04x5 FILLER_357_1040 ();
 b15zdnd11an1n16x5 FILLER_357_1054 ();
 b15zdnd11an1n08x5 FILLER_357_1070 ();
 b15zdnd00an1n02x5 FILLER_357_1078 ();
 b15zdnd00an1n01x5 FILLER_357_1080 ();
 b15zdnd11an1n64x5 FILLER_357_1087 ();
 b15zdnd11an1n64x5 FILLER_357_1151 ();
 b15zdnd11an1n64x5 FILLER_357_1215 ();
 b15zdnd11an1n32x5 FILLER_357_1279 ();
 b15zdnd11an1n16x5 FILLER_357_1311 ();
 b15zdnd11an1n04x5 FILLER_357_1327 ();
 b15zdnd00an1n02x5 FILLER_357_1331 ();
 b15zdnd00an1n01x5 FILLER_357_1333 ();
 b15zdnd11an1n04x5 FILLER_357_1346 ();
 b15zdnd11an1n04x5 FILLER_357_1378 ();
 b15zdnd00an1n01x5 FILLER_357_1382 ();
 b15zdnd11an1n32x5 FILLER_357_1389 ();
 b15zdnd11an1n04x5 FILLER_357_1421 ();
 b15zdnd00an1n01x5 FILLER_357_1425 ();
 b15zdnd11an1n08x5 FILLER_357_1438 ();
 b15zdnd11an1n04x5 FILLER_357_1446 ();
 b15zdnd00an1n02x5 FILLER_357_1450 ();
 b15zdnd00an1n01x5 FILLER_357_1452 ();
 b15zdnd11an1n08x5 FILLER_357_1465 ();
 b15zdnd11an1n04x5 FILLER_357_1473 ();
 b15zdnd00an1n02x5 FILLER_357_1477 ();
 b15zdnd00an1n01x5 FILLER_357_1479 ();
 b15zdnd11an1n32x5 FILLER_357_1486 ();
 b15zdnd11an1n08x5 FILLER_357_1518 ();
 b15zdnd11an1n08x5 FILLER_357_1532 ();
 b15zdnd11an1n04x5 FILLER_357_1540 ();
 b15zdnd00an1n02x5 FILLER_357_1544 ();
 b15zdnd11an1n64x5 FILLER_357_1552 ();
 b15zdnd11an1n16x5 FILLER_357_1616 ();
 b15zdnd11an1n04x5 FILLER_357_1632 ();
 b15zdnd00an1n02x5 FILLER_357_1636 ();
 b15zdnd11an1n32x5 FILLER_357_1642 ();
 b15zdnd00an1n02x5 FILLER_357_1674 ();
 b15zdnd00an1n01x5 FILLER_357_1676 ();
 b15zdnd11an1n32x5 FILLER_357_1687 ();
 b15zdnd11an1n64x5 FILLER_357_1735 ();
 b15zdnd11an1n16x5 FILLER_357_1799 ();
 b15zdnd11an1n08x5 FILLER_357_1815 ();
 b15zdnd00an1n01x5 FILLER_357_1823 ();
 b15zdnd11an1n16x5 FILLER_357_1830 ();
 b15zdnd11an1n08x5 FILLER_357_1846 ();
 b15zdnd11an1n16x5 FILLER_357_1860 ();
 b15zdnd11an1n08x5 FILLER_357_1876 ();
 b15zdnd00an1n02x5 FILLER_357_1884 ();
 b15zdnd11an1n64x5 FILLER_357_1891 ();
 b15zdnd11an1n32x5 FILLER_357_1955 ();
 b15zdnd11an1n16x5 FILLER_357_1987 ();
 b15zdnd11an1n04x5 FILLER_357_2003 ();
 b15zdnd11an1n32x5 FILLER_357_2012 ();
 b15zdnd11an1n08x5 FILLER_357_2044 ();
 b15zdnd00an1n02x5 FILLER_357_2052 ();
 b15zdnd00an1n01x5 FILLER_357_2054 ();
 b15zdnd11an1n04x5 FILLER_357_2060 ();
 b15zdnd11an1n16x5 FILLER_357_2073 ();
 b15zdnd11an1n04x5 FILLER_357_2089 ();
 b15zdnd11an1n32x5 FILLER_357_2099 ();
 b15zdnd00an1n02x5 FILLER_357_2131 ();
 b15zdnd00an1n01x5 FILLER_357_2133 ();
 b15zdnd11an1n16x5 FILLER_357_2142 ();
 b15zdnd11an1n04x5 FILLER_357_2158 ();
 b15zdnd11an1n08x5 FILLER_357_2167 ();
 b15zdnd11an1n04x5 FILLER_357_2175 ();
 b15zdnd00an1n01x5 FILLER_357_2179 ();
 b15zdnd11an1n64x5 FILLER_357_2186 ();
 b15zdnd11an1n32x5 FILLER_357_2250 ();
 b15zdnd00an1n02x5 FILLER_357_2282 ();
 b15zdnd11an1n64x5 FILLER_358_8 ();
 b15zdnd11an1n64x5 FILLER_358_72 ();
 b15zdnd11an1n64x5 FILLER_358_136 ();
 b15zdnd11an1n64x5 FILLER_358_200 ();
 b15zdnd11an1n08x5 FILLER_358_264 ();
 b15zdnd00an1n02x5 FILLER_358_272 ();
 b15zdnd00an1n01x5 FILLER_358_274 ();
 b15zdnd11an1n64x5 FILLER_358_280 ();
 b15zdnd11an1n64x5 FILLER_358_344 ();
 b15zdnd11an1n64x5 FILLER_358_408 ();
 b15zdnd11an1n64x5 FILLER_358_472 ();
 b15zdnd11an1n32x5 FILLER_358_536 ();
 b15zdnd11an1n16x5 FILLER_358_568 ();
 b15zdnd11an1n04x5 FILLER_358_584 ();
 b15zdnd00an1n01x5 FILLER_358_588 ();
 b15zdnd11an1n32x5 FILLER_358_593 ();
 b15zdnd11an1n16x5 FILLER_358_625 ();
 b15zdnd11an1n08x5 FILLER_358_641 ();
 b15zdnd11an1n04x5 FILLER_358_649 ();
 b15zdnd11an1n32x5 FILLER_358_667 ();
 b15zdnd11an1n16x5 FILLER_358_699 ();
 b15zdnd00an1n02x5 FILLER_358_715 ();
 b15zdnd00an1n01x5 FILLER_358_717 ();
 b15zdnd11an1n32x5 FILLER_358_726 ();
 b15zdnd00an1n02x5 FILLER_358_758 ();
 b15zdnd00an1n01x5 FILLER_358_760 ();
 b15zdnd11an1n16x5 FILLER_358_773 ();
 b15zdnd11an1n04x5 FILLER_358_802 ();
 b15zdnd11an1n32x5 FILLER_358_811 ();
 b15zdnd00an1n02x5 FILLER_358_843 ();
 b15zdnd11an1n16x5 FILLER_358_854 ();
 b15zdnd11an1n08x5 FILLER_358_870 ();
 b15zdnd11an1n04x5 FILLER_358_878 ();
 b15zdnd00an1n02x5 FILLER_358_882 ();
 b15zdnd00an1n01x5 FILLER_358_884 ();
 b15zdnd11an1n16x5 FILLER_358_897 ();
 b15zdnd11an1n08x5 FILLER_358_913 ();
 b15zdnd11an1n04x5 FILLER_358_921 ();
 b15zdnd00an1n01x5 FILLER_358_925 ();
 b15zdnd11an1n04x5 FILLER_358_946 ();
 b15zdnd11an1n08x5 FILLER_358_959 ();
 b15zdnd00an1n01x5 FILLER_358_967 ();
 b15zdnd11an1n32x5 FILLER_358_975 ();
 b15zdnd11an1n04x5 FILLER_358_1007 ();
 b15zdnd00an1n02x5 FILLER_358_1011 ();
 b15zdnd11an1n16x5 FILLER_358_1019 ();
 b15zdnd11an1n08x5 FILLER_358_1035 ();
 b15zdnd11an1n04x5 FILLER_358_1043 ();
 b15zdnd00an1n01x5 FILLER_358_1047 ();
 b15zdnd11an1n32x5 FILLER_358_1055 ();
 b15zdnd11an1n08x5 FILLER_358_1087 ();
 b15zdnd11an1n04x5 FILLER_358_1095 ();
 b15zdnd00an1n01x5 FILLER_358_1099 ();
 b15zdnd11an1n04x5 FILLER_358_1111 ();
 b15zdnd11an1n04x5 FILLER_358_1131 ();
 b15zdnd00an1n01x5 FILLER_358_1135 ();
 b15zdnd11an1n64x5 FILLER_358_1152 ();
 b15zdnd11an1n32x5 FILLER_358_1216 ();
 b15zdnd11an1n08x5 FILLER_358_1248 ();
 b15zdnd11an1n04x5 FILLER_358_1256 ();
 b15zdnd00an1n02x5 FILLER_358_1260 ();
 b15zdnd00an1n01x5 FILLER_358_1262 ();
 b15zdnd11an1n32x5 FILLER_358_1279 ();
 b15zdnd11an1n16x5 FILLER_358_1311 ();
 b15zdnd11an1n04x5 FILLER_358_1327 ();
 b15zdnd00an1n01x5 FILLER_358_1331 ();
 b15zdnd11an1n32x5 FILLER_358_1336 ();
 b15zdnd11an1n16x5 FILLER_358_1368 ();
 b15zdnd11an1n04x5 FILLER_358_1384 ();
 b15zdnd00an1n02x5 FILLER_358_1388 ();
 b15zdnd11an1n08x5 FILLER_358_1395 ();
 b15zdnd11an1n04x5 FILLER_358_1403 ();
 b15zdnd00an1n02x5 FILLER_358_1407 ();
 b15zdnd00an1n01x5 FILLER_358_1409 ();
 b15zdnd11an1n08x5 FILLER_358_1417 ();
 b15zdnd00an1n02x5 FILLER_358_1425 ();
 b15zdnd11an1n32x5 FILLER_358_1441 ();
 b15zdnd11an1n08x5 FILLER_358_1473 ();
 b15zdnd11an1n04x5 FILLER_358_1481 ();
 b15zdnd00an1n01x5 FILLER_358_1485 ();
 b15zdnd11an1n32x5 FILLER_358_1498 ();
 b15zdnd11an1n08x5 FILLER_358_1535 ();
 b15zdnd11an1n04x5 FILLER_358_1543 ();
 b15zdnd00an1n01x5 FILLER_358_1547 ();
 b15zdnd11an1n08x5 FILLER_358_1564 ();
 b15zdnd11an1n04x5 FILLER_358_1572 ();
 b15zdnd00an1n02x5 FILLER_358_1576 ();
 b15zdnd00an1n01x5 FILLER_358_1578 ();
 b15zdnd11an1n32x5 FILLER_358_1584 ();
 b15zdnd11an1n04x5 FILLER_358_1616 ();
 b15zdnd00an1n02x5 FILLER_358_1620 ();
 b15zdnd11an1n16x5 FILLER_358_1627 ();
 b15zdnd11an1n04x5 FILLER_358_1648 ();
 b15zdnd11an1n04x5 FILLER_358_1669 ();
 b15zdnd11an1n64x5 FILLER_358_1690 ();
 b15zdnd11an1n32x5 FILLER_358_1754 ();
 b15zdnd11an1n16x5 FILLER_358_1786 ();
 b15zdnd11an1n08x5 FILLER_358_1802 ();
 b15zdnd11an1n04x5 FILLER_358_1810 ();
 b15zdnd00an1n02x5 FILLER_358_1814 ();
 b15zdnd11an1n08x5 FILLER_358_1821 ();
 b15zdnd11an1n04x5 FILLER_358_1829 ();
 b15zdnd00an1n02x5 FILLER_358_1833 ();
 b15zdnd11an1n08x5 FILLER_358_1845 ();
 b15zdnd11an1n04x5 FILLER_358_1853 ();
 b15zdnd00an1n01x5 FILLER_358_1857 ();
 b15zdnd11an1n16x5 FILLER_358_1867 ();
 b15zdnd11an1n04x5 FILLER_358_1883 ();
 b15zdnd00an1n02x5 FILLER_358_1887 ();
 b15zdnd11an1n08x5 FILLER_358_1901 ();
 b15zdnd00an1n02x5 FILLER_358_1909 ();
 b15zdnd11an1n32x5 FILLER_358_1924 ();
 b15zdnd11an1n08x5 FILLER_358_1956 ();
 b15zdnd11an1n04x5 FILLER_358_1964 ();
 b15zdnd00an1n02x5 FILLER_358_1968 ();
 b15zdnd00an1n01x5 FILLER_358_1970 ();
 b15zdnd11an1n32x5 FILLER_358_1976 ();
 b15zdnd11an1n04x5 FILLER_358_2008 ();
 b15zdnd00an1n02x5 FILLER_358_2012 ();
 b15zdnd11an1n16x5 FILLER_358_2019 ();
 b15zdnd11an1n04x5 FILLER_358_2035 ();
 b15zdnd00an1n02x5 FILLER_358_2039 ();
 b15zdnd11an1n16x5 FILLER_358_2062 ();
 b15zdnd11an1n08x5 FILLER_358_2078 ();
 b15zdnd11an1n04x5 FILLER_358_2086 ();
 b15zdnd00an1n02x5 FILLER_358_2090 ();
 b15zdnd11an1n04x5 FILLER_358_2112 ();
 b15zdnd00an1n02x5 FILLER_358_2116 ();
 b15zdnd11an1n04x5 FILLER_358_2131 ();
 b15zdnd11an1n08x5 FILLER_358_2140 ();
 b15zdnd11an1n04x5 FILLER_358_2148 ();
 b15zdnd00an1n02x5 FILLER_358_2152 ();
 b15zdnd11an1n32x5 FILLER_358_2162 ();
 b15zdnd11an1n16x5 FILLER_358_2194 ();
 b15zdnd00an1n02x5 FILLER_358_2210 ();
 b15zdnd00an1n01x5 FILLER_358_2212 ();
 b15zdnd11an1n04x5 FILLER_358_2229 ();
 b15zdnd11an1n08x5 FILLER_358_2264 ();
 b15zdnd11an1n04x5 FILLER_358_2272 ();
 b15zdnd11an1n64x5 FILLER_359_0 ();
 b15zdnd11an1n64x5 FILLER_359_64 ();
 b15zdnd11an1n64x5 FILLER_359_128 ();
 b15zdnd11an1n16x5 FILLER_359_192 ();
 b15zdnd11an1n08x5 FILLER_359_208 ();
 b15zdnd00an1n02x5 FILLER_359_216 ();
 b15zdnd00an1n01x5 FILLER_359_218 ();
 b15zdnd11an1n04x5 FILLER_359_250 ();
 b15zdnd11an1n04x5 FILLER_359_258 ();
 b15zdnd11an1n08x5 FILLER_359_268 ();
 b15zdnd00an1n02x5 FILLER_359_276 ();
 b15zdnd00an1n01x5 FILLER_359_278 ();
 b15zdnd11an1n08x5 FILLER_359_294 ();
 b15zdnd00an1n01x5 FILLER_359_302 ();
 b15zdnd11an1n08x5 FILLER_359_313 ();
 b15zdnd00an1n02x5 FILLER_359_321 ();
 b15zdnd00an1n01x5 FILLER_359_323 ();
 b15zdnd11an1n32x5 FILLER_359_331 ();
 b15zdnd11an1n08x5 FILLER_359_363 ();
 b15zdnd00an1n02x5 FILLER_359_371 ();
 b15zdnd00an1n01x5 FILLER_359_373 ();
 b15zdnd11an1n08x5 FILLER_359_390 ();
 b15zdnd11an1n04x5 FILLER_359_398 ();
 b15zdnd00an1n02x5 FILLER_359_402 ();
 b15zdnd00an1n01x5 FILLER_359_404 ();
 b15zdnd11an1n08x5 FILLER_359_425 ();
 b15zdnd11an1n04x5 FILLER_359_433 ();
 b15zdnd11an1n32x5 FILLER_359_443 ();
 b15zdnd11an1n16x5 FILLER_359_475 ();
 b15zdnd00an1n02x5 FILLER_359_491 ();
 b15zdnd11an1n04x5 FILLER_359_497 ();
 b15zdnd11an1n08x5 FILLER_359_515 ();
 b15zdnd11an1n04x5 FILLER_359_523 ();
 b15zdnd00an1n02x5 FILLER_359_527 ();
 b15zdnd11an1n32x5 FILLER_359_560 ();
 b15zdnd00an1n02x5 FILLER_359_592 ();
 b15zdnd11an1n32x5 FILLER_359_620 ();
 b15zdnd00an1n02x5 FILLER_359_652 ();
 b15zdnd11an1n08x5 FILLER_359_679 ();
 b15zdnd11an1n04x5 FILLER_359_687 ();
 b15zdnd00an1n01x5 FILLER_359_691 ();
 b15zdnd11an1n16x5 FILLER_359_698 ();
 b15zdnd11an1n04x5 FILLER_359_714 ();
 b15zdnd00an1n01x5 FILLER_359_718 ();
 b15zdnd11an1n32x5 FILLER_359_726 ();
 b15zdnd11an1n04x5 FILLER_359_758 ();
 b15zdnd00an1n02x5 FILLER_359_762 ();
 b15zdnd11an1n08x5 FILLER_359_774 ();
 b15zdnd00an1n02x5 FILLER_359_782 ();
 b15zdnd11an1n64x5 FILLER_359_796 ();
 b15zdnd11an1n32x5 FILLER_359_860 ();
 b15zdnd11an1n16x5 FILLER_359_892 ();
 b15zdnd11an1n04x5 FILLER_359_908 ();
 b15zdnd00an1n02x5 FILLER_359_912 ();
 b15zdnd00an1n01x5 FILLER_359_914 ();
 b15zdnd11an1n32x5 FILLER_359_921 ();
 b15zdnd00an1n01x5 FILLER_359_953 ();
 b15zdnd11an1n04x5 FILLER_359_958 ();
 b15zdnd00an1n02x5 FILLER_359_962 ();
 b15zdnd11an1n32x5 FILLER_359_969 ();
 b15zdnd11an1n08x5 FILLER_359_1001 ();
 b15zdnd11an1n16x5 FILLER_359_1014 ();
 b15zdnd00an1n02x5 FILLER_359_1030 ();
 b15zdnd00an1n01x5 FILLER_359_1032 ();
 b15zdnd11an1n08x5 FILLER_359_1073 ();
 b15zdnd11an1n16x5 FILLER_359_1092 ();
 b15zdnd11an1n08x5 FILLER_359_1108 ();
 b15zdnd11an1n04x5 FILLER_359_1116 ();
 b15zdnd00an1n02x5 FILLER_359_1120 ();
 b15zdnd00an1n01x5 FILLER_359_1122 ();
 b15zdnd11an1n08x5 FILLER_359_1128 ();
 b15zdnd11an1n04x5 FILLER_359_1142 ();
 b15zdnd11an1n04x5 FILLER_359_1172 ();
 b15zdnd11an1n64x5 FILLER_359_1185 ();
 b15zdnd11an1n16x5 FILLER_359_1249 ();
 b15zdnd00an1n02x5 FILLER_359_1265 ();
 b15zdnd11an1n04x5 FILLER_359_1273 ();
 b15zdnd11an1n16x5 FILLER_359_1295 ();
 b15zdnd00an1n02x5 FILLER_359_1311 ();
 b15zdnd00an1n01x5 FILLER_359_1313 ();
 b15zdnd11an1n04x5 FILLER_359_1323 ();
 b15zdnd11an1n16x5 FILLER_359_1332 ();
 b15zdnd11an1n08x5 FILLER_359_1348 ();
 b15zdnd11an1n04x5 FILLER_359_1356 ();
 b15zdnd11an1n08x5 FILLER_359_1370 ();
 b15zdnd11an1n04x5 FILLER_359_1378 ();
 b15zdnd11an1n16x5 FILLER_359_1388 ();
 b15zdnd11an1n04x5 FILLER_359_1404 ();
 b15zdnd11an1n08x5 FILLER_359_1418 ();
 b15zdnd11an1n04x5 FILLER_359_1426 ();
 b15zdnd11an1n16x5 FILLER_359_1435 ();
 b15zdnd11an1n04x5 FILLER_359_1451 ();
 b15zdnd11an1n04x5 FILLER_359_1459 ();
 b15zdnd11an1n64x5 FILLER_359_1470 ();
 b15zdnd11an1n16x5 FILLER_359_1534 ();
 b15zdnd11an1n08x5 FILLER_359_1550 ();
 b15zdnd00an1n02x5 FILLER_359_1558 ();
 b15zdnd11an1n16x5 FILLER_359_1572 ();
 b15zdnd11an1n04x5 FILLER_359_1588 ();
 b15zdnd00an1n01x5 FILLER_359_1592 ();
 b15zdnd11an1n16x5 FILLER_359_1602 ();
 b15zdnd00an1n02x5 FILLER_359_1618 ();
 b15zdnd00an1n01x5 FILLER_359_1620 ();
 b15zdnd11an1n32x5 FILLER_359_1627 ();
 b15zdnd11an1n16x5 FILLER_359_1659 ();
 b15zdnd11an1n08x5 FILLER_359_1675 ();
 b15zdnd11an1n16x5 FILLER_359_1688 ();
 b15zdnd11an1n04x5 FILLER_359_1704 ();
 b15zdnd11an1n04x5 FILLER_359_1714 ();
 b15zdnd00an1n02x5 FILLER_359_1718 ();
 b15zdnd00an1n01x5 FILLER_359_1720 ();
 b15zdnd11an1n08x5 FILLER_359_1733 ();
 b15zdnd00an1n01x5 FILLER_359_1741 ();
 b15zdnd11an1n64x5 FILLER_359_1750 ();
 b15zdnd00an1n02x5 FILLER_359_1814 ();
 b15zdnd00an1n01x5 FILLER_359_1816 ();
 b15zdnd11an1n08x5 FILLER_359_1823 ();
 b15zdnd11an1n32x5 FILLER_359_1837 ();
 b15zdnd11an1n16x5 FILLER_359_1869 ();
 b15zdnd11an1n04x5 FILLER_359_1885 ();
 b15zdnd00an1n02x5 FILLER_359_1889 ();
 b15zdnd11an1n08x5 FILLER_359_1895 ();
 b15zdnd11an1n04x5 FILLER_359_1903 ();
 b15zdnd00an1n02x5 FILLER_359_1907 ();
 b15zdnd00an1n01x5 FILLER_359_1909 ();
 b15zdnd11an1n04x5 FILLER_359_1920 ();
 b15zdnd11an1n08x5 FILLER_359_1934 ();
 b15zdnd11an1n04x5 FILLER_359_1942 ();
 b15zdnd00an1n02x5 FILLER_359_1946 ();
 b15zdnd11an1n04x5 FILLER_359_1955 ();
 b15zdnd11an1n08x5 FILLER_359_1963 ();
 b15zdnd00an1n02x5 FILLER_359_1971 ();
 b15zdnd11an1n16x5 FILLER_359_1983 ();
 b15zdnd11an1n08x5 FILLER_359_2020 ();
 b15zdnd11an1n04x5 FILLER_359_2028 ();
 b15zdnd00an1n02x5 FILLER_359_2032 ();
 b15zdnd11an1n08x5 FILLER_359_2040 ();
 b15zdnd11an1n04x5 FILLER_359_2048 ();
 b15zdnd00an1n02x5 FILLER_359_2052 ();
 b15zdnd11an1n32x5 FILLER_359_2059 ();
 b15zdnd11an1n04x5 FILLER_359_2098 ();
 b15zdnd11an1n16x5 FILLER_359_2107 ();
 b15zdnd00an1n01x5 FILLER_359_2123 ();
 b15zdnd11an1n04x5 FILLER_359_2132 ();
 b15zdnd00an1n02x5 FILLER_359_2136 ();
 b15zdnd11an1n32x5 FILLER_359_2143 ();
 b15zdnd11an1n16x5 FILLER_359_2175 ();
 b15zdnd11an1n04x5 FILLER_359_2196 ();
 b15zdnd11an1n64x5 FILLER_359_2212 ();
 b15zdnd11an1n08x5 FILLER_359_2276 ();
 b15zdnd11an1n64x5 FILLER_360_8 ();
 b15zdnd11an1n64x5 FILLER_360_72 ();
 b15zdnd11an1n64x5 FILLER_360_136 ();
 b15zdnd11an1n32x5 FILLER_360_200 ();
 b15zdnd11an1n16x5 FILLER_360_232 ();
 b15zdnd00an1n02x5 FILLER_360_248 ();
 b15zdnd00an1n01x5 FILLER_360_250 ();
 b15zdnd11an1n16x5 FILLER_360_265 ();
 b15zdnd11an1n08x5 FILLER_360_281 ();
 b15zdnd00an1n02x5 FILLER_360_289 ();
 b15zdnd00an1n01x5 FILLER_360_291 ();
 b15zdnd11an1n04x5 FILLER_360_312 ();
 b15zdnd11an1n16x5 FILLER_360_323 ();
 b15zdnd11an1n08x5 FILLER_360_339 ();
 b15zdnd11an1n04x5 FILLER_360_347 ();
 b15zdnd00an1n02x5 FILLER_360_351 ();
 b15zdnd11an1n16x5 FILLER_360_360 ();
 b15zdnd11an1n08x5 FILLER_360_391 ();
 b15zdnd00an1n02x5 FILLER_360_399 ();
 b15zdnd00an1n01x5 FILLER_360_401 ();
 b15zdnd11an1n04x5 FILLER_360_407 ();
 b15zdnd11an1n16x5 FILLER_360_420 ();
 b15zdnd11an1n04x5 FILLER_360_436 ();
 b15zdnd11an1n08x5 FILLER_360_446 ();
 b15zdnd00an1n01x5 FILLER_360_454 ();
 b15zdnd11an1n16x5 FILLER_360_470 ();
 b15zdnd00an1n01x5 FILLER_360_486 ();
 b15zdnd11an1n32x5 FILLER_360_496 ();
 b15zdnd11an1n16x5 FILLER_360_528 ();
 b15zdnd00an1n01x5 FILLER_360_544 ();
 b15zdnd11an1n32x5 FILLER_360_549 ();
 b15zdnd11an1n04x5 FILLER_360_581 ();
 b15zdnd00an1n01x5 FILLER_360_585 ();
 b15zdnd11an1n04x5 FILLER_360_592 ();
 b15zdnd11an1n32x5 FILLER_360_616 ();
 b15zdnd11an1n04x5 FILLER_360_648 ();
 b15zdnd00an1n02x5 FILLER_360_652 ();
 b15zdnd00an1n01x5 FILLER_360_654 ();
 b15zdnd11an1n32x5 FILLER_360_662 ();
 b15zdnd11an1n08x5 FILLER_360_694 ();
 b15zdnd00an1n02x5 FILLER_360_702 ();
 b15zdnd00an1n02x5 FILLER_360_716 ();
 b15zdnd11an1n08x5 FILLER_360_726 ();
 b15zdnd00an1n01x5 FILLER_360_734 ();
 b15zdnd11an1n16x5 FILLER_360_746 ();
 b15zdnd11an1n08x5 FILLER_360_762 ();
 b15zdnd00an1n01x5 FILLER_360_770 ();
 b15zdnd11an1n16x5 FILLER_360_775 ();
 b15zdnd11an1n08x5 FILLER_360_791 ();
 b15zdnd11an1n04x5 FILLER_360_799 ();
 b15zdnd00an1n02x5 FILLER_360_803 ();
 b15zdnd11an1n32x5 FILLER_360_815 ();
 b15zdnd11an1n08x5 FILLER_360_847 ();
 b15zdnd11an1n04x5 FILLER_360_855 ();
 b15zdnd00an1n01x5 FILLER_360_859 ();
 b15zdnd11an1n32x5 FILLER_360_865 ();
 b15zdnd11an1n16x5 FILLER_360_897 ();
 b15zdnd00an1n01x5 FILLER_360_913 ();
 b15zdnd11an1n04x5 FILLER_360_926 ();
 b15zdnd11an1n08x5 FILLER_360_938 ();
 b15zdnd11an1n04x5 FILLER_360_946 ();
 b15zdnd00an1n02x5 FILLER_360_950 ();
 b15zdnd00an1n01x5 FILLER_360_952 ();
 b15zdnd11an1n64x5 FILLER_360_959 ();
 b15zdnd11an1n64x5 FILLER_360_1023 ();
 b15zdnd11an1n64x5 FILLER_360_1087 ();
 b15zdnd11an1n04x5 FILLER_360_1151 ();
 b15zdnd00an1n02x5 FILLER_360_1155 ();
 b15zdnd00an1n01x5 FILLER_360_1157 ();
 b15zdnd11an1n08x5 FILLER_360_1168 ();
 b15zdnd00an1n01x5 FILLER_360_1176 ();
 b15zdnd11an1n64x5 FILLER_360_1187 ();
 b15zdnd11an1n32x5 FILLER_360_1251 ();
 b15zdnd11an1n16x5 FILLER_360_1283 ();
 b15zdnd11an1n08x5 FILLER_360_1299 ();
 b15zdnd11an1n04x5 FILLER_360_1307 ();
 b15zdnd00an1n02x5 FILLER_360_1311 ();
 b15zdnd11an1n04x5 FILLER_360_1329 ();
 b15zdnd00an1n01x5 FILLER_360_1333 ();
 b15zdnd11an1n16x5 FILLER_360_1342 ();
 b15zdnd11an1n08x5 FILLER_360_1358 ();
 b15zdnd00an1n01x5 FILLER_360_1366 ();
 b15zdnd11an1n04x5 FILLER_360_1380 ();
 b15zdnd11an1n32x5 FILLER_360_1390 ();
 b15zdnd11an1n16x5 FILLER_360_1422 ();
 b15zdnd11an1n08x5 FILLER_360_1438 ();
 b15zdnd11an1n04x5 FILLER_360_1446 ();
 b15zdnd11an1n16x5 FILLER_360_1457 ();
 b15zdnd11an1n08x5 FILLER_360_1473 ();
 b15zdnd11an1n04x5 FILLER_360_1481 ();
 b15zdnd00an1n02x5 FILLER_360_1485 ();
 b15zdnd00an1n01x5 FILLER_360_1487 ();
 b15zdnd11an1n04x5 FILLER_360_1492 ();
 b15zdnd11an1n32x5 FILLER_360_1502 ();
 b15zdnd11an1n16x5 FILLER_360_1534 ();
 b15zdnd11an1n08x5 FILLER_360_1550 ();
 b15zdnd00an1n02x5 FILLER_360_1558 ();
 b15zdnd11an1n04x5 FILLER_360_1569 ();
 b15zdnd11an1n32x5 FILLER_360_1584 ();
 b15zdnd11an1n08x5 FILLER_360_1616 ();
 b15zdnd00an1n01x5 FILLER_360_1624 ();
 b15zdnd11an1n64x5 FILLER_360_1634 ();
 b15zdnd11an1n16x5 FILLER_360_1698 ();
 b15zdnd11an1n08x5 FILLER_360_1714 ();
 b15zdnd00an1n02x5 FILLER_360_1722 ();
 b15zdnd11an1n64x5 FILLER_360_1748 ();
 b15zdnd11an1n08x5 FILLER_360_1812 ();
 b15zdnd11an1n04x5 FILLER_360_1820 ();
 b15zdnd00an1n02x5 FILLER_360_1824 ();
 b15zdnd00an1n01x5 FILLER_360_1826 ();
 b15zdnd11an1n32x5 FILLER_360_1853 ();
 b15zdnd11an1n04x5 FILLER_360_1885 ();
 b15zdnd11an1n32x5 FILLER_360_1893 ();
 b15zdnd00an1n02x5 FILLER_360_1925 ();
 b15zdnd11an1n04x5 FILLER_360_1947 ();
 b15zdnd00an1n01x5 FILLER_360_1951 ();
 b15zdnd11an1n04x5 FILLER_360_1966 ();
 b15zdnd00an1n02x5 FILLER_360_1970 ();
 b15zdnd11an1n04x5 FILLER_360_1978 ();
 b15zdnd00an1n02x5 FILLER_360_1982 ();
 b15zdnd11an1n04x5 FILLER_360_1995 ();
 b15zdnd00an1n02x5 FILLER_360_1999 ();
 b15zdnd11an1n04x5 FILLER_360_2011 ();
 b15zdnd11an1n08x5 FILLER_360_2021 ();
 b15zdnd11an1n04x5 FILLER_360_2029 ();
 b15zdnd00an1n02x5 FILLER_360_2033 ();
 b15zdnd00an1n01x5 FILLER_360_2035 ();
 b15zdnd11an1n64x5 FILLER_360_2044 ();
 b15zdnd11an1n32x5 FILLER_360_2108 ();
 b15zdnd11an1n08x5 FILLER_360_2140 ();
 b15zdnd11an1n04x5 FILLER_360_2148 ();
 b15zdnd00an1n02x5 FILLER_360_2152 ();
 b15zdnd11an1n04x5 FILLER_360_2162 ();
 b15zdnd00an1n02x5 FILLER_360_2166 ();
 b15zdnd11an1n04x5 FILLER_360_2174 ();
 b15zdnd11an1n64x5 FILLER_360_2204 ();
 b15zdnd11an1n08x5 FILLER_360_2268 ();
 b15zdnd11an1n64x5 FILLER_361_0 ();
 b15zdnd11an1n64x5 FILLER_361_64 ();
 b15zdnd11an1n64x5 FILLER_361_128 ();
 b15zdnd11an1n16x5 FILLER_361_192 ();
 b15zdnd11an1n08x5 FILLER_361_208 ();
 b15zdnd00an1n01x5 FILLER_361_216 ();
 b15zdnd11an1n16x5 FILLER_361_233 ();
 b15zdnd00an1n02x5 FILLER_361_249 ();
 b15zdnd00an1n01x5 FILLER_361_251 ();
 b15zdnd11an1n32x5 FILLER_361_258 ();
 b15zdnd11an1n08x5 FILLER_361_290 ();
 b15zdnd11an1n04x5 FILLER_361_298 ();
 b15zdnd00an1n01x5 FILLER_361_302 ();
 b15zdnd11an1n16x5 FILLER_361_308 ();
 b15zdnd11an1n08x5 FILLER_361_324 ();
 b15zdnd11an1n04x5 FILLER_361_332 ();
 b15zdnd00an1n02x5 FILLER_361_336 ();
 b15zdnd00an1n01x5 FILLER_361_338 ();
 b15zdnd11an1n04x5 FILLER_361_353 ();
 b15zdnd11an1n08x5 FILLER_361_361 ();
 b15zdnd11an1n04x5 FILLER_361_369 ();
 b15zdnd11an1n08x5 FILLER_361_380 ();
 b15zdnd11an1n04x5 FILLER_361_388 ();
 b15zdnd11an1n64x5 FILLER_361_396 ();
 b15zdnd11an1n04x5 FILLER_361_460 ();
 b15zdnd00an1n02x5 FILLER_361_464 ();
 b15zdnd00an1n01x5 FILLER_361_466 ();
 b15zdnd11an1n16x5 FILLER_361_481 ();
 b15zdnd00an1n01x5 FILLER_361_497 ();
 b15zdnd11an1n16x5 FILLER_361_507 ();
 b15zdnd11an1n08x5 FILLER_361_523 ();
 b15zdnd00an1n02x5 FILLER_361_531 ();
 b15zdnd11an1n04x5 FILLER_361_537 ();
 b15zdnd00an1n01x5 FILLER_361_541 ();
 b15zdnd11an1n16x5 FILLER_361_556 ();
 b15zdnd11an1n08x5 FILLER_361_572 ();
 b15zdnd11an1n04x5 FILLER_361_580 ();
 b15zdnd00an1n01x5 FILLER_361_584 ();
 b15zdnd11an1n04x5 FILLER_361_601 ();
 b15zdnd11an1n32x5 FILLER_361_625 ();
 b15zdnd11an1n16x5 FILLER_361_657 ();
 b15zdnd11an1n04x5 FILLER_361_673 ();
 b15zdnd00an1n01x5 FILLER_361_677 ();
 b15zdnd11an1n16x5 FILLER_361_689 ();
 b15zdnd11an1n04x5 FILLER_361_705 ();
 b15zdnd11an1n32x5 FILLER_361_713 ();
 b15zdnd11an1n16x5 FILLER_361_745 ();
 b15zdnd11an1n16x5 FILLER_361_773 ();
 b15zdnd11an1n04x5 FILLER_361_789 ();
 b15zdnd00an1n01x5 FILLER_361_793 ();
 b15zdnd11an1n16x5 FILLER_361_801 ();
 b15zdnd11an1n04x5 FILLER_361_817 ();
 b15zdnd00an1n01x5 FILLER_361_821 ();
 b15zdnd11an1n16x5 FILLER_361_827 ();
 b15zdnd11an1n08x5 FILLER_361_843 ();
 b15zdnd00an1n02x5 FILLER_361_851 ();
 b15zdnd00an1n01x5 FILLER_361_853 ();
 b15zdnd11an1n32x5 FILLER_361_861 ();
 b15zdnd11an1n16x5 FILLER_361_899 ();
 b15zdnd00an1n01x5 FILLER_361_915 ();
 b15zdnd11an1n64x5 FILLER_361_922 ();
 b15zdnd11an1n64x5 FILLER_361_986 ();
 b15zdnd11an1n16x5 FILLER_361_1050 ();
 b15zdnd11an1n08x5 FILLER_361_1066 ();
 b15zdnd00an1n01x5 FILLER_361_1074 ();
 b15zdnd11an1n04x5 FILLER_361_1085 ();
 b15zdnd11an1n04x5 FILLER_361_1094 ();
 b15zdnd11an1n16x5 FILLER_361_1107 ();
 b15zdnd11an1n04x5 FILLER_361_1123 ();
 b15zdnd11an1n64x5 FILLER_361_1139 ();
 b15zdnd11an1n64x5 FILLER_361_1203 ();
 b15zdnd11an1n64x5 FILLER_361_1267 ();
 b15zdnd00an1n02x5 FILLER_361_1331 ();
 b15zdnd11an1n08x5 FILLER_361_1359 ();
 b15zdnd00an1n02x5 FILLER_361_1367 ();
 b15zdnd11an1n64x5 FILLER_361_1375 ();
 b15zdnd11an1n32x5 FILLER_361_1439 ();
 b15zdnd11an1n16x5 FILLER_361_1471 ();
 b15zdnd11an1n04x5 FILLER_361_1487 ();
 b15zdnd00an1n02x5 FILLER_361_1491 ();
 b15zdnd00an1n01x5 FILLER_361_1493 ();
 b15zdnd11an1n32x5 FILLER_361_1506 ();
 b15zdnd00an1n01x5 FILLER_361_1538 ();
 b15zdnd11an1n16x5 FILLER_361_1546 ();
 b15zdnd11an1n08x5 FILLER_361_1562 ();
 b15zdnd11an1n64x5 FILLER_361_1577 ();
 b15zdnd11an1n08x5 FILLER_361_1641 ();
 b15zdnd11an1n04x5 FILLER_361_1649 ();
 b15zdnd00an1n02x5 FILLER_361_1653 ();
 b15zdnd11an1n32x5 FILLER_361_1660 ();
 b15zdnd11an1n08x5 FILLER_361_1692 ();
 b15zdnd11an1n04x5 FILLER_361_1700 ();
 b15zdnd11an1n64x5 FILLER_361_1720 ();
 b15zdnd11an1n64x5 FILLER_361_1784 ();
 b15zdnd00an1n02x5 FILLER_361_1848 ();
 b15zdnd00an1n01x5 FILLER_361_1850 ();
 b15zdnd11an1n04x5 FILLER_361_1857 ();
 b15zdnd11an1n16x5 FILLER_361_1875 ();
 b15zdnd00an1n02x5 FILLER_361_1891 ();
 b15zdnd00an1n01x5 FILLER_361_1893 ();
 b15zdnd11an1n64x5 FILLER_361_1900 ();
 b15zdnd11an1n32x5 FILLER_361_1964 ();
 b15zdnd11an1n16x5 FILLER_361_1996 ();
 b15zdnd00an1n02x5 FILLER_361_2012 ();
 b15zdnd00an1n01x5 FILLER_361_2014 ();
 b15zdnd11an1n64x5 FILLER_361_2020 ();
 b15zdnd11an1n32x5 FILLER_361_2084 ();
 b15zdnd11an1n16x5 FILLER_361_2116 ();
 b15zdnd11an1n04x5 FILLER_361_2132 ();
 b15zdnd00an1n01x5 FILLER_361_2136 ();
 b15zdnd11an1n04x5 FILLER_361_2145 ();
 b15zdnd00an1n02x5 FILLER_361_2149 ();
 b15zdnd00an1n01x5 FILLER_361_2151 ();
 b15zdnd11an1n08x5 FILLER_361_2167 ();
 b15zdnd11an1n64x5 FILLER_361_2183 ();
 b15zdnd11an1n32x5 FILLER_361_2247 ();
 b15zdnd11an1n04x5 FILLER_361_2279 ();
 b15zdnd00an1n01x5 FILLER_361_2283 ();
 b15zdnd11an1n64x5 FILLER_362_8 ();
 b15zdnd11an1n64x5 FILLER_362_72 ();
 b15zdnd11an1n64x5 FILLER_362_136 ();
 b15zdnd11an1n32x5 FILLER_362_200 ();
 b15zdnd00an1n01x5 FILLER_362_232 ();
 b15zdnd11an1n04x5 FILLER_362_249 ();
 b15zdnd11an1n16x5 FILLER_362_271 ();
 b15zdnd11an1n04x5 FILLER_362_287 ();
 b15zdnd00an1n01x5 FILLER_362_291 ();
 b15zdnd11an1n16x5 FILLER_362_305 ();
 b15zdnd00an1n02x5 FILLER_362_321 ();
 b15zdnd11an1n64x5 FILLER_362_333 ();
 b15zdnd11an1n16x5 FILLER_362_397 ();
 b15zdnd11an1n04x5 FILLER_362_413 ();
 b15zdnd00an1n01x5 FILLER_362_417 ();
 b15zdnd11an1n16x5 FILLER_362_426 ();
 b15zdnd11an1n08x5 FILLER_362_447 ();
 b15zdnd11an1n04x5 FILLER_362_455 ();
 b15zdnd00an1n02x5 FILLER_362_459 ();
 b15zdnd00an1n01x5 FILLER_362_461 ();
 b15zdnd11an1n16x5 FILLER_362_468 ();
 b15zdnd11an1n08x5 FILLER_362_484 ();
 b15zdnd00an1n02x5 FILLER_362_492 ();
 b15zdnd11an1n04x5 FILLER_362_499 ();
 b15zdnd11an1n64x5 FILLER_362_513 ();
 b15zdnd11an1n16x5 FILLER_362_577 ();
 b15zdnd11an1n32x5 FILLER_362_597 ();
 b15zdnd11an1n08x5 FILLER_362_629 ();
 b15zdnd11an1n04x5 FILLER_362_637 ();
 b15zdnd11an1n08x5 FILLER_362_649 ();
 b15zdnd11an1n04x5 FILLER_362_657 ();
 b15zdnd00an1n01x5 FILLER_362_661 ();
 b15zdnd11an1n16x5 FILLER_362_667 ();
 b15zdnd11an1n08x5 FILLER_362_683 ();
 b15zdnd11an1n04x5 FILLER_362_691 ();
 b15zdnd00an1n01x5 FILLER_362_695 ();
 b15zdnd11an1n08x5 FILLER_362_700 ();
 b15zdnd00an1n02x5 FILLER_362_708 ();
 b15zdnd00an1n01x5 FILLER_362_710 ();
 b15zdnd00an1n02x5 FILLER_362_716 ();
 b15zdnd11an1n64x5 FILLER_362_726 ();
 b15zdnd00an1n01x5 FILLER_362_790 ();
 b15zdnd11an1n16x5 FILLER_362_796 ();
 b15zdnd11an1n08x5 FILLER_362_812 ();
 b15zdnd00an1n02x5 FILLER_362_820 ();
 b15zdnd00an1n01x5 FILLER_362_822 ();
 b15zdnd11an1n16x5 FILLER_362_835 ();
 b15zdnd11an1n04x5 FILLER_362_851 ();
 b15zdnd00an1n02x5 FILLER_362_855 ();
 b15zdnd11an1n16x5 FILLER_362_869 ();
 b15zdnd11an1n08x5 FILLER_362_885 ();
 b15zdnd00an1n02x5 FILLER_362_893 ();
 b15zdnd11an1n16x5 FILLER_362_899 ();
 b15zdnd11an1n64x5 FILLER_362_919 ();
 b15zdnd11an1n64x5 FILLER_362_983 ();
 b15zdnd11an1n08x5 FILLER_362_1047 ();
 b15zdnd11an1n04x5 FILLER_362_1055 ();
 b15zdnd00an1n02x5 FILLER_362_1059 ();
 b15zdnd00an1n01x5 FILLER_362_1061 ();
 b15zdnd11an1n08x5 FILLER_362_1067 ();
 b15zdnd00an1n02x5 FILLER_362_1075 ();
 b15zdnd11an1n64x5 FILLER_362_1084 ();
 b15zdnd11an1n64x5 FILLER_362_1148 ();
 b15zdnd11an1n64x5 FILLER_362_1212 ();
 b15zdnd11an1n64x5 FILLER_362_1276 ();
 b15zdnd11an1n64x5 FILLER_362_1340 ();
 b15zdnd11an1n64x5 FILLER_362_1404 ();
 b15zdnd11an1n16x5 FILLER_362_1468 ();
 b15zdnd11an1n04x5 FILLER_362_1484 ();
 b15zdnd00an1n02x5 FILLER_362_1488 ();
 b15zdnd11an1n64x5 FILLER_362_1494 ();
 b15zdnd11an1n64x5 FILLER_362_1558 ();
 b15zdnd11an1n08x5 FILLER_362_1622 ();
 b15zdnd11an1n04x5 FILLER_362_1630 ();
 b15zdnd00an1n02x5 FILLER_362_1634 ();
 b15zdnd00an1n01x5 FILLER_362_1636 ();
 b15zdnd11an1n04x5 FILLER_362_1650 ();
 b15zdnd11an1n08x5 FILLER_362_1663 ();
 b15zdnd11an1n04x5 FILLER_362_1671 ();
 b15zdnd11an1n32x5 FILLER_362_1687 ();
 b15zdnd11an1n08x5 FILLER_362_1719 ();
 b15zdnd11an1n04x5 FILLER_362_1727 ();
 b15zdnd11an1n08x5 FILLER_362_1735 ();
 b15zdnd00an1n01x5 FILLER_362_1743 ();
 b15zdnd11an1n64x5 FILLER_362_1754 ();
 b15zdnd11an1n08x5 FILLER_362_1818 ();
 b15zdnd00an1n01x5 FILLER_362_1826 ();
 b15zdnd11an1n32x5 FILLER_362_1837 ();
 b15zdnd11an1n16x5 FILLER_362_1869 ();
 b15zdnd11an1n04x5 FILLER_362_1885 ();
 b15zdnd11an1n64x5 FILLER_362_1896 ();
 b15zdnd11an1n64x5 FILLER_362_1960 ();
 b15zdnd11an1n64x5 FILLER_362_2024 ();
 b15zdnd11an1n32x5 FILLER_362_2088 ();
 b15zdnd11an1n04x5 FILLER_362_2120 ();
 b15zdnd00an1n02x5 FILLER_362_2124 ();
 b15zdnd11an1n08x5 FILLER_362_2145 ();
 b15zdnd00an1n01x5 FILLER_362_2153 ();
 b15zdnd11an1n32x5 FILLER_362_2162 ();
 b15zdnd11an1n16x5 FILLER_362_2194 ();
 b15zdnd00an1n02x5 FILLER_362_2210 ();
 b15zdnd11an1n32x5 FILLER_362_2224 ();
 b15zdnd11an1n16x5 FILLER_362_2256 ();
 b15zdnd11an1n04x5 FILLER_362_2272 ();
 b15zdnd11an1n64x5 FILLER_363_0 ();
 b15zdnd11an1n64x5 FILLER_363_64 ();
 b15zdnd11an1n64x5 FILLER_363_128 ();
 b15zdnd11an1n64x5 FILLER_363_192 ();
 b15zdnd11an1n08x5 FILLER_363_256 ();
 b15zdnd11an1n04x5 FILLER_363_264 ();
 b15zdnd11an1n32x5 FILLER_363_283 ();
 b15zdnd11an1n16x5 FILLER_363_315 ();
 b15zdnd11an1n08x5 FILLER_363_331 ();
 b15zdnd00an1n01x5 FILLER_363_339 ();
 b15zdnd11an1n16x5 FILLER_363_352 ();
 b15zdnd00an1n02x5 FILLER_363_368 ();
 b15zdnd11an1n04x5 FILLER_363_376 ();
 b15zdnd00an1n02x5 FILLER_363_380 ();
 b15zdnd00an1n01x5 FILLER_363_382 ();
 b15zdnd11an1n16x5 FILLER_363_389 ();
 b15zdnd11an1n08x5 FILLER_363_405 ();
 b15zdnd11an1n04x5 FILLER_363_413 ();
 b15zdnd00an1n02x5 FILLER_363_417 ();
 b15zdnd00an1n01x5 FILLER_363_419 ();
 b15zdnd11an1n16x5 FILLER_363_424 ();
 b15zdnd00an1n01x5 FILLER_363_440 ();
 b15zdnd11an1n08x5 FILLER_363_447 ();
 b15zdnd11an1n04x5 FILLER_363_455 ();
 b15zdnd00an1n01x5 FILLER_363_459 ();
 b15zdnd11an1n64x5 FILLER_363_465 ();
 b15zdnd11an1n08x5 FILLER_363_529 ();
 b15zdnd11an1n16x5 FILLER_363_562 ();
 b15zdnd11an1n04x5 FILLER_363_578 ();
 b15zdnd00an1n02x5 FILLER_363_582 ();
 b15zdnd00an1n01x5 FILLER_363_584 ();
 b15zdnd11an1n32x5 FILLER_363_591 ();
 b15zdnd11an1n16x5 FILLER_363_623 ();
 b15zdnd11an1n08x5 FILLER_363_639 ();
 b15zdnd11an1n04x5 FILLER_363_647 ();
 b15zdnd11an1n04x5 FILLER_363_656 ();
 b15zdnd00an1n02x5 FILLER_363_660 ();
 b15zdnd11an1n16x5 FILLER_363_669 ();
 b15zdnd11an1n32x5 FILLER_363_692 ();
 b15zdnd00an1n01x5 FILLER_363_724 ();
 b15zdnd11an1n32x5 FILLER_363_735 ();
 b15zdnd11an1n08x5 FILLER_363_767 ();
 b15zdnd00an1n01x5 FILLER_363_775 ();
 b15zdnd11an1n04x5 FILLER_363_782 ();
 b15zdnd00an1n02x5 FILLER_363_786 ();
 b15zdnd00an1n01x5 FILLER_363_788 ();
 b15zdnd11an1n16x5 FILLER_363_799 ();
 b15zdnd11an1n08x5 FILLER_363_815 ();
 b15zdnd00an1n01x5 FILLER_363_823 ();
 b15zdnd11an1n32x5 FILLER_363_836 ();
 b15zdnd11an1n16x5 FILLER_363_868 ();
 b15zdnd11an1n04x5 FILLER_363_884 ();
 b15zdnd11an1n04x5 FILLER_363_897 ();
 b15zdnd11an1n32x5 FILLER_363_906 ();
 b15zdnd11an1n16x5 FILLER_363_938 ();
 b15zdnd11an1n08x5 FILLER_363_954 ();
 b15zdnd11an1n32x5 FILLER_363_966 ();
 b15zdnd00an1n01x5 FILLER_363_998 ();
 b15zdnd11an1n04x5 FILLER_363_1004 ();
 b15zdnd11an1n16x5 FILLER_363_1017 ();
 b15zdnd00an1n01x5 FILLER_363_1033 ();
 b15zdnd11an1n08x5 FILLER_363_1045 ();
 b15zdnd11an1n04x5 FILLER_363_1053 ();
 b15zdnd00an1n02x5 FILLER_363_1057 ();
 b15zdnd00an1n01x5 FILLER_363_1059 ();
 b15zdnd11an1n32x5 FILLER_363_1076 ();
 b15zdnd11an1n16x5 FILLER_363_1108 ();
 b15zdnd11an1n08x5 FILLER_363_1124 ();
 b15zdnd00an1n01x5 FILLER_363_1132 ();
 b15zdnd11an1n64x5 FILLER_363_1138 ();
 b15zdnd11an1n64x5 FILLER_363_1202 ();
 b15zdnd11an1n08x5 FILLER_363_1266 ();
 b15zdnd11an1n04x5 FILLER_363_1274 ();
 b15zdnd00an1n02x5 FILLER_363_1278 ();
 b15zdnd11an1n04x5 FILLER_363_1298 ();
 b15zdnd11an1n04x5 FILLER_363_1306 ();
 b15zdnd11an1n04x5 FILLER_363_1323 ();
 b15zdnd11an1n64x5 FILLER_363_1339 ();
 b15zdnd11an1n04x5 FILLER_363_1403 ();
 b15zdnd11an1n64x5 FILLER_363_1412 ();
 b15zdnd11an1n08x5 FILLER_363_1476 ();
 b15zdnd00an1n02x5 FILLER_363_1484 ();
 b15zdnd00an1n01x5 FILLER_363_1486 ();
 b15zdnd11an1n32x5 FILLER_363_1494 ();
 b15zdnd11an1n04x5 FILLER_363_1526 ();
 b15zdnd00an1n02x5 FILLER_363_1530 ();
 b15zdnd11an1n64x5 FILLER_363_1542 ();
 b15zdnd11an1n08x5 FILLER_363_1606 ();
 b15zdnd00an1n01x5 FILLER_363_1614 ();
 b15zdnd11an1n04x5 FILLER_363_1621 ();
 b15zdnd11an1n04x5 FILLER_363_1631 ();
 b15zdnd00an1n02x5 FILLER_363_1635 ();
 b15zdnd11an1n64x5 FILLER_363_1658 ();
 b15zdnd11an1n04x5 FILLER_363_1722 ();
 b15zdnd00an1n02x5 FILLER_363_1726 ();
 b15zdnd00an1n01x5 FILLER_363_1728 ();
 b15zdnd11an1n64x5 FILLER_363_1742 ();
 b15zdnd11an1n08x5 FILLER_363_1806 ();
 b15zdnd11an1n04x5 FILLER_363_1814 ();
 b15zdnd11an1n16x5 FILLER_363_1827 ();
 b15zdnd11an1n08x5 FILLER_363_1843 ();
 b15zdnd00an1n02x5 FILLER_363_1851 ();
 b15zdnd00an1n01x5 FILLER_363_1853 ();
 b15zdnd11an1n64x5 FILLER_363_1870 ();
 b15zdnd11an1n08x5 FILLER_363_1934 ();
 b15zdnd11an1n04x5 FILLER_363_1942 ();
 b15zdnd00an1n02x5 FILLER_363_1946 ();
 b15zdnd00an1n01x5 FILLER_363_1948 ();
 b15zdnd11an1n64x5 FILLER_363_1954 ();
 b15zdnd11an1n32x5 FILLER_363_2018 ();
 b15zdnd11an1n16x5 FILLER_363_2050 ();
 b15zdnd11an1n08x5 FILLER_363_2066 ();
 b15zdnd11an1n04x5 FILLER_363_2074 ();
 b15zdnd00an1n02x5 FILLER_363_2078 ();
 b15zdnd00an1n01x5 FILLER_363_2080 ();
 b15zdnd11an1n64x5 FILLER_363_2087 ();
 b15zdnd11an1n64x5 FILLER_363_2151 ();
 b15zdnd11an1n64x5 FILLER_363_2215 ();
 b15zdnd11an1n04x5 FILLER_363_2279 ();
 b15zdnd00an1n01x5 FILLER_363_2283 ();
 b15zdnd11an1n64x5 FILLER_364_8 ();
 b15zdnd11an1n64x5 FILLER_364_72 ();
 b15zdnd11an1n64x5 FILLER_364_136 ();
 b15zdnd11an1n16x5 FILLER_364_200 ();
 b15zdnd11an1n32x5 FILLER_364_247 ();
 b15zdnd11an1n04x5 FILLER_364_279 ();
 b15zdnd11an1n16x5 FILLER_364_292 ();
 b15zdnd11an1n08x5 FILLER_364_308 ();
 b15zdnd11an1n04x5 FILLER_364_316 ();
 b15zdnd00an1n02x5 FILLER_364_320 ();
 b15zdnd11an1n16x5 FILLER_364_327 ();
 b15zdnd11an1n08x5 FILLER_364_343 ();
 b15zdnd11an1n04x5 FILLER_364_351 ();
 b15zdnd00an1n02x5 FILLER_364_355 ();
 b15zdnd00an1n01x5 FILLER_364_357 ();
 b15zdnd11an1n04x5 FILLER_364_378 ();
 b15zdnd11an1n32x5 FILLER_364_389 ();
 b15zdnd11an1n16x5 FILLER_364_421 ();
 b15zdnd11an1n04x5 FILLER_364_437 ();
 b15zdnd00an1n02x5 FILLER_364_441 ();
 b15zdnd11an1n64x5 FILLER_364_449 ();
 b15zdnd11an1n64x5 FILLER_364_513 ();
 b15zdnd11an1n64x5 FILLER_364_577 ();
 b15zdnd00an1n01x5 FILLER_364_641 ();
 b15zdnd11an1n64x5 FILLER_364_648 ();
 b15zdnd11an1n04x5 FILLER_364_712 ();
 b15zdnd00an1n02x5 FILLER_364_716 ();
 b15zdnd11an1n08x5 FILLER_364_726 ();
 b15zdnd11an1n04x5 FILLER_364_734 ();
 b15zdnd00an1n02x5 FILLER_364_738 ();
 b15zdnd00an1n01x5 FILLER_364_740 ();
 b15zdnd11an1n04x5 FILLER_364_751 ();
 b15zdnd11an1n32x5 FILLER_364_767 ();
 b15zdnd11an1n16x5 FILLER_364_799 ();
 b15zdnd11an1n04x5 FILLER_364_815 ();
 b15zdnd00an1n02x5 FILLER_364_819 ();
 b15zdnd11an1n08x5 FILLER_364_842 ();
 b15zdnd11an1n04x5 FILLER_364_850 ();
 b15zdnd00an1n02x5 FILLER_364_854 ();
 b15zdnd00an1n01x5 FILLER_364_856 ();
 b15zdnd11an1n64x5 FILLER_364_869 ();
 b15zdnd11an1n16x5 FILLER_364_933 ();
 b15zdnd11an1n08x5 FILLER_364_949 ();
 b15zdnd11an1n04x5 FILLER_364_957 ();
 b15zdnd00an1n01x5 FILLER_364_961 ();
 b15zdnd11an1n32x5 FILLER_364_974 ();
 b15zdnd00an1n01x5 FILLER_364_1006 ();
 b15zdnd11an1n08x5 FILLER_364_1027 ();
 b15zdnd00an1n02x5 FILLER_364_1035 ();
 b15zdnd11an1n04x5 FILLER_364_1045 ();
 b15zdnd11an1n32x5 FILLER_364_1054 ();
 b15zdnd11an1n16x5 FILLER_364_1086 ();
 b15zdnd11an1n08x5 FILLER_364_1102 ();
 b15zdnd11an1n04x5 FILLER_364_1110 ();
 b15zdnd00an1n02x5 FILLER_364_1114 ();
 b15zdnd11an1n04x5 FILLER_364_1128 ();
 b15zdnd11an1n16x5 FILLER_364_1140 ();
 b15zdnd11an1n04x5 FILLER_364_1156 ();
 b15zdnd00an1n02x5 FILLER_364_1160 ();
 b15zdnd11an1n04x5 FILLER_364_1172 ();
 b15zdnd11an1n04x5 FILLER_364_1183 ();
 b15zdnd00an1n02x5 FILLER_364_1187 ();
 b15zdnd11an1n64x5 FILLER_364_1201 ();
 b15zdnd11an1n32x5 FILLER_364_1265 ();
 b15zdnd11an1n08x5 FILLER_364_1297 ();
 b15zdnd11an1n04x5 FILLER_364_1305 ();
 b15zdnd00an1n01x5 FILLER_364_1309 ();
 b15zdnd11an1n08x5 FILLER_364_1322 ();
 b15zdnd11an1n04x5 FILLER_364_1330 ();
 b15zdnd11an1n16x5 FILLER_364_1341 ();
 b15zdnd11an1n04x5 FILLER_364_1357 ();
 b15zdnd00an1n01x5 FILLER_364_1361 ();
 b15zdnd11an1n16x5 FILLER_364_1366 ();
 b15zdnd11an1n04x5 FILLER_364_1382 ();
 b15zdnd11an1n16x5 FILLER_364_1392 ();
 b15zdnd11an1n04x5 FILLER_364_1415 ();
 b15zdnd00an1n02x5 FILLER_364_1419 ();
 b15zdnd11an1n16x5 FILLER_364_1427 ();
 b15zdnd11an1n08x5 FILLER_364_1443 ();
 b15zdnd11an1n04x5 FILLER_364_1451 ();
 b15zdnd00an1n01x5 FILLER_364_1455 ();
 b15zdnd11an1n16x5 FILLER_364_1463 ();
 b15zdnd11an1n04x5 FILLER_364_1479 ();
 b15zdnd00an1n02x5 FILLER_364_1483 ();
 b15zdnd00an1n01x5 FILLER_364_1485 ();
 b15zdnd11an1n32x5 FILLER_364_1492 ();
 b15zdnd11an1n16x5 FILLER_364_1524 ();
 b15zdnd11an1n04x5 FILLER_364_1540 ();
 b15zdnd00an1n02x5 FILLER_364_1544 ();
 b15zdnd11an1n64x5 FILLER_364_1556 ();
 b15zdnd00an1n02x5 FILLER_364_1620 ();
 b15zdnd00an1n01x5 FILLER_364_1622 ();
 b15zdnd11an1n16x5 FILLER_364_1632 ();
 b15zdnd11an1n08x5 FILLER_364_1648 ();
 b15zdnd11an1n32x5 FILLER_364_1673 ();
 b15zdnd11an1n16x5 FILLER_364_1705 ();
 b15zdnd11an1n04x5 FILLER_364_1721 ();
 b15zdnd00an1n02x5 FILLER_364_1725 ();
 b15zdnd11an1n04x5 FILLER_364_1742 ();
 b15zdnd00an1n02x5 FILLER_364_1746 ();
 b15zdnd11an1n32x5 FILLER_364_1768 ();
 b15zdnd11an1n08x5 FILLER_364_1800 ();
 b15zdnd00an1n01x5 FILLER_364_1808 ();
 b15zdnd11an1n32x5 FILLER_364_1816 ();
 b15zdnd11an1n04x5 FILLER_364_1848 ();
 b15zdnd11an1n04x5 FILLER_364_1860 ();
 b15zdnd00an1n02x5 FILLER_364_1864 ();
 b15zdnd00an1n01x5 FILLER_364_1866 ();
 b15zdnd11an1n08x5 FILLER_364_1873 ();
 b15zdnd11an1n04x5 FILLER_364_1881 ();
 b15zdnd00an1n02x5 FILLER_364_1885 ();
 b15zdnd00an1n01x5 FILLER_364_1887 ();
 b15zdnd11an1n32x5 FILLER_364_1898 ();
 b15zdnd11an1n16x5 FILLER_364_1930 ();
 b15zdnd11an1n04x5 FILLER_364_1946 ();
 b15zdnd11an1n04x5 FILLER_364_1960 ();
 b15zdnd11an1n32x5 FILLER_364_1975 ();
 b15zdnd11an1n04x5 FILLER_364_2007 ();
 b15zdnd00an1n02x5 FILLER_364_2011 ();
 b15zdnd11an1n08x5 FILLER_364_2018 ();
 b15zdnd11an1n04x5 FILLER_364_2026 ();
 b15zdnd00an1n01x5 FILLER_364_2030 ();
 b15zdnd11an1n16x5 FILLER_364_2043 ();
 b15zdnd11an1n04x5 FILLER_364_2059 ();
 b15zdnd11an1n04x5 FILLER_364_2069 ();
 b15zdnd11an1n16x5 FILLER_364_2083 ();
 b15zdnd00an1n02x5 FILLER_364_2099 ();
 b15zdnd11an1n16x5 FILLER_364_2117 ();
 b15zdnd11an1n08x5 FILLER_364_2133 ();
 b15zdnd11an1n04x5 FILLER_364_2141 ();
 b15zdnd00an1n02x5 FILLER_364_2152 ();
 b15zdnd11an1n32x5 FILLER_364_2162 ();
 b15zdnd11an1n08x5 FILLER_364_2194 ();
 b15zdnd00an1n01x5 FILLER_364_2202 ();
 b15zdnd11an1n08x5 FILLER_364_2208 ();
 b15zdnd00an1n01x5 FILLER_364_2216 ();
 b15zdnd11an1n04x5 FILLER_364_2227 ();
 b15zdnd11an1n32x5 FILLER_364_2237 ();
 b15zdnd11an1n04x5 FILLER_364_2269 ();
 b15zdnd00an1n02x5 FILLER_364_2273 ();
 b15zdnd00an1n01x5 FILLER_364_2275 ();
 b15zdnd11an1n64x5 FILLER_365_0 ();
 b15zdnd11an1n64x5 FILLER_365_64 ();
 b15zdnd11an1n64x5 FILLER_365_128 ();
 b15zdnd11an1n32x5 FILLER_365_192 ();
 b15zdnd11an1n04x5 FILLER_365_224 ();
 b15zdnd11an1n08x5 FILLER_365_237 ();
 b15zdnd11an1n04x5 FILLER_365_245 ();
 b15zdnd00an1n01x5 FILLER_365_249 ();
 b15zdnd11an1n08x5 FILLER_365_255 ();
 b15zdnd11an1n04x5 FILLER_365_263 ();
 b15zdnd00an1n01x5 FILLER_365_267 ();
 b15zdnd11an1n16x5 FILLER_365_275 ();
 b15zdnd11an1n04x5 FILLER_365_296 ();
 b15zdnd11an1n04x5 FILLER_365_307 ();
 b15zdnd11an1n04x5 FILLER_365_316 ();
 b15zdnd11an1n32x5 FILLER_365_324 ();
 b15zdnd11an1n16x5 FILLER_365_356 ();
 b15zdnd11an1n08x5 FILLER_365_372 ();
 b15zdnd11an1n04x5 FILLER_365_380 ();
 b15zdnd11an1n16x5 FILLER_365_389 ();
 b15zdnd00an1n01x5 FILLER_365_405 ();
 b15zdnd11an1n32x5 FILLER_365_412 ();
 b15zdnd11an1n32x5 FILLER_365_460 ();
 b15zdnd11an1n04x5 FILLER_365_492 ();
 b15zdnd00an1n02x5 FILLER_365_496 ();
 b15zdnd11an1n04x5 FILLER_365_503 ();
 b15zdnd11an1n08x5 FILLER_365_511 ();
 b15zdnd00an1n01x5 FILLER_365_519 ();
 b15zdnd11an1n04x5 FILLER_365_533 ();
 b15zdnd11an1n04x5 FILLER_365_541 ();
 b15zdnd00an1n02x5 FILLER_365_545 ();
 b15zdnd00an1n01x5 FILLER_365_547 ();
 b15zdnd11an1n16x5 FILLER_365_552 ();
 b15zdnd11an1n64x5 FILLER_365_582 ();
 b15zdnd11an1n32x5 FILLER_365_646 ();
 b15zdnd11an1n16x5 FILLER_365_678 ();
 b15zdnd11an1n08x5 FILLER_365_694 ();
 b15zdnd11an1n04x5 FILLER_365_702 ();
 b15zdnd11an1n16x5 FILLER_365_725 ();
 b15zdnd11an1n04x5 FILLER_365_741 ();
 b15zdnd00an1n02x5 FILLER_365_745 ();
 b15zdnd11an1n08x5 FILLER_365_768 ();
 b15zdnd00an1n01x5 FILLER_365_776 ();
 b15zdnd11an1n08x5 FILLER_365_790 ();
 b15zdnd00an1n02x5 FILLER_365_798 ();
 b15zdnd11an1n64x5 FILLER_365_804 ();
 b15zdnd11an1n08x5 FILLER_365_868 ();
 b15zdnd11an1n04x5 FILLER_365_876 ();
 b15zdnd00an1n01x5 FILLER_365_880 ();
 b15zdnd11an1n32x5 FILLER_365_886 ();
 b15zdnd11an1n04x5 FILLER_365_918 ();
 b15zdnd11an1n32x5 FILLER_365_931 ();
 b15zdnd00an1n02x5 FILLER_365_963 ();
 b15zdnd00an1n01x5 FILLER_365_965 ();
 b15zdnd11an1n04x5 FILLER_365_972 ();
 b15zdnd11an1n16x5 FILLER_365_982 ();
 b15zdnd11an1n04x5 FILLER_365_998 ();
 b15zdnd00an1n01x5 FILLER_365_1002 ();
 b15zdnd11an1n64x5 FILLER_365_1010 ();
 b15zdnd11an1n32x5 FILLER_365_1074 ();
 b15zdnd11an1n08x5 FILLER_365_1106 ();
 b15zdnd11an1n04x5 FILLER_365_1114 ();
 b15zdnd00an1n02x5 FILLER_365_1118 ();
 b15zdnd11an1n16x5 FILLER_365_1134 ();
 b15zdnd11an1n08x5 FILLER_365_1150 ();
 b15zdnd00an1n02x5 FILLER_365_1158 ();
 b15zdnd11an1n64x5 FILLER_365_1180 ();
 b15zdnd11an1n64x5 FILLER_365_1244 ();
 b15zdnd11an1n16x5 FILLER_365_1334 ();
 b15zdnd11an1n04x5 FILLER_365_1350 ();
 b15zdnd00an1n02x5 FILLER_365_1354 ();
 b15zdnd11an1n16x5 FILLER_365_1370 ();
 b15zdnd11an1n04x5 FILLER_365_1386 ();
 b15zdnd11an1n16x5 FILLER_365_1394 ();
 b15zdnd11an1n04x5 FILLER_365_1410 ();
 b15zdnd00an1n02x5 FILLER_365_1414 ();
 b15zdnd11an1n16x5 FILLER_365_1422 ();
 b15zdnd11an1n08x5 FILLER_365_1438 ();
 b15zdnd11an1n04x5 FILLER_365_1446 ();
 b15zdnd11an1n64x5 FILLER_365_1461 ();
 b15zdnd11an1n16x5 FILLER_365_1525 ();
 b15zdnd11an1n04x5 FILLER_365_1541 ();
 b15zdnd11an1n32x5 FILLER_365_1554 ();
 b15zdnd11an1n04x5 FILLER_365_1586 ();
 b15zdnd11an1n04x5 FILLER_365_1595 ();
 b15zdnd11an1n16x5 FILLER_365_1605 ();
 b15zdnd11an1n08x5 FILLER_365_1621 ();
 b15zdnd00an1n01x5 FILLER_365_1629 ();
 b15zdnd11an1n08x5 FILLER_365_1646 ();
 b15zdnd00an1n01x5 FILLER_365_1654 ();
 b15zdnd11an1n16x5 FILLER_365_1681 ();
 b15zdnd11an1n08x5 FILLER_365_1707 ();
 b15zdnd00an1n01x5 FILLER_365_1715 ();
 b15zdnd11an1n64x5 FILLER_365_1732 ();
 b15zdnd11an1n16x5 FILLER_365_1796 ();
 b15zdnd11an1n04x5 FILLER_365_1812 ();
 b15zdnd11an1n08x5 FILLER_365_1824 ();
 b15zdnd11an1n04x5 FILLER_365_1832 ();
 b15zdnd00an1n01x5 FILLER_365_1836 ();
 b15zdnd11an1n04x5 FILLER_365_1841 ();
 b15zdnd11an1n04x5 FILLER_365_1852 ();
 b15zdnd00an1n01x5 FILLER_365_1856 ();
 b15zdnd11an1n64x5 FILLER_365_1862 ();
 b15zdnd11an1n04x5 FILLER_365_1926 ();
 b15zdnd11an1n16x5 FILLER_365_1935 ();
 b15zdnd00an1n01x5 FILLER_365_1951 ();
 b15zdnd11an1n16x5 FILLER_365_1957 ();
 b15zdnd11an1n08x5 FILLER_365_1973 ();
 b15zdnd00an1n01x5 FILLER_365_1981 ();
 b15zdnd11an1n16x5 FILLER_365_1988 ();
 b15zdnd00an1n02x5 FILLER_365_2004 ();
 b15zdnd00an1n01x5 FILLER_365_2006 ();
 b15zdnd11an1n04x5 FILLER_365_2022 ();
 b15zdnd11an1n32x5 FILLER_365_2038 ();
 b15zdnd11an1n16x5 FILLER_365_2070 ();
 b15zdnd11an1n08x5 FILLER_365_2086 ();
 b15zdnd11an1n04x5 FILLER_365_2094 ();
 b15zdnd00an1n02x5 FILLER_365_2098 ();
 b15zdnd00an1n01x5 FILLER_365_2100 ();
 b15zdnd11an1n64x5 FILLER_365_2110 ();
 b15zdnd11an1n16x5 FILLER_365_2174 ();
 b15zdnd00an1n02x5 FILLER_365_2190 ();
 b15zdnd00an1n01x5 FILLER_365_2192 ();
 b15zdnd11an1n04x5 FILLER_365_2199 ();
 b15zdnd11an1n08x5 FILLER_365_2213 ();
 b15zdnd11an1n04x5 FILLER_365_2221 ();
 b15zdnd00an1n01x5 FILLER_365_2225 ();
 b15zdnd11an1n32x5 FILLER_365_2246 ();
 b15zdnd11an1n04x5 FILLER_365_2278 ();
 b15zdnd00an1n02x5 FILLER_365_2282 ();
 b15zdnd11an1n64x5 FILLER_366_8 ();
 b15zdnd11an1n64x5 FILLER_366_72 ();
 b15zdnd11an1n64x5 FILLER_366_136 ();
 b15zdnd11an1n32x5 FILLER_366_200 ();
 b15zdnd00an1n02x5 FILLER_366_232 ();
 b15zdnd00an1n01x5 FILLER_366_234 ();
 b15zdnd11an1n04x5 FILLER_366_252 ();
 b15zdnd11an1n64x5 FILLER_366_260 ();
 b15zdnd11an1n32x5 FILLER_366_324 ();
 b15zdnd11an1n16x5 FILLER_366_356 ();
 b15zdnd11an1n08x5 FILLER_366_372 ();
 b15zdnd00an1n02x5 FILLER_366_380 ();
 b15zdnd11an1n16x5 FILLER_366_394 ();
 b15zdnd11an1n64x5 FILLER_366_422 ();
 b15zdnd11an1n04x5 FILLER_366_486 ();
 b15zdnd00an1n02x5 FILLER_366_490 ();
 b15zdnd00an1n01x5 FILLER_366_492 ();
 b15zdnd11an1n32x5 FILLER_366_498 ();
 b15zdnd11an1n04x5 FILLER_366_530 ();
 b15zdnd00an1n01x5 FILLER_366_534 ();
 b15zdnd11an1n32x5 FILLER_366_561 ();
 b15zdnd00an1n02x5 FILLER_366_593 ();
 b15zdnd11an1n16x5 FILLER_366_627 ();
 b15zdnd11an1n04x5 FILLER_366_650 ();
 b15zdnd11an1n04x5 FILLER_366_659 ();
 b15zdnd00an1n02x5 FILLER_366_663 ();
 b15zdnd11an1n32x5 FILLER_366_675 ();
 b15zdnd11an1n08x5 FILLER_366_707 ();
 b15zdnd00an1n02x5 FILLER_366_715 ();
 b15zdnd00an1n01x5 FILLER_366_717 ();
 b15zdnd11an1n64x5 FILLER_366_726 ();
 b15zdnd11an1n32x5 FILLER_366_790 ();
 b15zdnd11an1n04x5 FILLER_366_822 ();
 b15zdnd00an1n02x5 FILLER_366_826 ();
 b15zdnd11an1n64x5 FILLER_366_832 ();
 b15zdnd11an1n64x5 FILLER_366_896 ();
 b15zdnd11an1n08x5 FILLER_366_960 ();
 b15zdnd11an1n64x5 FILLER_366_974 ();
 b15zdnd00an1n01x5 FILLER_366_1038 ();
 b15zdnd11an1n16x5 FILLER_366_1047 ();
 b15zdnd00an1n01x5 FILLER_366_1063 ();
 b15zdnd11an1n04x5 FILLER_366_1072 ();
 b15zdnd11an1n64x5 FILLER_366_1083 ();
 b15zdnd00an1n02x5 FILLER_366_1147 ();
 b15zdnd11an1n04x5 FILLER_366_1157 ();
 b15zdnd11an1n08x5 FILLER_366_1168 ();
 b15zdnd11an1n04x5 FILLER_366_1176 ();
 b15zdnd00an1n02x5 FILLER_366_1180 ();
 b15zdnd00an1n01x5 FILLER_366_1182 ();
 b15zdnd11an1n64x5 FILLER_366_1192 ();
 b15zdnd11an1n64x5 FILLER_366_1256 ();
 b15zdnd11an1n04x5 FILLER_366_1328 ();
 b15zdnd00an1n02x5 FILLER_366_1332 ();
 b15zdnd11an1n04x5 FILLER_366_1350 ();
 b15zdnd11an1n32x5 FILLER_366_1368 ();
 b15zdnd00an1n02x5 FILLER_366_1400 ();
 b15zdnd00an1n01x5 FILLER_366_1402 ();
 b15zdnd11an1n04x5 FILLER_366_1410 ();
 b15zdnd11an1n16x5 FILLER_366_1430 ();
 b15zdnd00an1n02x5 FILLER_366_1446 ();
 b15zdnd11an1n04x5 FILLER_366_1453 ();
 b15zdnd11an1n16x5 FILLER_366_1464 ();
 b15zdnd11an1n08x5 FILLER_366_1480 ();
 b15zdnd11an1n04x5 FILLER_366_1488 ();
 b15zdnd00an1n01x5 FILLER_366_1492 ();
 b15zdnd11an1n04x5 FILLER_366_1501 ();
 b15zdnd11an1n08x5 FILLER_366_1511 ();
 b15zdnd11an1n04x5 FILLER_366_1519 ();
 b15zdnd11an1n04x5 FILLER_366_1533 ();
 b15zdnd11an1n04x5 FILLER_366_1541 ();
 b15zdnd11an1n04x5 FILLER_366_1550 ();
 b15zdnd11an1n16x5 FILLER_366_1560 ();
 b15zdnd00an1n02x5 FILLER_366_1576 ();
 b15zdnd00an1n01x5 FILLER_366_1578 ();
 b15zdnd11an1n04x5 FILLER_366_1591 ();
 b15zdnd11an1n04x5 FILLER_366_1602 ();
 b15zdnd11an1n16x5 FILLER_366_1610 ();
 b15zdnd11an1n04x5 FILLER_366_1626 ();
 b15zdnd00an1n02x5 FILLER_366_1630 ();
 b15zdnd11an1n16x5 FILLER_366_1638 ();
 b15zdnd11an1n08x5 FILLER_366_1654 ();
 b15zdnd11an1n04x5 FILLER_366_1662 ();
 b15zdnd00an1n02x5 FILLER_366_1666 ();
 b15zdnd00an1n01x5 FILLER_366_1668 ();
 b15zdnd11an1n64x5 FILLER_366_1675 ();
 b15zdnd11an1n64x5 FILLER_366_1739 ();
 b15zdnd11an1n32x5 FILLER_366_1803 ();
 b15zdnd11an1n08x5 FILLER_366_1835 ();
 b15zdnd00an1n02x5 FILLER_366_1843 ();
 b15zdnd00an1n01x5 FILLER_366_1845 ();
 b15zdnd11an1n16x5 FILLER_366_1858 ();
 b15zdnd00an1n02x5 FILLER_366_1874 ();
 b15zdnd11an1n16x5 FILLER_366_1881 ();
 b15zdnd11an1n04x5 FILLER_366_1897 ();
 b15zdnd00an1n01x5 FILLER_366_1901 ();
 b15zdnd11an1n08x5 FILLER_366_1912 ();
 b15zdnd00an1n02x5 FILLER_366_1920 ();
 b15zdnd11an1n08x5 FILLER_366_1934 ();
 b15zdnd00an1n01x5 FILLER_366_1942 ();
 b15zdnd11an1n04x5 FILLER_366_1948 ();
 b15zdnd11an1n04x5 FILLER_366_1961 ();
 b15zdnd11an1n64x5 FILLER_366_1970 ();
 b15zdnd11an1n64x5 FILLER_366_2034 ();
 b15zdnd11an1n04x5 FILLER_366_2098 ();
 b15zdnd00an1n01x5 FILLER_366_2102 ();
 b15zdnd11an1n04x5 FILLER_366_2109 ();
 b15zdnd11an1n04x5 FILLER_366_2121 ();
 b15zdnd11an1n04x5 FILLER_366_2136 ();
 b15zdnd00an1n02x5 FILLER_366_2152 ();
 b15zdnd00an1n02x5 FILLER_366_2162 ();
 b15zdnd11an1n08x5 FILLER_366_2168 ();
 b15zdnd11an1n04x5 FILLER_366_2176 ();
 b15zdnd00an1n02x5 FILLER_366_2180 ();
 b15zdnd11an1n04x5 FILLER_366_2198 ();
 b15zdnd00an1n02x5 FILLER_366_2202 ();
 b15zdnd00an1n01x5 FILLER_366_2204 ();
 b15zdnd11an1n04x5 FILLER_366_2212 ();
 b15zdnd00an1n01x5 FILLER_366_2216 ();
 b15zdnd11an1n32x5 FILLER_366_2222 ();
 b15zdnd11an1n16x5 FILLER_366_2254 ();
 b15zdnd11an1n04x5 FILLER_366_2270 ();
 b15zdnd00an1n02x5 FILLER_366_2274 ();
 b15zdnd11an1n64x5 FILLER_367_0 ();
 b15zdnd11an1n64x5 FILLER_367_64 ();
 b15zdnd11an1n64x5 FILLER_367_128 ();
 b15zdnd11an1n16x5 FILLER_367_192 ();
 b15zdnd11an1n04x5 FILLER_367_208 ();
 b15zdnd11an1n64x5 FILLER_367_230 ();
 b15zdnd11an1n64x5 FILLER_367_294 ();
 b15zdnd11an1n64x5 FILLER_367_358 ();
 b15zdnd11an1n32x5 FILLER_367_422 ();
 b15zdnd11an1n08x5 FILLER_367_454 ();
 b15zdnd11an1n04x5 FILLER_367_462 ();
 b15zdnd00an1n02x5 FILLER_367_466 ();
 b15zdnd11an1n08x5 FILLER_367_472 ();
 b15zdnd00an1n01x5 FILLER_367_480 ();
 b15zdnd11an1n08x5 FILLER_367_488 ();
 b15zdnd00an1n02x5 FILLER_367_496 ();
 b15zdnd00an1n01x5 FILLER_367_498 ();
 b15zdnd11an1n32x5 FILLER_367_506 ();
 b15zdnd11an1n08x5 FILLER_367_538 ();
 b15zdnd11an1n04x5 FILLER_367_546 ();
 b15zdnd00an1n02x5 FILLER_367_550 ();
 b15zdnd00an1n01x5 FILLER_367_552 ();
 b15zdnd11an1n64x5 FILLER_367_558 ();
 b15zdnd11an1n16x5 FILLER_367_622 ();
 b15zdnd11an1n16x5 FILLER_367_643 ();
 b15zdnd00an1n02x5 FILLER_367_659 ();
 b15zdnd00an1n01x5 FILLER_367_661 ();
 b15zdnd11an1n08x5 FILLER_367_667 ();
 b15zdnd11an1n04x5 FILLER_367_685 ();
 b15zdnd11an1n04x5 FILLER_367_705 ();
 b15zdnd11an1n64x5 FILLER_367_714 ();
 b15zdnd11an1n08x5 FILLER_367_778 ();
 b15zdnd11an1n04x5 FILLER_367_786 ();
 b15zdnd00an1n02x5 FILLER_367_790 ();
 b15zdnd00an1n01x5 FILLER_367_792 ();
 b15zdnd11an1n16x5 FILLER_367_805 ();
 b15zdnd11an1n04x5 FILLER_367_821 ();
 b15zdnd00an1n02x5 FILLER_367_825 ();
 b15zdnd11an1n08x5 FILLER_367_836 ();
 b15zdnd11an1n04x5 FILLER_367_858 ();
 b15zdnd11an1n16x5 FILLER_367_867 ();
 b15zdnd11an1n04x5 FILLER_367_883 ();
 b15zdnd00an1n01x5 FILLER_367_887 ();
 b15zdnd11an1n04x5 FILLER_367_900 ();
 b15zdnd11an1n04x5 FILLER_367_910 ();
 b15zdnd00an1n01x5 FILLER_367_914 ();
 b15zdnd11an1n04x5 FILLER_367_925 ();
 b15zdnd11an1n64x5 FILLER_367_942 ();
 b15zdnd11an1n16x5 FILLER_367_1012 ();
 b15zdnd11an1n04x5 FILLER_367_1039 ();
 b15zdnd00an1n02x5 FILLER_367_1043 ();
 b15zdnd11an1n16x5 FILLER_367_1049 ();
 b15zdnd11an1n08x5 FILLER_367_1065 ();
 b15zdnd11an1n04x5 FILLER_367_1073 ();
 b15zdnd11an1n08x5 FILLER_367_1102 ();
 b15zdnd00an1n02x5 FILLER_367_1110 ();
 b15zdnd11an1n32x5 FILLER_367_1119 ();
 b15zdnd11an1n16x5 FILLER_367_1151 ();
 b15zdnd11an1n08x5 FILLER_367_1175 ();
 b15zdnd11an1n04x5 FILLER_367_1183 ();
 b15zdnd00an1n01x5 FILLER_367_1187 ();
 b15zdnd11an1n64x5 FILLER_367_1196 ();
 b15zdnd11an1n32x5 FILLER_367_1260 ();
 b15zdnd11an1n16x5 FILLER_367_1292 ();
 b15zdnd11an1n08x5 FILLER_367_1308 ();
 b15zdnd00an1n02x5 FILLER_367_1316 ();
 b15zdnd11an1n04x5 FILLER_367_1325 ();
 b15zdnd00an1n02x5 FILLER_367_1329 ();
 b15zdnd11an1n32x5 FILLER_367_1344 ();
 b15zdnd11an1n16x5 FILLER_367_1376 ();
 b15zdnd11an1n04x5 FILLER_367_1392 ();
 b15zdnd00an1n02x5 FILLER_367_1396 ();
 b15zdnd11an1n32x5 FILLER_367_1406 ();
 b15zdnd11an1n16x5 FILLER_367_1438 ();
 b15zdnd00an1n02x5 FILLER_367_1454 ();
 b15zdnd00an1n01x5 FILLER_367_1456 ();
 b15zdnd11an1n04x5 FILLER_367_1462 ();
 b15zdnd11an1n08x5 FILLER_367_1472 ();
 b15zdnd11an1n04x5 FILLER_367_1480 ();
 b15zdnd00an1n01x5 FILLER_367_1484 ();
 b15zdnd11an1n08x5 FILLER_367_1495 ();
 b15zdnd00an1n01x5 FILLER_367_1503 ();
 b15zdnd11an1n64x5 FILLER_367_1511 ();
 b15zdnd11an1n64x5 FILLER_367_1575 ();
 b15zdnd11an1n64x5 FILLER_367_1639 ();
 b15zdnd11an1n16x5 FILLER_367_1703 ();
 b15zdnd11an1n08x5 FILLER_367_1719 ();
 b15zdnd11an1n04x5 FILLER_367_1727 ();
 b15zdnd00an1n01x5 FILLER_367_1731 ();
 b15zdnd11an1n64x5 FILLER_367_1742 ();
 b15zdnd11an1n04x5 FILLER_367_1806 ();
 b15zdnd00an1n02x5 FILLER_367_1810 ();
 b15zdnd00an1n01x5 FILLER_367_1812 ();
 b15zdnd11an1n32x5 FILLER_367_1818 ();
 b15zdnd11an1n32x5 FILLER_367_1860 ();
 b15zdnd11an1n16x5 FILLER_367_1892 ();
 b15zdnd11an1n08x5 FILLER_367_1908 ();
 b15zdnd00an1n02x5 FILLER_367_1916 ();
 b15zdnd11an1n32x5 FILLER_367_1928 ();
 b15zdnd11an1n16x5 FILLER_367_1960 ();
 b15zdnd11an1n16x5 FILLER_367_1981 ();
 b15zdnd11an1n08x5 FILLER_367_1997 ();
 b15zdnd11an1n16x5 FILLER_367_2015 ();
 b15zdnd11an1n04x5 FILLER_367_2031 ();
 b15zdnd11an1n16x5 FILLER_367_2042 ();
 b15zdnd11an1n08x5 FILLER_367_2058 ();
 b15zdnd11an1n04x5 FILLER_367_2066 ();
 b15zdnd00an1n01x5 FILLER_367_2070 ();
 b15zdnd11an1n32x5 FILLER_367_2077 ();
 b15zdnd11an1n16x5 FILLER_367_2109 ();
 b15zdnd11an1n04x5 FILLER_367_2125 ();
 b15zdnd11an1n08x5 FILLER_367_2134 ();
 b15zdnd00an1n01x5 FILLER_367_2142 ();
 b15zdnd11an1n64x5 FILLER_367_2147 ();
 b15zdnd11an1n64x5 FILLER_367_2217 ();
 b15zdnd00an1n02x5 FILLER_367_2281 ();
 b15zdnd00an1n01x5 FILLER_367_2283 ();
 b15zdnd11an1n64x5 FILLER_368_8 ();
 b15zdnd11an1n64x5 FILLER_368_72 ();
 b15zdnd11an1n64x5 FILLER_368_136 ();
 b15zdnd11an1n16x5 FILLER_368_200 ();
 b15zdnd11an1n08x5 FILLER_368_216 ();
 b15zdnd00an1n01x5 FILLER_368_224 ();
 b15zdnd11an1n16x5 FILLER_368_241 ();
 b15zdnd11an1n64x5 FILLER_368_273 ();
 b15zdnd11an1n16x5 FILLER_368_337 ();
 b15zdnd11an1n32x5 FILLER_368_363 ();
 b15zdnd11an1n16x5 FILLER_368_395 ();
 b15zdnd11an1n08x5 FILLER_368_411 ();
 b15zdnd11an1n16x5 FILLER_368_428 ();
 b15zdnd11an1n08x5 FILLER_368_444 ();
 b15zdnd11an1n04x5 FILLER_368_452 ();
 b15zdnd11an1n16x5 FILLER_368_463 ();
 b15zdnd11an1n08x5 FILLER_368_479 ();
 b15zdnd00an1n01x5 FILLER_368_487 ();
 b15zdnd11an1n32x5 FILLER_368_494 ();
 b15zdnd11an1n16x5 FILLER_368_526 ();
 b15zdnd11an1n08x5 FILLER_368_542 ();
 b15zdnd11an1n04x5 FILLER_368_550 ();
 b15zdnd00an1n02x5 FILLER_368_554 ();
 b15zdnd11an1n64x5 FILLER_368_569 ();
 b15zdnd11an1n32x5 FILLER_368_633 ();
 b15zdnd11an1n16x5 FILLER_368_665 ();
 b15zdnd11an1n08x5 FILLER_368_681 ();
 b15zdnd11an1n04x5 FILLER_368_689 ();
 b15zdnd00an1n01x5 FILLER_368_693 ();
 b15zdnd11an1n08x5 FILLER_368_705 ();
 b15zdnd11an1n04x5 FILLER_368_713 ();
 b15zdnd00an1n01x5 FILLER_368_717 ();
 b15zdnd11an1n04x5 FILLER_368_726 ();
 b15zdnd00an1n02x5 FILLER_368_730 ();
 b15zdnd11an1n16x5 FILLER_368_737 ();
 b15zdnd00an1n02x5 FILLER_368_753 ();
 b15zdnd00an1n01x5 FILLER_368_755 ();
 b15zdnd11an1n04x5 FILLER_368_787 ();
 b15zdnd11an1n32x5 FILLER_368_799 ();
 b15zdnd11an1n16x5 FILLER_368_831 ();
 b15zdnd11an1n08x5 FILLER_368_847 ();
 b15zdnd11an1n04x5 FILLER_368_855 ();
 b15zdnd00an1n01x5 FILLER_368_859 ();
 b15zdnd11an1n04x5 FILLER_368_872 ();
 b15zdnd11an1n04x5 FILLER_368_897 ();
 b15zdnd11an1n16x5 FILLER_368_912 ();
 b15zdnd11an1n04x5 FILLER_368_928 ();
 b15zdnd00an1n02x5 FILLER_368_932 ();
 b15zdnd00an1n01x5 FILLER_368_934 ();
 b15zdnd11an1n08x5 FILLER_368_949 ();
 b15zdnd11an1n04x5 FILLER_368_963 ();
 b15zdnd11an1n32x5 FILLER_368_972 ();
 b15zdnd00an1n01x5 FILLER_368_1004 ();
 b15zdnd11an1n64x5 FILLER_368_1010 ();
 b15zdnd00an1n02x5 FILLER_368_1074 ();
 b15zdnd11an1n04x5 FILLER_368_1086 ();
 b15zdnd00an1n02x5 FILLER_368_1090 ();
 b15zdnd11an1n08x5 FILLER_368_1108 ();
 b15zdnd11an1n32x5 FILLER_368_1128 ();
 b15zdnd11an1n08x5 FILLER_368_1160 ();
 b15zdnd00an1n01x5 FILLER_368_1168 ();
 b15zdnd11an1n04x5 FILLER_368_1181 ();
 b15zdnd00an1n01x5 FILLER_368_1185 ();
 b15zdnd11an1n04x5 FILLER_368_1198 ();
 b15zdnd11an1n64x5 FILLER_368_1207 ();
 b15zdnd11an1n08x5 FILLER_368_1271 ();
 b15zdnd00an1n02x5 FILLER_368_1279 ();
 b15zdnd11an1n04x5 FILLER_368_1297 ();
 b15zdnd11an1n16x5 FILLER_368_1309 ();
 b15zdnd11an1n04x5 FILLER_368_1325 ();
 b15zdnd00an1n02x5 FILLER_368_1329 ();
 b15zdnd11an1n32x5 FILLER_368_1337 ();
 b15zdnd11an1n04x5 FILLER_368_1369 ();
 b15zdnd00an1n02x5 FILLER_368_1373 ();
 b15zdnd00an1n01x5 FILLER_368_1375 ();
 b15zdnd11an1n04x5 FILLER_368_1385 ();
 b15zdnd11an1n64x5 FILLER_368_1393 ();
 b15zdnd11an1n64x5 FILLER_368_1457 ();
 b15zdnd11an1n64x5 FILLER_368_1521 ();
 b15zdnd11an1n64x5 FILLER_368_1585 ();
 b15zdnd11an1n32x5 FILLER_368_1649 ();
 b15zdnd11an1n08x5 FILLER_368_1681 ();
 b15zdnd00an1n02x5 FILLER_368_1689 ();
 b15zdnd11an1n08x5 FILLER_368_1707 ();
 b15zdnd00an1n02x5 FILLER_368_1715 ();
 b15zdnd00an1n01x5 FILLER_368_1717 ();
 b15zdnd11an1n64x5 FILLER_368_1739 ();
 b15zdnd11an1n64x5 FILLER_368_1803 ();
 b15zdnd11an1n32x5 FILLER_368_1867 ();
 b15zdnd11an1n08x5 FILLER_368_1899 ();
 b15zdnd11an1n04x5 FILLER_368_1907 ();
 b15zdnd00an1n01x5 FILLER_368_1911 ();
 b15zdnd11an1n04x5 FILLER_368_1922 ();
 b15zdnd11an1n64x5 FILLER_368_1931 ();
 b15zdnd11an1n32x5 FILLER_368_1995 ();
 b15zdnd11an1n08x5 FILLER_368_2027 ();
 b15zdnd11an1n08x5 FILLER_368_2041 ();
 b15zdnd11an1n04x5 FILLER_368_2049 ();
 b15zdnd00an1n02x5 FILLER_368_2053 ();
 b15zdnd00an1n01x5 FILLER_368_2055 ();
 b15zdnd11an1n04x5 FILLER_368_2062 ();
 b15zdnd11an1n64x5 FILLER_368_2070 ();
 b15zdnd11an1n16x5 FILLER_368_2134 ();
 b15zdnd11an1n04x5 FILLER_368_2150 ();
 b15zdnd11an1n32x5 FILLER_368_2162 ();
 b15zdnd11an1n04x5 FILLER_368_2210 ();
 b15zdnd11an1n32x5 FILLER_368_2225 ();
 b15zdnd11an1n16x5 FILLER_368_2257 ();
 b15zdnd00an1n02x5 FILLER_368_2273 ();
 b15zdnd00an1n01x5 FILLER_368_2275 ();
 b15zdnd11an1n64x5 FILLER_369_0 ();
 b15zdnd11an1n64x5 FILLER_369_64 ();
 b15zdnd11an1n64x5 FILLER_369_128 ();
 b15zdnd11an1n16x5 FILLER_369_192 ();
 b15zdnd11an1n04x5 FILLER_369_208 ();
 b15zdnd00an1n01x5 FILLER_369_212 ();
 b15zdnd11an1n32x5 FILLER_369_238 ();
 b15zdnd11an1n04x5 FILLER_369_270 ();
 b15zdnd00an1n01x5 FILLER_369_274 ();
 b15zdnd11an1n16x5 FILLER_369_298 ();
 b15zdnd11an1n08x5 FILLER_369_326 ();
 b15zdnd11an1n04x5 FILLER_369_362 ();
 b15zdnd00an1n02x5 FILLER_369_366 ();
 b15zdnd00an1n01x5 FILLER_369_368 ();
 b15zdnd11an1n16x5 FILLER_369_383 ();
 b15zdnd00an1n02x5 FILLER_369_399 ();
 b15zdnd11an1n04x5 FILLER_369_413 ();
 b15zdnd00an1n01x5 FILLER_369_417 ();
 b15zdnd11an1n16x5 FILLER_369_424 ();
 b15zdnd11an1n08x5 FILLER_369_440 ();
 b15zdnd00an1n02x5 FILLER_369_448 ();
 b15zdnd00an1n01x5 FILLER_369_450 ();
 b15zdnd11an1n64x5 FILLER_369_464 ();
 b15zdnd11an1n16x5 FILLER_369_528 ();
 b15zdnd11an1n64x5 FILLER_369_562 ();
 b15zdnd11an1n16x5 FILLER_369_626 ();
 b15zdnd11an1n08x5 FILLER_369_642 ();
 b15zdnd00an1n02x5 FILLER_369_650 ();
 b15zdnd00an1n01x5 FILLER_369_652 ();
 b15zdnd11an1n16x5 FILLER_369_657 ();
 b15zdnd11an1n04x5 FILLER_369_673 ();
 b15zdnd00an1n02x5 FILLER_369_677 ();
 b15zdnd00an1n01x5 FILLER_369_679 ();
 b15zdnd11an1n08x5 FILLER_369_692 ();
 b15zdnd11an1n16x5 FILLER_369_706 ();
 b15zdnd11an1n08x5 FILLER_369_722 ();
 b15zdnd11an1n16x5 FILLER_369_737 ();
 b15zdnd00an1n02x5 FILLER_369_753 ();
 b15zdnd11an1n16x5 FILLER_369_768 ();
 b15zdnd11an1n04x5 FILLER_369_784 ();
 b15zdnd00an1n01x5 FILLER_369_788 ();
 b15zdnd11an1n64x5 FILLER_369_810 ();
 b15zdnd11an1n64x5 FILLER_369_874 ();
 b15zdnd11an1n64x5 FILLER_369_938 ();
 b15zdnd11an1n08x5 FILLER_369_1002 ();
 b15zdnd11an1n04x5 FILLER_369_1010 ();
 b15zdnd00an1n02x5 FILLER_369_1014 ();
 b15zdnd00an1n01x5 FILLER_369_1016 ();
 b15zdnd11an1n32x5 FILLER_369_1025 ();
 b15zdnd11an1n08x5 FILLER_369_1057 ();
 b15zdnd11an1n04x5 FILLER_369_1065 ();
 b15zdnd00an1n02x5 FILLER_369_1069 ();
 b15zdnd00an1n01x5 FILLER_369_1071 ();
 b15zdnd11an1n16x5 FILLER_369_1080 ();
 b15zdnd00an1n02x5 FILLER_369_1096 ();
 b15zdnd11an1n16x5 FILLER_369_1110 ();
 b15zdnd11an1n08x5 FILLER_369_1126 ();
 b15zdnd00an1n01x5 FILLER_369_1134 ();
 b15zdnd11an1n32x5 FILLER_369_1139 ();
 b15zdnd11an1n16x5 FILLER_369_1171 ();
 b15zdnd11an1n04x5 FILLER_369_1187 ();
 b15zdnd11an1n64x5 FILLER_369_1198 ();
 b15zdnd11an1n64x5 FILLER_369_1262 ();
 b15zdnd11an1n32x5 FILLER_369_1326 ();
 b15zdnd11an1n16x5 FILLER_369_1358 ();
 b15zdnd11an1n08x5 FILLER_369_1374 ();
 b15zdnd11an1n04x5 FILLER_369_1382 ();
 b15zdnd11an1n16x5 FILLER_369_1400 ();
 b15zdnd00an1n02x5 FILLER_369_1416 ();
 b15zdnd00an1n01x5 FILLER_369_1418 ();
 b15zdnd11an1n64x5 FILLER_369_1434 ();
 b15zdnd11an1n08x5 FILLER_369_1498 ();
 b15zdnd11an1n04x5 FILLER_369_1506 ();
 b15zdnd11an1n64x5 FILLER_369_1519 ();
 b15zdnd11an1n32x5 FILLER_369_1583 ();
 b15zdnd11an1n04x5 FILLER_369_1615 ();
 b15zdnd00an1n01x5 FILLER_369_1619 ();
 b15zdnd11an1n04x5 FILLER_369_1630 ();
 b15zdnd00an1n01x5 FILLER_369_1634 ();
 b15zdnd11an1n04x5 FILLER_369_1643 ();
 b15zdnd11an1n32x5 FILLER_369_1652 ();
 b15zdnd11an1n04x5 FILLER_369_1684 ();
 b15zdnd11an1n16x5 FILLER_369_1704 ();
 b15zdnd11an1n04x5 FILLER_369_1720 ();
 b15zdnd11an1n64x5 FILLER_369_1733 ();
 b15zdnd11an1n16x5 FILLER_369_1797 ();
 b15zdnd11an1n08x5 FILLER_369_1827 ();
 b15zdnd11an1n64x5 FILLER_369_1847 ();
 b15zdnd11an1n64x5 FILLER_369_1911 ();
 b15zdnd11an1n64x5 FILLER_369_1975 ();
 b15zdnd11an1n16x5 FILLER_369_2039 ();
 b15zdnd11an1n08x5 FILLER_369_2055 ();
 b15zdnd11an1n04x5 FILLER_369_2063 ();
 b15zdnd00an1n02x5 FILLER_369_2067 ();
 b15zdnd00an1n01x5 FILLER_369_2069 ();
 b15zdnd11an1n16x5 FILLER_369_2076 ();
 b15zdnd00an1n01x5 FILLER_369_2092 ();
 b15zdnd11an1n08x5 FILLER_369_2114 ();
 b15zdnd00an1n01x5 FILLER_369_2122 ();
 b15zdnd11an1n64x5 FILLER_369_2127 ();
 b15zdnd11an1n64x5 FILLER_369_2191 ();
 b15zdnd11an1n16x5 FILLER_369_2255 ();
 b15zdnd11an1n08x5 FILLER_369_2271 ();
 b15zdnd11an1n04x5 FILLER_369_2279 ();
 b15zdnd00an1n01x5 FILLER_369_2283 ();
 b15zdnd11an1n64x5 FILLER_370_8 ();
 b15zdnd11an1n64x5 FILLER_370_72 ();
 b15zdnd11an1n64x5 FILLER_370_136 ();
 b15zdnd11an1n32x5 FILLER_370_200 ();
 b15zdnd11an1n08x5 FILLER_370_232 ();
 b15zdnd11an1n08x5 FILLER_370_246 ();
 b15zdnd11an1n04x5 FILLER_370_254 ();
 b15zdnd00an1n01x5 FILLER_370_258 ();
 b15zdnd11an1n16x5 FILLER_370_271 ();
 b15zdnd11an1n04x5 FILLER_370_312 ();
 b15zdnd11an1n08x5 FILLER_370_340 ();
 b15zdnd00an1n02x5 FILLER_370_348 ();
 b15zdnd11an1n32x5 FILLER_370_356 ();
 b15zdnd00an1n01x5 FILLER_370_388 ();
 b15zdnd11an1n08x5 FILLER_370_395 ();
 b15zdnd11an1n04x5 FILLER_370_403 ();
 b15zdnd11an1n08x5 FILLER_370_416 ();
 b15zdnd11an1n04x5 FILLER_370_424 ();
 b15zdnd00an1n01x5 FILLER_370_428 ();
 b15zdnd11an1n64x5 FILLER_370_436 ();
 b15zdnd11an1n04x5 FILLER_370_500 ();
 b15zdnd11an1n04x5 FILLER_370_512 ();
 b15zdnd11an1n32x5 FILLER_370_528 ();
 b15zdnd11an1n16x5 FILLER_370_560 ();
 b15zdnd11an1n04x5 FILLER_370_576 ();
 b15zdnd00an1n02x5 FILLER_370_580 ();
 b15zdnd11an1n64x5 FILLER_370_592 ();
 b15zdnd11an1n32x5 FILLER_370_662 ();
 b15zdnd11an1n16x5 FILLER_370_694 ();
 b15zdnd11an1n08x5 FILLER_370_710 ();
 b15zdnd11an1n32x5 FILLER_370_726 ();
 b15zdnd00an1n01x5 FILLER_370_758 ();
 b15zdnd11an1n64x5 FILLER_370_764 ();
 b15zdnd11an1n04x5 FILLER_370_828 ();
 b15zdnd00an1n02x5 FILLER_370_832 ();
 b15zdnd00an1n01x5 FILLER_370_834 ();
 b15zdnd11an1n16x5 FILLER_370_839 ();
 b15zdnd11an1n08x5 FILLER_370_855 ();
 b15zdnd00an1n02x5 FILLER_370_863 ();
 b15zdnd00an1n01x5 FILLER_370_865 ();
 b15zdnd11an1n64x5 FILLER_370_880 ();
 b15zdnd11an1n64x5 FILLER_370_944 ();
 b15zdnd11an1n16x5 FILLER_370_1008 ();
 b15zdnd11an1n04x5 FILLER_370_1024 ();
 b15zdnd00an1n02x5 FILLER_370_1028 ();
 b15zdnd00an1n01x5 FILLER_370_1030 ();
 b15zdnd11an1n16x5 FILLER_370_1043 ();
 b15zdnd11an1n08x5 FILLER_370_1059 ();
 b15zdnd00an1n01x5 FILLER_370_1067 ();
 b15zdnd11an1n64x5 FILLER_370_1080 ();
 b15zdnd11an1n04x5 FILLER_370_1144 ();
 b15zdnd11an1n64x5 FILLER_370_1169 ();
 b15zdnd11an1n32x5 FILLER_370_1233 ();
 b15zdnd11an1n16x5 FILLER_370_1265 ();
 b15zdnd11an1n04x5 FILLER_370_1281 ();
 b15zdnd00an1n02x5 FILLER_370_1285 ();
 b15zdnd11an1n16x5 FILLER_370_1294 ();
 b15zdnd00an1n01x5 FILLER_370_1310 ();
 b15zdnd11an1n08x5 FILLER_370_1323 ();
 b15zdnd11an1n04x5 FILLER_370_1331 ();
 b15zdnd00an1n02x5 FILLER_370_1335 ();
 b15zdnd11an1n04x5 FILLER_370_1343 ();
 b15zdnd11an1n32x5 FILLER_370_1359 ();
 b15zdnd11an1n04x5 FILLER_370_1391 ();
 b15zdnd00an1n02x5 FILLER_370_1395 ();
 b15zdnd11an1n08x5 FILLER_370_1405 ();
 b15zdnd11an1n04x5 FILLER_370_1413 ();
 b15zdnd00an1n02x5 FILLER_370_1417 ();
 b15zdnd11an1n08x5 FILLER_370_1430 ();
 b15zdnd00an1n02x5 FILLER_370_1438 ();
 b15zdnd00an1n01x5 FILLER_370_1440 ();
 b15zdnd11an1n16x5 FILLER_370_1455 ();
 b15zdnd11an1n04x5 FILLER_370_1471 ();
 b15zdnd00an1n02x5 FILLER_370_1475 ();
 b15zdnd11an1n32x5 FILLER_370_1483 ();
 b15zdnd11an1n16x5 FILLER_370_1515 ();
 b15zdnd11an1n08x5 FILLER_370_1531 ();
 b15zdnd11an1n04x5 FILLER_370_1539 ();
 b15zdnd00an1n02x5 FILLER_370_1543 ();
 b15zdnd00an1n01x5 FILLER_370_1545 ();
 b15zdnd11an1n16x5 FILLER_370_1551 ();
 b15zdnd11an1n08x5 FILLER_370_1567 ();
 b15zdnd00an1n01x5 FILLER_370_1575 ();
 b15zdnd11an1n32x5 FILLER_370_1587 ();
 b15zdnd00an1n02x5 FILLER_370_1619 ();
 b15zdnd00an1n01x5 FILLER_370_1621 ();
 b15zdnd11an1n04x5 FILLER_370_1628 ();
 b15zdnd11an1n08x5 FILLER_370_1639 ();
 b15zdnd00an1n01x5 FILLER_370_1647 ();
 b15zdnd11an1n04x5 FILLER_370_1653 ();
 b15zdnd00an1n02x5 FILLER_370_1657 ();
 b15zdnd00an1n01x5 FILLER_370_1659 ();
 b15zdnd11an1n16x5 FILLER_370_1664 ();
 b15zdnd11an1n08x5 FILLER_370_1680 ();
 b15zdnd11an1n04x5 FILLER_370_1688 ();
 b15zdnd11an1n16x5 FILLER_370_1696 ();
 b15zdnd11an1n04x5 FILLER_370_1712 ();
 b15zdnd00an1n02x5 FILLER_370_1716 ();
 b15zdnd00an1n01x5 FILLER_370_1718 ();
 b15zdnd11an1n64x5 FILLER_370_1737 ();
 b15zdnd11an1n32x5 FILLER_370_1801 ();
 b15zdnd11an1n16x5 FILLER_370_1833 ();
 b15zdnd11an1n16x5 FILLER_370_1855 ();
 b15zdnd11an1n08x5 FILLER_370_1871 ();
 b15zdnd11an1n04x5 FILLER_370_1879 ();
 b15zdnd00an1n01x5 FILLER_370_1883 ();
 b15zdnd11an1n64x5 FILLER_370_1893 ();
 b15zdnd00an1n02x5 FILLER_370_1957 ();
 b15zdnd00an1n01x5 FILLER_370_1959 ();
 b15zdnd11an1n04x5 FILLER_370_1974 ();
 b15zdnd11an1n32x5 FILLER_370_1984 ();
 b15zdnd11an1n64x5 FILLER_370_2022 ();
 b15zdnd11an1n32x5 FILLER_370_2086 ();
 b15zdnd11an1n04x5 FILLER_370_2118 ();
 b15zdnd00an1n01x5 FILLER_370_2122 ();
 b15zdnd11an1n08x5 FILLER_370_2133 ();
 b15zdnd11an1n04x5 FILLER_370_2141 ();
 b15zdnd00an1n02x5 FILLER_370_2145 ();
 b15zdnd00an1n01x5 FILLER_370_2147 ();
 b15zdnd00an1n02x5 FILLER_370_2152 ();
 b15zdnd11an1n16x5 FILLER_370_2162 ();
 b15zdnd00an1n02x5 FILLER_370_2178 ();
 b15zdnd11an1n08x5 FILLER_370_2185 ();
 b15zdnd11an1n04x5 FILLER_370_2193 ();
 b15zdnd00an1n01x5 FILLER_370_2197 ();
 b15zdnd11an1n64x5 FILLER_370_2203 ();
 b15zdnd11an1n08x5 FILLER_370_2267 ();
 b15zdnd00an1n01x5 FILLER_370_2275 ();
 b15zdnd11an1n64x5 FILLER_371_0 ();
 b15zdnd11an1n64x5 FILLER_371_64 ();
 b15zdnd11an1n64x5 FILLER_371_128 ();
 b15zdnd11an1n32x5 FILLER_371_192 ();
 b15zdnd11an1n08x5 FILLER_371_224 ();
 b15zdnd00an1n02x5 FILLER_371_232 ();
 b15zdnd00an1n01x5 FILLER_371_234 ();
 b15zdnd11an1n04x5 FILLER_371_252 ();
 b15zdnd11an1n16x5 FILLER_371_275 ();
 b15zdnd11an1n08x5 FILLER_371_291 ();
 b15zdnd11an1n04x5 FILLER_371_299 ();
 b15zdnd00an1n01x5 FILLER_371_303 ();
 b15zdnd11an1n16x5 FILLER_371_318 ();
 b15zdnd11an1n16x5 FILLER_371_344 ();
 b15zdnd11an1n08x5 FILLER_371_360 ();
 b15zdnd00an1n02x5 FILLER_371_368 ();
 b15zdnd11an1n04x5 FILLER_371_376 ();
 b15zdnd11an1n64x5 FILLER_371_391 ();
 b15zdnd11an1n08x5 FILLER_371_455 ();
 b15zdnd11an1n04x5 FILLER_371_463 ();
 b15zdnd00an1n01x5 FILLER_371_467 ();
 b15zdnd11an1n08x5 FILLER_371_477 ();
 b15zdnd11an1n04x5 FILLER_371_485 ();
 b15zdnd00an1n01x5 FILLER_371_489 ();
 b15zdnd11an1n04x5 FILLER_371_496 ();
 b15zdnd11an1n16x5 FILLER_371_505 ();
 b15zdnd11an1n08x5 FILLER_371_521 ();
 b15zdnd11an1n04x5 FILLER_371_529 ();
 b15zdnd11an1n04x5 FILLER_371_537 ();
 b15zdnd11an1n08x5 FILLER_371_553 ();
 b15zdnd00an1n02x5 FILLER_371_561 ();
 b15zdnd00an1n01x5 FILLER_371_563 ();
 b15zdnd11an1n04x5 FILLER_371_582 ();
 b15zdnd11an1n64x5 FILLER_371_598 ();
 b15zdnd11an1n32x5 FILLER_371_662 ();
 b15zdnd11an1n04x5 FILLER_371_694 ();
 b15zdnd11an1n16x5 FILLER_371_707 ();
 b15zdnd11an1n04x5 FILLER_371_723 ();
 b15zdnd00an1n02x5 FILLER_371_727 ();
 b15zdnd11an1n04x5 FILLER_371_734 ();
 b15zdnd11an1n64x5 FILLER_371_746 ();
 b15zdnd11an1n16x5 FILLER_371_810 ();
 b15zdnd00an1n01x5 FILLER_371_826 ();
 b15zdnd11an1n16x5 FILLER_371_838 ();
 b15zdnd11an1n04x5 FILLER_371_854 ();
 b15zdnd00an1n02x5 FILLER_371_858 ();
 b15zdnd00an1n01x5 FILLER_371_860 ();
 b15zdnd11an1n64x5 FILLER_371_869 ();
 b15zdnd11an1n32x5 FILLER_371_933 ();
 b15zdnd11an1n04x5 FILLER_371_965 ();
 b15zdnd00an1n02x5 FILLER_371_969 ();
 b15zdnd00an1n01x5 FILLER_371_971 ();
 b15zdnd11an1n16x5 FILLER_371_978 ();
 b15zdnd11an1n08x5 FILLER_371_994 ();
 b15zdnd11an1n04x5 FILLER_371_1002 ();
 b15zdnd00an1n02x5 FILLER_371_1006 ();
 b15zdnd00an1n01x5 FILLER_371_1008 ();
 b15zdnd11an1n08x5 FILLER_371_1015 ();
 b15zdnd11an1n04x5 FILLER_371_1023 ();
 b15zdnd11an1n16x5 FILLER_371_1041 ();
 b15zdnd11an1n04x5 FILLER_371_1057 ();
 b15zdnd00an1n02x5 FILLER_371_1061 ();
 b15zdnd11an1n32x5 FILLER_371_1076 ();
 b15zdnd11an1n16x5 FILLER_371_1108 ();
 b15zdnd11an1n04x5 FILLER_371_1124 ();
 b15zdnd00an1n02x5 FILLER_371_1128 ();
 b15zdnd11an1n08x5 FILLER_371_1160 ();
 b15zdnd00an1n02x5 FILLER_371_1168 ();
 b15zdnd00an1n01x5 FILLER_371_1170 ();
 b15zdnd11an1n64x5 FILLER_371_1178 ();
 b15zdnd11an1n64x5 FILLER_371_1242 ();
 b15zdnd11an1n08x5 FILLER_371_1306 ();
 b15zdnd11an1n04x5 FILLER_371_1314 ();
 b15zdnd00an1n01x5 FILLER_371_1318 ();
 b15zdnd11an1n04x5 FILLER_371_1329 ();
 b15zdnd11an1n16x5 FILLER_371_1349 ();
 b15zdnd11an1n08x5 FILLER_371_1365 ();
 b15zdnd00an1n02x5 FILLER_371_1373 ();
 b15zdnd00an1n01x5 FILLER_371_1375 ();
 b15zdnd11an1n32x5 FILLER_371_1383 ();
 b15zdnd00an1n02x5 FILLER_371_1415 ();
 b15zdnd11an1n04x5 FILLER_371_1422 ();
 b15zdnd11an1n32x5 FILLER_371_1433 ();
 b15zdnd11an1n08x5 FILLER_371_1465 ();
 b15zdnd11an1n04x5 FILLER_371_1473 ();
 b15zdnd00an1n02x5 FILLER_371_1477 ();
 b15zdnd11an1n32x5 FILLER_371_1484 ();
 b15zdnd11an1n04x5 FILLER_371_1516 ();
 b15zdnd00an1n02x5 FILLER_371_1520 ();
 b15zdnd00an1n01x5 FILLER_371_1522 ();
 b15zdnd11an1n04x5 FILLER_371_1535 ();
 b15zdnd11an1n16x5 FILLER_371_1569 ();
 b15zdnd11an1n04x5 FILLER_371_1589 ();
 b15zdnd11an1n08x5 FILLER_371_1608 ();
 b15zdnd11an1n04x5 FILLER_371_1616 ();
 b15zdnd00an1n01x5 FILLER_371_1620 ();
 b15zdnd11an1n32x5 FILLER_371_1625 ();
 b15zdnd11an1n16x5 FILLER_371_1657 ();
 b15zdnd11an1n08x5 FILLER_371_1673 ();
 b15zdnd00an1n02x5 FILLER_371_1681 ();
 b15zdnd00an1n01x5 FILLER_371_1683 ();
 b15zdnd11an1n16x5 FILLER_371_1693 ();
 b15zdnd11an1n08x5 FILLER_371_1709 ();
 b15zdnd11an1n04x5 FILLER_371_1717 ();
 b15zdnd11an1n64x5 FILLER_371_1730 ();
 b15zdnd11an1n32x5 FILLER_371_1794 ();
 b15zdnd11an1n16x5 FILLER_371_1826 ();
 b15zdnd11an1n04x5 FILLER_371_1842 ();
 b15zdnd00an1n02x5 FILLER_371_1846 ();
 b15zdnd00an1n01x5 FILLER_371_1848 ();
 b15zdnd11an1n08x5 FILLER_371_1855 ();
 b15zdnd00an1n02x5 FILLER_371_1863 ();
 b15zdnd00an1n01x5 FILLER_371_1865 ();
 b15zdnd11an1n04x5 FILLER_371_1880 ();
 b15zdnd11an1n32x5 FILLER_371_1888 ();
 b15zdnd00an1n02x5 FILLER_371_1920 ();
 b15zdnd00an1n01x5 FILLER_371_1922 ();
 b15zdnd11an1n16x5 FILLER_371_1929 ();
 b15zdnd00an1n02x5 FILLER_371_1945 ();
 b15zdnd00an1n01x5 FILLER_371_1947 ();
 b15zdnd11an1n32x5 FILLER_371_1953 ();
 b15zdnd11an1n16x5 FILLER_371_1985 ();
 b15zdnd11an1n04x5 FILLER_371_2001 ();
 b15zdnd00an1n02x5 FILLER_371_2005 ();
 b15zdnd00an1n01x5 FILLER_371_2007 ();
 b15zdnd11an1n04x5 FILLER_371_2012 ();
 b15zdnd11an1n32x5 FILLER_371_2022 ();
 b15zdnd11an1n16x5 FILLER_371_2054 ();
 b15zdnd00an1n02x5 FILLER_371_2070 ();
 b15zdnd00an1n01x5 FILLER_371_2072 ();
 b15zdnd11an1n16x5 FILLER_371_2081 ();
 b15zdnd11an1n08x5 FILLER_371_2097 ();
 b15zdnd00an1n01x5 FILLER_371_2105 ();
 b15zdnd11an1n64x5 FILLER_371_2113 ();
 b15zdnd11an1n64x5 FILLER_371_2177 ();
 b15zdnd11an1n32x5 FILLER_371_2241 ();
 b15zdnd11an1n08x5 FILLER_371_2273 ();
 b15zdnd00an1n02x5 FILLER_371_2281 ();
 b15zdnd00an1n01x5 FILLER_371_2283 ();
 b15zdnd11an1n64x5 FILLER_372_8 ();
 b15zdnd11an1n64x5 FILLER_372_72 ();
 b15zdnd11an1n64x5 FILLER_372_136 ();
 b15zdnd11an1n32x5 FILLER_372_200 ();
 b15zdnd11an1n04x5 FILLER_372_232 ();
 b15zdnd11an1n64x5 FILLER_372_240 ();
 b15zdnd11an1n16x5 FILLER_372_304 ();
 b15zdnd00an1n02x5 FILLER_372_320 ();
 b15zdnd11an1n04x5 FILLER_372_334 ();
 b15zdnd11an1n16x5 FILLER_372_347 ();
 b15zdnd11an1n08x5 FILLER_372_363 ();
 b15zdnd11an1n08x5 FILLER_372_376 ();
 b15zdnd11an1n04x5 FILLER_372_384 ();
 b15zdnd00an1n01x5 FILLER_372_388 ();
 b15zdnd11an1n32x5 FILLER_372_394 ();
 b15zdnd11an1n16x5 FILLER_372_432 ();
 b15zdnd11an1n08x5 FILLER_372_448 ();
 b15zdnd11an1n64x5 FILLER_372_472 ();
 b15zdnd11an1n04x5 FILLER_372_536 ();
 b15zdnd00an1n02x5 FILLER_372_540 ();
 b15zdnd11an1n32x5 FILLER_372_548 ();
 b15zdnd11an1n08x5 FILLER_372_580 ();
 b15zdnd00an1n01x5 FILLER_372_588 ();
 b15zdnd11an1n64x5 FILLER_372_598 ();
 b15zdnd00an1n01x5 FILLER_372_662 ();
 b15zdnd11an1n04x5 FILLER_372_677 ();
 b15zdnd11an1n16x5 FILLER_372_693 ();
 b15zdnd11an1n08x5 FILLER_372_709 ();
 b15zdnd00an1n01x5 FILLER_372_717 ();
 b15zdnd11an1n64x5 FILLER_372_726 ();
 b15zdnd11an1n32x5 FILLER_372_790 ();
 b15zdnd00an1n02x5 FILLER_372_822 ();
 b15zdnd11an1n64x5 FILLER_372_830 ();
 b15zdnd11an1n16x5 FILLER_372_894 ();
 b15zdnd11an1n08x5 FILLER_372_910 ();
 b15zdnd11an1n04x5 FILLER_372_918 ();
 b15zdnd00an1n01x5 FILLER_372_922 ();
 b15zdnd11an1n32x5 FILLER_372_935 ();
 b15zdnd11an1n04x5 FILLER_372_967 ();
 b15zdnd11an1n16x5 FILLER_372_980 ();
 b15zdnd11an1n04x5 FILLER_372_996 ();
 b15zdnd00an1n02x5 FILLER_372_1000 ();
 b15zdnd11an1n16x5 FILLER_372_1019 ();
 b15zdnd00an1n01x5 FILLER_372_1035 ();
 b15zdnd11an1n08x5 FILLER_372_1043 ();
 b15zdnd11an1n04x5 FILLER_372_1051 ();
 b15zdnd00an1n02x5 FILLER_372_1055 ();
 b15zdnd00an1n01x5 FILLER_372_1057 ();
 b15zdnd11an1n32x5 FILLER_372_1072 ();
 b15zdnd11an1n16x5 FILLER_372_1104 ();
 b15zdnd11an1n04x5 FILLER_372_1126 ();
 b15zdnd00an1n01x5 FILLER_372_1130 ();
 b15zdnd11an1n08x5 FILLER_372_1140 ();
 b15zdnd11an1n04x5 FILLER_372_1148 ();
 b15zdnd00an1n02x5 FILLER_372_1152 ();
 b15zdnd11an1n08x5 FILLER_372_1160 ();
 b15zdnd11an1n04x5 FILLER_372_1168 ();
 b15zdnd11an1n64x5 FILLER_372_1186 ();
 b15zdnd11an1n16x5 FILLER_372_1250 ();
 b15zdnd00an1n01x5 FILLER_372_1266 ();
 b15zdnd11an1n04x5 FILLER_372_1290 ();
 b15zdnd11an1n04x5 FILLER_372_1312 ();
 b15zdnd11an1n32x5 FILLER_372_1324 ();
 b15zdnd11an1n16x5 FILLER_372_1356 ();
 b15zdnd11an1n08x5 FILLER_372_1372 ();
 b15zdnd00an1n01x5 FILLER_372_1380 ();
 b15zdnd11an1n16x5 FILLER_372_1388 ();
 b15zdnd11an1n04x5 FILLER_372_1414 ();
 b15zdnd00an1n02x5 FILLER_372_1418 ();
 b15zdnd00an1n01x5 FILLER_372_1420 ();
 b15zdnd11an1n16x5 FILLER_372_1426 ();
 b15zdnd11an1n04x5 FILLER_372_1442 ();
 b15zdnd00an1n01x5 FILLER_372_1446 ();
 b15zdnd11an1n16x5 FILLER_372_1455 ();
 b15zdnd11an1n08x5 FILLER_372_1471 ();
 b15zdnd11an1n32x5 FILLER_372_1486 ();
 b15zdnd00an1n02x5 FILLER_372_1518 ();
 b15zdnd00an1n01x5 FILLER_372_1520 ();
 b15zdnd11an1n16x5 FILLER_372_1528 ();
 b15zdnd11an1n04x5 FILLER_372_1544 ();
 b15zdnd00an1n02x5 FILLER_372_1548 ();
 b15zdnd00an1n01x5 FILLER_372_1550 ();
 b15zdnd11an1n08x5 FILLER_372_1557 ();
 b15zdnd11an1n04x5 FILLER_372_1565 ();
 b15zdnd00an1n02x5 FILLER_372_1569 ();
 b15zdnd11an1n04x5 FILLER_372_1578 ();
 b15zdnd11an1n64x5 FILLER_372_1589 ();
 b15zdnd11an1n16x5 FILLER_372_1653 ();
 b15zdnd00an1n02x5 FILLER_372_1669 ();
 b15zdnd11an1n04x5 FILLER_372_1687 ();
 b15zdnd11an1n64x5 FILLER_372_1700 ();
 b15zdnd11an1n32x5 FILLER_372_1764 ();
 b15zdnd11an1n16x5 FILLER_372_1796 ();
 b15zdnd11an1n08x5 FILLER_372_1812 ();
 b15zdnd11an1n04x5 FILLER_372_1820 ();
 b15zdnd00an1n02x5 FILLER_372_1824 ();
 b15zdnd11an1n04x5 FILLER_372_1830 ();
 b15zdnd11an1n04x5 FILLER_372_1846 ();
 b15zdnd11an1n08x5 FILLER_372_1858 ();
 b15zdnd11an1n04x5 FILLER_372_1866 ();
 b15zdnd00an1n02x5 FILLER_372_1870 ();
 b15zdnd00an1n01x5 FILLER_372_1872 ();
 b15zdnd11an1n08x5 FILLER_372_1879 ();
 b15zdnd11an1n04x5 FILLER_372_1887 ();
 b15zdnd00an1n01x5 FILLER_372_1891 ();
 b15zdnd11an1n16x5 FILLER_372_1896 ();
 b15zdnd11an1n04x5 FILLER_372_1912 ();
 b15zdnd00an1n02x5 FILLER_372_1916 ();
 b15zdnd00an1n01x5 FILLER_372_1918 ();
 b15zdnd11an1n04x5 FILLER_372_1931 ();
 b15zdnd11an1n08x5 FILLER_372_1940 ();
 b15zdnd11an1n04x5 FILLER_372_1948 ();
 b15zdnd11an1n04x5 FILLER_372_1958 ();
 b15zdnd11an1n16x5 FILLER_372_1967 ();
 b15zdnd11an1n04x5 FILLER_372_1988 ();
 b15zdnd11an1n08x5 FILLER_372_1997 ();
 b15zdnd11an1n04x5 FILLER_372_2005 ();
 b15zdnd11an1n16x5 FILLER_372_2016 ();
 b15zdnd11an1n08x5 FILLER_372_2032 ();
 b15zdnd00an1n02x5 FILLER_372_2040 ();
 b15zdnd11an1n32x5 FILLER_372_2046 ();
 b15zdnd11an1n04x5 FILLER_372_2078 ();
 b15zdnd00an1n02x5 FILLER_372_2082 ();
 b15zdnd00an1n01x5 FILLER_372_2084 ();
 b15zdnd11an1n04x5 FILLER_372_2095 ();
 b15zdnd00an1n02x5 FILLER_372_2099 ();
 b15zdnd00an1n01x5 FILLER_372_2101 ();
 b15zdnd11an1n04x5 FILLER_372_2114 ();
 b15zdnd11an1n16x5 FILLER_372_2134 ();
 b15zdnd11an1n04x5 FILLER_372_2150 ();
 b15zdnd11an1n04x5 FILLER_372_2162 ();
 b15zdnd00an1n02x5 FILLER_372_2166 ();
 b15zdnd00an1n01x5 FILLER_372_2168 ();
 b15zdnd11an1n08x5 FILLER_372_2185 ();
 b15zdnd00an1n01x5 FILLER_372_2193 ();
 b15zdnd11an1n04x5 FILLER_372_2200 ();
 b15zdnd11an1n04x5 FILLER_372_2210 ();
 b15zdnd00an1n02x5 FILLER_372_2214 ();
 b15zdnd11an1n32x5 FILLER_372_2228 ();
 b15zdnd11an1n16x5 FILLER_372_2260 ();
 b15zdnd11an1n64x5 FILLER_373_0 ();
 b15zdnd11an1n64x5 FILLER_373_64 ();
 b15zdnd11an1n64x5 FILLER_373_128 ();
 b15zdnd11an1n64x5 FILLER_373_192 ();
 b15zdnd11an1n04x5 FILLER_373_256 ();
 b15zdnd11an1n64x5 FILLER_373_278 ();
 b15zdnd11an1n16x5 FILLER_373_342 ();
 b15zdnd11an1n08x5 FILLER_373_358 ();
 b15zdnd11an1n04x5 FILLER_373_366 ();
 b15zdnd00an1n02x5 FILLER_373_370 ();
 b15zdnd11an1n32x5 FILLER_373_379 ();
 b15zdnd11an1n08x5 FILLER_373_411 ();
 b15zdnd00an1n01x5 FILLER_373_419 ();
 b15zdnd11an1n04x5 FILLER_373_429 ();
 b15zdnd00an1n01x5 FILLER_373_433 ();
 b15zdnd11an1n08x5 FILLER_373_447 ();
 b15zdnd11an1n04x5 FILLER_373_455 ();
 b15zdnd00an1n02x5 FILLER_373_459 ();
 b15zdnd00an1n01x5 FILLER_373_461 ();
 b15zdnd11an1n08x5 FILLER_373_468 ();
 b15zdnd11an1n04x5 FILLER_373_476 ();
 b15zdnd00an1n01x5 FILLER_373_480 ();
 b15zdnd11an1n64x5 FILLER_373_497 ();
 b15zdnd11an1n64x5 FILLER_373_561 ();
 b15zdnd11an1n32x5 FILLER_373_625 ();
 b15zdnd11an1n08x5 FILLER_373_657 ();
 b15zdnd11an1n08x5 FILLER_373_679 ();
 b15zdnd00an1n02x5 FILLER_373_687 ();
 b15zdnd00an1n01x5 FILLER_373_689 ();
 b15zdnd11an1n32x5 FILLER_373_708 ();
 b15zdnd11an1n16x5 FILLER_373_740 ();
 b15zdnd11an1n08x5 FILLER_373_756 ();
 b15zdnd00an1n01x5 FILLER_373_764 ();
 b15zdnd11an1n04x5 FILLER_373_772 ();
 b15zdnd11an1n04x5 FILLER_373_786 ();
 b15zdnd11an1n16x5 FILLER_373_803 ();
 b15zdnd11an1n04x5 FILLER_373_819 ();
 b15zdnd00an1n02x5 FILLER_373_823 ();
 b15zdnd00an1n01x5 FILLER_373_825 ();
 b15zdnd11an1n32x5 FILLER_373_832 ();
 b15zdnd11an1n08x5 FILLER_373_864 ();
 b15zdnd00an1n01x5 FILLER_373_872 ();
 b15zdnd11an1n16x5 FILLER_373_885 ();
 b15zdnd11an1n04x5 FILLER_373_901 ();
 b15zdnd11an1n04x5 FILLER_373_917 ();
 b15zdnd00an1n01x5 FILLER_373_921 ();
 b15zdnd11an1n04x5 FILLER_373_943 ();
 b15zdnd11an1n32x5 FILLER_373_959 ();
 b15zdnd11an1n16x5 FILLER_373_991 ();
 b15zdnd11an1n08x5 FILLER_373_1007 ();
 b15zdnd00an1n01x5 FILLER_373_1015 ();
 b15zdnd11an1n64x5 FILLER_373_1023 ();
 b15zdnd11an1n64x5 FILLER_373_1087 ();
 b15zdnd11an1n16x5 FILLER_373_1151 ();
 b15zdnd11an1n04x5 FILLER_373_1167 ();
 b15zdnd00an1n02x5 FILLER_373_1171 ();
 b15zdnd00an1n01x5 FILLER_373_1173 ();
 b15zdnd11an1n64x5 FILLER_373_1181 ();
 b15zdnd11an1n64x5 FILLER_373_1245 ();
 b15zdnd11an1n32x5 FILLER_373_1309 ();
 b15zdnd11an1n08x5 FILLER_373_1341 ();
 b15zdnd11an1n04x5 FILLER_373_1349 ();
 b15zdnd00an1n02x5 FILLER_373_1353 ();
 b15zdnd00an1n01x5 FILLER_373_1355 ();
 b15zdnd11an1n04x5 FILLER_373_1368 ();
 b15zdnd11an1n64x5 FILLER_373_1385 ();
 b15zdnd11an1n32x5 FILLER_373_1449 ();
 b15zdnd11an1n04x5 FILLER_373_1481 ();
 b15zdnd00an1n01x5 FILLER_373_1485 ();
 b15zdnd11an1n08x5 FILLER_373_1492 ();
 b15zdnd11an1n04x5 FILLER_373_1500 ();
 b15zdnd11an1n04x5 FILLER_373_1510 ();
 b15zdnd11an1n64x5 FILLER_373_1518 ();
 b15zdnd11an1n64x5 FILLER_373_1582 ();
 b15zdnd11an1n32x5 FILLER_373_1646 ();
 b15zdnd11an1n16x5 FILLER_373_1678 ();
 b15zdnd11an1n04x5 FILLER_373_1694 ();
 b15zdnd11an1n64x5 FILLER_373_1714 ();
 b15zdnd11an1n32x5 FILLER_373_1778 ();
 b15zdnd11an1n08x5 FILLER_373_1810 ();
 b15zdnd00an1n02x5 FILLER_373_1818 ();
 b15zdnd11an1n16x5 FILLER_373_1832 ();
 b15zdnd11an1n08x5 FILLER_373_1848 ();
 b15zdnd11an1n04x5 FILLER_373_1856 ();
 b15zdnd00an1n01x5 FILLER_373_1860 ();
 b15zdnd11an1n16x5 FILLER_373_1873 ();
 b15zdnd00an1n02x5 FILLER_373_1889 ();
 b15zdnd00an1n01x5 FILLER_373_1891 ();
 b15zdnd11an1n08x5 FILLER_373_1905 ();
 b15zdnd11an1n04x5 FILLER_373_1913 ();
 b15zdnd00an1n02x5 FILLER_373_1917 ();
 b15zdnd00an1n01x5 FILLER_373_1919 ();
 b15zdnd11an1n04x5 FILLER_373_1926 ();
 b15zdnd11an1n16x5 FILLER_373_1936 ();
 b15zdnd11an1n04x5 FILLER_373_1952 ();
 b15zdnd11an1n32x5 FILLER_373_1960 ();
 b15zdnd11an1n16x5 FILLER_373_1992 ();
 b15zdnd11an1n04x5 FILLER_373_2008 ();
 b15zdnd00an1n02x5 FILLER_373_2012 ();
 b15zdnd11an1n08x5 FILLER_373_2026 ();
 b15zdnd00an1n02x5 FILLER_373_2034 ();
 b15zdnd11an1n32x5 FILLER_373_2046 ();
 b15zdnd11an1n16x5 FILLER_373_2078 ();
 b15zdnd11an1n08x5 FILLER_373_2094 ();
 b15zdnd11an1n04x5 FILLER_373_2102 ();
 b15zdnd00an1n01x5 FILLER_373_2106 ();
 b15zdnd11an1n04x5 FILLER_373_2114 ();
 b15zdnd11an1n32x5 FILLER_373_2128 ();
 b15zdnd11an1n08x5 FILLER_373_2160 ();
 b15zdnd00an1n01x5 FILLER_373_2168 ();
 b15zdnd11an1n16x5 FILLER_373_2185 ();
 b15zdnd11an1n08x5 FILLER_373_2201 ();
 b15zdnd11an1n04x5 FILLER_373_2209 ();
 b15zdnd11an1n32x5 FILLER_373_2231 ();
 b15zdnd11an1n16x5 FILLER_373_2263 ();
 b15zdnd11an1n04x5 FILLER_373_2279 ();
 b15zdnd00an1n01x5 FILLER_373_2283 ();
 b15zdnd11an1n64x5 FILLER_374_8 ();
 b15zdnd11an1n64x5 FILLER_374_72 ();
 b15zdnd11an1n64x5 FILLER_374_136 ();
 b15zdnd11an1n16x5 FILLER_374_200 ();
 b15zdnd00an1n01x5 FILLER_374_216 ();
 b15zdnd11an1n64x5 FILLER_374_235 ();
 b15zdnd11an1n08x5 FILLER_374_299 ();
 b15zdnd11an1n64x5 FILLER_374_316 ();
 b15zdnd11an1n64x5 FILLER_374_380 ();
 b15zdnd00an1n01x5 FILLER_374_444 ();
 b15zdnd11an1n64x5 FILLER_374_450 ();
 b15zdnd11an1n16x5 FILLER_374_514 ();
 b15zdnd11an1n08x5 FILLER_374_530 ();
 b15zdnd00an1n02x5 FILLER_374_538 ();
 b15zdnd11an1n64x5 FILLER_374_547 ();
 b15zdnd11an1n32x5 FILLER_374_611 ();
 b15zdnd11an1n04x5 FILLER_374_650 ();
 b15zdnd11an1n32x5 FILLER_374_658 ();
 b15zdnd11an1n04x5 FILLER_374_690 ();
 b15zdnd00an1n02x5 FILLER_374_694 ();
 b15zdnd00an1n01x5 FILLER_374_696 ();
 b15zdnd11an1n04x5 FILLER_374_706 ();
 b15zdnd00an1n02x5 FILLER_374_716 ();
 b15zdnd11an1n16x5 FILLER_374_726 ();
 b15zdnd11an1n08x5 FILLER_374_742 ();
 b15zdnd11an1n04x5 FILLER_374_758 ();
 b15zdnd11an1n08x5 FILLER_374_768 ();
 b15zdnd00an1n01x5 FILLER_374_776 ();
 b15zdnd11an1n04x5 FILLER_374_786 ();
 b15zdnd11an1n16x5 FILLER_374_806 ();
 b15zdnd11an1n04x5 FILLER_374_822 ();
 b15zdnd11an1n32x5 FILLER_374_832 ();
 b15zdnd11an1n08x5 FILLER_374_864 ();
 b15zdnd11an1n04x5 FILLER_374_878 ();
 b15zdnd11an1n04x5 FILLER_374_889 ();
 b15zdnd11an1n04x5 FILLER_374_901 ();
 b15zdnd11an1n04x5 FILLER_374_926 ();
 b15zdnd11an1n16x5 FILLER_374_936 ();
 b15zdnd11an1n08x5 FILLER_374_952 ();
 b15zdnd11an1n04x5 FILLER_374_960 ();
 b15zdnd00an1n02x5 FILLER_374_964 ();
 b15zdnd00an1n01x5 FILLER_374_966 ();
 b15zdnd11an1n32x5 FILLER_374_973 ();
 b15zdnd11an1n04x5 FILLER_374_1005 ();
 b15zdnd00an1n01x5 FILLER_374_1009 ();
 b15zdnd11an1n08x5 FILLER_374_1022 ();
 b15zdnd00an1n02x5 FILLER_374_1030 ();
 b15zdnd00an1n01x5 FILLER_374_1032 ();
 b15zdnd11an1n16x5 FILLER_374_1037 ();
 b15zdnd11an1n04x5 FILLER_374_1053 ();
 b15zdnd00an1n02x5 FILLER_374_1057 ();
 b15zdnd00an1n01x5 FILLER_374_1059 ();
 b15zdnd11an1n16x5 FILLER_374_1074 ();
 b15zdnd11an1n04x5 FILLER_374_1095 ();
 b15zdnd00an1n01x5 FILLER_374_1099 ();
 b15zdnd11an1n64x5 FILLER_374_1106 ();
 b15zdnd11an1n08x5 FILLER_374_1170 ();
 b15zdnd11an1n04x5 FILLER_374_1178 ();
 b15zdnd00an1n01x5 FILLER_374_1182 ();
 b15zdnd11an1n64x5 FILLER_374_1199 ();
 b15zdnd11an1n64x5 FILLER_374_1263 ();
 b15zdnd11an1n64x5 FILLER_374_1347 ();
 b15zdnd11an1n64x5 FILLER_374_1411 ();
 b15zdnd11an1n04x5 FILLER_374_1475 ();
 b15zdnd00an1n02x5 FILLER_374_1479 ();
 b15zdnd11an1n16x5 FILLER_374_1488 ();
 b15zdnd11an1n64x5 FILLER_374_1510 ();
 b15zdnd11an1n08x5 FILLER_374_1574 ();
 b15zdnd11an1n04x5 FILLER_374_1582 ();
 b15zdnd00an1n01x5 FILLER_374_1586 ();
 b15zdnd11an1n16x5 FILLER_374_1599 ();
 b15zdnd00an1n02x5 FILLER_374_1615 ();
 b15zdnd00an1n01x5 FILLER_374_1617 ();
 b15zdnd11an1n64x5 FILLER_374_1629 ();
 b15zdnd11an1n64x5 FILLER_374_1693 ();
 b15zdnd11an1n64x5 FILLER_374_1757 ();
 b15zdnd11an1n32x5 FILLER_374_1821 ();
 b15zdnd11an1n08x5 FILLER_374_1853 ();
 b15zdnd11an1n04x5 FILLER_374_1861 ();
 b15zdnd11an1n16x5 FILLER_374_1871 ();
 b15zdnd11an1n64x5 FILLER_374_1903 ();
 b15zdnd11an1n64x5 FILLER_374_1967 ();
 b15zdnd11an1n04x5 FILLER_374_2031 ();
 b15zdnd00an1n02x5 FILLER_374_2035 ();
 b15zdnd00an1n01x5 FILLER_374_2037 ();
 b15zdnd11an1n04x5 FILLER_374_2043 ();
 b15zdnd11an1n64x5 FILLER_374_2056 ();
 b15zdnd00an1n01x5 FILLER_374_2120 ();
 b15zdnd11an1n16x5 FILLER_374_2135 ();
 b15zdnd00an1n02x5 FILLER_374_2151 ();
 b15zdnd00an1n01x5 FILLER_374_2153 ();
 b15zdnd11an1n16x5 FILLER_374_2162 ();
 b15zdnd11an1n08x5 FILLER_374_2178 ();
 b15zdnd11an1n64x5 FILLER_374_2202 ();
 b15zdnd11an1n08x5 FILLER_374_2266 ();
 b15zdnd00an1n02x5 FILLER_374_2274 ();
 b15zdnd11an1n64x5 FILLER_375_0 ();
 b15zdnd11an1n64x5 FILLER_375_64 ();
 b15zdnd11an1n64x5 FILLER_375_128 ();
 b15zdnd11an1n64x5 FILLER_375_192 ();
 b15zdnd11an1n16x5 FILLER_375_256 ();
 b15zdnd11an1n08x5 FILLER_375_272 ();
 b15zdnd11an1n64x5 FILLER_375_298 ();
 b15zdnd11an1n08x5 FILLER_375_362 ();
 b15zdnd11an1n04x5 FILLER_375_370 ();
 b15zdnd11an1n32x5 FILLER_375_388 ();
 b15zdnd11an1n04x5 FILLER_375_420 ();
 b15zdnd00an1n02x5 FILLER_375_424 ();
 b15zdnd00an1n01x5 FILLER_375_426 ();
 b15zdnd11an1n64x5 FILLER_375_433 ();
 b15zdnd00an1n02x5 FILLER_375_497 ();
 b15zdnd11an1n32x5 FILLER_375_505 ();
 b15zdnd11an1n16x5 FILLER_375_537 ();
 b15zdnd11an1n16x5 FILLER_375_560 ();
 b15zdnd11an1n08x5 FILLER_375_576 ();
 b15zdnd11an1n04x5 FILLER_375_584 ();
 b15zdnd11an1n32x5 FILLER_375_598 ();
 b15zdnd11an1n08x5 FILLER_375_630 ();
 b15zdnd00an1n02x5 FILLER_375_638 ();
 b15zdnd11an1n08x5 FILLER_375_656 ();
 b15zdnd11an1n04x5 FILLER_375_664 ();
 b15zdnd11an1n08x5 FILLER_375_680 ();
 b15zdnd11an1n04x5 FILLER_375_688 ();
 b15zdnd00an1n02x5 FILLER_375_692 ();
 b15zdnd11an1n04x5 FILLER_375_708 ();
 b15zdnd00an1n01x5 FILLER_375_712 ();
 b15zdnd11an1n64x5 FILLER_375_717 ();
 b15zdnd11an1n64x5 FILLER_375_781 ();
 b15zdnd00an1n02x5 FILLER_375_845 ();
 b15zdnd11an1n32x5 FILLER_375_854 ();
 b15zdnd11an1n16x5 FILLER_375_886 ();
 b15zdnd11an1n08x5 FILLER_375_902 ();
 b15zdnd00an1n01x5 FILLER_375_910 ();
 b15zdnd11an1n64x5 FILLER_375_915 ();
 b15zdnd11an1n16x5 FILLER_375_979 ();
 b15zdnd11an1n08x5 FILLER_375_995 ();
 b15zdnd11an1n04x5 FILLER_375_1003 ();
 b15zdnd00an1n02x5 FILLER_375_1007 ();
 b15zdnd11an1n08x5 FILLER_375_1016 ();
 b15zdnd11an1n04x5 FILLER_375_1024 ();
 b15zdnd00an1n01x5 FILLER_375_1028 ();
 b15zdnd11an1n16x5 FILLER_375_1045 ();
 b15zdnd00an1n01x5 FILLER_375_1061 ();
 b15zdnd11an1n16x5 FILLER_375_1071 ();
 b15zdnd00an1n01x5 FILLER_375_1087 ();
 b15zdnd11an1n32x5 FILLER_375_1093 ();
 b15zdnd11an1n16x5 FILLER_375_1125 ();
 b15zdnd11an1n04x5 FILLER_375_1141 ();
 b15zdnd00an1n02x5 FILLER_375_1145 ();
 b15zdnd00an1n01x5 FILLER_375_1147 ();
 b15zdnd11an1n64x5 FILLER_375_1164 ();
 b15zdnd11an1n64x5 FILLER_375_1228 ();
 b15zdnd11an1n32x5 FILLER_375_1292 ();
 b15zdnd00an1n02x5 FILLER_375_1324 ();
 b15zdnd00an1n01x5 FILLER_375_1326 ();
 b15zdnd11an1n64x5 FILLER_375_1339 ();
 b15zdnd11an1n32x5 FILLER_375_1403 ();
 b15zdnd00an1n01x5 FILLER_375_1435 ();
 b15zdnd11an1n32x5 FILLER_375_1447 ();
 b15zdnd11an1n16x5 FILLER_375_1479 ();
 b15zdnd11an1n08x5 FILLER_375_1495 ();
 b15zdnd00an1n02x5 FILLER_375_1503 ();
 b15zdnd11an1n64x5 FILLER_375_1514 ();
 b15zdnd11an1n32x5 FILLER_375_1578 ();
 b15zdnd11an1n04x5 FILLER_375_1610 ();
 b15zdnd11an1n04x5 FILLER_375_1624 ();
 b15zdnd00an1n01x5 FILLER_375_1628 ();
 b15zdnd11an1n04x5 FILLER_375_1634 ();
 b15zdnd11an1n16x5 FILLER_375_1644 ();
 b15zdnd11an1n08x5 FILLER_375_1660 ();
 b15zdnd00an1n02x5 FILLER_375_1668 ();
 b15zdnd00an1n01x5 FILLER_375_1670 ();
 b15zdnd11an1n08x5 FILLER_375_1677 ();
 b15zdnd11an1n04x5 FILLER_375_1685 ();
 b15zdnd00an1n02x5 FILLER_375_1689 ();
 b15zdnd11an1n04x5 FILLER_375_1712 ();
 b15zdnd11an1n64x5 FILLER_375_1732 ();
 b15zdnd11an1n32x5 FILLER_375_1796 ();
 b15zdnd11an1n16x5 FILLER_375_1842 ();
 b15zdnd11an1n04x5 FILLER_375_1858 ();
 b15zdnd00an1n02x5 FILLER_375_1862 ();
 b15zdnd00an1n01x5 FILLER_375_1864 ();
 b15zdnd11an1n32x5 FILLER_375_1870 ();
 b15zdnd11an1n08x5 FILLER_375_1902 ();
 b15zdnd11an1n04x5 FILLER_375_1910 ();
 b15zdnd00an1n02x5 FILLER_375_1914 ();
 b15zdnd00an1n01x5 FILLER_375_1916 ();
 b15zdnd11an1n64x5 FILLER_375_1921 ();
 b15zdnd11an1n64x5 FILLER_375_1985 ();
 b15zdnd11an1n64x5 FILLER_375_2049 ();
 b15zdnd11an1n64x5 FILLER_375_2113 ();
 b15zdnd11an1n64x5 FILLER_375_2177 ();
 b15zdnd11an1n32x5 FILLER_375_2241 ();
 b15zdnd11an1n08x5 FILLER_375_2273 ();
 b15zdnd00an1n02x5 FILLER_375_2281 ();
 b15zdnd00an1n01x5 FILLER_375_2283 ();
 b15zdnd11an1n64x5 FILLER_376_8 ();
 b15zdnd11an1n64x5 FILLER_376_72 ();
 b15zdnd11an1n64x5 FILLER_376_136 ();
 b15zdnd11an1n32x5 FILLER_376_200 ();
 b15zdnd11an1n04x5 FILLER_376_232 ();
 b15zdnd00an1n02x5 FILLER_376_236 ();
 b15zdnd11an1n04x5 FILLER_376_250 ();
 b15zdnd11an1n04x5 FILLER_376_261 ();
 b15zdnd11an1n08x5 FILLER_376_277 ();
 b15zdnd11an1n04x5 FILLER_376_285 ();
 b15zdnd11an1n08x5 FILLER_376_296 ();
 b15zdnd11an1n04x5 FILLER_376_304 ();
 b15zdnd00an1n01x5 FILLER_376_308 ();
 b15zdnd11an1n32x5 FILLER_376_314 ();
 b15zdnd11an1n16x5 FILLER_376_346 ();
 b15zdnd11an1n04x5 FILLER_376_362 ();
 b15zdnd00an1n02x5 FILLER_376_366 ();
 b15zdnd00an1n01x5 FILLER_376_368 ();
 b15zdnd11an1n04x5 FILLER_376_381 ();
 b15zdnd11an1n04x5 FILLER_376_397 ();
 b15zdnd11an1n16x5 FILLER_376_411 ();
 b15zdnd11an1n08x5 FILLER_376_427 ();
 b15zdnd11an1n04x5 FILLER_376_450 ();
 b15zdnd11an1n04x5 FILLER_376_466 ();
 b15zdnd00an1n01x5 FILLER_376_470 ();
 b15zdnd11an1n32x5 FILLER_376_477 ();
 b15zdnd11an1n08x5 FILLER_376_509 ();
 b15zdnd11an1n16x5 FILLER_376_523 ();
 b15zdnd11an1n08x5 FILLER_376_549 ();
 b15zdnd11an1n08x5 FILLER_376_564 ();
 b15zdnd00an1n01x5 FILLER_376_572 ();
 b15zdnd11an1n64x5 FILLER_376_589 ();
 b15zdnd11an1n08x5 FILLER_376_653 ();
 b15zdnd00an1n02x5 FILLER_376_661 ();
 b15zdnd00an1n01x5 FILLER_376_663 ();
 b15zdnd11an1n16x5 FILLER_376_684 ();
 b15zdnd11an1n04x5 FILLER_376_700 ();
 b15zdnd11an1n04x5 FILLER_376_714 ();
 b15zdnd11an1n64x5 FILLER_376_726 ();
 b15zdnd11an1n32x5 FILLER_376_790 ();
 b15zdnd11an1n08x5 FILLER_376_838 ();
 b15zdnd11an1n04x5 FILLER_376_846 ();
 b15zdnd00an1n01x5 FILLER_376_850 ();
 b15zdnd11an1n64x5 FILLER_376_866 ();
 b15zdnd11an1n64x5 FILLER_376_930 ();
 b15zdnd11an1n16x5 FILLER_376_994 ();
 b15zdnd11an1n16x5 FILLER_376_1015 ();
 b15zdnd00an1n02x5 FILLER_376_1031 ();
 b15zdnd11an1n64x5 FILLER_376_1041 ();
 b15zdnd11an1n64x5 FILLER_376_1105 ();
 b15zdnd11an1n64x5 FILLER_376_1169 ();
 b15zdnd11an1n64x5 FILLER_376_1233 ();
 b15zdnd11an1n16x5 FILLER_376_1297 ();
 b15zdnd00an1n02x5 FILLER_376_1313 ();
 b15zdnd00an1n01x5 FILLER_376_1315 ();
 b15zdnd11an1n16x5 FILLER_376_1326 ();
 b15zdnd11an1n32x5 FILLER_376_1353 ();
 b15zdnd11an1n16x5 FILLER_376_1385 ();
 b15zdnd11an1n08x5 FILLER_376_1401 ();
 b15zdnd11an1n64x5 FILLER_376_1425 ();
 b15zdnd11an1n64x5 FILLER_376_1489 ();
 b15zdnd11an1n16x5 FILLER_376_1553 ();
 b15zdnd00an1n01x5 FILLER_376_1569 ();
 b15zdnd11an1n08x5 FILLER_376_1575 ();
 b15zdnd00an1n02x5 FILLER_376_1583 ();
 b15zdnd11an1n08x5 FILLER_376_1597 ();
 b15zdnd11an1n04x5 FILLER_376_1605 ();
 b15zdnd00an1n02x5 FILLER_376_1609 ();
 b15zdnd00an1n01x5 FILLER_376_1611 ();
 b15zdnd11an1n16x5 FILLER_376_1617 ();
 b15zdnd11an1n08x5 FILLER_376_1633 ();
 b15zdnd11an1n04x5 FILLER_376_1641 ();
 b15zdnd00an1n01x5 FILLER_376_1645 ();
 b15zdnd11an1n16x5 FILLER_376_1652 ();
 b15zdnd00an1n02x5 FILLER_376_1668 ();
 b15zdnd11an1n08x5 FILLER_376_1678 ();
 b15zdnd00an1n02x5 FILLER_376_1686 ();
 b15zdnd11an1n16x5 FILLER_376_1693 ();
 b15zdnd00an1n02x5 FILLER_376_1709 ();
 b15zdnd11an1n64x5 FILLER_376_1727 ();
 b15zdnd11an1n64x5 FILLER_376_1791 ();
 b15zdnd11an1n16x5 FILLER_376_1855 ();
 b15zdnd11an1n04x5 FILLER_376_1871 ();
 b15zdnd11an1n08x5 FILLER_376_1881 ();
 b15zdnd00an1n02x5 FILLER_376_1889 ();
 b15zdnd00an1n01x5 FILLER_376_1891 ();
 b15zdnd11an1n64x5 FILLER_376_1897 ();
 b15zdnd11an1n16x5 FILLER_376_1961 ();
 b15zdnd11an1n08x5 FILLER_376_1977 ();
 b15zdnd11an1n04x5 FILLER_376_1985 ();
 b15zdnd11an1n64x5 FILLER_376_1999 ();
 b15zdnd11an1n16x5 FILLER_376_2063 ();
 b15zdnd11an1n08x5 FILLER_376_2079 ();
 b15zdnd11an1n04x5 FILLER_376_2087 ();
 b15zdnd00an1n01x5 FILLER_376_2091 ();
 b15zdnd11an1n04x5 FILLER_376_2097 ();
 b15zdnd11an1n32x5 FILLER_376_2107 ();
 b15zdnd00an1n01x5 FILLER_376_2139 ();
 b15zdnd11an1n08x5 FILLER_376_2144 ();
 b15zdnd00an1n02x5 FILLER_376_2152 ();
 b15zdnd00an1n02x5 FILLER_376_2162 ();
 b15zdnd00an1n01x5 FILLER_376_2164 ();
 b15zdnd11an1n16x5 FILLER_376_2183 ();
 b15zdnd00an1n02x5 FILLER_376_2199 ();
 b15zdnd11an1n32x5 FILLER_376_2219 ();
 b15zdnd11an1n16x5 FILLER_376_2251 ();
 b15zdnd11an1n08x5 FILLER_376_2267 ();
 b15zdnd00an1n01x5 FILLER_376_2275 ();
 b15zdnd11an1n64x5 FILLER_377_0 ();
 b15zdnd11an1n64x5 FILLER_377_64 ();
 b15zdnd11an1n64x5 FILLER_377_128 ();
 b15zdnd11an1n32x5 FILLER_377_192 ();
 b15zdnd11an1n16x5 FILLER_377_224 ();
 b15zdnd00an1n02x5 FILLER_377_240 ();
 b15zdnd11an1n32x5 FILLER_377_260 ();
 b15zdnd11an1n16x5 FILLER_377_292 ();
 b15zdnd11an1n04x5 FILLER_377_308 ();
 b15zdnd11an1n04x5 FILLER_377_317 ();
 b15zdnd00an1n02x5 FILLER_377_321 ();
 b15zdnd00an1n01x5 FILLER_377_323 ();
 b15zdnd11an1n08x5 FILLER_377_332 ();
 b15zdnd00an1n02x5 FILLER_377_340 ();
 b15zdnd11an1n08x5 FILLER_377_354 ();
 b15zdnd11an1n04x5 FILLER_377_362 ();
 b15zdnd00an1n01x5 FILLER_377_366 ();
 b15zdnd11an1n16x5 FILLER_377_391 ();
 b15zdnd11an1n08x5 FILLER_377_407 ();
 b15zdnd00an1n02x5 FILLER_377_415 ();
 b15zdnd00an1n01x5 FILLER_377_417 ();
 b15zdnd11an1n08x5 FILLER_377_425 ();
 b15zdnd00an1n02x5 FILLER_377_433 ();
 b15zdnd00an1n01x5 FILLER_377_435 ();
 b15zdnd11an1n16x5 FILLER_377_450 ();
 b15zdnd11an1n08x5 FILLER_377_466 ();
 b15zdnd00an1n02x5 FILLER_377_474 ();
 b15zdnd11an1n04x5 FILLER_377_491 ();
 b15zdnd00an1n02x5 FILLER_377_495 ();
 b15zdnd00an1n01x5 FILLER_377_497 ();
 b15zdnd11an1n32x5 FILLER_377_504 ();
 b15zdnd11an1n08x5 FILLER_377_536 ();
 b15zdnd00an1n02x5 FILLER_377_544 ();
 b15zdnd00an1n01x5 FILLER_377_546 ();
 b15zdnd11an1n04x5 FILLER_377_552 ();
 b15zdnd00an1n02x5 FILLER_377_556 ();
 b15zdnd11an1n64x5 FILLER_377_567 ();
 b15zdnd11an1n64x5 FILLER_377_631 ();
 b15zdnd11an1n64x5 FILLER_377_695 ();
 b15zdnd11an1n04x5 FILLER_377_759 ();
 b15zdnd11an1n32x5 FILLER_377_778 ();
 b15zdnd11an1n08x5 FILLER_377_810 ();
 b15zdnd11an1n04x5 FILLER_377_818 ();
 b15zdnd00an1n02x5 FILLER_377_822 ();
 b15zdnd11an1n64x5 FILLER_377_829 ();
 b15zdnd11an1n32x5 FILLER_377_893 ();
 b15zdnd00an1n02x5 FILLER_377_925 ();
 b15zdnd11an1n64x5 FILLER_377_941 ();
 b15zdnd11an1n32x5 FILLER_377_1005 ();
 b15zdnd00an1n02x5 FILLER_377_1037 ();
 b15zdnd00an1n01x5 FILLER_377_1039 ();
 b15zdnd11an1n64x5 FILLER_377_1056 ();
 b15zdnd11an1n16x5 FILLER_377_1120 ();
 b15zdnd00an1n01x5 FILLER_377_1136 ();
 b15zdnd11an1n64x5 FILLER_377_1153 ();
 b15zdnd11an1n64x5 FILLER_377_1217 ();
 b15zdnd11an1n32x5 FILLER_377_1281 ();
 b15zdnd00an1n02x5 FILLER_377_1313 ();
 b15zdnd00an1n01x5 FILLER_377_1315 ();
 b15zdnd11an1n08x5 FILLER_377_1332 ();
 b15zdnd00an1n02x5 FILLER_377_1340 ();
 b15zdnd00an1n01x5 FILLER_377_1342 ();
 b15zdnd11an1n08x5 FILLER_377_1351 ();
 b15zdnd11an1n04x5 FILLER_377_1359 ();
 b15zdnd11an1n04x5 FILLER_377_1371 ();
 b15zdnd11an1n32x5 FILLER_377_1381 ();
 b15zdnd11an1n04x5 FILLER_377_1413 ();
 b15zdnd00an1n02x5 FILLER_377_1417 ();
 b15zdnd11an1n08x5 FILLER_377_1427 ();
 b15zdnd11an1n04x5 FILLER_377_1435 ();
 b15zdnd00an1n02x5 FILLER_377_1439 ();
 b15zdnd11an1n04x5 FILLER_377_1448 ();
 b15zdnd11an1n08x5 FILLER_377_1457 ();
 b15zdnd00an1n02x5 FILLER_377_1465 ();
 b15zdnd00an1n01x5 FILLER_377_1467 ();
 b15zdnd11an1n32x5 FILLER_377_1480 ();
 b15zdnd00an1n01x5 FILLER_377_1512 ();
 b15zdnd11an1n16x5 FILLER_377_1529 ();
 b15zdnd00an1n01x5 FILLER_377_1545 ();
 b15zdnd11an1n04x5 FILLER_377_1554 ();
 b15zdnd11an1n16x5 FILLER_377_1564 ();
 b15zdnd11an1n08x5 FILLER_377_1580 ();
 b15zdnd11an1n32x5 FILLER_377_1594 ();
 b15zdnd11an1n16x5 FILLER_377_1626 ();
 b15zdnd11an1n04x5 FILLER_377_1642 ();
 b15zdnd00an1n02x5 FILLER_377_1646 ();
 b15zdnd11an1n16x5 FILLER_377_1660 ();
 b15zdnd00an1n02x5 FILLER_377_1676 ();
 b15zdnd11an1n64x5 FILLER_377_1696 ();
 b15zdnd11an1n64x5 FILLER_377_1760 ();
 b15zdnd11an1n04x5 FILLER_377_1840 ();
 b15zdnd11an1n16x5 FILLER_377_1856 ();
 b15zdnd11an1n04x5 FILLER_377_1872 ();
 b15zdnd00an1n01x5 FILLER_377_1876 ();
 b15zdnd11an1n08x5 FILLER_377_1883 ();
 b15zdnd00an1n02x5 FILLER_377_1891 ();
 b15zdnd11an1n04x5 FILLER_377_1900 ();
 b15zdnd11an1n16x5 FILLER_377_1909 ();
 b15zdnd11an1n08x5 FILLER_377_1925 ();
 b15zdnd00an1n01x5 FILLER_377_1933 ();
 b15zdnd11an1n08x5 FILLER_377_1942 ();
 b15zdnd00an1n02x5 FILLER_377_1950 ();
 b15zdnd11an1n04x5 FILLER_377_1978 ();
 b15zdnd00an1n01x5 FILLER_377_1982 ();
 b15zdnd11an1n04x5 FILLER_377_1989 ();
 b15zdnd11an1n04x5 FILLER_377_2002 ();
 b15zdnd11an1n04x5 FILLER_377_2025 ();
 b15zdnd11an1n16x5 FILLER_377_2050 ();
 b15zdnd11an1n08x5 FILLER_377_2066 ();
 b15zdnd00an1n02x5 FILLER_377_2074 ();
 b15zdnd11an1n32x5 FILLER_377_2087 ();
 b15zdnd00an1n01x5 FILLER_377_2119 ();
 b15zdnd11an1n08x5 FILLER_377_2126 ();
 b15zdnd11an1n04x5 FILLER_377_2134 ();
 b15zdnd11an1n16x5 FILLER_377_2148 ();
 b15zdnd11an1n04x5 FILLER_377_2164 ();
 b15zdnd00an1n02x5 FILLER_377_2168 ();
 b15zdnd11an1n64x5 FILLER_377_2186 ();
 b15zdnd11an1n32x5 FILLER_377_2250 ();
 b15zdnd00an1n02x5 FILLER_377_2282 ();
 b15zdnd11an1n64x5 FILLER_378_8 ();
 b15zdnd11an1n64x5 FILLER_378_72 ();
 b15zdnd11an1n64x5 FILLER_378_136 ();
 b15zdnd11an1n32x5 FILLER_378_200 ();
 b15zdnd11an1n08x5 FILLER_378_232 ();
 b15zdnd11an1n04x5 FILLER_378_240 ();
 b15zdnd00an1n02x5 FILLER_378_244 ();
 b15zdnd00an1n01x5 FILLER_378_246 ();
 b15zdnd11an1n32x5 FILLER_378_265 ();
 b15zdnd11an1n04x5 FILLER_378_297 ();
 b15zdnd11an1n08x5 FILLER_378_322 ();
 b15zdnd11an1n04x5 FILLER_378_330 ();
 b15zdnd00an1n01x5 FILLER_378_334 ();
 b15zdnd11an1n08x5 FILLER_378_356 ();
 b15zdnd11an1n04x5 FILLER_378_364 ();
 b15zdnd00an1n02x5 FILLER_378_368 ();
 b15zdnd00an1n01x5 FILLER_378_370 ();
 b15zdnd11an1n04x5 FILLER_378_379 ();
 b15zdnd00an1n02x5 FILLER_378_383 ();
 b15zdnd00an1n01x5 FILLER_378_385 ();
 b15zdnd11an1n64x5 FILLER_378_390 ();
 b15zdnd11an1n08x5 FILLER_378_454 ();
 b15zdnd11an1n04x5 FILLER_378_462 ();
 b15zdnd00an1n01x5 FILLER_378_466 ();
 b15zdnd11an1n32x5 FILLER_378_485 ();
 b15zdnd11an1n16x5 FILLER_378_517 ();
 b15zdnd11an1n08x5 FILLER_378_533 ();
 b15zdnd11an1n04x5 FILLER_378_541 ();
 b15zdnd00an1n02x5 FILLER_378_545 ();
 b15zdnd00an1n01x5 FILLER_378_547 ();
 b15zdnd11an1n64x5 FILLER_378_555 ();
 b15zdnd11an1n32x5 FILLER_378_619 ();
 b15zdnd11an1n16x5 FILLER_378_651 ();
 b15zdnd00an1n01x5 FILLER_378_667 ();
 b15zdnd11an1n04x5 FILLER_378_678 ();
 b15zdnd11an1n16x5 FILLER_378_687 ();
 b15zdnd11an1n04x5 FILLER_378_703 ();
 b15zdnd00an1n02x5 FILLER_378_707 ();
 b15zdnd00an1n01x5 FILLER_378_709 ();
 b15zdnd00an1n02x5 FILLER_378_716 ();
 b15zdnd11an1n08x5 FILLER_378_726 ();
 b15zdnd00an1n02x5 FILLER_378_734 ();
 b15zdnd00an1n01x5 FILLER_378_736 ();
 b15zdnd11an1n04x5 FILLER_378_752 ();
 b15zdnd11an1n32x5 FILLER_378_765 ();
 b15zdnd11an1n16x5 FILLER_378_808 ();
 b15zdnd11an1n08x5 FILLER_378_824 ();
 b15zdnd00an1n02x5 FILLER_378_832 ();
 b15zdnd00an1n01x5 FILLER_378_834 ();
 b15zdnd11an1n64x5 FILLER_378_845 ();
 b15zdnd11an1n16x5 FILLER_378_909 ();
 b15zdnd11an1n08x5 FILLER_378_925 ();
 b15zdnd11an1n04x5 FILLER_378_941 ();
 b15zdnd11an1n04x5 FILLER_378_956 ();
 b15zdnd00an1n02x5 FILLER_378_960 ();
 b15zdnd11an1n64x5 FILLER_378_967 ();
 b15zdnd00an1n01x5 FILLER_378_1031 ();
 b15zdnd11an1n64x5 FILLER_378_1048 ();
 b15zdnd11an1n32x5 FILLER_378_1112 ();
 b15zdnd00an1n02x5 FILLER_378_1144 ();
 b15zdnd00an1n01x5 FILLER_378_1146 ();
 b15zdnd11an1n64x5 FILLER_378_1159 ();
 b15zdnd11an1n64x5 FILLER_378_1223 ();
 b15zdnd11an1n16x5 FILLER_378_1287 ();
 b15zdnd11an1n04x5 FILLER_378_1303 ();
 b15zdnd00an1n02x5 FILLER_378_1307 ();
 b15zdnd11an1n16x5 FILLER_378_1325 ();
 b15zdnd00an1n02x5 FILLER_378_1341 ();
 b15zdnd00an1n01x5 FILLER_378_1343 ();
 b15zdnd11an1n04x5 FILLER_378_1348 ();
 b15zdnd11an1n16x5 FILLER_378_1360 ();
 b15zdnd11an1n16x5 FILLER_378_1380 ();
 b15zdnd11an1n04x5 FILLER_378_1396 ();
 b15zdnd00an1n02x5 FILLER_378_1400 ();
 b15zdnd00an1n01x5 FILLER_378_1402 ();
 b15zdnd11an1n04x5 FILLER_378_1418 ();
 b15zdnd11an1n32x5 FILLER_378_1438 ();
 b15zdnd11an1n04x5 FILLER_378_1470 ();
 b15zdnd11an1n16x5 FILLER_378_1481 ();
 b15zdnd11an1n08x5 FILLER_378_1497 ();
 b15zdnd11an1n04x5 FILLER_378_1505 ();
 b15zdnd00an1n01x5 FILLER_378_1509 ();
 b15zdnd11an1n04x5 FILLER_378_1531 ();
 b15zdnd11an1n64x5 FILLER_378_1541 ();
 b15zdnd11an1n64x5 FILLER_378_1605 ();
 b15zdnd11an1n64x5 FILLER_378_1669 ();
 b15zdnd11an1n64x5 FILLER_378_1733 ();
 b15zdnd11an1n32x5 FILLER_378_1797 ();
 b15zdnd11an1n16x5 FILLER_378_1829 ();
 b15zdnd11an1n04x5 FILLER_378_1845 ();
 b15zdnd00an1n02x5 FILLER_378_1849 ();
 b15zdnd11an1n32x5 FILLER_378_1863 ();
 b15zdnd11an1n16x5 FILLER_378_1900 ();
 b15zdnd11an1n08x5 FILLER_378_1916 ();
 b15zdnd11an1n04x5 FILLER_378_1924 ();
 b15zdnd00an1n02x5 FILLER_378_1928 ();
 b15zdnd00an1n01x5 FILLER_378_1930 ();
 b15zdnd11an1n04x5 FILLER_378_1945 ();
 b15zdnd00an1n02x5 FILLER_378_1949 ();
 b15zdnd11an1n08x5 FILLER_378_1965 ();
 b15zdnd11an1n04x5 FILLER_378_1973 ();
 b15zdnd11an1n32x5 FILLER_378_1982 ();
 b15zdnd11an1n08x5 FILLER_378_2014 ();
 b15zdnd00an1n01x5 FILLER_378_2022 ();
 b15zdnd11an1n04x5 FILLER_378_2033 ();
 b15zdnd00an1n02x5 FILLER_378_2037 ();
 b15zdnd00an1n01x5 FILLER_378_2039 ();
 b15zdnd11an1n16x5 FILLER_378_2044 ();
 b15zdnd11an1n08x5 FILLER_378_2060 ();
 b15zdnd00an1n02x5 FILLER_378_2068 ();
 b15zdnd11an1n04x5 FILLER_378_2075 ();
 b15zdnd11an1n08x5 FILLER_378_2088 ();
 b15zdnd11an1n04x5 FILLER_378_2096 ();
 b15zdnd00an1n02x5 FILLER_378_2100 ();
 b15zdnd00an1n01x5 FILLER_378_2102 ();
 b15zdnd11an1n04x5 FILLER_378_2124 ();
 b15zdnd11an1n04x5 FILLER_378_2148 ();
 b15zdnd00an1n02x5 FILLER_378_2152 ();
 b15zdnd00an1n02x5 FILLER_378_2162 ();
 b15zdnd00an1n01x5 FILLER_378_2164 ();
 b15zdnd11an1n08x5 FILLER_378_2181 ();
 b15zdnd11an1n64x5 FILLER_378_2205 ();
 b15zdnd11an1n04x5 FILLER_378_2269 ();
 b15zdnd00an1n02x5 FILLER_378_2273 ();
 b15zdnd00an1n01x5 FILLER_378_2275 ();
 b15zdnd11an1n64x5 FILLER_379_0 ();
 b15zdnd11an1n64x5 FILLER_379_64 ();
 b15zdnd11an1n64x5 FILLER_379_128 ();
 b15zdnd11an1n64x5 FILLER_379_192 ();
 b15zdnd11an1n16x5 FILLER_379_256 ();
 b15zdnd11an1n04x5 FILLER_379_272 ();
 b15zdnd00an1n01x5 FILLER_379_276 ();
 b15zdnd11an1n16x5 FILLER_379_297 ();
 b15zdnd00an1n02x5 FILLER_379_313 ();
 b15zdnd11an1n08x5 FILLER_379_325 ();
 b15zdnd00an1n02x5 FILLER_379_333 ();
 b15zdnd00an1n01x5 FILLER_379_335 ();
 b15zdnd11an1n04x5 FILLER_379_341 ();
 b15zdnd11an1n64x5 FILLER_379_351 ();
 b15zdnd11an1n16x5 FILLER_379_415 ();
 b15zdnd11an1n04x5 FILLER_379_431 ();
 b15zdnd00an1n02x5 FILLER_379_435 ();
 b15zdnd00an1n01x5 FILLER_379_437 ();
 b15zdnd11an1n04x5 FILLER_379_445 ();
 b15zdnd11an1n16x5 FILLER_379_454 ();
 b15zdnd00an1n01x5 FILLER_379_470 ();
 b15zdnd11an1n32x5 FILLER_379_478 ();
 b15zdnd11an1n32x5 FILLER_379_520 ();
 b15zdnd11an1n08x5 FILLER_379_552 ();
 b15zdnd11an1n32x5 FILLER_379_570 ();
 b15zdnd11an1n16x5 FILLER_379_602 ();
 b15zdnd11an1n08x5 FILLER_379_618 ();
 b15zdnd11an1n04x5 FILLER_379_626 ();
 b15zdnd11an1n16x5 FILLER_379_654 ();
 b15zdnd00an1n02x5 FILLER_379_670 ();
 b15zdnd11an1n04x5 FILLER_379_677 ();
 b15zdnd11an1n04x5 FILLER_379_685 ();
 b15zdnd11an1n32x5 FILLER_379_705 ();
 b15zdnd11an1n08x5 FILLER_379_737 ();
 b15zdnd11an1n04x5 FILLER_379_745 ();
 b15zdnd11an1n16x5 FILLER_379_754 ();
 b15zdnd11an1n04x5 FILLER_379_770 ();
 b15zdnd11an1n16x5 FILLER_379_778 ();
 b15zdnd11an1n08x5 FILLER_379_794 ();
 b15zdnd11an1n04x5 FILLER_379_802 ();
 b15zdnd11an1n08x5 FILLER_379_817 ();
 b15zdnd00an1n02x5 FILLER_379_825 ();
 b15zdnd11an1n16x5 FILLER_379_838 ();
 b15zdnd00an1n02x5 FILLER_379_854 ();
 b15zdnd11an1n04x5 FILLER_379_865 ();
 b15zdnd11an1n04x5 FILLER_379_874 ();
 b15zdnd00an1n02x5 FILLER_379_878 ();
 b15zdnd11an1n04x5 FILLER_379_890 ();
 b15zdnd11an1n04x5 FILLER_379_898 ();
 b15zdnd00an1n01x5 FILLER_379_902 ();
 b15zdnd11an1n08x5 FILLER_379_909 ();
 b15zdnd00an1n01x5 FILLER_379_917 ();
 b15zdnd11an1n16x5 FILLER_379_928 ();
 b15zdnd00an1n01x5 FILLER_379_944 ();
 b15zdnd11an1n04x5 FILLER_379_952 ();
 b15zdnd00an1n01x5 FILLER_379_956 ();
 b15zdnd11an1n08x5 FILLER_379_978 ();
 b15zdnd11an1n08x5 FILLER_379_999 ();
 b15zdnd11an1n04x5 FILLER_379_1007 ();
 b15zdnd00an1n02x5 FILLER_379_1011 ();
 b15zdnd00an1n01x5 FILLER_379_1013 ();
 b15zdnd11an1n08x5 FILLER_379_1018 ();
 b15zdnd11an1n04x5 FILLER_379_1026 ();
 b15zdnd11an1n16x5 FILLER_379_1038 ();
 b15zdnd11an1n08x5 FILLER_379_1054 ();
 b15zdnd00an1n02x5 FILLER_379_1062 ();
 b15zdnd00an1n01x5 FILLER_379_1064 ();
 b15zdnd11an1n04x5 FILLER_379_1077 ();
 b15zdnd00an1n02x5 FILLER_379_1081 ();
 b15zdnd11an1n08x5 FILLER_379_1091 ();
 b15zdnd11an1n04x5 FILLER_379_1099 ();
 b15zdnd11an1n16x5 FILLER_379_1119 ();
 b15zdnd11an1n04x5 FILLER_379_1141 ();
 b15zdnd11an1n08x5 FILLER_379_1161 ();
 b15zdnd11an1n04x5 FILLER_379_1169 ();
 b15zdnd11an1n64x5 FILLER_379_1205 ();
 b15zdnd11an1n64x5 FILLER_379_1269 ();
 b15zdnd00an1n02x5 FILLER_379_1333 ();
 b15zdnd11an1n32x5 FILLER_379_1351 ();
 b15zdnd11an1n08x5 FILLER_379_1383 ();
 b15zdnd11an1n04x5 FILLER_379_1391 ();
 b15zdnd00an1n01x5 FILLER_379_1395 ();
 b15zdnd11an1n16x5 FILLER_379_1401 ();
 b15zdnd11an1n32x5 FILLER_379_1425 ();
 b15zdnd11an1n08x5 FILLER_379_1457 ();
 b15zdnd11an1n04x5 FILLER_379_1465 ();
 b15zdnd00an1n02x5 FILLER_379_1469 ();
 b15zdnd11an1n04x5 FILLER_379_1479 ();
 b15zdnd11an1n64x5 FILLER_379_1488 ();
 b15zdnd11an1n32x5 FILLER_379_1552 ();
 b15zdnd11an1n04x5 FILLER_379_1584 ();
 b15zdnd00an1n02x5 FILLER_379_1588 ();
 b15zdnd00an1n01x5 FILLER_379_1590 ();
 b15zdnd11an1n04x5 FILLER_379_1601 ();
 b15zdnd11an1n16x5 FILLER_379_1617 ();
 b15zdnd11an1n08x5 FILLER_379_1633 ();
 b15zdnd11an1n04x5 FILLER_379_1641 ();
 b15zdnd00an1n02x5 FILLER_379_1645 ();
 b15zdnd00an1n01x5 FILLER_379_1647 ();
 b15zdnd11an1n32x5 FILLER_379_1661 ();
 b15zdnd11an1n04x5 FILLER_379_1693 ();
 b15zdnd00an1n01x5 FILLER_379_1697 ();
 b15zdnd11an1n64x5 FILLER_379_1716 ();
 b15zdnd11an1n64x5 FILLER_379_1780 ();
 b15zdnd11an1n64x5 FILLER_379_1844 ();
 b15zdnd11an1n64x5 FILLER_379_1908 ();
 b15zdnd11an1n64x5 FILLER_379_1972 ();
 b15zdnd11an1n04x5 FILLER_379_2036 ();
 b15zdnd00an1n01x5 FILLER_379_2040 ();
 b15zdnd11an1n32x5 FILLER_379_2049 ();
 b15zdnd11an1n04x5 FILLER_379_2081 ();
 b15zdnd11an1n04x5 FILLER_379_2091 ();
 b15zdnd11an1n64x5 FILLER_379_2101 ();
 b15zdnd11an1n32x5 FILLER_379_2165 ();
 b15zdnd00an1n01x5 FILLER_379_2197 ();
 b15zdnd11an1n08x5 FILLER_379_2214 ();
 b15zdnd00an1n02x5 FILLER_379_2222 ();
 b15zdnd00an1n01x5 FILLER_379_2224 ();
 b15zdnd11an1n32x5 FILLER_379_2239 ();
 b15zdnd11an1n08x5 FILLER_379_2271 ();
 b15zdnd11an1n04x5 FILLER_379_2279 ();
 b15zdnd00an1n01x5 FILLER_379_2283 ();
 b15zdnd11an1n64x5 FILLER_380_8 ();
 b15zdnd11an1n64x5 FILLER_380_72 ();
 b15zdnd11an1n64x5 FILLER_380_136 ();
 b15zdnd11an1n64x5 FILLER_380_200 ();
 b15zdnd11an1n08x5 FILLER_380_264 ();
 b15zdnd11an1n64x5 FILLER_380_288 ();
 b15zdnd11an1n32x5 FILLER_380_352 ();
 b15zdnd11an1n08x5 FILLER_380_384 ();
 b15zdnd11an1n04x5 FILLER_380_392 ();
 b15zdnd11an1n32x5 FILLER_380_404 ();
 b15zdnd11an1n04x5 FILLER_380_436 ();
 b15zdnd00an1n01x5 FILLER_380_440 ();
 b15zdnd11an1n64x5 FILLER_380_445 ();
 b15zdnd11an1n16x5 FILLER_380_509 ();
 b15zdnd00an1n02x5 FILLER_380_525 ();
 b15zdnd00an1n01x5 FILLER_380_527 ();
 b15zdnd11an1n16x5 FILLER_380_532 ();
 b15zdnd11an1n08x5 FILLER_380_548 ();
 b15zdnd11an1n04x5 FILLER_380_556 ();
 b15zdnd00an1n01x5 FILLER_380_560 ();
 b15zdnd11an1n64x5 FILLER_380_573 ();
 b15zdnd11an1n08x5 FILLER_380_637 ();
 b15zdnd00an1n01x5 FILLER_380_645 ();
 b15zdnd11an1n32x5 FILLER_380_658 ();
 b15zdnd11an1n08x5 FILLER_380_690 ();
 b15zdnd11an1n04x5 FILLER_380_698 ();
 b15zdnd11an1n08x5 FILLER_380_706 ();
 b15zdnd11an1n04x5 FILLER_380_714 ();
 b15zdnd11an1n64x5 FILLER_380_726 ();
 b15zdnd00an1n02x5 FILLER_380_790 ();
 b15zdnd11an1n16x5 FILLER_380_801 ();
 b15zdnd11an1n08x5 FILLER_380_817 ();
 b15zdnd11an1n04x5 FILLER_380_830 ();
 b15zdnd11an1n32x5 FILLER_380_839 ();
 b15zdnd11an1n04x5 FILLER_380_878 ();
 b15zdnd11an1n64x5 FILLER_380_887 ();
 b15zdnd11an1n16x5 FILLER_380_951 ();
 b15zdnd00an1n02x5 FILLER_380_967 ();
 b15zdnd00an1n01x5 FILLER_380_969 ();
 b15zdnd11an1n08x5 FILLER_380_980 ();
 b15zdnd00an1n02x5 FILLER_380_988 ();
 b15zdnd00an1n01x5 FILLER_380_990 ();
 b15zdnd11an1n04x5 FILLER_380_998 ();
 b15zdnd11an1n08x5 FILLER_380_1007 ();
 b15zdnd00an1n01x5 FILLER_380_1015 ();
 b15zdnd11an1n04x5 FILLER_380_1040 ();
 b15zdnd11an1n04x5 FILLER_380_1048 ();
 b15zdnd11an1n16x5 FILLER_380_1068 ();
 b15zdnd11an1n08x5 FILLER_380_1084 ();
 b15zdnd00an1n02x5 FILLER_380_1092 ();
 b15zdnd00an1n01x5 FILLER_380_1094 ();
 b15zdnd11an1n04x5 FILLER_380_1119 ();
 b15zdnd11an1n16x5 FILLER_380_1139 ();
 b15zdnd11an1n04x5 FILLER_380_1155 ();
 b15zdnd00an1n02x5 FILLER_380_1159 ();
 b15zdnd00an1n01x5 FILLER_380_1161 ();
 b15zdnd11an1n64x5 FILLER_380_1178 ();
 b15zdnd11an1n64x5 FILLER_380_1242 ();
 b15zdnd11an1n64x5 FILLER_380_1306 ();
 b15zdnd11an1n64x5 FILLER_380_1370 ();
 b15zdnd11an1n32x5 FILLER_380_1434 ();
 b15zdnd11an1n04x5 FILLER_380_1466 ();
 b15zdnd00an1n01x5 FILLER_380_1470 ();
 b15zdnd11an1n32x5 FILLER_380_1476 ();
 b15zdnd11an1n64x5 FILLER_380_1514 ();
 b15zdnd11an1n04x5 FILLER_380_1578 ();
 b15zdnd00an1n01x5 FILLER_380_1582 ();
 b15zdnd11an1n32x5 FILLER_380_1589 ();
 b15zdnd11an1n16x5 FILLER_380_1621 ();
 b15zdnd11an1n08x5 FILLER_380_1637 ();
 b15zdnd00an1n02x5 FILLER_380_1645 ();
 b15zdnd00an1n01x5 FILLER_380_1647 ();
 b15zdnd11an1n32x5 FILLER_380_1655 ();
 b15zdnd11an1n04x5 FILLER_380_1687 ();
 b15zdnd00an1n02x5 FILLER_380_1691 ();
 b15zdnd00an1n01x5 FILLER_380_1693 ();
 b15zdnd11an1n64x5 FILLER_380_1726 ();
 b15zdnd11an1n32x5 FILLER_380_1790 ();
 b15zdnd11an1n04x5 FILLER_380_1822 ();
 b15zdnd00an1n02x5 FILLER_380_1826 ();
 b15zdnd00an1n01x5 FILLER_380_1828 ();
 b15zdnd11an1n04x5 FILLER_380_1845 ();
 b15zdnd11an1n08x5 FILLER_380_1867 ();
 b15zdnd00an1n01x5 FILLER_380_1875 ();
 b15zdnd11an1n04x5 FILLER_380_1885 ();
 b15zdnd00an1n01x5 FILLER_380_1889 ();
 b15zdnd11an1n32x5 FILLER_380_1896 ();
 b15zdnd11an1n16x5 FILLER_380_1928 ();
 b15zdnd00an1n02x5 FILLER_380_1944 ();
 b15zdnd00an1n01x5 FILLER_380_1946 ();
 b15zdnd11an1n32x5 FILLER_380_1960 ();
 b15zdnd11an1n08x5 FILLER_380_1992 ();
 b15zdnd11an1n32x5 FILLER_380_2006 ();
 b15zdnd11an1n04x5 FILLER_380_2038 ();
 b15zdnd00an1n01x5 FILLER_380_2042 ();
 b15zdnd11an1n64x5 FILLER_380_2048 ();
 b15zdnd11an1n32x5 FILLER_380_2112 ();
 b15zdnd11an1n08x5 FILLER_380_2144 ();
 b15zdnd00an1n02x5 FILLER_380_2152 ();
 b15zdnd00an1n02x5 FILLER_380_2162 ();
 b15zdnd11an1n16x5 FILLER_380_2185 ();
 b15zdnd11an1n04x5 FILLER_380_2201 ();
 b15zdnd11an1n32x5 FILLER_380_2223 ();
 b15zdnd11an1n16x5 FILLER_380_2255 ();
 b15zdnd11an1n04x5 FILLER_380_2271 ();
 b15zdnd00an1n01x5 FILLER_380_2275 ();
 b15zdnd11an1n64x5 FILLER_381_0 ();
 b15zdnd11an1n64x5 FILLER_381_64 ();
 b15zdnd11an1n64x5 FILLER_381_128 ();
 b15zdnd11an1n64x5 FILLER_381_192 ();
 b15zdnd11an1n32x5 FILLER_381_256 ();
 b15zdnd11an1n16x5 FILLER_381_288 ();
 b15zdnd00an1n01x5 FILLER_381_304 ();
 b15zdnd11an1n08x5 FILLER_381_321 ();
 b15zdnd00an1n02x5 FILLER_381_329 ();
 b15zdnd00an1n01x5 FILLER_381_331 ();
 b15zdnd11an1n16x5 FILLER_381_352 ();
 b15zdnd00an1n02x5 FILLER_381_368 ();
 b15zdnd11an1n08x5 FILLER_381_382 ();
 b15zdnd11an1n04x5 FILLER_381_390 ();
 b15zdnd00an1n01x5 FILLER_381_394 ();
 b15zdnd11an1n04x5 FILLER_381_405 ();
 b15zdnd00an1n01x5 FILLER_381_409 ();
 b15zdnd11an1n08x5 FILLER_381_422 ();
 b15zdnd00an1n02x5 FILLER_381_430 ();
 b15zdnd00an1n01x5 FILLER_381_432 ();
 b15zdnd11an1n16x5 FILLER_381_447 ();
 b15zdnd11an1n04x5 FILLER_381_463 ();
 b15zdnd00an1n01x5 FILLER_381_467 ();
 b15zdnd11an1n16x5 FILLER_381_473 ();
 b15zdnd11an1n08x5 FILLER_381_489 ();
 b15zdnd11an1n04x5 FILLER_381_497 ();
 b15zdnd00an1n02x5 FILLER_381_501 ();
 b15zdnd11an1n08x5 FILLER_381_512 ();
 b15zdnd11an1n04x5 FILLER_381_520 ();
 b15zdnd00an1n01x5 FILLER_381_524 ();
 b15zdnd11an1n08x5 FILLER_381_532 ();
 b15zdnd00an1n01x5 FILLER_381_540 ();
 b15zdnd11an1n04x5 FILLER_381_553 ();
 b15zdnd11an1n16x5 FILLER_381_565 ();
 b15zdnd11an1n32x5 FILLER_381_597 ();
 b15zdnd11an1n04x5 FILLER_381_645 ();
 b15zdnd11an1n16x5 FILLER_381_667 ();
 b15zdnd11an1n08x5 FILLER_381_683 ();
 b15zdnd00an1n02x5 FILLER_381_691 ();
 b15zdnd00an1n01x5 FILLER_381_693 ();
 b15zdnd11an1n16x5 FILLER_381_700 ();
 b15zdnd00an1n02x5 FILLER_381_716 ();
 b15zdnd00an1n01x5 FILLER_381_718 ();
 b15zdnd11an1n64x5 FILLER_381_725 ();
 b15zdnd11an1n64x5 FILLER_381_789 ();
 b15zdnd11an1n32x5 FILLER_381_853 ();
 b15zdnd11an1n08x5 FILLER_381_885 ();
 b15zdnd11an1n04x5 FILLER_381_893 ();
 b15zdnd00an1n02x5 FILLER_381_897 ();
 b15zdnd11an1n64x5 FILLER_381_907 ();
 b15zdnd11an1n16x5 FILLER_381_971 ();
 b15zdnd11an1n04x5 FILLER_381_987 ();
 b15zdnd11an1n04x5 FILLER_381_997 ();
 b15zdnd11an1n16x5 FILLER_381_1005 ();
 b15zdnd11an1n04x5 FILLER_381_1021 ();
 b15zdnd00an1n02x5 FILLER_381_1025 ();
 b15zdnd11an1n32x5 FILLER_381_1039 ();
 b15zdnd11an1n08x5 FILLER_381_1071 ();
 b15zdnd11an1n64x5 FILLER_381_1095 ();
 b15zdnd11an1n64x5 FILLER_381_1159 ();
 b15zdnd11an1n64x5 FILLER_381_1223 ();
 b15zdnd11an1n64x5 FILLER_381_1287 ();
 b15zdnd11an1n32x5 FILLER_381_1351 ();
 b15zdnd00an1n02x5 FILLER_381_1383 ();
 b15zdnd11an1n64x5 FILLER_381_1399 ();
 b15zdnd11an1n04x5 FILLER_381_1463 ();
 b15zdnd00an1n02x5 FILLER_381_1467 ();
 b15zdnd00an1n01x5 FILLER_381_1469 ();
 b15zdnd11an1n16x5 FILLER_381_1474 ();
 b15zdnd11an1n08x5 FILLER_381_1490 ();
 b15zdnd00an1n01x5 FILLER_381_1498 ();
 b15zdnd11an1n04x5 FILLER_381_1505 ();
 b15zdnd11an1n16x5 FILLER_381_1513 ();
 b15zdnd00an1n02x5 FILLER_381_1529 ();
 b15zdnd11an1n32x5 FILLER_381_1536 ();
 b15zdnd11an1n16x5 FILLER_381_1568 ();
 b15zdnd00an1n01x5 FILLER_381_1584 ();
 b15zdnd11an1n16x5 FILLER_381_1598 ();
 b15zdnd11an1n04x5 FILLER_381_1614 ();
 b15zdnd00an1n02x5 FILLER_381_1618 ();
 b15zdnd11an1n16x5 FILLER_381_1626 ();
 b15zdnd11an1n04x5 FILLER_381_1642 ();
 b15zdnd00an1n02x5 FILLER_381_1646 ();
 b15zdnd11an1n08x5 FILLER_381_1655 ();
 b15zdnd11an1n04x5 FILLER_381_1663 ();
 b15zdnd00an1n02x5 FILLER_381_1667 ();
 b15zdnd00an1n01x5 FILLER_381_1669 ();
 b15zdnd11an1n04x5 FILLER_381_1688 ();
 b15zdnd00an1n02x5 FILLER_381_1692 ();
 b15zdnd00an1n01x5 FILLER_381_1694 ();
 b15zdnd11an1n04x5 FILLER_381_1707 ();
 b15zdnd11an1n64x5 FILLER_381_1728 ();
 b15zdnd11an1n32x5 FILLER_381_1792 ();
 b15zdnd11an1n16x5 FILLER_381_1824 ();
 b15zdnd11an1n08x5 FILLER_381_1840 ();
 b15zdnd00an1n02x5 FILLER_381_1848 ();
 b15zdnd00an1n01x5 FILLER_381_1850 ();
 b15zdnd11an1n08x5 FILLER_381_1857 ();
 b15zdnd00an1n02x5 FILLER_381_1865 ();
 b15zdnd11an1n04x5 FILLER_381_1873 ();
 b15zdnd11an1n64x5 FILLER_381_1889 ();
 b15zdnd11an1n16x5 FILLER_381_1953 ();
 b15zdnd00an1n01x5 FILLER_381_1969 ();
 b15zdnd11an1n16x5 FILLER_381_1976 ();
 b15zdnd00an1n02x5 FILLER_381_1992 ();
 b15zdnd11an1n04x5 FILLER_381_1999 ();
 b15zdnd11an1n64x5 FILLER_381_2009 ();
 b15zdnd11an1n16x5 FILLER_381_2073 ();
 b15zdnd11an1n04x5 FILLER_381_2089 ();
 b15zdnd00an1n01x5 FILLER_381_2093 ();
 b15zdnd11an1n16x5 FILLER_381_2104 ();
 b15zdnd11an1n08x5 FILLER_381_2120 ();
 b15zdnd00an1n02x5 FILLER_381_2128 ();
 b15zdnd11an1n64x5 FILLER_381_2135 ();
 b15zdnd11an1n64x5 FILLER_381_2199 ();
 b15zdnd11an1n16x5 FILLER_381_2263 ();
 b15zdnd11an1n04x5 FILLER_381_2279 ();
 b15zdnd00an1n01x5 FILLER_381_2283 ();
 b15zdnd11an1n64x5 FILLER_382_8 ();
 b15zdnd11an1n64x5 FILLER_382_72 ();
 b15zdnd11an1n64x5 FILLER_382_136 ();
 b15zdnd11an1n64x5 FILLER_382_200 ();
 b15zdnd11an1n64x5 FILLER_382_264 ();
 b15zdnd11an1n64x5 FILLER_382_328 ();
 b15zdnd11an1n08x5 FILLER_382_392 ();
 b15zdnd11an1n16x5 FILLER_382_406 ();
 b15zdnd11an1n04x5 FILLER_382_422 ();
 b15zdnd00an1n02x5 FILLER_382_426 ();
 b15zdnd00an1n01x5 FILLER_382_428 ();
 b15zdnd11an1n04x5 FILLER_382_436 ();
 b15zdnd11an1n32x5 FILLER_382_444 ();
 b15zdnd11an1n16x5 FILLER_382_476 ();
 b15zdnd11an1n08x5 FILLER_382_515 ();
 b15zdnd00an1n02x5 FILLER_382_523 ();
 b15zdnd00an1n01x5 FILLER_382_525 ();
 b15zdnd11an1n16x5 FILLER_382_530 ();
 b15zdnd11an1n08x5 FILLER_382_546 ();
 b15zdnd00an1n01x5 FILLER_382_554 ();
 b15zdnd11an1n64x5 FILLER_382_567 ();
 b15zdnd11an1n08x5 FILLER_382_631 ();
 b15zdnd11an1n04x5 FILLER_382_639 ();
 b15zdnd00an1n01x5 FILLER_382_643 ();
 b15zdnd11an1n04x5 FILLER_382_666 ();
 b15zdnd00an1n02x5 FILLER_382_670 ();
 b15zdnd00an1n01x5 FILLER_382_672 ();
 b15zdnd11an1n32x5 FILLER_382_685 ();
 b15zdnd00an1n01x5 FILLER_382_717 ();
 b15zdnd11an1n64x5 FILLER_382_726 ();
 b15zdnd11an1n04x5 FILLER_382_790 ();
 b15zdnd00an1n01x5 FILLER_382_794 ();
 b15zdnd11an1n64x5 FILLER_382_805 ();
 b15zdnd11an1n64x5 FILLER_382_869 ();
 b15zdnd11an1n64x5 FILLER_382_933 ();
 b15zdnd11an1n32x5 FILLER_382_997 ();
 b15zdnd11an1n08x5 FILLER_382_1029 ();
 b15zdnd11an1n04x5 FILLER_382_1037 ();
 b15zdnd11an1n64x5 FILLER_382_1053 ();
 b15zdnd11an1n08x5 FILLER_382_1117 ();
 b15zdnd11an1n64x5 FILLER_382_1146 ();
 b15zdnd11an1n64x5 FILLER_382_1210 ();
 b15zdnd11an1n32x5 FILLER_382_1274 ();
 b15zdnd11an1n08x5 FILLER_382_1306 ();
 b15zdnd11an1n04x5 FILLER_382_1314 ();
 b15zdnd00an1n01x5 FILLER_382_1318 ();
 b15zdnd11an1n04x5 FILLER_382_1333 ();
 b15zdnd11an1n32x5 FILLER_382_1353 ();
 b15zdnd11an1n08x5 FILLER_382_1385 ();
 b15zdnd00an1n02x5 FILLER_382_1393 ();
 b15zdnd11an1n16x5 FILLER_382_1400 ();
 b15zdnd11an1n04x5 FILLER_382_1416 ();
 b15zdnd00an1n02x5 FILLER_382_1420 ();
 b15zdnd11an1n16x5 FILLER_382_1430 ();
 b15zdnd11an1n04x5 FILLER_382_1446 ();
 b15zdnd00an1n02x5 FILLER_382_1450 ();
 b15zdnd00an1n01x5 FILLER_382_1452 ();
 b15zdnd11an1n04x5 FILLER_382_1469 ();
 b15zdnd11an1n32x5 FILLER_382_1478 ();
 b15zdnd11an1n32x5 FILLER_382_1520 ();
 b15zdnd11an1n16x5 FILLER_382_1552 ();
 b15zdnd11an1n08x5 FILLER_382_1568 ();
 b15zdnd00an1n02x5 FILLER_382_1576 ();
 b15zdnd11an1n32x5 FILLER_382_1594 ();
 b15zdnd11an1n64x5 FILLER_382_1631 ();
 b15zdnd11an1n64x5 FILLER_382_1695 ();
 b15zdnd11an1n32x5 FILLER_382_1759 ();
 b15zdnd11an1n16x5 FILLER_382_1791 ();
 b15zdnd00an1n02x5 FILLER_382_1807 ();
 b15zdnd11an1n64x5 FILLER_382_1825 ();
 b15zdnd11an1n04x5 FILLER_382_1889 ();
 b15zdnd11an1n16x5 FILLER_382_1908 ();
 b15zdnd00an1n02x5 FILLER_382_1924 ();
 b15zdnd00an1n01x5 FILLER_382_1926 ();
 b15zdnd11an1n32x5 FILLER_382_1931 ();
 b15zdnd11an1n04x5 FILLER_382_1963 ();
 b15zdnd11an1n16x5 FILLER_382_1979 ();
 b15zdnd11an1n08x5 FILLER_382_1995 ();
 b15zdnd11an1n16x5 FILLER_382_2017 ();
 b15zdnd00an1n01x5 FILLER_382_2033 ();
 b15zdnd11an1n64x5 FILLER_382_2046 ();
 b15zdnd11an1n16x5 FILLER_382_2110 ();
 b15zdnd11an1n04x5 FILLER_382_2126 ();
 b15zdnd00an1n01x5 FILLER_382_2130 ();
 b15zdnd11an1n08x5 FILLER_382_2141 ();
 b15zdnd11an1n04x5 FILLER_382_2149 ();
 b15zdnd00an1n01x5 FILLER_382_2153 ();
 b15zdnd11an1n16x5 FILLER_382_2162 ();
 b15zdnd11an1n04x5 FILLER_382_2178 ();
 b15zdnd00an1n01x5 FILLER_382_2182 ();
 b15zdnd11an1n04x5 FILLER_382_2215 ();
 b15zdnd11an1n32x5 FILLER_382_2236 ();
 b15zdnd11an1n08x5 FILLER_382_2268 ();
 b15zdnd11an1n64x5 FILLER_383_0 ();
 b15zdnd11an1n64x5 FILLER_383_64 ();
 b15zdnd11an1n64x5 FILLER_383_128 ();
 b15zdnd11an1n64x5 FILLER_383_192 ();
 b15zdnd11an1n64x5 FILLER_383_256 ();
 b15zdnd11an1n64x5 FILLER_383_320 ();
 b15zdnd11an1n64x5 FILLER_383_384 ();
 b15zdnd11an1n32x5 FILLER_383_448 ();
 b15zdnd11an1n16x5 FILLER_383_480 ();
 b15zdnd11an1n04x5 FILLER_383_496 ();
 b15zdnd00an1n02x5 FILLER_383_500 ();
 b15zdnd00an1n01x5 FILLER_383_502 ();
 b15zdnd11an1n64x5 FILLER_383_508 ();
 b15zdnd11an1n64x5 FILLER_383_572 ();
 b15zdnd11an1n16x5 FILLER_383_636 ();
 b15zdnd11an1n08x5 FILLER_383_652 ();
 b15zdnd00an1n01x5 FILLER_383_660 ();
 b15zdnd11an1n16x5 FILLER_383_684 ();
 b15zdnd11an1n08x5 FILLER_383_700 ();
 b15zdnd00an1n02x5 FILLER_383_708 ();
 b15zdnd11an1n08x5 FILLER_383_717 ();
 b15zdnd11an1n04x5 FILLER_383_725 ();
 b15zdnd00an1n02x5 FILLER_383_729 ();
 b15zdnd11an1n04x5 FILLER_383_737 ();
 b15zdnd00an1n02x5 FILLER_383_741 ();
 b15zdnd00an1n01x5 FILLER_383_743 ();
 b15zdnd11an1n04x5 FILLER_383_750 ();
 b15zdnd11an1n16x5 FILLER_383_770 ();
 b15zdnd11an1n08x5 FILLER_383_786 ();
 b15zdnd00an1n02x5 FILLER_383_794 ();
 b15zdnd00an1n01x5 FILLER_383_796 ();
 b15zdnd11an1n64x5 FILLER_383_803 ();
 b15zdnd11an1n04x5 FILLER_383_867 ();
 b15zdnd11an1n64x5 FILLER_383_878 ();
 b15zdnd11an1n64x5 FILLER_383_942 ();
 b15zdnd11an1n32x5 FILLER_383_1006 ();
 b15zdnd11an1n08x5 FILLER_383_1038 ();
 b15zdnd11an1n64x5 FILLER_383_1061 ();
 b15zdnd11an1n08x5 FILLER_383_1125 ();
 b15zdnd00an1n01x5 FILLER_383_1133 ();
 b15zdnd11an1n04x5 FILLER_383_1143 ();
 b15zdnd00an1n02x5 FILLER_383_1147 ();
 b15zdnd00an1n01x5 FILLER_383_1149 ();
 b15zdnd11an1n64x5 FILLER_383_1173 ();
 b15zdnd11an1n64x5 FILLER_383_1237 ();
 b15zdnd11an1n32x5 FILLER_383_1301 ();
 b15zdnd11an1n04x5 FILLER_383_1333 ();
 b15zdnd00an1n01x5 FILLER_383_1337 ();
 b15zdnd11an1n04x5 FILLER_383_1344 ();
 b15zdnd11an1n08x5 FILLER_383_1358 ();
 b15zdnd00an1n02x5 FILLER_383_1366 ();
 b15zdnd11an1n16x5 FILLER_383_1384 ();
 b15zdnd11an1n08x5 FILLER_383_1400 ();
 b15zdnd00an1n02x5 FILLER_383_1408 ();
 b15zdnd11an1n04x5 FILLER_383_1416 ();
 b15zdnd00an1n02x5 FILLER_383_1420 ();
 b15zdnd11an1n32x5 FILLER_383_1434 ();
 b15zdnd11an1n08x5 FILLER_383_1466 ();
 b15zdnd11an1n16x5 FILLER_383_1480 ();
 b15zdnd11an1n08x5 FILLER_383_1496 ();
 b15zdnd11an1n04x5 FILLER_383_1504 ();
 b15zdnd00an1n02x5 FILLER_383_1508 ();
 b15zdnd00an1n01x5 FILLER_383_1510 ();
 b15zdnd11an1n16x5 FILLER_383_1517 ();
 b15zdnd11an1n08x5 FILLER_383_1533 ();
 b15zdnd00an1n02x5 FILLER_383_1541 ();
 b15zdnd00an1n01x5 FILLER_383_1543 ();
 b15zdnd11an1n16x5 FILLER_383_1555 ();
 b15zdnd11an1n08x5 FILLER_383_1571 ();
 b15zdnd11an1n04x5 FILLER_383_1579 ();
 b15zdnd00an1n02x5 FILLER_383_1583 ();
 b15zdnd11an1n32x5 FILLER_383_1591 ();
 b15zdnd11an1n16x5 FILLER_383_1623 ();
 b15zdnd11an1n08x5 FILLER_383_1639 ();
 b15zdnd11an1n04x5 FILLER_383_1647 ();
 b15zdnd00an1n02x5 FILLER_383_1651 ();
 b15zdnd00an1n01x5 FILLER_383_1653 ();
 b15zdnd11an1n04x5 FILLER_383_1672 ();
 b15zdnd11an1n64x5 FILLER_383_1707 ();
 b15zdnd11an1n64x5 FILLER_383_1771 ();
 b15zdnd00an1n02x5 FILLER_383_1835 ();
 b15zdnd00an1n01x5 FILLER_383_1837 ();
 b15zdnd11an1n04x5 FILLER_383_1854 ();
 b15zdnd11an1n08x5 FILLER_383_1874 ();
 b15zdnd11an1n04x5 FILLER_383_1882 ();
 b15zdnd00an1n02x5 FILLER_383_1886 ();
 b15zdnd00an1n01x5 FILLER_383_1888 ();
 b15zdnd11an1n32x5 FILLER_383_1896 ();
 b15zdnd11an1n08x5 FILLER_383_1928 ();
 b15zdnd00an1n01x5 FILLER_383_1936 ();
 b15zdnd11an1n64x5 FILLER_383_1942 ();
 b15zdnd11an1n16x5 FILLER_383_2006 ();
 b15zdnd11an1n08x5 FILLER_383_2022 ();
 b15zdnd11an1n04x5 FILLER_383_2030 ();
 b15zdnd00an1n02x5 FILLER_383_2034 ();
 b15zdnd11an1n04x5 FILLER_383_2045 ();
 b15zdnd00an1n02x5 FILLER_383_2049 ();
 b15zdnd11an1n08x5 FILLER_383_2058 ();
 b15zdnd00an1n01x5 FILLER_383_2066 ();
 b15zdnd11an1n08x5 FILLER_383_2071 ();
 b15zdnd11an1n04x5 FILLER_383_2079 ();
 b15zdnd11an1n32x5 FILLER_383_2091 ();
 b15zdnd11an1n04x5 FILLER_383_2123 ();
 b15zdnd11an1n32x5 FILLER_383_2132 ();
 b15zdnd11an1n04x5 FILLER_383_2164 ();
 b15zdnd11an1n04x5 FILLER_383_2184 ();
 b15zdnd11an1n64x5 FILLER_383_2204 ();
 b15zdnd11an1n16x5 FILLER_383_2268 ();
 b15zdnd11an1n64x5 FILLER_384_8 ();
 b15zdnd11an1n64x5 FILLER_384_72 ();
 b15zdnd11an1n64x5 FILLER_384_136 ();
 b15zdnd11an1n64x5 FILLER_384_200 ();
 b15zdnd11an1n64x5 FILLER_384_264 ();
 b15zdnd11an1n64x5 FILLER_384_328 ();
 b15zdnd11an1n64x5 FILLER_384_392 ();
 b15zdnd11an1n64x5 FILLER_384_456 ();
 b15zdnd11an1n64x5 FILLER_384_520 ();
 b15zdnd11an1n64x5 FILLER_384_584 ();
 b15zdnd11an1n16x5 FILLER_384_648 ();
 b15zdnd11an1n04x5 FILLER_384_664 ();
 b15zdnd00an1n01x5 FILLER_384_668 ();
 b15zdnd11an1n32x5 FILLER_384_685 ();
 b15zdnd00an1n01x5 FILLER_384_717 ();
 b15zdnd11an1n08x5 FILLER_384_726 ();
 b15zdnd00an1n02x5 FILLER_384_734 ();
 b15zdnd11an1n04x5 FILLER_384_754 ();
 b15zdnd11an1n16x5 FILLER_384_762 ();
 b15zdnd11an1n08x5 FILLER_384_778 ();
 b15zdnd11an1n04x5 FILLER_384_786 ();
 b15zdnd00an1n01x5 FILLER_384_790 ();
 b15zdnd11an1n32x5 FILLER_384_803 ();
 b15zdnd11an1n08x5 FILLER_384_835 ();
 b15zdnd00an1n01x5 FILLER_384_843 ();
 b15zdnd11an1n64x5 FILLER_384_854 ();
 b15zdnd11an1n32x5 FILLER_384_918 ();
 b15zdnd11an1n04x5 FILLER_384_950 ();
 b15zdnd00an1n02x5 FILLER_384_954 ();
 b15zdnd11an1n64x5 FILLER_384_966 ();
 b15zdnd11an1n16x5 FILLER_384_1030 ();
 b15zdnd11an1n04x5 FILLER_384_1046 ();
 b15zdnd00an1n01x5 FILLER_384_1050 ();
 b15zdnd11an1n32x5 FILLER_384_1055 ();
 b15zdnd11an1n16x5 FILLER_384_1087 ();
 b15zdnd00an1n01x5 FILLER_384_1103 ();
 b15zdnd11an1n16x5 FILLER_384_1120 ();
 b15zdnd11an1n08x5 FILLER_384_1136 ();
 b15zdnd00an1n01x5 FILLER_384_1144 ();
 b15zdnd11an1n64x5 FILLER_384_1153 ();
 b15zdnd11an1n64x5 FILLER_384_1217 ();
 b15zdnd11an1n32x5 FILLER_384_1281 ();
 b15zdnd11an1n08x5 FILLER_384_1333 ();
 b15zdnd00an1n02x5 FILLER_384_1341 ();
 b15zdnd11an1n08x5 FILLER_384_1353 ();
 b15zdnd11an1n04x5 FILLER_384_1361 ();
 b15zdnd11an1n32x5 FILLER_384_1372 ();
 b15zdnd11an1n16x5 FILLER_384_1404 ();
 b15zdnd00an1n02x5 FILLER_384_1420 ();
 b15zdnd11an1n16x5 FILLER_384_1428 ();
 b15zdnd11an1n08x5 FILLER_384_1444 ();
 b15zdnd11an1n04x5 FILLER_384_1452 ();
 b15zdnd00an1n02x5 FILLER_384_1456 ();
 b15zdnd00an1n01x5 FILLER_384_1458 ();
 b15zdnd11an1n04x5 FILLER_384_1475 ();
 b15zdnd00an1n01x5 FILLER_384_1479 ();
 b15zdnd11an1n16x5 FILLER_384_1484 ();
 b15zdnd11an1n08x5 FILLER_384_1500 ();
 b15zdnd11an1n04x5 FILLER_384_1508 ();
 b15zdnd00an1n02x5 FILLER_384_1512 ();
 b15zdnd00an1n01x5 FILLER_384_1514 ();
 b15zdnd11an1n04x5 FILLER_384_1522 ();
 b15zdnd11an1n04x5 FILLER_384_1531 ();
 b15zdnd00an1n01x5 FILLER_384_1535 ();
 b15zdnd11an1n64x5 FILLER_384_1545 ();
 b15zdnd11an1n08x5 FILLER_384_1609 ();
 b15zdnd11an1n04x5 FILLER_384_1617 ();
 b15zdnd00an1n01x5 FILLER_384_1621 ();
 b15zdnd11an1n16x5 FILLER_384_1627 ();
 b15zdnd11an1n64x5 FILLER_384_1651 ();
 b15zdnd11an1n64x5 FILLER_384_1715 ();
 b15zdnd11an1n64x5 FILLER_384_1779 ();
 b15zdnd11an1n32x5 FILLER_384_1843 ();
 b15zdnd11an1n08x5 FILLER_384_1875 ();
 b15zdnd00an1n01x5 FILLER_384_1883 ();
 b15zdnd11an1n64x5 FILLER_384_1896 ();
 b15zdnd11an1n08x5 FILLER_384_1960 ();
 b15zdnd11an1n16x5 FILLER_384_1972 ();
 b15zdnd00an1n02x5 FILLER_384_1988 ();
 b15zdnd00an1n01x5 FILLER_384_1990 ();
 b15zdnd11an1n64x5 FILLER_384_1997 ();
 b15zdnd11an1n04x5 FILLER_384_2061 ();
 b15zdnd00an1n02x5 FILLER_384_2065 ();
 b15zdnd11an1n32x5 FILLER_384_2075 ();
 b15zdnd11an1n16x5 FILLER_384_2107 ();
 b15zdnd11an1n04x5 FILLER_384_2123 ();
 b15zdnd00an1n02x5 FILLER_384_2127 ();
 b15zdnd00an1n01x5 FILLER_384_2129 ();
 b15zdnd11an1n16x5 FILLER_384_2137 ();
 b15zdnd00an1n01x5 FILLER_384_2153 ();
 b15zdnd11an1n08x5 FILLER_384_2162 ();
 b15zdnd11an1n04x5 FILLER_384_2170 ();
 b15zdnd11an1n08x5 FILLER_384_2192 ();
 b15zdnd00an1n01x5 FILLER_384_2200 ();
 b15zdnd11an1n32x5 FILLER_384_2225 ();
 b15zdnd11an1n16x5 FILLER_384_2257 ();
 b15zdnd00an1n02x5 FILLER_384_2273 ();
 b15zdnd00an1n01x5 FILLER_384_2275 ();
 b15zdnd11an1n64x5 FILLER_385_0 ();
 b15zdnd11an1n64x5 FILLER_385_64 ();
 b15zdnd11an1n64x5 FILLER_385_128 ();
 b15zdnd11an1n64x5 FILLER_385_192 ();
 b15zdnd11an1n64x5 FILLER_385_256 ();
 b15zdnd11an1n64x5 FILLER_385_320 ();
 b15zdnd11an1n64x5 FILLER_385_384 ();
 b15zdnd11an1n64x5 FILLER_385_448 ();
 b15zdnd11an1n64x5 FILLER_385_512 ();
 b15zdnd11an1n64x5 FILLER_385_576 ();
 b15zdnd11an1n04x5 FILLER_385_640 ();
 b15zdnd11an1n08x5 FILLER_385_660 ();
 b15zdnd11an1n08x5 FILLER_385_676 ();
 b15zdnd11an1n04x5 FILLER_385_684 ();
 b15zdnd11an1n16x5 FILLER_385_694 ();
 b15zdnd11an1n04x5 FILLER_385_710 ();
 b15zdnd00an1n02x5 FILLER_385_714 ();
 b15zdnd11an1n16x5 FILLER_385_720 ();
 b15zdnd11an1n08x5 FILLER_385_736 ();
 b15zdnd00an1n02x5 FILLER_385_744 ();
 b15zdnd11an1n04x5 FILLER_385_750 ();
 b15zdnd11an1n04x5 FILLER_385_767 ();
 b15zdnd00an1n02x5 FILLER_385_771 ();
 b15zdnd11an1n08x5 FILLER_385_783 ();
 b15zdnd11an1n04x5 FILLER_385_791 ();
 b15zdnd00an1n02x5 FILLER_385_795 ();
 b15zdnd00an1n01x5 FILLER_385_797 ();
 b15zdnd11an1n08x5 FILLER_385_802 ();
 b15zdnd11an1n08x5 FILLER_385_819 ();
 b15zdnd11an1n04x5 FILLER_385_827 ();
 b15zdnd00an1n02x5 FILLER_385_831 ();
 b15zdnd00an1n01x5 FILLER_385_833 ();
 b15zdnd11an1n04x5 FILLER_385_850 ();
 b15zdnd11an1n16x5 FILLER_385_863 ();
 b15zdnd11an1n04x5 FILLER_385_893 ();
 b15zdnd00an1n02x5 FILLER_385_897 ();
 b15zdnd00an1n01x5 FILLER_385_899 ();
 b15zdnd11an1n04x5 FILLER_385_911 ();
 b15zdnd11an1n16x5 FILLER_385_921 ();
 b15zdnd11an1n08x5 FILLER_385_937 ();
 b15zdnd00an1n02x5 FILLER_385_945 ();
 b15zdnd11an1n08x5 FILLER_385_961 ();
 b15zdnd00an1n02x5 FILLER_385_969 ();
 b15zdnd11an1n04x5 FILLER_385_983 ();
 b15zdnd00an1n02x5 FILLER_385_987 ();
 b15zdnd11an1n08x5 FILLER_385_999 ();
 b15zdnd00an1n02x5 FILLER_385_1007 ();
 b15zdnd11an1n08x5 FILLER_385_1016 ();
 b15zdnd00an1n01x5 FILLER_385_1024 ();
 b15zdnd11an1n32x5 FILLER_385_1035 ();
 b15zdnd11an1n08x5 FILLER_385_1067 ();
 b15zdnd11an1n16x5 FILLER_385_1091 ();
 b15zdnd11an1n08x5 FILLER_385_1107 ();
 b15zdnd11an1n04x5 FILLER_385_1115 ();
 b15zdnd00an1n01x5 FILLER_385_1119 ();
 b15zdnd11an1n04x5 FILLER_385_1152 ();
 b15zdnd00an1n02x5 FILLER_385_1156 ();
 b15zdnd11an1n64x5 FILLER_385_1174 ();
 b15zdnd11an1n64x5 FILLER_385_1238 ();
 b15zdnd11an1n64x5 FILLER_385_1302 ();
 b15zdnd11an1n16x5 FILLER_385_1366 ();
 b15zdnd11an1n08x5 FILLER_385_1391 ();
 b15zdnd11an1n04x5 FILLER_385_1399 ();
 b15zdnd00an1n02x5 FILLER_385_1403 ();
 b15zdnd11an1n64x5 FILLER_385_1411 ();
 b15zdnd11an1n04x5 FILLER_385_1475 ();
 b15zdnd11an1n08x5 FILLER_385_1486 ();
 b15zdnd00an1n02x5 FILLER_385_1494 ();
 b15zdnd00an1n01x5 FILLER_385_1496 ();
 b15zdnd11an1n64x5 FILLER_385_1509 ();
 b15zdnd11an1n32x5 FILLER_385_1573 ();
 b15zdnd11an1n08x5 FILLER_385_1605 ();
 b15zdnd11an1n04x5 FILLER_385_1613 ();
 b15zdnd00an1n02x5 FILLER_385_1617 ();
 b15zdnd11an1n64x5 FILLER_385_1627 ();
 b15zdnd11an1n64x5 FILLER_385_1691 ();
 b15zdnd11an1n64x5 FILLER_385_1755 ();
 b15zdnd11an1n32x5 FILLER_385_1819 ();
 b15zdnd11an1n08x5 FILLER_385_1851 ();
 b15zdnd11an1n04x5 FILLER_385_1859 ();
 b15zdnd00an1n01x5 FILLER_385_1863 ();
 b15zdnd11an1n16x5 FILLER_385_1872 ();
 b15zdnd00an1n02x5 FILLER_385_1888 ();
 b15zdnd11an1n16x5 FILLER_385_1896 ();
 b15zdnd00an1n02x5 FILLER_385_1912 ();
 b15zdnd00an1n01x5 FILLER_385_1914 ();
 b15zdnd11an1n04x5 FILLER_385_1919 ();
 b15zdnd00an1n02x5 FILLER_385_1923 ();
 b15zdnd00an1n01x5 FILLER_385_1925 ();
 b15zdnd11an1n04x5 FILLER_385_1942 ();
 b15zdnd11an1n16x5 FILLER_385_1952 ();
 b15zdnd11an1n16x5 FILLER_385_1977 ();
 b15zdnd11an1n08x5 FILLER_385_1993 ();
 b15zdnd11an1n04x5 FILLER_385_2001 ();
 b15zdnd11an1n64x5 FILLER_385_2025 ();
 b15zdnd11an1n08x5 FILLER_385_2089 ();
 b15zdnd11an1n04x5 FILLER_385_2097 ();
 b15zdnd00an1n02x5 FILLER_385_2101 ();
 b15zdnd11an1n16x5 FILLER_385_2121 ();
 b15zdnd00an1n02x5 FILLER_385_2137 ();
 b15zdnd11an1n64x5 FILLER_385_2170 ();
 b15zdnd11an1n32x5 FILLER_385_2234 ();
 b15zdnd11an1n16x5 FILLER_385_2266 ();
 b15zdnd00an1n02x5 FILLER_385_2282 ();
 b15zdnd11an1n64x5 FILLER_386_8 ();
 b15zdnd11an1n64x5 FILLER_386_72 ();
 b15zdnd11an1n64x5 FILLER_386_136 ();
 b15zdnd11an1n64x5 FILLER_386_200 ();
 b15zdnd11an1n64x5 FILLER_386_264 ();
 b15zdnd11an1n64x5 FILLER_386_328 ();
 b15zdnd11an1n64x5 FILLER_386_392 ();
 b15zdnd11an1n64x5 FILLER_386_456 ();
 b15zdnd11an1n64x5 FILLER_386_520 ();
 b15zdnd11an1n32x5 FILLER_386_584 ();
 b15zdnd11an1n16x5 FILLER_386_616 ();
 b15zdnd11an1n08x5 FILLER_386_652 ();
 b15zdnd00an1n01x5 FILLER_386_660 ();
 b15zdnd11an1n04x5 FILLER_386_670 ();
 b15zdnd11an1n04x5 FILLER_386_686 ();
 b15zdnd11an1n08x5 FILLER_386_694 ();
 b15zdnd00an1n02x5 FILLER_386_702 ();
 b15zdnd00an1n02x5 FILLER_386_716 ();
 b15zdnd11an1n16x5 FILLER_386_726 ();
 b15zdnd11an1n04x5 FILLER_386_742 ();
 b15zdnd00an1n01x5 FILLER_386_746 ();
 b15zdnd11an1n04x5 FILLER_386_763 ();
 b15zdnd11an1n16x5 FILLER_386_786 ();
 b15zdnd11an1n04x5 FILLER_386_802 ();
 b15zdnd00an1n02x5 FILLER_386_806 ();
 b15zdnd11an1n08x5 FILLER_386_818 ();
 b15zdnd00an1n01x5 FILLER_386_826 ();
 b15zdnd11an1n04x5 FILLER_386_836 ();
 b15zdnd11an1n08x5 FILLER_386_846 ();
 b15zdnd11an1n04x5 FILLER_386_854 ();
 b15zdnd11an1n16x5 FILLER_386_871 ();
 b15zdnd11an1n08x5 FILLER_386_887 ();
 b15zdnd00an1n02x5 FILLER_386_895 ();
 b15zdnd00an1n01x5 FILLER_386_897 ();
 b15zdnd11an1n04x5 FILLER_386_903 ();
 b15zdnd11an1n08x5 FILLER_386_913 ();
 b15zdnd00an1n02x5 FILLER_386_921 ();
 b15zdnd11an1n08x5 FILLER_386_933 ();
 b15zdnd11an1n04x5 FILLER_386_941 ();
 b15zdnd11an1n08x5 FILLER_386_958 ();
 b15zdnd00an1n01x5 FILLER_386_966 ();
 b15zdnd11an1n04x5 FILLER_386_975 ();
 b15zdnd00an1n02x5 FILLER_386_979 ();
 b15zdnd11an1n32x5 FILLER_386_985 ();
 b15zdnd00an1n01x5 FILLER_386_1017 ();
 b15zdnd11an1n04x5 FILLER_386_1024 ();
 b15zdnd11an1n64x5 FILLER_386_1060 ();
 b15zdnd11an1n08x5 FILLER_386_1124 ();
 b15zdnd11an1n64x5 FILLER_386_1136 ();
 b15zdnd11an1n64x5 FILLER_386_1200 ();
 b15zdnd11an1n64x5 FILLER_386_1264 ();
 b15zdnd11an1n04x5 FILLER_386_1328 ();
 b15zdnd00an1n02x5 FILLER_386_1332 ();
 b15zdnd11an1n32x5 FILLER_386_1338 ();
 b15zdnd11an1n08x5 FILLER_386_1370 ();
 b15zdnd11an1n04x5 FILLER_386_1378 ();
 b15zdnd00an1n01x5 FILLER_386_1382 ();
 b15zdnd11an1n04x5 FILLER_386_1399 ();
 b15zdnd11an1n64x5 FILLER_386_1407 ();
 b15zdnd11an1n16x5 FILLER_386_1471 ();
 b15zdnd00an1n01x5 FILLER_386_1487 ();
 b15zdnd11an1n04x5 FILLER_386_1495 ();
 b15zdnd00an1n02x5 FILLER_386_1499 ();
 b15zdnd11an1n04x5 FILLER_386_1513 ();
 b15zdnd11an1n64x5 FILLER_386_1522 ();
 b15zdnd11an1n16x5 FILLER_386_1586 ();
 b15zdnd11an1n08x5 FILLER_386_1602 ();
 b15zdnd00an1n01x5 FILLER_386_1610 ();
 b15zdnd11an1n04x5 FILLER_386_1617 ();
 b15zdnd11an1n04x5 FILLER_386_1630 ();
 b15zdnd11an1n64x5 FILLER_386_1639 ();
 b15zdnd11an1n64x5 FILLER_386_1703 ();
 b15zdnd11an1n64x5 FILLER_386_1767 ();
 b15zdnd11an1n32x5 FILLER_386_1831 ();
 b15zdnd11an1n16x5 FILLER_386_1863 ();
 b15zdnd11an1n04x5 FILLER_386_1879 ();
 b15zdnd11an1n16x5 FILLER_386_1895 ();
 b15zdnd00an1n02x5 FILLER_386_1911 ();
 b15zdnd11an1n08x5 FILLER_386_1922 ();
 b15zdnd11an1n04x5 FILLER_386_1930 ();
 b15zdnd00an1n02x5 FILLER_386_1934 ();
 b15zdnd00an1n01x5 FILLER_386_1936 ();
 b15zdnd11an1n08x5 FILLER_386_1945 ();
 b15zdnd11an1n04x5 FILLER_386_1953 ();
 b15zdnd00an1n02x5 FILLER_386_1957 ();
 b15zdnd11an1n04x5 FILLER_386_1965 ();
 b15zdnd00an1n02x5 FILLER_386_1969 ();
 b15zdnd00an1n01x5 FILLER_386_1971 ();
 b15zdnd11an1n16x5 FILLER_386_1977 ();
 b15zdnd11an1n16x5 FILLER_386_2007 ();
 b15zdnd00an1n02x5 FILLER_386_2023 ();
 b15zdnd00an1n01x5 FILLER_386_2025 ();
 b15zdnd11an1n04x5 FILLER_386_2033 ();
 b15zdnd11an1n04x5 FILLER_386_2044 ();
 b15zdnd11an1n08x5 FILLER_386_2058 ();
 b15zdnd00an1n02x5 FILLER_386_2066 ();
 b15zdnd11an1n08x5 FILLER_386_2078 ();
 b15zdnd11an1n08x5 FILLER_386_2104 ();
 b15zdnd00an1n02x5 FILLER_386_2112 ();
 b15zdnd11an1n04x5 FILLER_386_2126 ();
 b15zdnd11an1n16x5 FILLER_386_2134 ();
 b15zdnd11an1n04x5 FILLER_386_2150 ();
 b15zdnd00an1n02x5 FILLER_386_2162 ();
 b15zdnd00an1n01x5 FILLER_386_2164 ();
 b15zdnd11an1n64x5 FILLER_386_2181 ();
 b15zdnd11an1n16x5 FILLER_386_2245 ();
 b15zdnd11an1n08x5 FILLER_386_2261 ();
 b15zdnd11an1n04x5 FILLER_386_2269 ();
 b15zdnd00an1n02x5 FILLER_386_2273 ();
 b15zdnd00an1n01x5 FILLER_386_2275 ();
 b15zdnd11an1n64x5 FILLER_387_0 ();
 b15zdnd11an1n64x5 FILLER_387_64 ();
 b15zdnd11an1n64x5 FILLER_387_128 ();
 b15zdnd11an1n64x5 FILLER_387_192 ();
 b15zdnd11an1n64x5 FILLER_387_256 ();
 b15zdnd11an1n64x5 FILLER_387_320 ();
 b15zdnd11an1n64x5 FILLER_387_384 ();
 b15zdnd11an1n64x5 FILLER_387_448 ();
 b15zdnd11an1n64x5 FILLER_387_512 ();
 b15zdnd11an1n64x5 FILLER_387_576 ();
 b15zdnd00an1n02x5 FILLER_387_640 ();
 b15zdnd00an1n01x5 FILLER_387_642 ();
 b15zdnd11an1n16x5 FILLER_387_657 ();
 b15zdnd11an1n04x5 FILLER_387_673 ();
 b15zdnd11an1n64x5 FILLER_387_681 ();
 b15zdnd11an1n32x5 FILLER_387_745 ();
 b15zdnd00an1n02x5 FILLER_387_777 ();
 b15zdnd00an1n01x5 FILLER_387_779 ();
 b15zdnd11an1n32x5 FILLER_387_784 ();
 b15zdnd11an1n04x5 FILLER_387_816 ();
 b15zdnd00an1n02x5 FILLER_387_820 ();
 b15zdnd11an1n32x5 FILLER_387_827 ();
 b15zdnd11an1n16x5 FILLER_387_859 ();
 b15zdnd11an1n08x5 FILLER_387_875 ();
 b15zdnd11an1n04x5 FILLER_387_883 ();
 b15zdnd00an1n02x5 FILLER_387_887 ();
 b15zdnd11an1n08x5 FILLER_387_893 ();
 b15zdnd00an1n02x5 FILLER_387_901 ();
 b15zdnd11an1n16x5 FILLER_387_910 ();
 b15zdnd11an1n08x5 FILLER_387_926 ();
 b15zdnd00an1n02x5 FILLER_387_934 ();
 b15zdnd00an1n01x5 FILLER_387_936 ();
 b15zdnd11an1n16x5 FILLER_387_941 ();
 b15zdnd11an1n08x5 FILLER_387_957 ();
 b15zdnd00an1n01x5 FILLER_387_965 ();
 b15zdnd11an1n32x5 FILLER_387_974 ();
 b15zdnd11an1n16x5 FILLER_387_1006 ();
 b15zdnd11an1n04x5 FILLER_387_1022 ();
 b15zdnd00an1n02x5 FILLER_387_1026 ();
 b15zdnd11an1n32x5 FILLER_387_1049 ();
 b15zdnd11an1n08x5 FILLER_387_1081 ();
 b15zdnd11an1n04x5 FILLER_387_1089 ();
 b15zdnd00an1n02x5 FILLER_387_1093 ();
 b15zdnd00an1n01x5 FILLER_387_1095 ();
 b15zdnd11an1n64x5 FILLER_387_1100 ();
 b15zdnd11an1n32x5 FILLER_387_1164 ();
 b15zdnd11an1n08x5 FILLER_387_1196 ();
 b15zdnd11an1n04x5 FILLER_387_1204 ();
 b15zdnd00an1n02x5 FILLER_387_1208 ();
 b15zdnd11an1n64x5 FILLER_387_1214 ();
 b15zdnd11an1n64x5 FILLER_387_1278 ();
 b15zdnd11an1n64x5 FILLER_387_1342 ();
 b15zdnd11an1n08x5 FILLER_387_1406 ();
 b15zdnd11an1n64x5 FILLER_387_1418 ();
 b15zdnd11an1n64x5 FILLER_387_1482 ();
 b15zdnd11an1n64x5 FILLER_387_1546 ();
 b15zdnd11an1n64x5 FILLER_387_1610 ();
 b15zdnd11an1n64x5 FILLER_387_1674 ();
 b15zdnd11an1n64x5 FILLER_387_1738 ();
 b15zdnd11an1n64x5 FILLER_387_1802 ();
 b15zdnd11an1n16x5 FILLER_387_1866 ();
 b15zdnd11an1n08x5 FILLER_387_1882 ();
 b15zdnd11an1n04x5 FILLER_387_1890 ();
 b15zdnd00an1n01x5 FILLER_387_1894 ();
 b15zdnd11an1n64x5 FILLER_387_1899 ();
 b15zdnd11an1n16x5 FILLER_387_1963 ();
 b15zdnd11an1n08x5 FILLER_387_1979 ();
 b15zdnd11an1n04x5 FILLER_387_1987 ();
 b15zdnd11an1n08x5 FILLER_387_2003 ();
 b15zdnd11an1n04x5 FILLER_387_2011 ();
 b15zdnd00an1n02x5 FILLER_387_2015 ();
 b15zdnd11an1n64x5 FILLER_387_2029 ();
 b15zdnd11an1n32x5 FILLER_387_2093 ();
 b15zdnd11an1n08x5 FILLER_387_2125 ();
 b15zdnd11an1n04x5 FILLER_387_2133 ();
 b15zdnd00an1n02x5 FILLER_387_2137 ();
 b15zdnd00an1n01x5 FILLER_387_2139 ();
 b15zdnd11an1n64x5 FILLER_387_2156 ();
 b15zdnd11an1n64x5 FILLER_387_2220 ();
 b15zdnd11an1n64x5 FILLER_388_8 ();
 b15zdnd11an1n64x5 FILLER_388_72 ();
 b15zdnd11an1n64x5 FILLER_388_136 ();
 b15zdnd11an1n64x5 FILLER_388_200 ();
 b15zdnd11an1n64x5 FILLER_388_264 ();
 b15zdnd11an1n64x5 FILLER_388_328 ();
 b15zdnd11an1n64x5 FILLER_388_392 ();
 b15zdnd11an1n64x5 FILLER_388_456 ();
 b15zdnd11an1n64x5 FILLER_388_520 ();
 b15zdnd11an1n64x5 FILLER_388_584 ();
 b15zdnd11an1n64x5 FILLER_388_648 ();
 b15zdnd11an1n04x5 FILLER_388_712 ();
 b15zdnd00an1n02x5 FILLER_388_716 ();
 b15zdnd11an1n64x5 FILLER_388_726 ();
 b15zdnd11an1n64x5 FILLER_388_790 ();
 b15zdnd11an1n32x5 FILLER_388_854 ();
 b15zdnd11an1n16x5 FILLER_388_886 ();
 b15zdnd11an1n04x5 FILLER_388_902 ();
 b15zdnd00an1n02x5 FILLER_388_906 ();
 b15zdnd00an1n01x5 FILLER_388_908 ();
 b15zdnd11an1n32x5 FILLER_388_916 ();
 b15zdnd11an1n16x5 FILLER_388_954 ();
 b15zdnd11an1n04x5 FILLER_388_970 ();
 b15zdnd00an1n02x5 FILLER_388_974 ();
 b15zdnd00an1n01x5 FILLER_388_976 ();
 b15zdnd11an1n16x5 FILLER_388_981 ();
 b15zdnd11an1n04x5 FILLER_388_1001 ();
 b15zdnd11an1n16x5 FILLER_388_1010 ();
 b15zdnd11an1n04x5 FILLER_388_1026 ();
 b15zdnd11an1n32x5 FILLER_388_1034 ();
 b15zdnd11an1n32x5 FILLER_388_1070 ();
 b15zdnd11an1n16x5 FILLER_388_1102 ();
 b15zdnd11an1n08x5 FILLER_388_1118 ();
 b15zdnd11an1n04x5 FILLER_388_1131 ();
 b15zdnd11an1n16x5 FILLER_388_1141 ();
 b15zdnd11an1n04x5 FILLER_388_1157 ();
 b15zdnd00an1n01x5 FILLER_388_1161 ();
 b15zdnd11an1n32x5 FILLER_388_1167 ();
 b15zdnd11an1n08x5 FILLER_388_1199 ();
 b15zdnd11an1n64x5 FILLER_388_1212 ();
 b15zdnd11an1n32x5 FILLER_388_1276 ();
 b15zdnd11an1n16x5 FILLER_388_1308 ();
 b15zdnd11an1n08x5 FILLER_388_1324 ();
 b15zdnd11an1n04x5 FILLER_388_1332 ();
 b15zdnd11an1n64x5 FILLER_388_1340 ();
 b15zdnd11an1n08x5 FILLER_388_1404 ();
 b15zdnd11an1n16x5 FILLER_388_1416 ();
 b15zdnd11an1n64x5 FILLER_388_1437 ();
 b15zdnd11an1n64x5 FILLER_388_1501 ();
 b15zdnd11an1n64x5 FILLER_388_1565 ();
 b15zdnd11an1n64x5 FILLER_388_1629 ();
 b15zdnd11an1n64x5 FILLER_388_1693 ();
 b15zdnd11an1n64x5 FILLER_388_1757 ();
 b15zdnd11an1n64x5 FILLER_388_1821 ();
 b15zdnd11an1n64x5 FILLER_388_1885 ();
 b15zdnd11an1n64x5 FILLER_388_1949 ();
 b15zdnd11an1n64x5 FILLER_388_2013 ();
 b15zdnd11an1n64x5 FILLER_388_2077 ();
 b15zdnd11an1n08x5 FILLER_388_2141 ();
 b15zdnd11an1n04x5 FILLER_388_2149 ();
 b15zdnd00an1n01x5 FILLER_388_2153 ();
 b15zdnd11an1n64x5 FILLER_388_2162 ();
 b15zdnd11an1n32x5 FILLER_388_2226 ();
 b15zdnd11an1n16x5 FILLER_388_2258 ();
 b15zdnd00an1n02x5 FILLER_388_2274 ();
 b15zdnd11an1n64x5 FILLER_389_0 ();
 b15zdnd11an1n64x5 FILLER_389_64 ();
 b15zdnd11an1n64x5 FILLER_389_128 ();
 b15zdnd11an1n64x5 FILLER_389_192 ();
 b15zdnd11an1n64x5 FILLER_389_256 ();
 b15zdnd11an1n64x5 FILLER_389_320 ();
 b15zdnd11an1n64x5 FILLER_389_384 ();
 b15zdnd11an1n64x5 FILLER_389_448 ();
 b15zdnd11an1n64x5 FILLER_389_512 ();
 b15zdnd11an1n64x5 FILLER_389_576 ();
 b15zdnd11an1n64x5 FILLER_389_640 ();
 b15zdnd11an1n64x5 FILLER_389_704 ();
 b15zdnd11an1n64x5 FILLER_389_768 ();
 b15zdnd11an1n08x5 FILLER_389_832 ();
 b15zdnd11an1n04x5 FILLER_389_840 ();
 b15zdnd11an1n16x5 FILLER_389_849 ();
 b15zdnd00an1n01x5 FILLER_389_865 ();
 b15zdnd11an1n08x5 FILLER_389_871 ();
 b15zdnd11an1n04x5 FILLER_389_879 ();
 b15zdnd11an1n04x5 FILLER_389_889 ();
 b15zdnd11an1n04x5 FILLER_389_898 ();
 b15zdnd11an1n16x5 FILLER_389_907 ();
 b15zdnd00an1n02x5 FILLER_389_923 ();
 b15zdnd11an1n04x5 FILLER_389_930 ();
 b15zdnd11an1n04x5 FILLER_389_939 ();
 b15zdnd11an1n08x5 FILLER_389_948 ();
 b15zdnd00an1n02x5 FILLER_389_956 ();
 b15zdnd11an1n04x5 FILLER_389_963 ();
 b15zdnd11an1n16x5 FILLER_389_971 ();
 b15zdnd00an1n02x5 FILLER_389_987 ();
 b15zdnd11an1n04x5 FILLER_389_993 ();
 b15zdnd00an1n02x5 FILLER_389_997 ();
 b15zdnd11an1n16x5 FILLER_389_1003 ();
 b15zdnd11an1n04x5 FILLER_389_1019 ();
 b15zdnd00an1n02x5 FILLER_389_1023 ();
 b15zdnd11an1n08x5 FILLER_389_1029 ();
 b15zdnd11an1n04x5 FILLER_389_1037 ();
 b15zdnd11an1n16x5 FILLER_389_1045 ();
 b15zdnd11an1n04x5 FILLER_389_1061 ();
 b15zdnd00an1n02x5 FILLER_389_1065 ();
 b15zdnd00an1n01x5 FILLER_389_1067 ();
 b15zdnd11an1n04x5 FILLER_389_1072 ();
 b15zdnd11an1n04x5 FILLER_389_1082 ();
 b15zdnd11an1n04x5 FILLER_389_1090 ();
 b15zdnd00an1n01x5 FILLER_389_1094 ();
 b15zdnd11an1n08x5 FILLER_389_1099 ();
 b15zdnd11an1n04x5 FILLER_389_1107 ();
 b15zdnd00an1n02x5 FILLER_389_1111 ();
 b15zdnd11an1n04x5 FILLER_389_1117 ();
 b15zdnd11an1n04x5 FILLER_389_1126 ();
 b15zdnd00an1n01x5 FILLER_389_1130 ();
 b15zdnd11an1n04x5 FILLER_389_1136 ();
 b15zdnd11an1n16x5 FILLER_389_1145 ();
 b15zdnd11an1n04x5 FILLER_389_1166 ();
 b15zdnd00an1n02x5 FILLER_389_1170 ();
 b15zdnd00an1n01x5 FILLER_389_1172 ();
 b15zdnd11an1n16x5 FILLER_389_1178 ();
 b15zdnd11an1n08x5 FILLER_389_1194 ();
 b15zdnd00an1n02x5 FILLER_389_1202 ();
 b15zdnd00an1n01x5 FILLER_389_1204 ();
 b15zdnd11an1n08x5 FILLER_389_1210 ();
 b15zdnd11an1n04x5 FILLER_389_1223 ();
 b15zdnd11an1n08x5 FILLER_389_1232 ();
 b15zdnd11an1n04x5 FILLER_389_1240 ();
 b15zdnd00an1n02x5 FILLER_389_1244 ();
 b15zdnd00an1n01x5 FILLER_389_1246 ();
 b15zdnd11an1n16x5 FILLER_389_1252 ();
 b15zdnd11an1n08x5 FILLER_389_1268 ();
 b15zdnd11an1n04x5 FILLER_389_1276 ();
 b15zdnd00an1n02x5 FILLER_389_1280 ();
 b15zdnd11an1n04x5 FILLER_389_1286 ();
 b15zdnd11an1n04x5 FILLER_389_1295 ();
 b15zdnd00an1n02x5 FILLER_389_1299 ();
 b15zdnd00an1n01x5 FILLER_389_1301 ();
 b15zdnd11an1n32x5 FILLER_389_1307 ();
 b15zdnd00an1n02x5 FILLER_389_1339 ();
 b15zdnd11an1n16x5 FILLER_389_1347 ();
 b15zdnd11an1n08x5 FILLER_389_1363 ();
 b15zdnd00an1n02x5 FILLER_389_1371 ();
 b15zdnd00an1n01x5 FILLER_389_1373 ();
 b15zdnd11an1n08x5 FILLER_389_1379 ();
 b15zdnd11an1n04x5 FILLER_389_1387 ();
 b15zdnd11an1n32x5 FILLER_389_1396 ();
 b15zdnd11an1n04x5 FILLER_389_1428 ();
 b15zdnd00an1n01x5 FILLER_389_1432 ();
 b15zdnd11an1n16x5 FILLER_389_1437 ();
 b15zdnd00an1n02x5 FILLER_389_1453 ();
 b15zdnd00an1n01x5 FILLER_389_1455 ();
 b15zdnd11an1n04x5 FILLER_389_1460 ();
 b15zdnd11an1n16x5 FILLER_389_1469 ();
 b15zdnd00an1n02x5 FILLER_389_1485 ();
 b15zdnd11an1n64x5 FILLER_389_1491 ();
 b15zdnd11an1n64x5 FILLER_389_1555 ();
 b15zdnd11an1n64x5 FILLER_389_1619 ();
 b15zdnd11an1n64x5 FILLER_389_1683 ();
 b15zdnd11an1n64x5 FILLER_389_1747 ();
 b15zdnd11an1n64x5 FILLER_389_1811 ();
 b15zdnd11an1n64x5 FILLER_389_1875 ();
 b15zdnd11an1n64x5 FILLER_389_1939 ();
 b15zdnd11an1n64x5 FILLER_389_2003 ();
 b15zdnd11an1n64x5 FILLER_389_2067 ();
 b15zdnd11an1n64x5 FILLER_389_2131 ();
 b15zdnd11an1n64x5 FILLER_389_2195 ();
 b15zdnd11an1n16x5 FILLER_389_2259 ();
 b15zdnd11an1n08x5 FILLER_389_2275 ();
 b15zdnd00an1n01x5 FILLER_389_2283 ();
endmodule
