VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO Noise_injection_block_final_v11
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN Noise_injection_block_final_v11 0 0 ;
  SIZE 18.576 BY 189 ;
  SYMMETRY X Y R90 ;
  PIN Iout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m3 ;
        RECT 1.5995 188.9585 1.6435 189.0025 ;
    END
  END Iout
  PIN Random
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m4 ;
        RECT 0 188.691 0.3215 188.735 ;
    END
  END Random
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 1.868 0.044 1.912 ;
    END
  END S[0]
  PIN S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 129.308 0.044 129.352 ;
    END
  END S[10]
  PIN S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 18.532 129.308 18.576 129.352 ;
    END
  END S[11]
  PIN S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 144.428 0.044 144.472 ;
    END
  END S[12]
  PIN S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 158.468 0.044 158.512 ;
    END
  END S[13]
  PIN S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 176.828 0.044 176.872 ;
    END
  END S[14]
  PIN S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 18.532 176.828 18.576 176.872 ;
    END
  END S[15]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 15.908 0.044 15.952 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 34.268 0.044 34.312 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 18.532 34.268 18.576 34.312 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 49.388 0.044 49.432 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 63.428 0.044 63.472 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 81.788 0.044 81.832 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 18.532 81.788 18.576 81.832 ;
    END
  END S[7]
  PIN S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 96.908 0.044 96.952 ;
    END
  END S[8]
  PIN S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 110.948 0.044 110.992 ;
    END
  END S[9]
  PIN VB[0]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m6 ;
        RECT 0 0.0925 0.448 0.1825 ;
    END
  END VB[0]
  PIN VB[1]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m6 ;
        RECT 0 47.6125 0.25 47.7025 ;
    END
  END VB[1]
  PIN VB[2]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m6 ;
        RECT 0 95.1325 0.25 95.2225 ;
    END
  END VB[2]
  PIN VB[3]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m6 ;
        RECT 0 142.6525 0.358 142.7425 ;
    END
  END VB[3]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER m7 ;
        RECT 2.054 0.251 2.374 188.999 ;
    END
    PORT
      LAYER m7 ;
        RECT 17.3065 -0.0005 17.6265 188.999 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m7 ;
        RECT 1.315 0.251 1.635 188.9995 ;
    END
  END vss
  OBS
    LAYER m1 SPACING 0.04 ;
      RECT 0 0 18.576 189 ;
    LAYER m5 SPACING 0.046 ;
      RECT 0 188.831 18.576 189 ;
      RECT 0.4175 0 18.576 189 ;
      RECT 0 0 18.576 188.595 ;
    LAYER m2 ;
      RECT 7.0425 188.9015 11.5335 188.9915 ;
      RECT 11.4435 188.3735 11.5335 188.9915 ;
      RECT 7.0425 188.353 7.1325 188.9915 ;
      RECT 18.0285 -0.022 18.1885 0.022 ;
      RECT 18.0285 188.978 18.1885 189.022 ;
      RECT 0.3875 188.978 0.5475 189.022 ;
    LAYER m2 SPACING 0.046 ;
      RECT 0 0 18.576 189 ;
    LAYER m3 ;
      RECT 18.0865 -0.05 18.1305 189.05 ;
      RECT 17.721 -0.0005 17.765 188.9975 ;
      RECT 1.5995 36.49 1.6435 188.8585 ;
      RECT 0.811 -0.002 0.855 189 ;
      RECT 0.4455 0 0.4895 189.05 ;
    LAYER m3 SPACING 0.046 ;
      RECT 1.7235 0 18.576 189 ;
      RECT 0 0 1.5195 189 ;
      RECT 0 0 18.576 188.8785 ;
    LAYER m4 SPACING 0.046 ;
      RECT 1.7395 0 18.576 189 ;
      RECT 0.9015 0 18.576 188.8625 ;
      RECT 0 0 18.576 188.111 ;
    LAYER m6 ;
      RECT 17.787 34.268 18.432 34.312 ;
      RECT 17.825 81.788 18.432 81.832 ;
      RECT 17.825 129.308 18.432 129.352 ;
      RECT 17.8185 176.828 18.432 176.872 ;
      RECT 0.548 0.0925 7.1325 0.1825 ;
      RECT 0.35 47.6125 7.0425 47.7025 ;
      RECT 0.35 95.1325 7.0425 95.2225 ;
      RECT 0.458 142.6525 7.0425 142.7425 ;
      RECT 0.144 49.388 0.4255 49.432 ;
      RECT 0.144 176.828 0.425 176.872 ;
      RECT 0.144 63.428 0.3515 63.472 ;
      RECT 0.144 158.468 0.348 158.512 ;
      RECT 0.144 1.868 0.3475 1.912 ;
      RECT 0.144 15.908 0.3455 15.952 ;
      RECT 0.144 110.948 0.3455 110.992 ;
      RECT 0.144 144.428 0.344 144.472 ;
      RECT 0.144 81.788 0.343 81.832 ;
      RECT 0.144 129.308 0.3265 129.352 ;
      RECT 0.144 34.268 0.3225 34.312 ;
      RECT 0.144 96.908 0.3165 96.952 ;
    LAYER m6 SPACING 0.046 ;
      RECT 0 177.078 18.576 189 ;
      RECT 0.25 142.9485 18.326 189 ;
      RECT 0 158.718 18.576 176.622 ;
      RECT 0.564 129.558 18.576 176.622 ;
      RECT 0 144.678 18.576 158.262 ;
      RECT 0 142.9485 18.576 144.222 ;
      RECT 0 129.558 18.576 142.4465 ;
      RECT 0.25 95.4285 18.326 142.4465 ;
      RECT 0 111.198 18.576 129.102 ;
      RECT 0.456 82.038 18.576 129.102 ;
      RECT 0 97.158 18.576 110.742 ;
      RECT 0 95.4285 18.576 96.702 ;
      RECT 0 82.038 18.576 94.9265 ;
      RECT 0.25 47.9085 18.326 94.9265 ;
      RECT 0 63.678 18.576 81.582 ;
      RECT 0.456 34.518 18.576 81.582 ;
      RECT 0 49.638 18.576 63.222 ;
      RECT 0 47.9085 18.576 49.182 ;
      RECT 0 34.518 18.576 47.4065 ;
      RECT 0.25 0.3885 18.326 47.4065 ;
      RECT 0 16.158 18.576 34.062 ;
      RECT 0.654 0 18.576 34.062 ;
      RECT 0 2.118 18.576 15.702 ;
      RECT 0 0.3885 18.576 1.662 ;
    LAYER m7 SPACING 0.18 ;
      RECT 0 177.212 0.895 189 ;
      RECT 0.698 0.5225 0.895 189 ;
      RECT 0.384 143.0825 0.895 189 ;
      RECT 0 158.852 0.895 176.488 ;
      RECT 0 144.812 0.895 158.128 ;
      RECT 0 143.0825 0.895 144.088 ;
      RECT 0 129.692 0.895 142.3125 ;
      RECT 0.59 0.5225 0.895 142.3125 ;
      RECT 0.384 95.5625 0.895 142.3125 ;
      RECT 0 111.332 0.895 128.968 ;
      RECT 0 97.292 0.895 110.608 ;
      RECT 0 95.5625 0.895 96.568 ;
      RECT 0 82.172 0.895 94.7925 ;
      RECT 0.384 48.0425 0.895 94.7925 ;
      RECT 0 63.812 0.895 81.448 ;
      RECT 0 49.772 0.895 63.088 ;
      RECT 0 48.0425 0.895 49.048 ;
      RECT 0 34.652 0.895 47.2725 ;
      RECT 0.384 0.5225 0.895 47.2725 ;
      RECT 0 16.292 0.895 33.928 ;
      RECT 0 2.252 0.895 15.568 ;
      RECT 0 0.5225 0.895 1.528 ;
      RECT 18.0465 0 18.576 33.928 ;
      RECT 18.0465 34.652 18.576 81.448 ;
      RECT 18.0465 82.172 18.576 128.968 ;
      RECT 18.0465 129.692 18.576 176.488 ;
      RECT 18.0465 177.212 18.576 189 ;
      RECT 2.794 0 16.8865 189 ;
  END
END Noise_injection_block_final_v11

END LIBRARY
