module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire net11;
 wire net10;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire net9;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire net8;
 wire _189_;
 wire net7;
 wire net6;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire net5;
 wire _223_;
 wire net4;
 wire _225_;
 wire _226_;
 wire net3;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire net2;
 wire _247_;
 wire net1;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 b15inv000as1n03x5 _298_ (.a(\dpath.a_lt_b$in0[0] ),
    .o1(_035_));
 b15nand02aq1n06x5 _299_ (.a(_035_),
    .b(\dpath.a_lt_b$in1[0] ),
    .o1(_036_));
 b15inv040as1n02x5 _300_ (.a(_036_),
    .o1(_037_));
 b15norp02as1n02x5 _301_ (.a(_035_),
    .b(\dpath.a_lt_b$in1[0] ),
    .o1(_038_));
 b15nor002aq1n02x5 _302_ (.a(_037_),
    .b(_038_),
    .o1(_039_));
 b15inv040ah1n02x5 _303_ (.a(_039_),
    .o1(net37));
 b15nor004as1n02x5 _304_ (.a(\dpath.a_lt_b$in1[15] ),
    .b(\dpath.a_lt_b$in1[14] ),
    .c(\dpath.a_lt_b$in1[13] ),
    .d(\dpath.a_lt_b$in1[12] ),
    .o1(_040_));
 b15nor004an1n02x5 _305_ (.a(\dpath.a_lt_b$in1[11] ),
    .b(\dpath.a_lt_b$in1[10] ),
    .c(\dpath.a_lt_b$in1[9] ),
    .d(\dpath.a_lt_b$in1[8] ),
    .o1(_041_));
 b15nor004ah1n06x5 _306_ (.a(\dpath.a_lt_b$in1[7] ),
    .b(\dpath.a_lt_b$in1[6] ),
    .c(\dpath.a_lt_b$in1[5] ),
    .d(\dpath.a_lt_b$in1[4] ),
    .o1(_042_));
 b15nor004ah1n04x5 _307_ (.a(\dpath.a_lt_b$in1[0] ),
    .b(\dpath.a_lt_b$in1[3] ),
    .c(\dpath.a_lt_b$in1[2] ),
    .d(\dpath.a_lt_b$in1[1] ),
    .o1(_043_));
 b15nand04al1n06x5 _308_ (.a(_040_),
    .b(_041_),
    .c(_042_),
    .d(_043_),
    .o1(_044_));
 b15inv000as1n03x5 _309_ (.a(net34),
    .o1(_045_));
 b15nandp3ar1n02x5 _310_ (.a(_044_),
    .b(_045_),
    .c(\ctrl.state.out[2] ),
    .o1(_046_));
 b15ztpn00an1n08x5 PHY_12 ();
 b15ztpn00an1n08x5 PHY_11 ();
 b15nandp3ar1n02x5 _313_ (.a(_045_),
    .b(net36),
    .c(net33),
    .o1(_049_));
 b15nand02ar1n02x5 _314_ (.a(_046_),
    .b(_049_),
    .o1(_002_));
 b15nor002ah1n32x5 _315_ (.a(\ctrl.state.out[2] ),
    .b(net36),
    .o1(_050_));
 b15and002ar1n02x5 _316_ (.a(_050_),
    .b(\ctrl.state.out[1] ),
    .o(net53));
 b15nand02ar1n02x5 _317_ (.a(net53),
    .b(net35),
    .o1(_051_));
 b15inv020an1n40x5 _318_ (.a(net36),
    .o1(_052_));
 b15ztpn00an1n08x5 PHY_10 ();
 b15oai112aq1n04x5 _320_ (.a(_051_),
    .b(_045_),
    .c(_052_),
    .d(net33),
    .o1(_000_));
 b15nandp3ar1n02x5 _321_ (.a(_051_),
    .b(_045_),
    .c(\ctrl.state.out[1] ),
    .o1(_054_));
 b15inv000ah1n10x5 _322_ (.a(\ctrl.state.out[2] ),
    .o1(_055_));
 b15oai013ar1n02x5 _323_ (.a(_054_),
    .b(_044_),
    .c(net34),
    .d(_055_),
    .o1(_001_));
 b15inv040as1n02x5 _324_ (.a(\dpath.a_lt_b$in1[14] ),
    .o1(_056_));
 b15nand02aq1n02x5 _325_ (.a(_056_),
    .b(\dpath.a_lt_b$in0[14] ),
    .o1(_057_));
 b15inv000al1n02x5 _326_ (.a(_057_),
    .o1(_058_));
 b15nanb02al1n04x5 _327_ (.a(\dpath.a_lt_b$in1[13] ),
    .b(\dpath.a_lt_b$in0[13] ),
    .out0(_059_));
 b15nanb02ar1n02x5 _328_ (.a(\dpath.a_lt_b$in0[13] ),
    .b(\dpath.a_lt_b$in1[13] ),
    .out0(_060_));
 b15nandp2aq1n04x5 _329_ (.a(_059_),
    .b(_060_),
    .o1(_061_));
 b15inv000as1n03x5 _330_ (.a(\dpath.a_lt_b$in1[12] ),
    .o1(_062_));
 b15nand02ar1n02x5 _331_ (.a(_062_),
    .b(\dpath.a_lt_b$in0[12] ),
    .o1(_063_));
 b15oai012al1n02x5 _332_ (.a(_059_),
    .b(_061_),
    .c(_063_),
    .o1(_064_));
 b15inv040ah1n02x5 _333_ (.a(\dpath.a_lt_b$in0[11] ),
    .o1(_065_));
 b15norp02ar1n04x5 _334_ (.a(_065_),
    .b(\dpath.a_lt_b$in1[11] ),
    .o1(_066_));
 b15inv040ah1n02x5 _335_ (.a(\dpath.a_lt_b$in1[11] ),
    .o1(_067_));
 b15norp02ah1n02x5 _336_ (.a(_067_),
    .b(\dpath.a_lt_b$in0[11] ),
    .o1(_068_));
 b15inv000al1n02x5 _337_ (.a(_068_),
    .o1(_069_));
 b15inv040as1n02x5 _338_ (.a(\dpath.a_lt_b$in1[10] ),
    .o1(_070_));
 b15nandp2al1n02x5 _339_ (.a(_070_),
    .b(\dpath.a_lt_b$in0[10] ),
    .o1(_071_));
 b15inv000as1n02x5 _340_ (.a(_071_),
    .o1(_072_));
 b15aoi012ar1n02x5 _341_ (.a(_066_),
    .b(_069_),
    .c(_072_),
    .o1(_073_));
 b15norp02ah1n03x5 _342_ (.a(_066_),
    .b(_068_),
    .o1(_074_));
 b15inv000as1n03x5 _343_ (.a(_074_),
    .o1(_075_));
 b15nanb02an1n03x5 _344_ (.a(\dpath.a_lt_b$in0[10] ),
    .b(\dpath.a_lt_b$in1[10] ),
    .out0(_076_));
 b15nand02aq1n03x5 _345_ (.a(_076_),
    .b(_071_),
    .o1(_077_));
 b15nor002as1n04x5 _346_ (.a(_075_),
    .b(_077_),
    .o1(_078_));
 b15inv040ah1n02x5 _347_ (.a(\dpath.a_lt_b$in1[9] ),
    .o1(_079_));
 b15nandp2al1n02x5 _348_ (.a(_079_),
    .b(\dpath.a_lt_b$in0[9] ),
    .o1(_080_));
 b15norp02al1n04x5 _349_ (.a(_079_),
    .b(\dpath.a_lt_b$in0[9] ),
    .o1(_081_));
 b15cinv00as1n04x5 _350_ (.clk(\dpath.a_lt_b$in1[8] ),
    .clkout(_082_));
 b15nand02ah1n04x5 _351_ (.a(_082_),
    .b(\dpath.a_lt_b$in0[8] ),
    .o1(_083_));
 b15oai012al1n03x5 _352_ (.a(_080_),
    .b(_081_),
    .c(_083_),
    .o1(_084_));
 b15aob012ar1n02x5 _353_ (.a(_073_),
    .b(_078_),
    .c(_084_),
    .out0(_085_));
 b15inv020as1n05x5 _354_ (.a(\dpath.a_lt_b$in0[7] ),
    .o1(_086_));
 b15norp02ar1n02x5 _355_ (.a(_086_),
    .b(\dpath.a_lt_b$in1[7] ),
    .o1(_087_));
 b15inv000ah1n03x5 _356_ (.a(\dpath.a_lt_b$in0[6] ),
    .o1(_088_));
 b15norp02as1n02x5 _357_ (.a(_088_),
    .b(\dpath.a_lt_b$in1[6] ),
    .o1(_089_));
 b15nand02ar1n02x5 _358_ (.a(_086_),
    .b(\dpath.a_lt_b$in1[7] ),
    .o1(_090_));
 b15aoi012al1n02x5 _359_ (.a(_087_),
    .b(_089_),
    .c(_090_),
    .o1(_091_));
 b15inv000as1n03x5 _360_ (.a(\dpath.a_lt_b$in0[5] ),
    .o1(_092_));
 b15nor002al1n06x5 _361_ (.a(_092_),
    .b(\dpath.a_lt_b$in1[5] ),
    .o1(_093_));
 b15inv040ah1n03x5 _362_ (.a(\dpath.a_lt_b$in0[4] ),
    .o1(_094_));
 b15norp02aq1n02x5 _363_ (.a(_094_),
    .b(\dpath.a_lt_b$in1[4] ),
    .o1(_095_));
 b15nandp2al1n05x5 _364_ (.a(_092_),
    .b(\dpath.a_lt_b$in1[5] ),
    .o1(_096_));
 b15aoi012ar1n02x5 _365_ (.a(_093_),
    .b(_095_),
    .c(_096_),
    .o1(_097_));
 b15xor002ah1n04x5 _366_ (.a(_086_),
    .b(\dpath.a_lt_b$in1[7] ),
    .out0(_098_));
 b15xor002al1n06x5 _367_ (.a(_088_),
    .b(\dpath.a_lt_b$in1[6] ),
    .out0(_099_));
 b15nand02ar1n12x5 _368_ (.a(_098_),
    .b(_099_),
    .o1(_100_));
 b15oai012ah1n04x5 _369_ (.a(_091_),
    .b(_097_),
    .c(_100_),
    .o1(_101_));
 b15inv040ah1n03x5 _370_ (.a(\dpath.a_lt_b$in0[3] ),
    .o1(_102_));
 b15norp02an1n02x5 _371_ (.a(_102_),
    .b(\dpath.a_lt_b$in1[3] ),
    .o1(_103_));
 b15inv040as1n02x5 _372_ (.a(\dpath.a_lt_b$in0[2] ),
    .o1(_104_));
 b15nor002as1n02x5 _373_ (.a(_104_),
    .b(\dpath.a_lt_b$in1[2] ),
    .o1(_105_));
 b15nandp2ar1n02x5 _374_ (.a(_102_),
    .b(\dpath.a_lt_b$in1[3] ),
    .o1(_106_));
 b15aoi012al1n02x5 _375_ (.a(_103_),
    .b(_105_),
    .c(_106_),
    .o1(_107_));
 b15inv000as1n03x5 _376_ (.a(\dpath.a_lt_b$in0[1] ),
    .o1(_108_));
 b15qgbno2an1n05x5 _377_ (.o1(_109_),
    .a(_108_),
    .b(\dpath.a_lt_b$in1[1] ));
 b15nand02aq1n04x5 _378_ (.a(_108_),
    .b(\dpath.a_lt_b$in1[1] ),
    .o1(_110_));
 b15aoi012as1n06x5 _379_ (.a(_109_),
    .b(_036_),
    .c(_110_),
    .o1(_111_));
 b15xor002ar1n04x5 _380_ (.a(_102_),
    .b(\dpath.a_lt_b$in1[3] ),
    .out0(_112_));
 b15xor002ar1n03x5 _381_ (.a(_104_),
    .b(\dpath.a_lt_b$in1[2] ),
    .out0(_113_));
 b15nand02al1n04x5 _382_ (.a(_112_),
    .b(_113_),
    .o1(_114_));
 b15oai012as1n08x5 _383_ (.a(_107_),
    .b(_111_),
    .c(_114_),
    .o1(_115_));
 b15nanb02aq1n04x5 _384_ (.a(_093_),
    .b(_096_),
    .out0(_116_));
 b15inv000as1n02x5 _385_ (.a(_095_),
    .o1(_117_));
 b15nand02ah1n04x5 _386_ (.a(_094_),
    .b(\dpath.a_lt_b$in1[4] ),
    .o1(_118_));
 b15nand02al1n06x5 _387_ (.a(_117_),
    .b(_118_),
    .o1(_119_));
 b15norp03an1n04x5 _388_ (.a(_100_),
    .b(_116_),
    .c(_119_),
    .o1(_120_));
 b15aoi012an1n08x5 _389_ (.a(_101_),
    .b(_115_),
    .c(_120_),
    .o1(_121_));
 b15norp02ar1n04x5 _390_ (.a(_082_),
    .b(\dpath.a_lt_b$in0[8] ),
    .o1(_122_));
 b15nanb02ah1n04x5 _391_ (.a(_122_),
    .b(_083_),
    .out0(_123_));
 b15inv000an1n02x5 _392_ (.a(_080_),
    .o1(_124_));
 b15nor002al1n04x5 _393_ (.a(_124_),
    .b(_081_),
    .o1(_125_));
 b15nanb02al1n03x5 _394_ (.a(_123_),
    .b(_125_),
    .out0(_126_));
 b15nanb02an1n06x5 _395_ (.a(_126_),
    .b(_078_),
    .out0(_127_));
 b15oabi12aq1n06x5 _396_ (.a(_085_),
    .b(_121_),
    .c(_127_),
    .out0(_128_));
 b15norp02aq1n04x5 _397_ (.a(_062_),
    .b(\dpath.a_lt_b$in0[12] ),
    .o1(_129_));
 b15inv040an1n02x5 _398_ (.a(_063_),
    .o1(_130_));
 b15nor003aq1n04x5 _399_ (.a(_061_),
    .b(_129_),
    .c(_130_),
    .o1(_131_));
 b15aoi012al1n04x5 _400_ (.a(_064_),
    .b(_128_),
    .c(_131_),
    .o1(_132_));
 b15nanb02al1n03x5 _401_ (.a(\dpath.a_lt_b$in0[14] ),
    .b(\dpath.a_lt_b$in1[14] ),
    .out0(_133_));
 b15nand02an1n04x5 _402_ (.a(_133_),
    .b(_057_),
    .o1(_134_));
 b15oabi12an1n02x5 _403_ (.a(_058_),
    .b(_132_),
    .c(_134_),
    .out0(_135_));
 b15nanb02ar1n03x5 _404_ (.a(\dpath.a_lt_b$in0[15] ),
    .b(\dpath.a_lt_b$in1[15] ),
    .out0(_136_));
 b15inv000as1n02x5 _405_ (.a(\dpath.a_lt_b$in1[15] ),
    .o1(_137_));
 b15nand02ar1n02x5 _406_ (.a(_137_),
    .b(\dpath.a_lt_b$in0[15] ),
    .o1(_138_));
 b15nand02an1n04x5 _407_ (.a(_136_),
    .b(_138_),
    .o1(_139_));
 b15xor002ah1n02x5 _408_ (.a(_135_),
    .b(_139_),
    .out0(_140_));
 b15inv040ah1n02x5 _409_ (.a(_140_),
    .o1(net43));
 b15nonb02al1n03x5 _410_ (.a(_110_),
    .b(_109_),
    .out0(_141_));
 b15xor002an1n02x5 _411_ (.a(_141_),
    .b(_036_),
    .out0(net44));
 b15inv040ah1n02x5 _412_ (.a(_113_),
    .o1(_142_));
 b15xor002al1n02x5 _413_ (.a(_111_),
    .b(_142_),
    .out0(net45));
 b15oabi12an1n02x5 _414_ (.a(_105_),
    .b(_111_),
    .c(_142_),
    .out0(_143_));
 b15xor002an1n02x5 _415_ (.a(_143_),
    .b(_112_),
    .out0(net46));
 b15xnr002ar1n04x5 _416_ (.a(_115_),
    .b(_119_),
    .out0(net47));
 b15aob012ah1n04x5 _417_ (.a(_117_),
    .b(_115_),
    .c(_118_),
    .out0(_144_));
 b15xnr002as1n02x5 _418_ (.a(_144_),
    .b(_116_),
    .out0(net48));
 b15aoi012ar1n04x5 _419_ (.a(_093_),
    .b(_144_),
    .c(_096_),
    .o1(_145_));
 b15inv000al1n02x5 _420_ (.a(_099_),
    .o1(_146_));
 b15xor002an1n02x5 _421_ (.a(_145_),
    .b(_146_),
    .out0(net49));
 b15nonb02an1n02x5 _422_ (.a(\dpath.a_lt_b$in1[6] ),
    .b(\dpath.a_lt_b$in0[6] ),
    .out0(_147_));
 b15oabi12an1n02x5 _423_ (.a(_089_),
    .b(_145_),
    .c(_147_),
    .out0(_148_));
 b15xor002ah1n02x5 _424_ (.a(_148_),
    .b(_098_),
    .out0(net50));
 b15xor002al1n06x5 _425_ (.a(_121_),
    .b(_123_),
    .out0(net51));
 b15oai012aq1n03x5 _426_ (.a(_083_),
    .b(_121_),
    .c(_122_),
    .o1(_149_));
 b15xor002ah1n04x5 _427_ (.a(_149_),
    .b(_125_),
    .out0(net52));
 b15oabi12ah1n02x5 _428_ (.a(_084_),
    .b(_121_),
    .c(_126_),
    .out0(_150_));
 b15inv000al1n02x5 _429_ (.a(_077_),
    .o1(_151_));
 b15and002as1n02x5 _430_ (.a(_150_),
    .b(_151_),
    .o(_152_));
 b15norp02ar1n02x5 _431_ (.a(_150_),
    .b(_151_),
    .o1(_153_));
 b15nor002aq1n04x5 _432_ (.a(_152_),
    .b(_153_),
    .o1(net38));
 b15orn003ar1n02x5 _433_ (.a(_152_),
    .b(_072_),
    .c(_074_),
    .o(_154_));
 b15oai012al1n02x5 _434_ (.a(_074_),
    .b(_152_),
    .c(_072_),
    .o1(_155_));
 b15and002an1n02x5 _435_ (.a(_154_),
    .b(_155_),
    .o(net39));
 b15norp02ar1n02x5 _436_ (.a(_130_),
    .b(_129_),
    .o1(_156_));
 b15and002ar1n02x5 _437_ (.a(_128_),
    .b(_156_),
    .o(_157_));
 b15norp02ar1n02x5 _438_ (.a(_128_),
    .b(_156_),
    .o1(_158_));
 b15norp02an1n02x5 _439_ (.a(_157_),
    .b(_158_),
    .o1(net40));
 b15norp02ah1n02x5 _440_ (.a(_157_),
    .b(_130_),
    .o1(_159_));
 b15xor002al1n02x5 _441_ (.a(_159_),
    .b(_061_),
    .out0(net41));
 b15xor002an1n02x5 _442_ (.a(_132_),
    .b(_134_),
    .out0(net42));
 b15nor002ah1n03x5 _443_ (.a(_139_),
    .b(_134_),
    .o1(_160_));
 b15nandp2al1n05x5 _444_ (.a(_131_),
    .b(_160_),
    .o1(_161_));
 b15inv040ah1n02x5 _445_ (.a(_114_),
    .o1(_162_));
 b15nandp3ar1n03x5 _446_ (.a(_162_),
    .b(_039_),
    .c(_141_),
    .o1(_163_));
 b15norp02ar1n02x5 _447_ (.a(_116_),
    .b(_119_),
    .o1(_164_));
 b15nanb02an1n04x5 _448_ (.a(_100_),
    .b(_164_),
    .out0(_165_));
 b15nor004as1n06x5 _449_ (.a(_127_),
    .b(_161_),
    .c(_163_),
    .d(_165_),
    .o1(_166_));
 b15nor002ar1n02x5 _450_ (.a(_127_),
    .b(_161_),
    .o1(_167_));
 b15aoi012ar1n02x5 _451_ (.a(_109_),
    .b(_038_),
    .c(_110_),
    .o1(_168_));
 b15nand02ar1n02x5 _452_ (.a(_162_),
    .b(_168_),
    .o1(_169_));
 b15nand02ar1n02x5 _453_ (.a(_104_),
    .b(\dpath.a_lt_b$in1[2] ),
    .o1(_170_));
 b15oa0012ar1n02x5 _454_ (.a(_106_),
    .b(_103_),
    .c(_170_),
    .o(_171_));
 b15aoi012ar1n02x5 _455_ (.a(_165_),
    .b(_169_),
    .c(_171_),
    .o1(_172_));
 b15rm6013eh1n04x5 _456_ (.a(\dpath.a_lt_b$in1[7] ),
    .b(_086_),
    .c(_147_),
    .carryb(_173_));
 b15and002ar1n02x5 _457_ (.a(_118_),
    .b(_096_),
    .o(_174_));
 b15oai013al1n06x5 _458_ (.a(_173_),
    .b(_100_),
    .c(_174_),
    .d(_093_),
    .o1(_175_));
 b15oai012ar1n06x5 _459_ (.a(_167_),
    .b(_172_),
    .c(_175_),
    .o1(_176_));
 b15oai012as1n02x5 _460_ (.a(_136_),
    .b(_139_),
    .c(_133_),
    .o1(_177_));
 b15nanb02ar1n02x5 _461_ (.a(_129_),
    .b(_060_),
    .out0(_178_));
 b15qgbao4an1n05x5 _462_ (.o1(_179_),
    .a(_177_),
    .b(_059_),
    .c(_160_),
    .d(_178_));
 b15inv040ah1n02x5 _463_ (.a(_161_),
    .o1(_180_));
 b15aoi012ar1n02x5 _464_ (.a(_066_),
    .b(_069_),
    .c(_076_),
    .o1(_181_));
 b15oab012an1n02x5 _465_ (.a(_124_),
    .b(_122_),
    .c(_081_),
    .out0(_182_));
 b15aoai13ar1n04x5 _466_ (.a(_180_),
    .b(_181_),
    .c(_078_),
    .d(_182_),
    .o1(_183_));
 b15nand03an1n12x5 _467_ (.a(_176_),
    .b(_179_),
    .c(_183_),
    .o1(_184_));
 b15nanb02an1n24x5 _468_ (.a(_166_),
    .b(_184_),
    .out0(_185_));
 b15norp02as1n48x5 _469_ (.a(_185_),
    .b(_055_),
    .o1(_186_));
 b15norp02an1n32x5 _470_ (.a(_186_),
    .b(net36),
    .o1(_187_));
 b15ztpn00an1n08x5 PHY_9 ();
 b15nand02ar1n02x5 _472_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[0] ),
    .o1(_189_));
 b15ztpn00an1n08x5 PHY_8 ();
 b15ztpn00an1n08x5 PHY_7 ();
 b15nandp3ar1n02x5 _475_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[0] ),
    .c(_052_),
    .o1(_192_));
 b15nand02ar1n02x5 _476_ (.a(net36),
    .b(net1),
    .o1(_193_));
 b15nand03an1n04x5 _477_ (.a(_189_),
    .b(_192_),
    .c(_193_),
    .o1(_003_));
 b15nand02ar1n02x5 _478_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[1] ),
    .o1(_194_));
 b15nandp3ar1n02x5 _479_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[1] ),
    .c(_052_),
    .o1(_195_));
 b15nand02al1n02x5 _480_ (.a(net36),
    .b(net12),
    .o1(_196_));
 b15nandp3ar1n03x5 _481_ (.a(_194_),
    .b(_195_),
    .c(_196_),
    .o1(_004_));
 b15nand02ar1n02x5 _482_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[2] ),
    .o1(_197_));
 b15nandp3ar1n02x5 _483_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[2] ),
    .c(_052_),
    .o1(_198_));
 b15nand02ar1n02x5 _484_ (.a(net36),
    .b(net23),
    .o1(_199_));
 b15nandp3ah1n04x5 _485_ (.a(_197_),
    .b(_198_),
    .c(_199_),
    .o1(_005_));
 b15nand02ar1n02x5 _486_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[3] ),
    .o1(_200_));
 b15nandp3ar1n02x5 _487_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[3] ),
    .c(_052_),
    .o1(_201_));
 b15nandp2an1n02x5 _488_ (.a(net36),
    .b(net26),
    .o1(_202_));
 b15nand03an1n04x5 _489_ (.a(_200_),
    .b(_201_),
    .c(_202_),
    .o1(_006_));
 b15nand02ar1n02x5 _490_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[4] ),
    .o1(_203_));
 b15nandp2al1n02x5 _491_ (.a(_094_),
    .b(_052_),
    .o1(_204_));
 b15oai012al1n03x5 _492_ (.a(_204_),
    .b(_052_),
    .c(net27),
    .o1(_205_));
 b15oai012aq1n02x5 _493_ (.a(_203_),
    .b(_187_),
    .c(_205_),
    .o1(_007_));
 b15nand02ar1n02x5 _494_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[5] ),
    .o1(_206_));
 b15nandp3ar1n02x5 _495_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[5] ),
    .c(_052_),
    .o1(_207_));
 b15nand02ar1n02x5 _496_ (.a(net36),
    .b(net28),
    .o1(_208_));
 b15nand03an1n03x5 _497_ (.a(_206_),
    .b(_207_),
    .c(_208_),
    .o1(_008_));
 b15nand02ar1n02x5 _498_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[6] ),
    .o1(_209_));
 b15nandp3ar1n02x5 _499_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[6] ),
    .c(_052_),
    .o1(_210_));
 b15nand02ar1n02x5 _500_ (.a(net36),
    .b(net29),
    .o1(_211_));
 b15nand03an1n03x5 _501_ (.a(_209_),
    .b(_210_),
    .c(_211_),
    .o1(_009_));
 b15nand02ar1n02x5 _502_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[7] ),
    .o1(_212_));
 b15nandp3ar1n02x5 _503_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[7] ),
    .c(_052_),
    .o1(_213_));
 b15nand02ar1n02x5 _504_ (.a(net36),
    .b(net30),
    .o1(_214_));
 b15nand03ar1n04x5 _505_ (.a(_212_),
    .b(_213_),
    .c(_214_),
    .o1(_010_));
 b15nand02ar1n02x5 _506_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[8] ),
    .o1(_215_));
 b15nandp3ar1n02x5 _507_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[8] ),
    .c(_052_),
    .o1(_216_));
 b15nand02ar1n02x5 _508_ (.a(net36),
    .b(net31),
    .o1(_217_));
 b15nand03ar1n03x5 _509_ (.a(_215_),
    .b(_216_),
    .c(_217_),
    .o1(_011_));
 b15nand02ar1n02x5 _510_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[9] ),
    .o1(_218_));
 b15nandp3ar1n02x5 _511_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[9] ),
    .c(_052_),
    .o1(_219_));
 b15nand02ar1n02x5 _512_ (.a(net36),
    .b(net32),
    .o1(_220_));
 b15nandp3an1n02x5 _513_ (.a(_218_),
    .b(_219_),
    .c(_220_),
    .o1(_012_));
 b15nand02ar1n02x5 _514_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[10] ),
    .o1(_221_));
 b15ztpn00an1n08x5 PHY_6 ();
 b15nandp3ar1n02x5 _516_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[10] ),
    .c(_052_),
    .o1(_223_));
 b15ztpn00an1n08x5 PHY_5 ();
 b15nand02ar1n02x5 _518_ (.a(net36),
    .b(net2),
    .o1(_225_));
 b15nandp3ar1n02x5 _519_ (.a(_221_),
    .b(_223_),
    .c(_225_),
    .o1(_013_));
 b15nand02ar1n02x5 _520_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[11] ),
    .o1(_226_));
 b15ztpn00an1n08x5 PHY_4 ();
 b15nandp3ar1n02x5 _522_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[11] ),
    .c(_052_),
    .o1(_228_));
 b15nand02ar1n02x5 _523_ (.a(net36),
    .b(net3),
    .o1(_229_));
 b15nandp3ar1n02x5 _524_ (.a(_226_),
    .b(_228_),
    .c(_229_),
    .o1(_014_));
 b15nand02ar1n02x5 _525_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[12] ),
    .o1(_230_));
 b15nandp3ar1n02x5 _526_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[12] ),
    .c(_052_),
    .o1(_231_));
 b15nand02ar1n02x5 _527_ (.a(net36),
    .b(net4),
    .o1(_232_));
 b15nandp3an1n03x5 _528_ (.a(_230_),
    .b(_231_),
    .c(_232_),
    .o1(_015_));
 b15nand02ar1n02x5 _529_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[13] ),
    .o1(_233_));
 b15nandp3ar1n02x5 _530_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[13] ),
    .c(_052_),
    .o1(_234_));
 b15nand02ar1n02x5 _531_ (.a(net36),
    .b(net5),
    .o1(_235_));
 b15nand03ah1n04x5 _532_ (.a(_233_),
    .b(_234_),
    .c(_235_),
    .o1(_016_));
 b15nand02ar1n02x5 _533_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[14] ),
    .o1(_236_));
 b15nandp3ar1n02x5 _534_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[14] ),
    .c(_052_),
    .o1(_237_));
 b15nand02ar1n02x5 _535_ (.a(net36),
    .b(net6),
    .o1(_238_));
 b15nand03aq1n06x5 _536_ (.a(_236_),
    .b(_237_),
    .c(_238_),
    .o1(_017_));
 b15nand02ar1n02x5 _537_ (.a(_187_),
    .b(\dpath.a_lt_b$in1[15] ),
    .o1(_239_));
 b15nandp3ar1n02x5 _538_ (.a(_186_),
    .b(\dpath.a_lt_b$in0[15] ),
    .c(_052_),
    .o1(_240_));
 b15nand02ar1n02x5 _539_ (.a(net36),
    .b(net7),
    .o1(_241_));
 b15nandp3al1n02x5 _540_ (.a(_239_),
    .b(_240_),
    .c(_241_),
    .o1(_018_));
 b15nand03ar1n02x5 _541_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[0] ),
    .c(_052_),
    .o1(_242_));
 b15norp02an1n04x5 _542_ (.a(_055_),
    .b(net36),
    .o1(_243_));
 b15nand02an1n08x5 _543_ (.a(_185_),
    .b(_243_),
    .o1(_244_));
 b15inv000ah1n20x5 _544_ (.a(_244_),
    .o1(_245_));
 b15ztpn00an1n08x5 PHY_3 ();
 b15nand02ar1n02x5 _546_ (.a(_245_),
    .b(net37),
    .o1(_247_));
 b15ztpn00an1n08x5 PHY_2 ();
 b15aoi022ar1n02x5 _548_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[0] ),
    .c(net36),
    .d(net8),
    .o1(_249_));
 b15nand03ah1n06x5 _549_ (.a(_242_),
    .b(_247_),
    .c(_249_),
    .o1(_019_));
 b15nandp3an1n02x5 _550_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[1] ),
    .c(_052_),
    .o1(_250_));
 b15nandp2ar1n02x5 _551_ (.a(_245_),
    .b(net44),
    .o1(_251_));
 b15aoi022al1n02x5 _552_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[1] ),
    .c(net36),
    .d(net9),
    .o1(_252_));
 b15nand03ar1n08x5 _553_ (.a(_250_),
    .b(_251_),
    .c(_252_),
    .o1(_020_));
 b15ztpn00an1n08x5 PHY_1 ();
 b15nandp3ar1n02x5 _555_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[2] ),
    .c(_052_),
    .o1(_254_));
 b15nand02ar1n02x5 _556_ (.a(_245_),
    .b(net45),
    .o1(_255_));
 b15aoi022ar1n02x5 _557_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[2] ),
    .c(net36),
    .d(net10),
    .o1(_256_));
 b15nandp3ah1n04x5 _558_ (.a(_254_),
    .b(_255_),
    .c(_256_),
    .o1(_021_));
 b15nandp3ar1n02x5 _559_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[3] ),
    .c(_052_),
    .o1(_257_));
 b15nand02ar1n02x5 _560_ (.a(_245_),
    .b(net46),
    .o1(_258_));
 b15aoi022ar1n02x5 _561_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[3] ),
    .c(net36),
    .d(net11),
    .o1(_259_));
 b15nandp3aq1n03x5 _562_ (.a(_257_),
    .b(_258_),
    .c(_259_),
    .o1(_022_));
 b15nandp3ar1n02x5 _563_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[4] ),
    .c(_052_),
    .o1(_260_));
 b15nand02ar1n02x5 _564_ (.a(_245_),
    .b(net47),
    .o1(_261_));
 b15ztpn00an1n08x5 PHY_0 ();
 b15aoai13ar1n02x5 _566_ (.a(_204_),
    .b(_050_),
    .c(net36),
    .d(net13),
    .o1(_263_));
 b15nand03as1n03x5 _567_ (.a(_260_),
    .b(_261_),
    .c(_263_),
    .o1(_023_));
 b15nandp3ar1n02x5 _568_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[5] ),
    .c(_052_),
    .o1(_264_));
 b15nand02ar1n02x5 _569_ (.a(_245_),
    .b(net48),
    .o1(_265_));
 b15aoi022ar1n02x5 _570_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[5] ),
    .c(net36),
    .d(net14),
    .o1(_266_));
 b15nand03ar1n04x5 _571_ (.a(_264_),
    .b(_265_),
    .c(_266_),
    .o1(_024_));
 b15nandp3ar1n02x5 _572_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[6] ),
    .c(_052_),
    .o1(_267_));
 b15nand02ar1n02x5 _573_ (.a(_245_),
    .b(net49),
    .o1(_268_));
 b15aoi022ar1n02x5 _574_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[6] ),
    .c(net36),
    .d(net15),
    .o1(_269_));
 b15nandp3aq1n03x5 _575_ (.a(_267_),
    .b(_268_),
    .c(_269_),
    .o1(_025_));
 b15nand02ar1n02x5 _576_ (.a(net50),
    .b(_245_),
    .o1(_270_));
 b15nandp3ar1n02x5 _577_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[7] ),
    .c(_052_),
    .o1(_271_));
 b15aoi022ar1n02x5 _578_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[7] ),
    .c(net36),
    .d(net16),
    .o1(_272_));
 b15nand03al1n02x5 _579_ (.a(_270_),
    .b(_271_),
    .c(_272_),
    .o1(_026_));
 b15nandp3ar1n02x5 _580_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[8] ),
    .c(_052_),
    .o1(_273_));
 b15nand02ar1n02x5 _581_ (.a(_245_),
    .b(net51),
    .o1(_274_));
 b15aoi022ar1n02x5 _582_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[8] ),
    .c(net36),
    .d(net17),
    .o1(_275_));
 b15nand03ar1n03x5 _583_ (.a(_273_),
    .b(_274_),
    .c(_275_),
    .o1(_027_));
 b15nandp3ar1n02x5 _584_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[9] ),
    .c(_052_),
    .o1(_276_));
 b15nand02ar1n02x5 _585_ (.a(_245_),
    .b(net52),
    .o1(_277_));
 b15aoi022ar1n02x5 _586_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[9] ),
    .c(net36),
    .d(net18),
    .o1(_278_));
 b15nandp3ar1n02x5 _587_ (.a(_276_),
    .b(_277_),
    .c(_278_),
    .o1(_028_));
 b15nandp3ar1n02x5 _588_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[10] ),
    .c(_052_),
    .o1(_279_));
 b15nand02ar1n02x5 _589_ (.a(_245_),
    .b(net38),
    .o1(_280_));
 b15aoi022ar1n02x5 _590_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[10] ),
    .c(net36),
    .d(net19),
    .o1(_281_));
 b15nandp3ar1n02x5 _591_ (.a(_279_),
    .b(_280_),
    .c(_281_),
    .o1(_029_));
 b15nandp3ar1n02x5 _592_ (.a(_154_),
    .b(_245_),
    .c(_155_),
    .o1(_282_));
 b15aoi022ar1n02x5 _593_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[11] ),
    .c(net36),
    .d(net20),
    .o1(_283_));
 b15nano22ar1n02x5 _594_ (.a(\dpath.a_lt_b$in1[11] ),
    .b(_243_),
    .c(_185_),
    .out0(_284_));
 b15nonb02ar1n02x5 _595_ (.a(_283_),
    .b(_284_),
    .out0(_285_));
 b15nandp2al1n02x5 _596_ (.a(_282_),
    .b(_285_),
    .o1(_030_));
 b15nand03ar1n03x5 _597_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[12] ),
    .c(_052_),
    .o1(_286_));
 b15nand02ar1n02x5 _598_ (.a(_245_),
    .b(net40),
    .o1(_287_));
 b15aoi022ar1n02x5 _599_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[12] ),
    .c(net36),
    .d(net21),
    .o1(_288_));
 b15nand03ah1n06x5 _600_ (.a(_286_),
    .b(_287_),
    .c(_288_),
    .o1(_031_));
 b15nand02ar1n02x5 _601_ (.a(net41),
    .b(_245_),
    .o1(_289_));
 b15nandp3ar1n02x5 _602_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[13] ),
    .c(_052_),
    .o1(_290_));
 b15aoi022ar1n02x5 _603_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[13] ),
    .c(net36),
    .d(net22),
    .o1(_291_));
 b15nandp3ah1n03x5 _604_ (.a(_289_),
    .b(_290_),
    .c(_291_),
    .o1(_032_));
 b15nandp3ar1n02x5 _605_ (.a(_186_),
    .b(\dpath.a_lt_b$in1[14] ),
    .c(_052_),
    .o1(_292_));
 b15nand02ar1n02x5 _606_ (.a(_245_),
    .b(net42),
    .o1(_293_));
 b15aoi022al1n02x5 _607_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[14] ),
    .c(net36),
    .d(net24),
    .o1(_294_));
 b15nand03ar1n06x5 _608_ (.a(_292_),
    .b(_293_),
    .c(_294_),
    .o1(_033_));
 b15nona23ar1n02x5 _609_ (.a(_137_),
    .b(_166_),
    .c(_184_),
    .d(_243_),
    .out0(_295_));
 b15aoi022ar1n02x5 _610_ (.a(_050_),
    .b(\dpath.a_lt_b$in0[15] ),
    .c(net36),
    .d(net25),
    .o1(_296_));
 b15nand02ar1n02x5 _611_ (.a(_295_),
    .b(_296_),
    .o1(_297_));
 b15oabi12as1n02x5 _612_ (.a(_297_),
    .b(_140_),
    .c(_244_),
    .out0(_034_));
 b15fpn000hn1n04x5 _613_ (.clk(clknet_2_2__leaf_clk),
    .d(_000_),
    .o(net36));
 b15fpn000hn1n04x5 _614_ (.clk(clknet_2_3__leaf_clk),
    .d(_001_),
    .o(\ctrl.state.out[1] ));
 b15fpn000hn1n04x5 _615_ (.clk(clknet_2_3__leaf_clk),
    .d(_002_),
    .o(\ctrl.state.out[2] ));
 b15fpn000hn1n04x5 _616_ (.clk(clknet_2_3__leaf_clk),
    .d(_003_),
    .o(\dpath.a_lt_b$in1[0] ));
 b15fpn000hn1n04x5 _617_ (.clk(clknet_2_1__leaf_clk),
    .d(_004_),
    .o(\dpath.a_lt_b$in1[1] ));
 b15fpn000hn1n04x5 _618_ (.clk(clknet_2_1__leaf_clk),
    .d(_005_),
    .o(\dpath.a_lt_b$in1[2] ));
 b15fpn000hn1n04x5 _619_ (.clk(clknet_2_1__leaf_clk),
    .d(_006_),
    .o(\dpath.a_lt_b$in1[3] ));
 b15fpn000hn1n04x5 _620_ (.clk(clknet_2_0__leaf_clk),
    .d(_007_),
    .o(\dpath.a_lt_b$in1[4] ));
 b15fpn000hn1n04x5 _621_ (.clk(clknet_2_0__leaf_clk),
    .d(_008_),
    .o(\dpath.a_lt_b$in1[5] ));
 b15fpn000hn1n04x5 _622_ (.clk(clknet_2_0__leaf_clk),
    .d(_009_),
    .o(\dpath.a_lt_b$in1[6] ));
 b15fpn000hn1n04x5 _623_ (.clk(clknet_2_0__leaf_clk),
    .d(_010_),
    .o(\dpath.a_lt_b$in1[7] ));
 b15fpn000hn1n04x5 _624_ (.clk(clknet_2_0__leaf_clk),
    .d(_011_),
    .o(\dpath.a_lt_b$in1[8] ));
 b15fpn000hn1n04x5 _625_ (.clk(clknet_2_2__leaf_clk),
    .d(_012_),
    .o(\dpath.a_lt_b$in1[9] ));
 b15fpn000hn1n04x5 _626_ (.clk(clknet_2_2__leaf_clk),
    .d(_013_),
    .o(\dpath.a_lt_b$in1[10] ));
 b15fpn000hn1n04x5 _627_ (.clk(clknet_2_2__leaf_clk),
    .d(_014_),
    .o(\dpath.a_lt_b$in1[11] ));
 b15fpn000hn1n04x5 _628_ (.clk(clknet_2_3__leaf_clk),
    .d(_015_),
    .o(\dpath.a_lt_b$in1[12] ));
 b15fpn000hn1n04x5 _629_ (.clk(clknet_2_3__leaf_clk),
    .d(_016_),
    .o(\dpath.a_lt_b$in1[13] ));
 b15fpn000hn1n04x5 _630_ (.clk(clknet_2_2__leaf_clk),
    .d(_017_),
    .o(\dpath.a_lt_b$in1[14] ));
 b15fpn000hn1n04x5 _631_ (.clk(clknet_2_3__leaf_clk),
    .d(_018_),
    .o(\dpath.a_lt_b$in1[15] ));
 b15fpn000hn1n04x5 _632_ (.clk(clknet_2_1__leaf_clk),
    .d(_019_),
    .o(\dpath.a_lt_b$in0[0] ));
 b15fpn000hn1n04x5 _633_ (.clk(clknet_2_1__leaf_clk),
    .d(_020_),
    .o(\dpath.a_lt_b$in0[1] ));
 b15fpn000hn1n04x5 _634_ (.clk(clknet_2_1__leaf_clk),
    .d(_021_),
    .o(\dpath.a_lt_b$in0[2] ));
 b15fpn000hn1n04x5 _635_ (.clk(clknet_2_1__leaf_clk),
    .d(_022_),
    .o(\dpath.a_lt_b$in0[3] ));
 b15fpn000hn1n04x5 _636_ (.clk(clknet_2_1__leaf_clk),
    .d(_023_),
    .o(\dpath.a_lt_b$in0[4] ));
 b15fpn000hn1n04x5 _637_ (.clk(clknet_2_1__leaf_clk),
    .d(_024_),
    .o(\dpath.a_lt_b$in0[5] ));
 b15fpn000hn1n04x5 _638_ (.clk(clknet_2_0__leaf_clk),
    .d(_025_),
    .o(\dpath.a_lt_b$in0[6] ));
 b15fpn000hn1n04x5 _639_ (.clk(clknet_2_0__leaf_clk),
    .d(_026_),
    .o(\dpath.a_lt_b$in0[7] ));
 b15fpn000hn1n04x5 _640_ (.clk(clknet_2_1__leaf_clk),
    .d(_027_),
    .o(\dpath.a_lt_b$in0[8] ));
 b15fpn000hn1n04x5 _641_ (.clk(clknet_2_0__leaf_clk),
    .d(_028_),
    .o(\dpath.a_lt_b$in0[9] ));
 b15fpn000hn1n04x5 _642_ (.clk(clknet_2_2__leaf_clk),
    .d(_029_),
    .o(\dpath.a_lt_b$in0[10] ));
 b15fpn000hn1n04x5 _643_ (.clk(clknet_2_2__leaf_clk),
    .d(_030_),
    .o(\dpath.a_lt_b$in0[11] ));
 b15fpn000hn1n04x5 _644_ (.clk(clknet_2_3__leaf_clk),
    .d(_031_),
    .o(\dpath.a_lt_b$in0[12] ));
 b15fpn000hn1n04x5 _645_ (.clk(clknet_2_3__leaf_clk),
    .d(_032_),
    .o(\dpath.a_lt_b$in0[13] ));
 b15fpn000hn1n04x5 _646_ (.clk(clknet_2_3__leaf_clk),
    .d(_033_),
    .o(\dpath.a_lt_b$in0[14] ));
 b15fpn000hn1n04x5 _647_ (.clk(clknet_2_3__leaf_clk),
    .d(_034_),
    .o(\dpath.a_lt_b$in0[15] ));
 b15ztpn00an1n08x5 PHY_13 ();
 b15ztpn00an1n08x5 PHY_14 ();
 b15ztpn00an1n08x5 PHY_15 ();
 b15ztpn00an1n08x5 PHY_16 ();
 b15ztpn00an1n08x5 PHY_17 ();
 b15ztpn00an1n08x5 PHY_18 ();
 b15ztpn00an1n08x5 PHY_19 ();
 b15ztpn00an1n08x5 PHY_20 ();
 b15ztpn00an1n08x5 PHY_21 ();
 b15ztpn00an1n08x5 PHY_22 ();
 b15ztpn00an1n08x5 PHY_23 ();
 b15ztpn00an1n08x5 PHY_24 ();
 b15ztpn00an1n08x5 PHY_25 ();
 b15ztpn00an1n08x5 PHY_26 ();
 b15ztpn00an1n08x5 PHY_27 ();
 b15ztpn00an1n08x5 PHY_28 ();
 b15ztpn00an1n08x5 PHY_29 ();
 b15ztpn00an1n08x5 PHY_30 ();
 b15ztpn00an1n08x5 PHY_31 ();
 b15ztpn00an1n08x5 PHY_32 ();
 b15ztpn00an1n08x5 PHY_33 ();
 b15ztpn00an1n08x5 PHY_34 ();
 b15ztpn00an1n08x5 PHY_35 ();
 b15bfn000ar1n02x5 input1 (.a(req_msg[0]),
    .o(net1));
 b15bfn000ar1n02x5 input2 (.a(req_msg[10]),
    .o(net2));
 b15bfn000ar1n02x5 input3 (.a(req_msg[11]),
    .o(net3));
 b15bfn000ar1n02x5 input4 (.a(req_msg[12]),
    .o(net4));
 b15bfn000ar1n02x5 input5 (.a(req_msg[13]),
    .o(net5));
 b15bfn000ar1n02x5 input6 (.a(req_msg[14]),
    .o(net6));
 b15bfn000ar1n02x5 input7 (.a(req_msg[15]),
    .o(net7));
 b15bfn000ar1n02x5 input8 (.a(req_msg[16]),
    .o(net8));
 b15bfn000ar1n02x5 input9 (.a(req_msg[17]),
    .o(net9));
 b15bfn000ar1n02x5 input10 (.a(req_msg[18]),
    .o(net10));
 b15bfn000ar1n02x5 input11 (.a(req_msg[19]),
    .o(net11));
 b15bfn000ar1n02x5 input12 (.a(req_msg[1]),
    .o(net12));
 b15bfn000ar1n02x5 input13 (.a(req_msg[20]),
    .o(net13));
 b15bfn000ar1n02x5 input14 (.a(req_msg[21]),
    .o(net14));
 b15bfn000ar1n02x5 input15 (.a(req_msg[22]),
    .o(net15));
 b15bfn000ar1n02x5 input16 (.a(req_msg[23]),
    .o(net16));
 b15bfn000ar1n02x5 input17 (.a(req_msg[24]),
    .o(net17));
 b15bfn000ar1n02x5 input18 (.a(req_msg[25]),
    .o(net18));
 b15bfn000ar1n02x5 input19 (.a(req_msg[26]),
    .o(net19));
 b15bfn000ar1n02x5 input20 (.a(req_msg[27]),
    .o(net20));
 b15bfn000ar1n02x5 input21 (.a(req_msg[28]),
    .o(net21));
 b15bfn000ar1n02x5 input22 (.a(req_msg[29]),
    .o(net22));
 b15bfn000ar1n02x5 input23 (.a(req_msg[2]),
    .o(net23));
 b15bfn000ar1n02x5 input24 (.a(req_msg[30]),
    .o(net24));
 b15bfn000ar1n02x5 input25 (.a(req_msg[31]),
    .o(net25));
 b15bfn000ar1n02x5 input26 (.a(req_msg[3]),
    .o(net26));
 b15bfn000ar1n02x5 input27 (.a(req_msg[4]),
    .o(net27));
 b15bfn000ar1n02x5 input28 (.a(req_msg[5]),
    .o(net28));
 b15bfn000ar1n02x5 input29 (.a(req_msg[6]),
    .o(net29));
 b15bfn000ar1n02x5 input30 (.a(req_msg[7]),
    .o(net30));
 b15bfn000ar1n02x5 input31 (.a(req_msg[8]),
    .o(net31));
 b15bfn000ar1n02x5 input32 (.a(req_msg[9]),
    .o(net32));
 b15bfn000ar1n02x5 input33 (.a(req_val),
    .o(net33));
 b15bfn000ar1n02x5 input34 (.a(reset),
    .o(net34));
 b15bfn000ar1n02x5 input35 (.a(resp_rdy),
    .o(net35));
 b15bfn000al1n02x5 output36 (.a(net36),
    .o(req_rdy));
 b15bfn000al1n02x5 output37 (.a(net37),
    .o(resp_msg[0]));
 b15bfn000al1n02x5 output38 (.a(net38),
    .o(resp_msg[10]));
 b15bfn000al1n02x5 output39 (.a(net39),
    .o(resp_msg[11]));
 b15bfn000al1n02x5 output40 (.a(net40),
    .o(resp_msg[12]));
 b15bfn000al1n02x5 output41 (.a(net41),
    .o(resp_msg[13]));
 b15bfn000al1n02x5 output42 (.a(net42),
    .o(resp_msg[14]));
 b15bfn000al1n02x5 output43 (.a(net43),
    .o(resp_msg[15]));
 b15bfn000al1n02x5 output44 (.a(net44),
    .o(resp_msg[1]));
 b15bfn000al1n02x5 output45 (.a(net45),
    .o(resp_msg[2]));
 b15bfn000al1n02x5 output46 (.a(net46),
    .o(resp_msg[3]));
 b15bfn000al1n02x5 output47 (.a(net47),
    .o(resp_msg[4]));
 b15bfn000al1n02x5 output48 (.a(net48),
    .o(resp_msg[5]));
 b15bfn000al1n02x5 output49 (.a(net49),
    .o(resp_msg[6]));
 b15bfn000al1n02x5 output50 (.a(net50),
    .o(resp_msg[7]));
 b15bfn000al1n02x5 output51 (.a(net51),
    .o(resp_msg[8]));
 b15bfn000al1n02x5 output52 (.a(net52),
    .o(resp_msg[9]));
 b15bfn000al1n02x5 output53 (.a(net53),
    .o(resp_val));
 b15cbf000an1n16x5 clkbuf_0_clk (.clk(clk),
    .clkout(clknet_0_clk));
 b15cbf000an1n16x5 clkbuf_2_0__f_clk (.clk(clknet_0_clk),
    .clkout(clknet_2_0__leaf_clk));
 b15cbf000an1n16x5 clkbuf_2_1__f_clk (.clk(clknet_0_clk),
    .clkout(clknet_2_1__leaf_clk));
 b15cbf000an1n16x5 clkbuf_2_2__f_clk (.clk(clknet_0_clk),
    .clkout(clknet_2_2__leaf_clk));
 b15cbf000an1n16x5 clkbuf_2_3__f_clk (.clk(clknet_0_clk),
    .clkout(clknet_2_3__leaf_clk));
 b15zdnd11an1n08x5 FILLER_0_8 ();
 b15zdnd00an1n02x5 FILLER_0_16 ();
 b15zdnd00an1n01x5 FILLER_0_18 ();
 b15zdnd11an1n04x5 FILLER_0_23 ();
 b15zdnd11an1n04x5 FILLER_0_31 ();
 b15zdnd00an1n01x5 FILLER_0_35 ();
 b15zdnd11an1n08x5 FILLER_0_40 ();
 b15zdnd11an1n04x5 FILLER_0_48 ();
 b15zdnd00an1n01x5 FILLER_0_52 ();
 b15zdnd11an1n08x5 FILLER_0_57 ();
 b15zdnd11an1n04x5 FILLER_0_65 ();
 b15zdnd00an1n02x5 FILLER_0_69 ();
 b15zdnd11an1n04x5 FILLER_0_75 ();
 b15zdnd11an1n04x5 FILLER_0_83 ();
 b15zdnd11an1n04x5 FILLER_0_91 ();
 b15zdnd00an1n02x5 FILLER_0_95 ();
 b15zdnd11an1n04x5 FILLER_0_101 ();
 b15zdnd00an1n02x5 FILLER_0_105 ();
 b15zdnd00an1n01x5 FILLER_0_107 ();
 b15zdnd11an1n04x5 FILLER_0_112 ();
 b15zdnd00an1n01x5 FILLER_0_116 ();
 b15zdnd11an1n04x5 FILLER_0_121 ();
 b15zdnd00an1n02x5 FILLER_0_125 ();
 b15zdnd00an1n01x5 FILLER_0_127 ();
 b15zdnd11an1n08x5 FILLER_0_132 ();
 b15zdnd11an1n04x5 FILLER_0_140 ();
 b15zdnd00an1n02x5 FILLER_0_144 ();
 b15zdnd11an1n04x5 FILLER_0_150 ();
 b15zdnd11an1n04x5 FILLER_0_158 ();
 b15zdnd11an1n04x5 FILLER_0_166 ();
 b15zdnd11an1n04x5 FILLER_0_174 ();
 b15zdnd00an1n02x5 FILLER_0_178 ();
 b15zdnd00an1n01x5 FILLER_0_180 ();
 b15zdnd11an1n16x5 FILLER_0_185 ();
 b15zdnd11an1n04x5 FILLER_0_201 ();
 b15zdnd00an1n01x5 FILLER_0_205 ();
 b15zdnd11an1n16x5 FILLER_1_0 ();
 b15zdnd11an1n04x5 FILLER_1_20 ();
 b15zdnd11an1n08x5 FILLER_1_29 ();
 b15zdnd11an1n04x5 FILLER_1_41 ();
 b15zdnd00an1n01x5 FILLER_1_45 ();
 b15zdnd11an1n04x5 FILLER_1_51 ();
 b15zdnd11an1n08x5 FILLER_1_61 ();
 b15zdnd00an1n01x5 FILLER_1_69 ();
 b15zdnd11an1n08x5 FILLER_1_74 ();
 b15zdnd11an1n04x5 FILLER_1_82 ();
 b15zdnd00an1n02x5 FILLER_1_86 ();
 b15zdnd00an1n01x5 FILLER_1_88 ();
 b15zdnd11an1n04x5 FILLER_1_93 ();
 b15zdnd11an1n04x5 FILLER_1_101 ();
 b15zdnd11an1n04x5 FILLER_1_109 ();
 b15zdnd11an1n04x5 FILLER_1_119 ();
 b15zdnd11an1n32x5 FILLER_1_127 ();
 b15zdnd00an1n02x5 FILLER_1_159 ();
 b15zdnd11an1n04x5 FILLER_1_166 ();
 b15zdnd00an1n02x5 FILLER_1_170 ();
 b15zdnd00an1n01x5 FILLER_1_172 ();
 b15zdnd11an1n04x5 FILLER_1_179 ();
 b15zdnd11an1n04x5 FILLER_1_188 ();
 b15zdnd11an1n08x5 FILLER_1_196 ();
 b15zdnd11an1n04x5 FILLER_1_204 ();
 b15zdnd00an1n02x5 FILLER_1_212 ();
 b15zdnd11an1n08x5 FILLER_2_8 ();
 b15zdnd11an1n04x5 FILLER_2_16 ();
 b15zdnd00an1n02x5 FILLER_2_20 ();
 b15zdnd11an1n16x5 FILLER_2_27 ();
 b15zdnd00an1n02x5 FILLER_2_43 ();
 b15zdnd11an1n04x5 FILLER_2_50 ();
 b15zdnd11an1n04x5 FILLER_2_74 ();
 b15zdnd11an1n08x5 FILLER_2_83 ();
 b15zdnd11an1n04x5 FILLER_2_96 ();
 b15zdnd00an1n01x5 FILLER_2_100 ();
 b15zdnd11an1n04x5 FILLER_2_110 ();
 b15zdnd00an1n02x5 FILLER_2_114 ();
 b15zdnd00an1n01x5 FILLER_2_116 ();
 b15zdnd11an1n04x5 FILLER_2_122 ();
 b15zdnd11an1n16x5 FILLER_2_131 ();
 b15zdnd00an1n01x5 FILLER_2_147 ();
 b15zdnd11an1n04x5 FILLER_2_153 ();
 b15zdnd11an1n04x5 FILLER_2_166 ();
 b15zdnd11an1n08x5 FILLER_2_175 ();
 b15zdnd00an1n01x5 FILLER_2_183 ();
 b15zdnd00an1n02x5 FILLER_2_204 ();
 b15zdnd11an1n16x5 FILLER_3_0 ();
 b15zdnd11an1n04x5 FILLER_3_16 ();
 b15zdnd00an1n01x5 FILLER_3_20 ();
 b15zdnd11an1n32x5 FILLER_3_26 ();
 b15zdnd11an1n08x5 FILLER_3_58 ();
 b15zdnd00an1n02x5 FILLER_3_66 ();
 b15zdnd11an1n04x5 FILLER_3_72 ();
 b15zdnd11an1n08x5 FILLER_3_82 ();
 b15zdnd00an1n01x5 FILLER_3_90 ();
 b15zdnd11an1n04x5 FILLER_3_96 ();
 b15zdnd00an1n02x5 FILLER_3_100 ();
 b15zdnd11an1n04x5 FILLER_3_122 ();
 b15zdnd11an1n08x5 FILLER_3_146 ();
 b15zdnd11an1n04x5 FILLER_3_154 ();
 b15zdnd00an1n01x5 FILLER_3_158 ();
 b15zdnd11an1n08x5 FILLER_3_179 ();
 b15zdnd11an1n04x5 FILLER_3_187 ();
 b15zdnd00an1n01x5 FILLER_3_191 ();
 b15zdnd00an1n02x5 FILLER_3_212 ();
 b15zdnd11an1n04x5 FILLER_4_8 ();
 b15zdnd11an1n04x5 FILLER_4_16 ();
 b15zdnd11an1n32x5 FILLER_4_25 ();
 b15zdnd00an1n01x5 FILLER_4_57 ();
 b15zdnd11an1n16x5 FILLER_4_78 ();
 b15zdnd11an1n08x5 FILLER_4_94 ();
 b15zdnd11an1n04x5 FILLER_4_122 ();
 b15zdnd11an1n32x5 FILLER_4_146 ();
 b15zdnd11an1n16x5 FILLER_4_178 ();
 b15zdnd11an1n08x5 FILLER_4_194 ();
 b15zdnd11an1n04x5 FILLER_4_202 ();
 b15zdnd00an1n02x5 FILLER_5_0 ();
 b15zdnd00an1n01x5 FILLER_5_2 ();
 b15zdnd11an1n08x5 FILLER_5_7 ();
 b15zdnd11an1n04x5 FILLER_5_21 ();
 b15zdnd11an1n08x5 FILLER_5_28 ();
 b15zdnd00an1n02x5 FILLER_5_36 ();
 b15zdnd00an1n01x5 FILLER_5_38 ();
 b15zdnd11an1n08x5 FILLER_5_45 ();
 b15zdnd00an1n02x5 FILLER_5_53 ();
 b15zdnd11an1n32x5 FILLER_5_58 ();
 b15zdnd00an1n02x5 FILLER_5_90 ();
 b15zdnd11an1n64x5 FILLER_5_97 ();
 b15zdnd11an1n16x5 FILLER_5_161 ();
 b15zdnd11an1n04x5 FILLER_5_177 ();
 b15zdnd00an1n02x5 FILLER_5_181 ();
 b15zdnd11an1n08x5 FILLER_5_187 ();
 b15zdnd00an1n01x5 FILLER_5_195 ();
 b15zdnd11an1n08x5 FILLER_5_200 ();
 b15zdnd11an1n04x5 FILLER_5_208 ();
 b15zdnd00an1n02x5 FILLER_5_212 ();
 b15zdnd11an1n08x5 FILLER_6_8 ();
 b15zdnd11an1n04x5 FILLER_6_16 ();
 b15zdnd00an1n02x5 FILLER_6_20 ();
 b15zdnd00an1n01x5 FILLER_6_22 ();
 b15zdnd11an1n04x5 FILLER_6_27 ();
 b15zdnd11an1n04x5 FILLER_6_39 ();
 b15zdnd00an1n02x5 FILLER_6_43 ();
 b15zdnd00an1n01x5 FILLER_6_45 ();
 b15zdnd11an1n04x5 FILLER_6_54 ();
 b15zdnd11an1n04x5 FILLER_6_78 ();
 b15zdnd00an1n02x5 FILLER_6_82 ();
 b15zdnd00an1n01x5 FILLER_6_84 ();
 b15zdnd11an1n04x5 FILLER_6_89 ();
 b15zdnd11an1n16x5 FILLER_6_98 ();
 b15zdnd00an1n02x5 FILLER_6_114 ();
 b15zdnd00an1n01x5 FILLER_6_116 ();
 b15zdnd11an1n32x5 FILLER_6_137 ();
 b15zdnd11an1n32x5 FILLER_6_174 ();
 b15zdnd11an1n16x5 FILLER_7_0 ();
 b15zdnd11an1n08x5 FILLER_7_16 ();
 b15zdnd00an1n02x5 FILLER_7_24 ();
 b15zdnd11an1n04x5 FILLER_7_35 ();
 b15zdnd11an1n04x5 FILLER_7_51 ();
 b15zdnd11an1n04x5 FILLER_7_59 ();
 b15zdnd00an1n02x5 FILLER_7_63 ();
 b15zdnd00an1n01x5 FILLER_7_65 ();
 b15zdnd11an1n04x5 FILLER_7_86 ();
 b15zdnd11an1n32x5 FILLER_7_103 ();
 b15zdnd11an1n16x5 FILLER_7_135 ();
 b15zdnd11an1n08x5 FILLER_7_151 ();
 b15zdnd00an1n02x5 FILLER_7_159 ();
 b15zdnd00an1n01x5 FILLER_7_161 ();
 b15zdnd11an1n32x5 FILLER_7_182 ();
 b15zdnd00an1n02x5 FILLER_8_8 ();
 b15zdnd00an1n01x5 FILLER_8_10 ();
 b15zdnd11an1n04x5 FILLER_8_20 ();
 b15zdnd11an1n04x5 FILLER_8_39 ();
 b15zdnd11an1n04x5 FILLER_8_48 ();
 b15zdnd11an1n16x5 FILLER_8_56 ();
 b15zdnd00an1n01x5 FILLER_8_72 ();
 b15zdnd11an1n04x5 FILLER_8_82 ();
 b15zdnd11an1n32x5 FILLER_8_106 ();
 b15zdnd11an1n04x5 FILLER_8_138 ();
 b15zdnd00an1n02x5 FILLER_8_142 ();
 b15zdnd11an1n04x5 FILLER_8_164 ();
 b15zdnd00an1n01x5 FILLER_8_168 ();
 b15zdnd11an1n08x5 FILLER_8_174 ();
 b15zdnd00an1n02x5 FILLER_8_182 ();
 b15zdnd00an1n02x5 FILLER_8_204 ();
 b15zdnd00an1n02x5 FILLER_9_0 ();
 b15zdnd11an1n04x5 FILLER_9_6 ();
 b15zdnd11an1n08x5 FILLER_9_13 ();
 b15zdnd00an1n02x5 FILLER_9_21 ();
 b15zdnd00an1n01x5 FILLER_9_23 ();
 b15zdnd11an1n08x5 FILLER_9_32 ();
 b15zdnd00an1n02x5 FILLER_9_40 ();
 b15zdnd00an1n01x5 FILLER_9_42 ();
 b15zdnd11an1n16x5 FILLER_9_47 ();
 b15zdnd11an1n08x5 FILLER_9_63 ();
 b15zdnd11an1n04x5 FILLER_9_71 ();
 b15zdnd00an1n01x5 FILLER_9_75 ();
 b15zdnd11an1n04x5 FILLER_9_82 ();
 b15zdnd11an1n16x5 FILLER_9_106 ();
 b15zdnd11an1n04x5 FILLER_9_122 ();
 b15zdnd11an1n04x5 FILLER_9_146 ();
 b15zdnd11an1n08x5 FILLER_9_159 ();
 b15zdnd11an1n04x5 FILLER_9_167 ();
 b15zdnd11an1n16x5 FILLER_9_175 ();
 b15zdnd11an1n04x5 FILLER_9_191 ();
 b15zdnd00an1n01x5 FILLER_9_195 ();
 b15zdnd11an1n08x5 FILLER_9_200 ();
 b15zdnd11an1n04x5 FILLER_9_208 ();
 b15zdnd00an1n02x5 FILLER_9_212 ();
 b15zdnd00an1n02x5 FILLER_10_8 ();
 b15zdnd11an1n08x5 FILLER_10_14 ();
 b15zdnd11an1n08x5 FILLER_10_26 ();
 b15zdnd11an1n04x5 FILLER_10_39 ();
 b15zdnd11an1n04x5 FILLER_10_48 ();
 b15zdnd00an1n02x5 FILLER_10_52 ();
 b15zdnd00an1n01x5 FILLER_10_54 ();
 b15zdnd11an1n04x5 FILLER_10_75 ();
 b15zdnd11an1n04x5 FILLER_10_84 ();
 b15zdnd11an1n32x5 FILLER_10_92 ();
 b15zdnd11an1n16x5 FILLER_10_124 ();
 b15zdnd11an1n04x5 FILLER_10_140 ();
 b15zdnd11an1n08x5 FILLER_10_164 ();
 b15zdnd11an1n04x5 FILLER_10_172 ();
 b15zdnd11an1n04x5 FILLER_10_196 ();
 b15zdnd00an1n02x5 FILLER_10_204 ();
 b15zdnd11an1n16x5 FILLER_11_0 ();
 b15zdnd11an1n04x5 FILLER_11_21 ();
 b15zdnd11an1n04x5 FILLER_11_28 ();
 b15zdnd00an1n02x5 FILLER_11_32 ();
 b15zdnd11an1n08x5 FILLER_11_40 ();
 b15zdnd11an1n04x5 FILLER_11_48 ();
 b15zdnd11an1n16x5 FILLER_11_56 ();
 b15zdnd00an1n01x5 FILLER_11_72 ();
 b15zdnd11an1n64x5 FILLER_11_78 ();
 b15zdnd11an1n08x5 FILLER_11_142 ();
 b15zdnd11an1n04x5 FILLER_11_150 ();
 b15zdnd00an1n02x5 FILLER_11_154 ();
 b15zdnd00an1n01x5 FILLER_11_156 ();
 b15zdnd11an1n04x5 FILLER_11_166 ();
 b15zdnd11an1n04x5 FILLER_11_174 ();
 b15zdnd11an1n08x5 FILLER_11_198 ();
 b15zdnd11an1n04x5 FILLER_11_210 ();
 b15zdnd11an1n08x5 FILLER_12_8 ();
 b15zdnd11an1n04x5 FILLER_12_16 ();
 b15zdnd00an1n02x5 FILLER_12_20 ();
 b15zdnd11an1n04x5 FILLER_12_28 ();
 b15zdnd00an1n02x5 FILLER_12_32 ();
 b15zdnd11an1n08x5 FILLER_12_38 ();
 b15zdnd00an1n02x5 FILLER_12_46 ();
 b15zdnd11an1n08x5 FILLER_12_53 ();
 b15zdnd00an1n02x5 FILLER_12_61 ();
 b15zdnd11an1n64x5 FILLER_12_83 ();
 b15zdnd11an1n08x5 FILLER_12_147 ();
 b15zdnd11an1n04x5 FILLER_12_155 ();
 b15zdnd00an1n01x5 FILLER_12_159 ();
 b15zdnd11an1n04x5 FILLER_12_180 ();
 b15zdnd00an1n02x5 FILLER_12_204 ();
 b15zdnd11an1n16x5 FILLER_13_0 ();
 b15zdnd00an1n02x5 FILLER_13_16 ();
 b15zdnd00an1n01x5 FILLER_13_18 ();
 b15zdnd11an1n08x5 FILLER_13_25 ();
 b15zdnd00an1n02x5 FILLER_13_33 ();
 b15zdnd11an1n16x5 FILLER_13_44 ();
 b15zdnd00an1n02x5 FILLER_13_60 ();
 b15zdnd00an1n01x5 FILLER_13_62 ();
 b15zdnd11an1n04x5 FILLER_13_83 ();
 b15zdnd11an1n04x5 FILLER_13_107 ();
 b15zdnd11an1n04x5 FILLER_13_131 ();
 b15zdnd11an1n04x5 FILLER_13_155 ();
 b15zdnd11an1n08x5 FILLER_13_179 ();
 b15zdnd11an1n04x5 FILLER_13_187 ();
 b15zdnd00an1n01x5 FILLER_13_191 ();
 b15zdnd00an1n02x5 FILLER_13_212 ();
 b15zdnd11an1n08x5 FILLER_14_8 ();
 b15zdnd00an1n02x5 FILLER_14_16 ();
 b15zdnd11an1n04x5 FILLER_14_22 ();
 b15zdnd11an1n08x5 FILLER_14_30 ();
 b15zdnd00an1n02x5 FILLER_14_38 ();
 b15zdnd11an1n04x5 FILLER_14_45 ();
 b15zdnd11an1n04x5 FILLER_14_61 ();
 b15zdnd00an1n02x5 FILLER_14_65 ();
 b15zdnd00an1n01x5 FILLER_14_67 ();
 b15zdnd11an1n04x5 FILLER_14_88 ();
 b15zdnd11an1n32x5 FILLER_14_112 ();
 b15zdnd11an1n16x5 FILLER_14_144 ();
 b15zdnd11an1n08x5 FILLER_14_160 ();
 b15zdnd11an1n04x5 FILLER_14_188 ();
 b15zdnd11an1n04x5 FILLER_14_196 ();
 b15zdnd00an1n02x5 FILLER_14_204 ();
 b15zdnd00an1n02x5 FILLER_15_0 ();
 b15zdnd11an1n08x5 FILLER_15_6 ();
 b15zdnd11an1n04x5 FILLER_15_14 ();
 b15zdnd00an1n02x5 FILLER_15_18 ();
 b15zdnd00an1n01x5 FILLER_15_20 ();
 b15zdnd11an1n08x5 FILLER_15_25 ();
 b15zdnd00an1n02x5 FILLER_15_33 ();
 b15zdnd00an1n01x5 FILLER_15_35 ();
 b15zdnd11an1n04x5 FILLER_15_42 ();
 b15zdnd11an1n04x5 FILLER_15_51 ();
 b15zdnd11an1n08x5 FILLER_15_59 ();
 b15zdnd11an1n04x5 FILLER_15_67 ();
 b15zdnd11an1n04x5 FILLER_15_74 ();
 b15zdnd11an1n16x5 FILLER_15_83 ();
 b15zdnd11an1n04x5 FILLER_15_99 ();
 b15zdnd00an1n01x5 FILLER_15_103 ();
 b15zdnd11an1n04x5 FILLER_15_124 ();
 b15zdnd11an1n08x5 FILLER_15_132 ();
 b15zdnd11an1n04x5 FILLER_15_140 ();
 b15zdnd11an1n16x5 FILLER_15_150 ();
 b15zdnd11an1n04x5 FILLER_15_166 ();
 b15zdnd00an1n02x5 FILLER_15_170 ();
 b15zdnd00an1n01x5 FILLER_15_172 ();
 b15zdnd11an1n04x5 FILLER_15_178 ();
 b15zdnd00an1n02x5 FILLER_15_182 ();
 b15zdnd00an1n01x5 FILLER_15_184 ();
 b15zdnd11an1n04x5 FILLER_15_191 ();
 b15zdnd11an1n04x5 FILLER_15_200 ();
 b15zdnd11an1n04x5 FILLER_15_208 ();
 b15zdnd00an1n02x5 FILLER_15_212 ();
 b15zdnd11an1n04x5 FILLER_16_8 ();
 b15zdnd11an1n04x5 FILLER_16_19 ();
 b15zdnd00an1n01x5 FILLER_16_23 ();
 b15zdnd11an1n04x5 FILLER_16_35 ();
 b15zdnd11an1n04x5 FILLER_16_43 ();
 b15zdnd11an1n16x5 FILLER_16_54 ();
 b15zdnd11an1n04x5 FILLER_16_70 ();
 b15zdnd00an1n02x5 FILLER_16_74 ();
 b15zdnd00an1n01x5 FILLER_16_76 ();
 b15zdnd11an1n04x5 FILLER_16_81 ();
 b15zdnd11an1n08x5 FILLER_16_89 ();
 b15zdnd00an1n02x5 FILLER_16_97 ();
 b15zdnd11an1n16x5 FILLER_16_111 ();
 b15zdnd11an1n04x5 FILLER_16_127 ();
 b15zdnd11an1n08x5 FILLER_16_134 ();
 b15zdnd11an1n04x5 FILLER_16_142 ();
 b15zdnd11an1n04x5 FILLER_16_156 ();
 b15zdnd11an1n08x5 FILLER_16_166 ();
 b15zdnd11an1n04x5 FILLER_16_178 ();
 b15zdnd11an1n04x5 FILLER_16_187 ();
 b15zdnd00an1n01x5 FILLER_16_191 ();
 b15zdnd11an1n04x5 FILLER_16_200 ();
 b15zdnd00an1n02x5 FILLER_16_204 ();
 b15zdnd11an1n16x5 FILLER_17_0 ();
 b15zdnd00an1n01x5 FILLER_17_16 ();
 b15zdnd11an1n04x5 FILLER_17_22 ();
 b15zdnd11an1n04x5 FILLER_17_31 ();
 b15zdnd11an1n04x5 FILLER_17_40 ();
 b15zdnd11an1n32x5 FILLER_17_47 ();
 b15zdnd11an1n04x5 FILLER_17_79 ();
 b15zdnd11an1n04x5 FILLER_17_95 ();
 b15zdnd11an1n16x5 FILLER_17_102 ();
 b15zdnd11an1n08x5 FILLER_17_118 ();
 b15zdnd00an1n02x5 FILLER_17_126 ();
 b15zdnd11an1n32x5 FILLER_17_134 ();
 b15zdnd00an1n01x5 FILLER_17_166 ();
 b15zdnd11an1n04x5 FILLER_17_173 ();
 b15zdnd11an1n04x5 FILLER_17_181 ();
 b15zdnd11an1n04x5 FILLER_17_188 ();
 b15zdnd00an1n01x5 FILLER_17_192 ();
 b15zdnd11an1n16x5 FILLER_17_198 ();
 b15zdnd00an1n02x5 FILLER_18_8 ();
 b15zdnd11an1n04x5 FILLER_18_14 ();
 b15zdnd11an1n16x5 FILLER_18_22 ();
 b15zdnd11an1n04x5 FILLER_18_44 ();
 b15zdnd11an1n32x5 FILLER_18_54 ();
 b15zdnd11an1n04x5 FILLER_18_86 ();
 b15zdnd00an1n02x5 FILLER_18_90 ();
 b15zdnd11an1n04x5 FILLER_18_96 ();
 b15zdnd11an1n16x5 FILLER_18_104 ();
 b15zdnd00an1n02x5 FILLER_18_120 ();
 b15zdnd00an1n01x5 FILLER_18_122 ();
 b15zdnd11an1n16x5 FILLER_18_129 ();
 b15zdnd11an1n04x5 FILLER_18_145 ();
 b15zdnd11an1n08x5 FILLER_18_154 ();
 b15zdnd00an1n01x5 FILLER_18_162 ();
 b15zdnd11an1n16x5 FILLER_18_187 ();
 b15zdnd00an1n02x5 FILLER_18_203 ();
 b15zdnd00an1n01x5 FILLER_18_205 ();
 b15zdnd00an1n02x5 FILLER_19_0 ();
 b15zdnd11an1n04x5 FILLER_19_6 ();
 b15zdnd00an1n01x5 FILLER_19_10 ();
 b15zdnd11an1n04x5 FILLER_19_15 ();
 b15zdnd11an1n04x5 FILLER_19_36 ();
 b15zdnd11an1n04x5 FILLER_19_46 ();
 b15zdnd00an1n01x5 FILLER_19_50 ();
 b15zdnd11an1n08x5 FILLER_19_63 ();
 b15zdnd00an1n02x5 FILLER_19_71 ();
 b15zdnd00an1n01x5 FILLER_19_73 ();
 b15zdnd11an1n04x5 FILLER_19_80 ();
 b15zdnd11an1n04x5 FILLER_19_89 ();
 b15zdnd11an1n04x5 FILLER_19_98 ();
 b15zdnd11an1n08x5 FILLER_19_105 ();
 b15zdnd11an1n04x5 FILLER_19_113 ();
 b15zdnd00an1n01x5 FILLER_19_117 ();
 b15zdnd11an1n04x5 FILLER_19_122 ();
 b15zdnd11an1n08x5 FILLER_19_130 ();
 b15zdnd00an1n01x5 FILLER_19_138 ();
 b15zdnd11an1n04x5 FILLER_19_145 ();
 b15zdnd00an1n02x5 FILLER_19_149 ();
 b15zdnd00an1n01x5 FILLER_19_151 ();
 b15zdnd11an1n08x5 FILLER_19_156 ();
 b15zdnd00an1n01x5 FILLER_19_164 ();
 b15zdnd11an1n16x5 FILLER_19_171 ();
 b15zdnd11an1n04x5 FILLER_19_187 ();
 b15zdnd00an1n01x5 FILLER_19_191 ();
 b15zdnd11an1n16x5 FILLER_19_196 ();
 b15zdnd00an1n02x5 FILLER_19_212 ();
 b15zdnd11an1n32x5 FILLER_20_8 ();
 b15zdnd11an1n04x5 FILLER_20_40 ();
 b15zdnd00an1n02x5 FILLER_20_44 ();
 b15zdnd00an1n01x5 FILLER_20_46 ();
 b15zdnd11an1n04x5 FILLER_20_51 ();
 b15zdnd11an1n08x5 FILLER_20_61 ();
 b15zdnd11an1n04x5 FILLER_20_84 ();
 b15zdnd00an1n01x5 FILLER_20_88 ();
 b15zdnd11an1n04x5 FILLER_20_95 ();
 b15zdnd11an1n08x5 FILLER_20_105 ();
 b15zdnd11an1n04x5 FILLER_20_113 ();
 b15zdnd00an1n02x5 FILLER_20_117 ();
 b15zdnd00an1n01x5 FILLER_20_119 ();
 b15zdnd11an1n04x5 FILLER_20_125 ();
 b15zdnd11an1n08x5 FILLER_20_132 ();
 b15zdnd11an1n04x5 FILLER_20_145 ();
 b15zdnd00an1n01x5 FILLER_20_149 ();
 b15zdnd11an1n16x5 FILLER_20_155 ();
 b15zdnd11an1n04x5 FILLER_20_194 ();
 b15zdnd00an1n02x5 FILLER_20_203 ();
 b15zdnd00an1n01x5 FILLER_20_205 ();
 b15zdnd11an1n16x5 FILLER_21_0 ();
 b15zdnd11an1n04x5 FILLER_21_21 ();
 b15zdnd11an1n32x5 FILLER_21_30 ();
 b15zdnd11an1n16x5 FILLER_21_62 ();
 b15zdnd11an1n08x5 FILLER_21_78 ();
 b15zdnd11an1n04x5 FILLER_21_92 ();
 b15zdnd00an1n01x5 FILLER_21_96 ();
 b15zdnd11an1n08x5 FILLER_21_105 ();
 b15zdnd11an1n04x5 FILLER_21_113 ();
 b15zdnd00an1n02x5 FILLER_21_117 ();
 b15zdnd11an1n32x5 FILLER_21_122 ();
 b15zdnd11an1n08x5 FILLER_21_154 ();
 b15zdnd11an1n04x5 FILLER_21_162 ();
 b15zdnd11an1n04x5 FILLER_21_173 ();
 b15zdnd11an1n08x5 FILLER_21_181 ();
 b15zdnd11an1n04x5 FILLER_21_189 ();
 b15zdnd00an1n02x5 FILLER_21_193 ();
 b15zdnd11an1n04x5 FILLER_21_200 ();
 b15zdnd11an1n04x5 FILLER_21_208 ();
 b15zdnd00an1n02x5 FILLER_21_212 ();
 b15zdnd11an1n04x5 FILLER_22_8 ();
 b15zdnd11an1n32x5 FILLER_22_16 ();
 b15zdnd11an1n08x5 FILLER_22_48 ();
 b15zdnd00an1n02x5 FILLER_22_56 ();
 b15zdnd11an1n16x5 FILLER_22_62 ();
 b15zdnd11an1n04x5 FILLER_22_78 ();
 b15zdnd00an1n02x5 FILLER_22_82 ();
 b15zdnd00an1n01x5 FILLER_22_84 ();
 b15zdnd11an1n04x5 FILLER_22_93 ();
 b15zdnd00an1n02x5 FILLER_22_97 ();
 b15zdnd11an1n08x5 FILLER_22_105 ();
 b15zdnd11an1n04x5 FILLER_22_113 ();
 b15zdnd11an1n04x5 FILLER_22_123 ();
 b15zdnd11an1n04x5 FILLER_22_132 ();
 b15zdnd11an1n08x5 FILLER_22_139 ();
 b15zdnd11an1n04x5 FILLER_22_151 ();
 b15zdnd11an1n04x5 FILLER_22_158 ();
 b15zdnd11an1n16x5 FILLER_22_165 ();
 b15zdnd11an1n04x5 FILLER_22_189 ();
 b15zdnd11an1n04x5 FILLER_22_196 ();
 b15zdnd00an1n02x5 FILLER_22_204 ();
 b15zdnd00an1n02x5 FILLER_23_0 ();
 b15zdnd11an1n04x5 FILLER_23_6 ();
 b15zdnd11an1n04x5 FILLER_23_14 ();
 b15zdnd11an1n04x5 FILLER_23_24 ();
 b15zdnd11an1n04x5 FILLER_23_31 ();
 b15zdnd11an1n04x5 FILLER_23_39 ();
 b15zdnd11an1n08x5 FILLER_23_47 ();
 b15zdnd00an1n02x5 FILLER_23_55 ();
 b15zdnd00an1n01x5 FILLER_23_57 ();
 b15zdnd11an1n04x5 FILLER_23_64 ();
 b15zdnd11an1n16x5 FILLER_23_73 ();
 b15zdnd11an1n04x5 FILLER_23_89 ();
 b15zdnd00an1n02x5 FILLER_23_93 ();
 b15zdnd00an1n01x5 FILLER_23_95 ();
 b15zdnd11an1n08x5 FILLER_23_109 ();
 b15zdnd11an1n04x5 FILLER_23_117 ();
 b15zdnd00an1n02x5 FILLER_23_121 ();
 b15zdnd11an1n04x5 FILLER_23_128 ();
 b15zdnd00an1n01x5 FILLER_23_132 ();
 b15zdnd11an1n04x5 FILLER_23_136 ();
 b15zdnd00an1n02x5 FILLER_23_140 ();
 b15zdnd11an1n08x5 FILLER_23_146 ();
 b15zdnd11an1n04x5 FILLER_23_154 ();
 b15zdnd11an1n16x5 FILLER_23_162 ();
 b15zdnd11an1n04x5 FILLER_23_178 ();
 b15zdnd11an1n08x5 FILLER_23_186 ();
 b15zdnd11an1n08x5 FILLER_23_200 ();
 b15zdnd00an1n02x5 FILLER_23_212 ();
 b15zdnd00an1n02x5 FILLER_24_8 ();
 b15zdnd11an1n04x5 FILLER_24_19 ();
 b15zdnd11an1n04x5 FILLER_24_35 ();
 b15zdnd00an1n02x5 FILLER_24_39 ();
 b15zdnd00an1n01x5 FILLER_24_41 ();
 b15zdnd11an1n08x5 FILLER_24_50 ();
 b15zdnd00an1n01x5 FILLER_24_58 ();
 b15zdnd11an1n08x5 FILLER_24_64 ();
 b15zdnd00an1n01x5 FILLER_24_72 ();
 b15zdnd11an1n04x5 FILLER_24_83 ();
 b15zdnd00an1n02x5 FILLER_24_87 ();
 b15zdnd00an1n01x5 FILLER_24_89 ();
 b15zdnd11an1n08x5 FILLER_24_94 ();
 b15zdnd11an1n04x5 FILLER_24_102 ();
 b15zdnd00an1n02x5 FILLER_24_106 ();
 b15zdnd00an1n01x5 FILLER_24_108 ();
 b15zdnd11an1n04x5 FILLER_24_119 ();
 b15zdnd11an1n32x5 FILLER_24_126 ();
 b15zdnd11an1n08x5 FILLER_24_158 ();
 b15zdnd11an1n04x5 FILLER_24_166 ();
 b15zdnd00an1n02x5 FILLER_24_170 ();
 b15zdnd00an1n01x5 FILLER_24_172 ();
 b15zdnd11an1n04x5 FILLER_24_179 ();
 b15zdnd11an1n08x5 FILLER_24_190 ();
 b15zdnd00an1n02x5 FILLER_24_198 ();
 b15zdnd00an1n02x5 FILLER_24_204 ();
 b15zdnd11an1n16x5 FILLER_25_0 ();
 b15zdnd11an1n04x5 FILLER_25_16 ();
 b15zdnd11an1n04x5 FILLER_25_24 ();
 b15zdnd11an1n04x5 FILLER_25_32 ();
 b15zdnd00an1n02x5 FILLER_25_36 ();
 b15zdnd11an1n32x5 FILLER_25_43 ();
 b15zdnd11an1n04x5 FILLER_25_75 ();
 b15zdnd00an1n01x5 FILLER_25_79 ();
 b15zdnd11an1n16x5 FILLER_25_93 ();
 b15zdnd00an1n02x5 FILLER_25_109 ();
 b15zdnd00an1n01x5 FILLER_25_111 ();
 b15zdnd11an1n16x5 FILLER_25_123 ();
 b15zdnd00an1n01x5 FILLER_25_139 ();
 b15zdnd11an1n08x5 FILLER_25_144 ();
 b15zdnd11an1n04x5 FILLER_25_170 ();
 b15zdnd11an1n04x5 FILLER_25_182 ();
 b15zdnd11an1n04x5 FILLER_25_189 ();
 b15zdnd11an1n16x5 FILLER_25_198 ();
 b15zdnd11an1n08x5 FILLER_26_8 ();
 b15zdnd11an1n08x5 FILLER_26_24 ();
 b15zdnd00an1n01x5 FILLER_26_32 ();
 b15zdnd11an1n08x5 FILLER_26_43 ();
 b15zdnd00an1n02x5 FILLER_26_51 ();
 b15zdnd00an1n01x5 FILLER_26_53 ();
 b15zdnd11an1n16x5 FILLER_26_57 ();
 b15zdnd00an1n01x5 FILLER_26_73 ();
 b15zdnd11an1n16x5 FILLER_26_79 ();
 b15zdnd11an1n04x5 FILLER_26_95 ();
 b15zdnd00an1n02x5 FILLER_26_99 ();
 b15zdnd11an1n16x5 FILLER_26_106 ();
 b15zdnd11an1n08x5 FILLER_26_122 ();
 b15zdnd11an1n04x5 FILLER_26_130 ();
 b15zdnd00an1n02x5 FILLER_26_134 ();
 b15zdnd11an1n32x5 FILLER_26_141 ();
 b15zdnd00an1n02x5 FILLER_26_173 ();
 b15zdnd00an1n01x5 FILLER_26_175 ();
 b15zdnd11an1n04x5 FILLER_26_182 ();
 b15zdnd11an1n04x5 FILLER_26_190 ();
 b15zdnd00an1n02x5 FILLER_26_204 ();
 b15zdnd11an1n08x5 FILLER_27_0 ();
 b15zdnd00an1n02x5 FILLER_27_8 ();
 b15zdnd11an1n08x5 FILLER_27_14 ();
 b15zdnd00an1n02x5 FILLER_27_22 ();
 b15zdnd11an1n04x5 FILLER_27_27 ();
 b15zdnd00an1n02x5 FILLER_27_31 ();
 b15zdnd00an1n01x5 FILLER_27_33 ();
 b15zdnd11an1n16x5 FILLER_27_38 ();
 b15zdnd11an1n04x5 FILLER_27_54 ();
 b15zdnd00an1n01x5 FILLER_27_58 ();
 b15zdnd11an1n04x5 FILLER_27_63 ();
 b15zdnd11an1n08x5 FILLER_27_72 ();
 b15zdnd11an1n04x5 FILLER_27_80 ();
 b15zdnd00an1n01x5 FILLER_27_84 ();
 b15zdnd11an1n08x5 FILLER_27_89 ();
 b15zdnd11an1n04x5 FILLER_27_97 ();
 b15zdnd00an1n02x5 FILLER_27_101 ();
 b15zdnd11an1n16x5 FILLER_27_109 ();
 b15zdnd11an1n08x5 FILLER_27_125 ();
 b15zdnd00an1n02x5 FILLER_27_133 ();
 b15zdnd11an1n32x5 FILLER_27_140 ();
 b15zdnd11an1n08x5 FILLER_27_172 ();
 b15zdnd00an1n02x5 FILLER_27_180 ();
 b15zdnd11an1n04x5 FILLER_27_186 ();
 b15zdnd11an1n08x5 FILLER_27_194 ();
 b15zdnd11an1n04x5 FILLER_27_202 ();
 b15zdnd00an1n01x5 FILLER_27_206 ();
 b15zdnd00an1n02x5 FILLER_27_211 ();
 b15zdnd00an1n01x5 FILLER_27_213 ();
 b15zdnd11an1n04x5 FILLER_28_8 ();
 b15zdnd00an1n02x5 FILLER_28_12 ();
 b15zdnd11an1n08x5 FILLER_28_23 ();
 b15zdnd11an1n04x5 FILLER_28_41 ();
 b15zdnd11an1n08x5 FILLER_28_49 ();
 b15zdnd00an1n02x5 FILLER_28_57 ();
 b15zdnd00an1n01x5 FILLER_28_59 ();
 b15zdnd11an1n08x5 FILLER_28_65 ();
 b15zdnd00an1n02x5 FILLER_28_73 ();
 b15zdnd11an1n16x5 FILLER_28_80 ();
 b15zdnd11an1n04x5 FILLER_28_96 ();
 b15zdnd00an1n02x5 FILLER_28_100 ();
 b15zdnd11an1n16x5 FILLER_28_106 ();
 b15zdnd00an1n01x5 FILLER_28_122 ();
 b15zdnd11an1n04x5 FILLER_28_127 ();
 b15zdnd11an1n08x5 FILLER_28_140 ();
 b15zdnd11an1n04x5 FILLER_28_148 ();
 b15zdnd00an1n02x5 FILLER_28_152 ();
 b15zdnd00an1n01x5 FILLER_28_154 ();
 b15zdnd11an1n04x5 FILLER_28_171 ();
 b15zdnd11an1n08x5 FILLER_28_179 ();
 b15zdnd11an1n08x5 FILLER_28_195 ();
 b15zdnd00an1n02x5 FILLER_28_203 ();
 b15zdnd00an1n01x5 FILLER_28_205 ();
 b15zdnd00an1n02x5 FILLER_29_0 ();
 b15zdnd11an1n08x5 FILLER_29_6 ();
 b15zdnd00an1n01x5 FILLER_29_14 ();
 b15zdnd11an1n04x5 FILLER_29_19 ();
 b15zdnd11an1n04x5 FILLER_29_29 ();
 b15zdnd00an1n02x5 FILLER_29_33 ();
 b15zdnd11an1n08x5 FILLER_29_38 ();
 b15zdnd11an1n04x5 FILLER_29_46 ();
 b15zdnd00an1n02x5 FILLER_29_50 ();
 b15zdnd00an1n01x5 FILLER_29_52 ();
 b15zdnd11an1n04x5 FILLER_29_63 ();
 b15zdnd11an1n04x5 FILLER_29_73 ();
 b15zdnd11an1n04x5 FILLER_29_81 ();
 b15zdnd11an1n32x5 FILLER_29_88 ();
 b15zdnd11an1n04x5 FILLER_29_129 ();
 b15zdnd00an1n02x5 FILLER_29_133 ();
 b15zdnd11an1n04x5 FILLER_29_140 ();
 b15zdnd00an1n02x5 FILLER_29_144 ();
 b15zdnd00an1n01x5 FILLER_29_146 ();
 b15zdnd11an1n04x5 FILLER_29_151 ();
 b15zdnd00an1n01x5 FILLER_29_155 ();
 b15zdnd11an1n08x5 FILLER_29_162 ();
 b15zdnd00an1n02x5 FILLER_29_170 ();
 b15zdnd11an1n04x5 FILLER_29_177 ();
 b15zdnd11an1n04x5 FILLER_29_190 ();
 b15zdnd11an1n08x5 FILLER_29_200 ();
 b15zdnd11an1n04x5 FILLER_29_208 ();
 b15zdnd00an1n02x5 FILLER_29_212 ();
 b15zdnd11an1n08x5 FILLER_30_8 ();
 b15zdnd11an1n04x5 FILLER_30_16 ();
 b15zdnd00an1n02x5 FILLER_30_20 ();
 b15zdnd00an1n01x5 FILLER_30_22 ();
 b15zdnd11an1n32x5 FILLER_30_28 ();
 b15zdnd00an1n02x5 FILLER_30_60 ();
 b15zdnd11an1n04x5 FILLER_30_70 ();
 b15zdnd11an1n04x5 FILLER_30_77 ();
 b15zdnd11an1n04x5 FILLER_30_85 ();
 b15zdnd11an1n04x5 FILLER_30_93 ();
 b15zdnd11an1n08x5 FILLER_30_100 ();
 b15zdnd11an1n04x5 FILLER_30_108 ();
 b15zdnd00an1n01x5 FILLER_30_112 ();
 b15zdnd11an1n04x5 FILLER_30_117 ();
 b15zdnd00an1n01x5 FILLER_30_121 ();
 b15zdnd11an1n04x5 FILLER_30_125 ();
 b15zdnd11an1n04x5 FILLER_30_133 ();
 b15zdnd11an1n04x5 FILLER_30_141 ();
 b15zdnd11an1n08x5 FILLER_30_150 ();
 b15zdnd00an1n01x5 FILLER_30_158 ();
 b15zdnd11an1n16x5 FILLER_30_164 ();
 b15zdnd11an1n04x5 FILLER_30_180 ();
 b15zdnd00an1n02x5 FILLER_30_184 ();
 b15zdnd00an1n01x5 FILLER_30_186 ();
 b15zdnd11an1n04x5 FILLER_30_196 ();
 b15zdnd00an1n02x5 FILLER_30_204 ();
 b15zdnd00an1n02x5 FILLER_31_0 ();
 b15zdnd00an1n01x5 FILLER_31_2 ();
 b15zdnd11an1n16x5 FILLER_31_7 ();
 b15zdnd11an1n08x5 FILLER_31_29 ();
 b15zdnd11an1n16x5 FILLER_31_42 ();
 b15zdnd11an1n08x5 FILLER_31_58 ();
 b15zdnd00an1n01x5 FILLER_31_66 ();
 b15zdnd11an1n08x5 FILLER_31_76 ();
 b15zdnd11an1n04x5 FILLER_31_84 ();
 b15zdnd00an1n02x5 FILLER_31_88 ();
 b15zdnd11an1n08x5 FILLER_31_96 ();
 b15zdnd11an1n04x5 FILLER_31_104 ();
 b15zdnd00an1n02x5 FILLER_31_108 ();
 b15zdnd11an1n04x5 FILLER_31_115 ();
 b15zdnd11an1n04x5 FILLER_31_123 ();
 b15zdnd11an1n04x5 FILLER_31_131 ();
 b15zdnd11an1n32x5 FILLER_31_138 ();
 b15zdnd11an1n08x5 FILLER_31_170 ();
 b15zdnd11an1n04x5 FILLER_31_178 ();
 b15zdnd00an1n01x5 FILLER_31_182 ();
 b15zdnd11an1n04x5 FILLER_31_186 ();
 b15zdnd11an1n16x5 FILLER_31_194 ();
 b15zdnd11an1n04x5 FILLER_31_210 ();
 b15zdnd11an1n16x5 FILLER_32_8 ();
 b15zdnd11an1n04x5 FILLER_32_24 ();
 b15zdnd00an1n01x5 FILLER_32_28 ();
 b15zdnd11an1n04x5 FILLER_32_33 ();
 b15zdnd11an1n16x5 FILLER_32_43 ();
 b15zdnd11an1n04x5 FILLER_32_59 ();
 b15zdnd11an1n08x5 FILLER_32_68 ();
 b15zdnd11an1n04x5 FILLER_32_76 ();
 b15zdnd00an1n02x5 FILLER_32_80 ();
 b15zdnd11an1n04x5 FILLER_32_85 ();
 b15zdnd11an1n16x5 FILLER_32_94 ();
 b15zdnd00an1n01x5 FILLER_32_110 ();
 b15zdnd11an1n16x5 FILLER_32_115 ();
 b15zdnd11an1n04x5 FILLER_32_131 ();
 b15zdnd11an1n08x5 FILLER_32_144 ();
 b15zdnd11an1n04x5 FILLER_32_152 ();
 b15zdnd00an1n01x5 FILLER_32_156 ();
 b15zdnd11an1n04x5 FILLER_32_162 ();
 b15zdnd11an1n16x5 FILLER_32_170 ();
 b15zdnd11an1n04x5 FILLER_32_186 ();
 b15zdnd00an1n01x5 FILLER_32_190 ();
 b15zdnd11an1n04x5 FILLER_32_197 ();
 b15zdnd00an1n02x5 FILLER_32_204 ();
 b15zdnd11an1n16x5 FILLER_33_0 ();
 b15zdnd11an1n04x5 FILLER_33_16 ();
 b15zdnd00an1n02x5 FILLER_33_20 ();
 b15zdnd00an1n01x5 FILLER_33_22 ();
 b15zdnd11an1n04x5 FILLER_33_32 ();
 b15zdnd00an1n02x5 FILLER_33_36 ();
 b15zdnd11an1n04x5 FILLER_33_54 ();
 b15zdnd00an1n02x5 FILLER_33_58 ();
 b15zdnd00an1n01x5 FILLER_33_60 ();
 b15zdnd11an1n08x5 FILLER_33_71 ();
 b15zdnd00an1n02x5 FILLER_33_79 ();
 b15zdnd11an1n04x5 FILLER_33_85 ();
 b15zdnd11an1n08x5 FILLER_33_99 ();
 b15zdnd11an1n04x5 FILLER_33_107 ();
 b15zdnd00an1n02x5 FILLER_33_111 ();
 b15zdnd00an1n01x5 FILLER_33_113 ();
 b15zdnd11an1n04x5 FILLER_33_118 ();
 b15zdnd11an1n04x5 FILLER_33_132 ();
 b15zdnd11an1n08x5 FILLER_33_141 ();
 b15zdnd00an1n01x5 FILLER_33_149 ();
 b15zdnd11an1n08x5 FILLER_33_155 ();
 b15zdnd00an1n01x5 FILLER_33_163 ();
 b15zdnd11an1n04x5 FILLER_33_170 ();
 b15zdnd11an1n04x5 FILLER_33_179 ();
 b15zdnd00an1n02x5 FILLER_33_183 ();
 b15zdnd11an1n04x5 FILLER_33_189 ();
 b15zdnd11an1n04x5 FILLER_33_198 ();
 b15zdnd00an1n01x5 FILLER_33_202 ();
 b15zdnd11an1n04x5 FILLER_33_207 ();
 b15zdnd00an1n02x5 FILLER_33_211 ();
 b15zdnd00an1n01x5 FILLER_33_213 ();
 b15zdnd11an1n16x5 FILLER_34_8 ();
 b15zdnd11an1n04x5 FILLER_34_24 ();
 b15zdnd00an1n01x5 FILLER_34_28 ();
 b15zdnd11an1n04x5 FILLER_34_33 ();
 b15zdnd11an1n08x5 FILLER_34_41 ();
 b15zdnd11an1n04x5 FILLER_34_49 ();
 b15zdnd00an1n02x5 FILLER_34_53 ();
 b15zdnd11an1n04x5 FILLER_34_59 ();
 b15zdnd11an1n04x5 FILLER_34_67 ();
 b15zdnd11an1n16x5 FILLER_34_77 ();
 b15zdnd11an1n04x5 FILLER_34_99 ();
 b15zdnd11an1n04x5 FILLER_34_107 ();
 b15zdnd00an1n02x5 FILLER_34_111 ();
 b15zdnd00an1n01x5 FILLER_34_113 ();
 b15zdnd11an1n08x5 FILLER_34_118 ();
 b15zdnd11an1n04x5 FILLER_34_132 ();
 b15zdnd11an1n04x5 FILLER_34_140 ();
 b15zdnd11an1n04x5 FILLER_34_148 ();
 b15zdnd11an1n08x5 FILLER_34_158 ();
 b15zdnd00an1n02x5 FILLER_34_166 ();
 b15zdnd00an1n01x5 FILLER_34_168 ();
 b15zdnd11an1n08x5 FILLER_34_173 ();
 b15zdnd11an1n04x5 FILLER_34_181 ();
 b15zdnd00an1n01x5 FILLER_34_185 ();
 b15zdnd11an1n04x5 FILLER_34_196 ();
 b15zdnd00an1n02x5 FILLER_34_204 ();
 b15zdnd11an1n32x5 FILLER_35_0 ();
 b15zdnd11an1n16x5 FILLER_35_32 ();
 b15zdnd11an1n08x5 FILLER_35_48 ();
 b15zdnd11an1n04x5 FILLER_35_60 ();
 b15zdnd00an1n02x5 FILLER_35_64 ();
 b15zdnd11an1n04x5 FILLER_35_70 ();
 b15zdnd00an1n01x5 FILLER_35_74 ();
 b15zdnd11an1n04x5 FILLER_35_79 ();
 b15zdnd00an1n01x5 FILLER_35_83 ();
 b15zdnd11an1n04x5 FILLER_35_88 ();
 b15zdnd11an1n04x5 FILLER_35_96 ();
 b15zdnd00an1n01x5 FILLER_35_100 ();
 b15zdnd11an1n08x5 FILLER_35_105 ();
 b15zdnd11an1n04x5 FILLER_35_113 ();
 b15zdnd00an1n02x5 FILLER_35_117 ();
 b15zdnd11an1n04x5 FILLER_35_123 ();
 b15zdnd11an1n04x5 FILLER_35_131 ();
 b15zdnd00an1n02x5 FILLER_35_135 ();
 b15zdnd11an1n08x5 FILLER_35_141 ();
 b15zdnd00an1n02x5 FILLER_35_149 ();
 b15zdnd11an1n16x5 FILLER_35_155 ();
 b15zdnd11an1n16x5 FILLER_35_175 ();
 b15zdnd11an1n04x5 FILLER_35_191 ();
 b15zdnd00an1n01x5 FILLER_35_195 ();
 b15zdnd11an1n08x5 FILLER_35_200 ();
 b15zdnd11an1n04x5 FILLER_35_208 ();
 b15zdnd00an1n02x5 FILLER_35_212 ();
endmodule
