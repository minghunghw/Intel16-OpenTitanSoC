## ##############################################################################
## ## Intel Top Secret                                                         ##
## ##############################################################################
## ## Copyright © Intel Corporation.                                           ##
## ##                                                                          ##
## ## This is the property of Intel Corporation and may only be utilized       ##
## ## pursuant to a written Restricted Use Nondisclosure Agreement             ##
## ## with Intel Corporation.  It may not be used, reproduced, or              ##
## ## disclosed to others except in accordance with the terms and              ##
## ## conditions of such agreement.                                            ##
## ##                                                                          ##
## ## All products, processes, computer systems, dates, and figures            ##
## ## specified are preliminary based on current expectations, and are         ##
## ## subject to change without notice.                                        ##
## ##############################################################################
## ## Text_Tag % __Placeholder neutral1


VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO b15aboi22as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aboi22as1n02x3 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.3155 0.682 0.3595 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.3155 0.898 0.3595 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.702 0.202 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.4275 0.574 0.4715 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.373 0.142 0.417 ;
        RECT 0.722 0.4275 0.79 0.4715 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.398 0.202 0.466 0.246 ;
        RECT 0.83 0.048 0.898 0.092 ;
    END
  END vssx
END b15aboi22as1n02x3

MACRO b15aboi22as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aboi22as1n02x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 0.682 0.472 ;
        RECT 0.614 0.068 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.202 0.682 0.246 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.382 0.142 0.426 ;
        RECT 0.83 0.538 0.898 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.398 0.202 0.466 0.246 ;
        RECT 0.938 0.048 1.006 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.518 0.466 0.562 ;
    LAYER m1 ;
      RECT 0.29 0.518 0.722 0.562 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.428 1.026 0.472 ;
  END
END b15aboi22as1n02x5

MACRO b15aboi22as1n04x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aboi22as1n04x3 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.594 0.292 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.918 0.112 ;
        RECT 0.29 0.158 0.79 0.202 ;
        RECT 0.722 0.068 0.79 0.202 ;
        RECT 0.29 0.518 0.574 0.562 ;
        RECT 0.506 0.428 0.574 0.562 ;
        RECT 0.29 0.158 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.508 0.448 0.572 0.492 ;
        RECT 0.83 0.068 0.898 0.112 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.722 0.448 0.79 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
    LAYER v0 ;
      RECT 0.182 0.1575 0.25 0.2015 ;
      RECT 0.182 0.338 0.25 0.382 ;
  END
END b15aboi22as1n04x3

MACRO b15aboi22as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aboi22as1n04x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.574 0.382 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 0.682 0.472 ;
        RECT 0.614 0.068 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.2065 0.682 0.2505 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.398 0.203 0.466 0.247 ;
        RECT 0.938 0.048 1.006 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.518 0.722 0.562 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.428 1.026 0.472 ;
  END
END b15aboi22as1n04x5

MACRO b15aboi22as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aboi22as1n06x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.79 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.546 0.382 ;
        RECT 1.478 0.158 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.438 0.292 ;
        RECT 1.046 0.158 1.114 0.292 ;
      LAYER v0 ;
        RECT 1.262 0.248 1.33 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 1.566 0.112 ;
        RECT 1.154 0.158 1.438 0.202 ;
        RECT 1.37 0.068 1.438 0.202 ;
        RECT 1.154 0.068 1.222 0.202 ;
        RECT 0.938 0.068 1.222 0.112 ;
        RECT 0.398 0.428 1.006 0.472 ;
        RECT 0.938 0.068 1.006 0.472 ;
        RECT 0.398 0.158 1.006 0.202 ;
        RECT 0.398 0.068 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.4 0.088 0.464 0.132 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.068 1.114 0.112 ;
        RECT 1.478 0.068 1.546 0.112 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.493 0.142 0.537 ;
        RECT 1.154 0.538 1.222 0.582 ;
        RECT 1.37 0.538 1.438 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.518 1.046 0.562 ;
    LAYER v0 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.338 0.466 0.382 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.182 0.164 0.25 0.208 ;
      RECT 0.182 0.493 0.25 0.537 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.898 0.382 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.114 0.428 1.566 0.472 ;
  END
END b15aboi22as1n06x5

MACRO b15aboi22as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aboi22as1n08x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.79 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.546 0.382 ;
        RECT 1.478 0.158 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.438 0.292 ;
        RECT 1.046 0.158 1.114 0.292 ;
      LAYER v0 ;
        RECT 1.262 0.248 1.33 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 1.566 0.112 ;
        RECT 1.154 0.158 1.438 0.202 ;
        RECT 1.37 0.068 1.438 0.202 ;
        RECT 1.154 0.068 1.222 0.202 ;
        RECT 0.938 0.068 1.222 0.112 ;
        RECT 0.398 0.428 1.006 0.472 ;
        RECT 0.938 0.068 1.006 0.472 ;
        RECT 0.398 0.158 1.006 0.202 ;
        RECT 0.398 0.068 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.4 0.088 0.464 0.132 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.068 1.114 0.112 ;
        RECT 1.478 0.068 1.546 0.112 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.493 0.142 0.537 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.518 1.046 0.562 ;
    LAYER v0 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.338 0.466 0.382 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.182 0.164 0.25 0.208 ;
      RECT 0.182 0.493 0.25 0.537 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.898 0.382 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.114 0.428 1.566 0.472 ;
  END
END b15aboi22as1n08x5

MACRO b15aboi22as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aboi22as1n12x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.70571425 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.70571425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 1.222 0.292 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.338 2.086 0.382 ;
        RECT 2.018 0.158 2.086 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.338 1.654 0.382 ;
        RECT 1.91 0.338 1.978 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.248 1.978 0.292 ;
        RECT 1.37 0.248 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.478 0.248 1.546 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 2.106 0.112 ;
        RECT 0.506 0.158 1.978 0.202 ;
        RECT 1.91 0.068 1.978 0.202 ;
        RECT 0.486 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.472 ;
        RECT 0.506 0.068 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.508 0.088 0.572 0.132 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.018 0.068 2.086 0.112 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.518 1.37 0.562 ;
    LAYER v0 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.182 0.1595 0.25 0.2035 ;
      RECT 0.182 0.454 0.25 0.498 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 1.114 0.382 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.438 0.428 2.106 0.472 ;
  END
END b15aboi22as1n12x5

MACRO b15aboi22as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aboi22as1n16x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 1.438 0.382 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.338 2.518 0.382 ;
        RECT 2.45 0.158 2.518 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.338 1.762 0.382 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.342 0.338 2.41 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.248 2.41 0.292 ;
        RECT 1.586 0.158 1.654 0.292 ;
      LAYER v0 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.234 0.248 2.302 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11016 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.538 0.112 ;
        RECT 1.694 0.158 2.41 0.202 ;
        RECT 2.342 0.068 2.41 0.202 ;
        RECT 1.694 0.068 1.762 0.202 ;
        RECT 1.478 0.068 1.762 0.112 ;
        RECT 0.506 0.428 1.546 0.472 ;
        RECT 1.478 0.068 1.546 0.472 ;
        RECT 0.614 0.158 1.546 0.202 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.586 0.068 1.654 0.112 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.45 0.068 2.518 0.112 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.518 1.586 0.562 ;
    LAYER v0 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.454 0.25 0.498 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.25 0.338 0.29 0.382 ;
      RECT 0.074 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.382 ;
      RECT 0.358 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.292 ;
      RECT 0.574 0.248 1.33 0.292 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.654 0.428 2.538 0.472 ;
  END
END b15aboi22as1n16x5

MACRO b15aboi22as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aboi22as1n24x5 0 0 ;
  SIZE 3.564 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 1.978 0.382 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.338 3.49 0.382 ;
        RECT 3.422 0.158 3.49 0.382 ;
      LAYER v0 ;
        RECT 2.234 0.338 2.302 0.382 ;
        RECT 2.558 0.338 2.626 0.382 ;
        RECT 2.99 0.338 3.058 0.382 ;
        RECT 3.314 0.338 3.382 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.248 3.382 0.292 ;
        RECT 2.126 0.158 2.194 0.292 ;
      LAYER v0 ;
        RECT 2.342 0.248 2.41 0.292 ;
        RECT 2.774 0.248 2.842 0.292 ;
        RECT 3.206 0.248 3.274 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.15912 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.068 3.51 0.112 ;
        RECT 2.234 0.158 3.382 0.202 ;
        RECT 3.314 0.068 3.382 0.202 ;
        RECT 2.234 0.068 2.302 0.202 ;
        RECT 2.018 0.068 2.302 0.112 ;
        RECT 0.614 0.428 2.086 0.472 ;
        RECT 2.018 0.068 2.086 0.472 ;
        RECT 0.722 0.158 2.086 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 2.126 0.068 2.194 0.112 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.422 0.068 3.49 0.112 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.316 0.538 3.38 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.598 0.022 ;
        RECT 3.206 -0.022 3.274 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 3.208 0.048 3.272 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.518 2.126 0.562 ;
    LAYER v0 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.454 0.466 0.498 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.454 0.25 0.498 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.25 0.338 0.29 0.382 ;
      RECT 0.074 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.382 ;
      RECT 0.358 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.358 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.248 1.87 0.292 ;
      RECT 2.126 0.428 2.194 0.562 ;
      RECT 2.194 0.428 3.51 0.472 ;
  END
END b15aboi22as1n24x5

MACRO b15and002as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and002as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.383 0.466 0.427 ;
        RECT 0.398 0.178 0.466 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.473 0.358 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.383 0.25 0.427 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.472 ;
  END
END b15and002as1n02x5

MACRO b15and002as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and002as1n03x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.383 0.466 0.427 ;
        RECT 0.398 0.178 0.466 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.473 0.358 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.383 0.25 0.427 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.472 ;
  END
END b15and002as1n03x5

MACRO b15and002as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and002as1n04x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.2705 0.358 0.3145 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.372 0.466 0.416 ;
        RECT 0.398 0.178 0.466 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.4645 0.358 0.5085 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.372 0.25 0.416 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.472 ;
  END
END b15and002as1n04x5

MACRO b15and002as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and002as1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.378 0.292 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 1.4114285 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.408 0.682 0.452 ;
        RECT 0.614 0.1415 0.682 0.1855 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4785 0.25 0.5225 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.722 0.489 0.79 0.533 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.292 0.088 0.356 0.132 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.378 0.428 0.506 0.472 ;
      RECT 0.358 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.472 ;
  END
END b15and002as1n08x5

MACRO b15and002as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and002as1n12x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.396923 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.472 ;
        RECT 0.722 0.248 1.006 0.292 ;
        RECT 0.722 0.068 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.363 0.79 0.407 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.363 1.006 0.407 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.83 0.448 0.898 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.1135 0.25 0.1575 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.29 0.363 0.358 0.407 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.358 0.068 0.506 0.112 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.574 0.338 0.614 0.382 ;
      RECT 0.574 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.382 ;
  END
END b15and002as1n12x5

MACRO b15and002as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and002as1n16x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.562 ;
        RECT 0.938 0.338 1.222 0.382 ;
        RECT 0.938 0.158 1.006 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.4455 1.006 0.4895 ;
        RECT 0.938 0.1835 1.006 0.2275 ;
        RECT 1.154 0.4455 1.222 0.4895 ;
        RECT 1.154 0.1835 1.222 0.2275 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.093 0.574 0.137 ;
        RECT 0.83 0.093 0.898 0.137 ;
        RECT 1.046 0.093 1.114 0.137 ;
        RECT 1.262 0.093 1.33 0.137 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
    LAYER v0 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.614 0.1835 0.682 0.2275 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.1835 0.466 0.2275 ;
      RECT 0.29 0.1835 0.358 0.2275 ;
      RECT 0.182 0.068 0.25 0.112 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.1835 0.142 0.2275 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.358 0.428 0.83 0.472 ;
      RECT 0.83 0.248 0.898 0.472 ;
  END
END b15and002as1n16x5

MACRO b15and002as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and002as1n24x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5875925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.42734 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.898 0.382 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.654 0.382 ;
        RECT 1.586 0.158 1.654 0.382 ;
        RECT 0.938 0.158 1.654 0.202 ;
        RECT 1.478 0.338 1.546 0.562 ;
        RECT 1.262 0.338 1.33 0.562 ;
        RECT 1.046 0.338 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
    LAYER v0 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.228 0.248 0.272 ;
      RECT 0.076 0.1425 0.14 0.1865 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.158 0.79 0.202 ;
      RECT 0.142 0.068 0.466 0.112 ;
      RECT 0.142 0.428 0.938 0.472 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.006 0.248 1.546 0.292 ;
  END
END b15and002as1n24x5

MACRO b15and002as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and002as1n32x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63973075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.682 0.382 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.81 0.338 1.222 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.428 2.194 0.472 ;
        RECT 2.126 0.158 2.194 0.472 ;
        RECT 1.262 0.158 2.194 0.202 ;
        RECT 1.37 0.338 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.372 0.358 1.436 0.402 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
    LAYER v0 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 1.048 0.228 1.112 0.272 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.228 0.248 0.272 ;
      RECT 0.076 0.138 0.14 0.182 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 0.142 0.068 0.682 0.112 ;
      RECT 0.142 0.428 1.262 0.472 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.33 0.248 2.086 0.292 ;
  END
END b15and002as1n32x5

MACRO b15and003as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and003as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.113 0.358 0.157 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.506 0.203 0.574 0.247 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.398 -0.022 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END vssx
END b15and003as1n02x5

MACRO b15and003as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and003as1n03x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.506 0.158 0.574 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.398 0.048 0.466 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.448 0.142 0.492 ;
  END
END b15and003as1n03x5

MACRO b15and003as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and003as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.158 0.142 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.068 0.25 0.112 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.338 0.25 0.382 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.25 0.428 0.506 0.472 ;
      RECT 0.506 0.068 0.574 0.472 ;
      RECT 0.574 0.428 0.702 0.472 ;
      RECT 0.574 0.068 0.702 0.112 ;
  END
END b15and003as1n04x5

MACRO b15and003as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and003as1n08x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.23925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.23925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.23925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.466 0.358 0.51 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.938 0.518 1.006 0.562 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.938 0.068 1.006 0.112 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.473 0.142 0.517 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.398 0.518 0.614 0.562 ;
      RECT 0.142 0.068 0.614 0.112 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.428 0.722 0.472 ;
      RECT 0.682 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.472 ;
  END
END b15and003as1n08x5

MACRO b15and003as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and003as1n12x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.43712425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0171 LAYER m1 ;
      ANTENNAMAXAREACAR 0.50222225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 1.438 0.562 ;
        RECT 1.154 0.248 1.438 0.292 ;
        RECT 1.154 0.068 1.222 0.562 ;
      LAYER v0 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.262 0.518 1.33 0.562 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.722 -0.022 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.046 0.068 1.114 0.112 ;
        RECT 1.262 0.068 1.33 0.112 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.182 0.472 ;
    LAYER v0 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.506 0.112 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.428 1.046 0.472 ;
      RECT 1.046 0.248 1.114 0.472 ;
  END
END b15and003as1n12x5

MACRO b15and003as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and003as1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.9025 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.81 0.292 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.382 ;
        RECT 0.918 0.248 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.562 ;
        RECT 1.262 0.248 1.546 0.292 ;
        RECT 1.262 0.068 1.33 0.562 ;
      LAYER v0 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.37 0.518 1.438 0.562 ;
        RECT 1.586 0.518 1.654 0.562 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
      LAYER v0 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.37 0.068 1.438 0.112 ;
        RECT 1.586 0.068 1.654 0.112 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.898 0.112 ;
      RECT 0.506 0.158 1.222 0.202 ;
    LAYER v0 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.068 0.25 0.112 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.428 0.398 0.472 ;
      RECT 0.054 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.518 0.722 0.562 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.428 1.154 0.472 ;
      RECT 1.154 0.248 1.222 0.472 ;
  END
END b15and003as1n16x5

MACRO b15and003as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15and003as1n24x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.43757575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.35267975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.28915825 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 1.222 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.472 ;
        RECT 1.262 0.158 1.978 0.202 ;
        RECT 1.37 0.338 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.372 0.358 1.436 0.402 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
      LAYER v0 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.898 0.112 ;
      RECT 0.054 0.428 0.398 0.472 ;
    LAYER v0 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 1.048 0.178 1.112 0.222 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.832 0.178 0.896 0.222 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.068 0.25 0.112 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.158 0.898 0.292 ;
      RECT 0.898 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 0.054 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.428 1.262 0.472 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.33 0.248 1.87 0.292 ;
  END
END b15and003as1n24x5

MACRO b15andc04as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15andc04as1n02x3 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.3155 1.006 0.3595 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.3155 0.79 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 0.682 0.472 ;
        RECT 0.614 0.068 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.83 0.068 0.898 0.562 ;
    LAYER v0 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.068 0.378 0.112 ;
      RECT 0.898 0.068 1.026 0.112 ;
  END
END b15andc04as1n02x3

MACRO b15andc04as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15andc04as1n02x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.3155 1.006 0.3595 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.3155 0.79 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 0.682 0.472 ;
        RECT 0.614 0.068 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.83 0.068 0.898 0.562 ;
    LAYER v0 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.83 0.4575 0.898 0.5015 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.4575 0.25 0.5015 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.068 0.378 0.112 ;
      RECT 0.898 0.068 1.026 0.112 ;
  END
END b15andc04as1n02x5

MACRO b15andc04as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15andc04as1n03x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.3155 1.006 0.3595 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.3155 0.79 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 0.682 0.472 ;
        RECT 0.614 0.068 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.83 0.068 0.898 0.562 ;
    LAYER v0 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.83 0.4575 0.898 0.5015 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.4575 0.25 0.5015 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.068 0.378 0.112 ;
      RECT 0.898 0.068 1.026 0.112 ;
  END
END b15andc04as1n03x5

MACRO b15andc04as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15andc04as1n04x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.472 ;
        RECT 0.074 0.068 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.068 0.25 0.112 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.682 0.562 ;
        RECT 0.506 0.338 0.682 0.382 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.163 0.574 0.207 ;
        RECT 0.614 0.428 0.682 0.472 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.383 0.142 0.427 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 1.046 0.538 1.114 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.163 0.682 0.207 ;
        RECT 1.046 0.048 1.114 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.382 ;
    LAYER v0 ;
      RECT 0.938 0.448 1.006 0.492 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.182 0.383 0.25 0.427 ;
      RECT 0.076 0.178 0.14 0.222 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.292 ;
      RECT 0.142 0.248 0.182 0.292 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.562 ;
  END
END b15andc04as1n04x5

MACRO b15andc04as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15andc04as1n06x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.158 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.428 0.898 0.472 ;
        RECT 0.83 0.068 0.898 0.472 ;
        RECT 0.614 0.248 0.898 0.292 ;
        RECT 0.722 0.428 0.79 0.562 ;
        RECT 0.614 0.068 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 0.724 0.498 0.788 0.542 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.398 0.4505 0.466 0.4945 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.154 0.538 1.222 0.582 ;
        RECT 1.37 0.538 1.438 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.37 0.048 1.438 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.134 0.068 1.262 0.112 ;
    LAYER v0 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.4505 0.25 0.4945 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.466 0.338 0.79 0.382 ;
      RECT 1.262 0.068 1.33 0.562 ;
  END
END b15andc04as1n06x5

MACRO b15andc04as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15andc04as1n08x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.378 0.112 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.574 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.068 2.086 0.292 ;
        RECT 1.89 0.068 2.086 0.112 ;
      LAYER v0 ;
        RECT 1.91 0.068 1.978 0.112 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.338 2.194 0.382 ;
        RECT 2.126 0.158 2.194 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.338 1.87 0.382 ;
        RECT 2.018 0.338 2.086 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 1.438 0.292 ;
        RECT 1.37 0.158 1.438 0.292 ;
        RECT 1.046 0.158 1.114 0.292 ;
        RECT 0.938 0.248 1.006 0.472 ;
        RECT 0.83 0.158 0.898 0.292 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 0.832 0.178 0.896 0.222 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.048 0.178 1.112 0.222 ;
        RECT 1.372 0.178 1.436 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.694 0.538 1.762 0.582 ;
        RECT 1.91 0.538 1.978 0.582 ;
        RECT 2.126 0.538 2.194 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 1.478 0.048 1.546 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 2.126 0.048 2.194 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.518 1.154 0.562 ;
      RECT 1.586 0.158 1.654 0.472 ;
    LAYER v0 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.912 0.228 1.976 0.272 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.37 0.4575 1.438 0.5015 ;
      RECT 1.156 0.408 1.22 0.452 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.292 0.228 0.356 0.272 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.292 ;
      RECT 0.074 0.428 0.614 0.472 ;
      RECT 0.358 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.654 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.292 ;
      RECT 1.654 0.428 2.194 0.472 ;
  END
END b15andc04as1n08x5

MACRO b15andc04as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15andc04as1n12x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.248 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.293 2.194 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.248 2.626 0.562 ;
      LAYER v0 ;
        RECT 2.558 0.293 2.626 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07956 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.78666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 1.87 0.292 ;
        RECT 1.802 0.158 1.87 0.292 ;
        RECT 1.586 0.158 1.654 0.292 ;
        RECT 1.262 0.158 1.33 0.292 ;
        RECT 1.154 0.248 1.222 0.472 ;
        RECT 1.046 0.158 1.114 0.292 ;
        RECT 0.938 0.248 1.006 0.472 ;
        RECT 0.83 0.158 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.832 0.178 0.896 0.222 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.048 0.178 1.112 0.222 ;
        RECT 1.154 0.408 1.222 0.452 ;
        RECT 1.264 0.178 1.328 0.222 ;
        RECT 1.588 0.178 1.652 0.222 ;
        RECT 1.804 0.178 1.868 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.45 0.428 2.518 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.478 0.048 1.546 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 2.45 0.048 2.518 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.682 0.202 ;
      RECT 0.722 0.518 1.37 0.562 ;
      RECT 1.91 0.068 1.978 0.382 ;
      RECT 2.018 0.158 2.646 0.202 ;
    LAYER v0 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.4575 1.87 0.5015 ;
      RECT 1.586 0.4575 1.654 0.5015 ;
      RECT 1.372 0.408 1.436 0.452 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.378 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.978 0.068 2.322 0.112 ;
  END
END b15andc04as1n12x5

MACRO b15andc04as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15andc04as1n16x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.248 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.293 2.842 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.248 3.274 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.293 3.274 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11016 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 2.194 0.292 ;
        RECT 2.126 0.158 2.194 0.292 ;
        RECT 1.91 0.158 1.978 0.292 ;
        RECT 1.586 0.158 1.654 0.292 ;
        RECT 1.478 0.248 1.546 0.472 ;
        RECT 1.37 0.158 1.438 0.292 ;
        RECT 1.262 0.248 1.33 0.472 ;
        RECT 1.154 0.158 1.222 0.292 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.408 1.114 0.452 ;
        RECT 1.156 0.178 1.22 0.222 ;
        RECT 1.262 0.408 1.33 0.452 ;
        RECT 1.372 0.178 1.436 0.222 ;
        RECT 1.478 0.408 1.546 0.452 ;
        RECT 1.588 0.178 1.652 0.222 ;
        RECT 1.912 0.178 1.976 0.222 ;
        RECT 2.128 0.178 2.192 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 3.206 -0.022 3.274 0.112 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 1.478 0.048 1.546 0.092 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.99 0.048 3.058 0.092 ;
        RECT 3.206 0.048 3.274 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.702 0.202 ;
      RECT 0.83 0.518 1.694 0.562 ;
      RECT 2.45 0.068 2.518 0.472 ;
      RECT 2.558 0.158 3.274 0.202 ;
    LAYER v0 ;
      RECT 3.098 0.158 3.166 0.202 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.774 0.068 2.842 0.112 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.45 0.293 2.518 0.337 ;
      RECT 2.342 0.4575 2.41 0.5015 ;
      RECT 2.126 0.4575 2.194 0.5015 ;
      RECT 1.91 0.4575 1.978 0.5015 ;
      RECT 1.696 0.408 1.76 0.452 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.486 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.762 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.978 0.338 2.126 0.382 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.194 0.338 2.342 0.382 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.518 0.068 2.862 0.112 ;
  END
END b15andc04as1n16x5

MACRO b15ao0012as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0012as1n02x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.292 ;
        RECT 0.27 0.068 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0018 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.3835 0.574 0.4275 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.385 0.142 0.429 ;
        RECT 0.29 0.383 0.358 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.2025 0.142 0.2465 ;
        RECT 0.614 0.1155 0.682 0.1595 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.472 ;
    LAYER v0 ;
      RECT 0.722 0.203 0.79 0.247 ;
      RECT 0.722 0.383 0.79 0.427 ;
  END
END b15ao0012as1n02x5

MACRO b15ao0012as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0012as1n03x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 2.014 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.292 ;
        RECT 0.27 0.068 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0027 LAYER m1 ;
      ANTENNAMAXAREACAR 3.67333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.3835 0.574 0.4275 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.385 0.142 0.429 ;
        RECT 0.29 0.42 0.358 0.464 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.2025 0.142 0.2465 ;
        RECT 0.614 0.1155 0.682 0.1595 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.472 ;
    LAYER v0 ;
      RECT 0.722 0.203 0.79 0.247 ;
      RECT 0.722 0.383 0.79 0.427 ;
  END
END b15ao0012as1n03x5

MACRO b15ao0012as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0012as1n04x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.522639 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.03018525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.228 0.682 0.272 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.4005 0.79 0.4445 ;
        RECT 0.722 0.1405 0.79 0.1845 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.83 0.4005 0.898 0.4445 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.506 0.135 0.574 0.179 ;
        RECT 0.83 0.1405 0.898 0.1845 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.382 ;
    LAYER v0 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.398 0.135 0.466 0.179 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.076 0.498 0.14 0.542 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.574 0.472 ;
      RECT 0.398 0.518 0.614 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
  END
END b15ao0012as1n04x5

MACRO b15ao0012as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0012as1n06x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.574 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.4645 0.898 0.5085 ;
        RECT 0.83 0.101 0.898 0.145 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.722 0.4645 0.79 0.5085 ;
        RECT 0.938 0.4645 1.006 0.5085 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.722 0.101 0.79 0.145 ;
        RECT 0.938 0.101 1.006 0.145 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.202 ;
    LAYER v0 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.4 0.088 0.464 0.132 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.518 0.574 0.562 ;
      RECT 0.398 0.428 0.614 0.472 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
  END
END b15ao0012as1n06x5

MACRO b15ao0012as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0012as1n08x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.25076925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.25076925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.498 0.466 0.542 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.046 0.138 1.114 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.506 0.3675 0.574 0.4115 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.154 0.448 1.222 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
    LAYER v0 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.29 0.4055 0.358 0.4495 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.4055 0.25 0.4495 ;
    LAYER m1 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.358 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.562 ;
  END
END b15ao0012as1n08x5

MACRO b15ao0012as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0012as1n12x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.199375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.59916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.498 1.114 0.542 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.318 0.682 0.362 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4128395 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.574 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.472 ;
        RECT 1.262 0.248 1.546 0.292 ;
        RECT 1.262 0.068 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.408 1.33 0.452 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.478 0.408 1.546 0.452 ;
        RECT 1.478 0.138 1.546 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.154 0.408 1.222 0.452 ;
        RECT 1.37 0.408 1.438 0.452 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.37 0.138 1.438 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.074 0.428 1.006 0.472 ;
    LAYER v0 ;
      RECT 0.938 0.138 1.006 0.182 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.398 0.228 0.466 0.272 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.138 0.142 0.182 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.142 0.248 0.29 0.292 ;
      RECT 0.29 0.068 0.358 0.292 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
  END
END b15ao0012as1n12x5

MACRO b15ao0012as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0012as1n16x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.114 0.382 ;
        RECT 1.046 0.158 1.114 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.594 0.338 0.79 0.382 ;
        RECT 0.722 0.068 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4611965 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.068 1.654 0.562 ;
        RECT 1.37 0.338 1.654 0.382 ;
        RECT 1.37 0.068 1.438 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.474 1.438 0.518 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.474 1.654 0.518 ;
        RECT 1.586 0.138 1.654 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 1.262 0.474 1.33 0.518 ;
        RECT 1.478 0.474 1.546 0.518 ;
        RECT 1.694 0.474 1.762 0.518 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.83 0.1805 0.898 0.2245 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.694 0.138 1.762 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 0.054 0.428 1.026 0.472 ;
    LAYER v0 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.1805 1.006 0.2245 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.81 0.518 1.154 0.562 ;
      RECT 1.006 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.562 ;
  END
END b15ao0012as1n16x5

MACRO b15ao0012as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0012as1n24x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.97375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.29833325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.338 1.87 0.562 ;
      LAYER v0 ;
        RECT 1.802 0.443 1.87 0.487 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.222 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.574 0.382 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.158 2.518 0.472 ;
        RECT 2.018 0.338 2.518 0.382 ;
        RECT 2.234 0.158 2.302 0.472 ;
        RECT 2.018 0.158 2.086 0.472 ;
      LAYER v0 ;
        RECT 2.02 0.408 2.084 0.452 ;
        RECT 2.018 0.194 2.086 0.238 ;
        RECT 2.236 0.408 2.3 0.452 ;
        RECT 2.234 0.194 2.302 0.238 ;
        RECT 2.452 0.408 2.516 0.452 ;
        RECT 2.45 0.194 2.518 0.238 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.126 0.538 2.194 0.582 ;
        RECT 2.342 0.538 2.41 0.582 ;
        RECT 2.558 0.538 2.626 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 1.91 0.113 1.978 0.157 ;
        RECT 2.126 0.113 2.194 0.157 ;
        RECT 2.342 0.113 2.41 0.157 ;
        RECT 2.558 0.113 2.626 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.068 1.262 0.112 ;
      RECT 0.182 0.428 1.762 0.472 ;
    LAYER v0 ;
      RECT 1.694 0.138 1.762 0.182 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.138 1.33 0.182 ;
      RECT 1.048 0.178 1.112 0.222 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.832 0.178 0.896 0.222 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.158 0.898 0.292 ;
      RECT 0.898 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 1.262 0.068 1.33 0.292 ;
      RECT 1.33 0.248 1.694 0.292 ;
      RECT 1.694 0.068 1.762 0.292 ;
  END
END b15ao0012as1n24x5

MACRO b15ao0012as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0012as1n32x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.83916675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 1.220606 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.338 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.498 2.518 0.542 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57879625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57879625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 1.654 0.382 ;
        RECT 1.586 0.158 1.654 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.478 0.338 1.546 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57879625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57879625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.79 0.382 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11016 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.158 3.382 0.472 ;
        RECT 2.666 0.338 3.382 0.382 ;
        RECT 3.098 0.158 3.166 0.472 ;
        RECT 2.882 0.158 2.95 0.472 ;
        RECT 2.666 0.158 2.734 0.472 ;
      LAYER v0 ;
        RECT 2.668 0.408 2.732 0.452 ;
        RECT 2.666 0.194 2.734 0.238 ;
        RECT 2.884 0.408 2.948 0.452 ;
        RECT 2.882 0.194 2.95 0.238 ;
        RECT 3.1 0.408 3.164 0.452 ;
        RECT 3.098 0.194 3.166 0.238 ;
        RECT 3.316 0.408 3.38 0.452 ;
        RECT 3.314 0.194 3.382 0.238 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 2.558 0.498 2.626 0.542 ;
        RECT 2.774 0.4985 2.842 0.5425 ;
        RECT 2.99 0.4985 3.058 0.5425 ;
        RECT 3.206 0.493 3.274 0.537 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.99 -0.022 3.058 0.292 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.234 -0.022 2.302 0.292 ;
        RECT 2.018 -0.022 2.086 0.292 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.558 0.113 2.626 0.157 ;
        RECT 2.774 0.194 2.842 0.238 ;
        RECT 2.99 0.194 3.058 0.238 ;
        RECT 3.206 0.113 3.274 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.83 0.068 1.694 0.112 ;
      RECT 0.182 0.428 2.41 0.472 ;
    LAYER v0 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.48 0.178 1.544 0.222 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.264 0.178 1.328 0.222 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.048 0.178 1.112 0.222 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.832 0.178 0.896 0.222 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.158 0.898 0.292 ;
      RECT 0.898 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 1.114 0.248 1.262 0.292 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.33 0.248 1.478 0.292 ;
      RECT 1.478 0.158 1.546 0.292 ;
      RECT 1.694 0.068 1.762 0.382 ;
      RECT 1.762 0.338 2.342 0.382 ;
      RECT 2.342 0.068 2.41 0.382 ;
  END
END b15ao0012as1n32x5

MACRO b15ao0022as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0022as1n02x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
    LAYER v0 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.29 0.178 0.358 0.222 ;
      RECT 0.29 0.408 0.358 0.452 ;
      RECT 0.182 0.408 0.25 0.452 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.29 0.562 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.25 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.562 ;
  END
END b15ao0022as1n02x5

MACRO b15ao0022as1n03x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0022as1n03x3 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.113 0.466 0.157 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 0.83 0.181 0.898 0.225 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
        RECT 0.506 0.113 0.574 0.157 ;
        RECT 0.722 0.181 0.79 0.225 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.203 0.358 0.247 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
  END
END b15ao0022as1n03x3

MACRO b15ao0022as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0022as1n03x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.408 0.142 0.452 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.83 0.048 0.898 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.562 ;
    LAYER v0 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.4005 0.79 0.4445 ;
      RECT 0.614 0.1855 0.682 0.2295 ;
      RECT 0.614 0.4005 0.682 0.4445 ;
      RECT 0.29 0.383 0.358 0.427 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.358 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.682 0.518 0.918 0.562 ;
  END
END b15ao0022as1n03x5

MACRO b15ao0022as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0022as1n04x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.4555 0.898 0.4995 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
    LAYER v0 ;
      RECT 0.614 0.4505 0.682 0.4945 ;
      RECT 0.29 0.1805 0.358 0.2245 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.182 0.383 0.25 0.427 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.29 0.562 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.25 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.562 ;
  END
END b15ao0022as1n04x5

MACRO b15ao0022as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0022as1n06x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 1.006 0.292 ;
        RECT 0.722 0.158 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.466 1.114 0.51 ;
        RECT 1.046 0.138 1.114 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
      LAYER v0 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.938 0.466 1.006 0.51 ;
        RECT 1.154 0.466 1.222 0.51 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.428 0.398 0.472 ;
    LAYER v0 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.398 0.1525 0.466 0.1965 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.506 0.562 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.428 0.898 0.472 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 0.466 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.382 ;
      RECT 0.682 0.338 1.006 0.382 ;
  END
END b15ao0022as1n06x5

MACRO b15ao0022as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0022as1n08x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.562 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.338 1.654 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4055 0.25 0.4495 ;
        RECT 0.398 0.4055 0.466 0.4495 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.586 0.428 1.654 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.18 0.25 0.224 ;
        RECT 0.83 0.18 0.898 0.224 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.158 1.654 0.202 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.154 0.4055 1.222 0.4495 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.4055 1.006 0.4495 ;
      RECT 0.722 0.4055 0.79 0.4495 ;
      RECT 0.398 0.18 0.466 0.224 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.79 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.006 0.518 1.154 0.562 ;
      RECT 0.938 0.158 1.154 0.202 ;
      RECT 1.154 0.158 1.222 0.562 ;
  END
END b15ao0022as1n08x5

MACRO b15ao0022as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0022as1n12x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.574 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 1.114 0.292 ;
        RECT 1.046 0.158 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.222 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.068 1.654 0.562 ;
        RECT 1.37 0.338 1.654 0.382 ;
        RECT 1.37 0.068 1.438 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.454 1.438 0.498 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.454 1.654 0.498 ;
        RECT 1.586 0.138 1.654 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
      LAYER v0 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.202 ;
    LAYER v0 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.292 0.088 0.356 0.132 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.722 0.562 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.428 1.33 0.472 ;
      RECT 0.074 0.428 0.614 0.472 ;
      RECT 0.358 0.158 0.614 0.202 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 0.682 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.202 ;
      RECT 1.222 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.382 ;
  END
END b15ao0022as1n12x5

MACRO b15ao0022as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0022as1n16x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.79 0.292 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.574 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.438 0.292 ;
        RECT 0.938 0.158 1.006 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.262 0.248 1.33 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.338 1.762 0.472 ;
        RECT 1.046 0.338 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.478 0.338 1.546 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.338 2.194 0.382 ;
        RECT 2.126 0.158 2.194 0.382 ;
        RECT 1.694 0.158 2.194 0.202 ;
        RECT 2.018 0.338 2.086 0.562 ;
        RECT 1.802 0.338 1.87 0.562 ;
      LAYER v0 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.018 0.158 2.086 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
      LAYER v0 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.586 0.112 1.654 0.156 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.202 ;
    LAYER v0 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.292 0.088 0.356 0.132 ;
      RECT 0.182 0.518 0.25 0.562 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.518 0.722 0.562 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.428 1.654 0.472 ;
      RECT 0.054 0.428 0.614 0.472 ;
      RECT 0.358 0.158 0.614 0.202 ;
      RECT 0.614 0.338 0.682 0.472 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.682 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.114 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.292 ;
      RECT 1.546 0.248 2.086 0.292 ;
  END
END b15ao0022as1n16x5

MACRO b15ao0022as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0022as1n24x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.338 2.322 0.382 ;
        RECT 1.91 0.248 1.978 0.382 ;
      LAYER v0 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.234 0.338 2.302 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.248 2.95 0.472 ;
        RECT 2.558 0.248 2.95 0.292 ;
      LAYER v0 ;
        RECT 2.666 0.248 2.734 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.674 0.382 ;
        RECT 0.83 0.338 0.898 0.562 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.87 0.382 ;
        RECT 0.938 0.248 1.87 0.292 ;
        RECT 0.938 0.158 1.006 0.292 ;
      LAYER v0 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.694 0.248 1.762 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.79 0.202 ;
        RECT 0.614 0.338 0.682 0.562 ;
        RECT 0.074 0.338 0.682 0.382 ;
        RECT 0.398 0.338 0.466 0.562 ;
        RECT 0.29 0.158 0.358 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.938 0.428 1.91 0.472 ;
      RECT 1.998 0.068 2.342 0.112 ;
    LAYER v0 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.882 0.518 2.95 0.562 ;
      RECT 2.776 0.358 2.84 0.402 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.45 0.518 2.518 0.562 ;
      RECT 2.342 0.248 2.41 0.292 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
    LAYER m1 ;
      RECT 0.486 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.114 0.158 2.234 0.202 ;
      RECT 2.234 0.158 2.302 0.292 ;
      RECT 2.106 0.428 2.45 0.472 ;
      RECT 2.302 0.248 2.45 0.292 ;
      RECT 2.45 0.248 2.518 0.472 ;
      RECT 2.518 0.428 2.774 0.472 ;
      RECT 2.774 0.338 2.842 0.472 ;
      RECT 1.91 0.428 1.978 0.562 ;
      RECT 1.978 0.518 2.97 0.562 ;
      RECT 2.342 0.068 2.41 0.202 ;
      RECT 2.41 0.158 2.97 0.202 ;
  END
END b15ao0022as1n24x5

MACRO b15ao0022as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ao0022as1n32x5 0 0 ;
  SIZE 4.104 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.338 3.186 0.382 ;
        RECT 2.558 0.248 2.626 0.382 ;
      LAYER v0 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 2.882 0.338 2.95 0.382 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.248 4.03 0.472 ;
        RECT 3.51 0.248 4.03 0.292 ;
      LAYER v0 ;
        RECT 3.53 0.248 3.598 0.292 ;
        RECT 3.746 0.248 3.814 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 2.322 0.382 ;
        RECT 1.046 0.338 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
        RECT 2.234 0.338 2.302 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.248 2.518 0.382 ;
        RECT 1.154 0.248 2.518 0.292 ;
        RECT 1.154 0.158 1.222 0.292 ;
      LAYER v0 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.586 0.248 1.654 0.292 ;
        RECT 1.91 0.248 1.978 0.292 ;
        RECT 2.126 0.248 2.194 0.292 ;
        RECT 2.342 0.248 2.41 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 1.006 0.202 ;
        RECT 0.074 0.428 0.898 0.472 ;
        RECT 0.83 0.338 0.898 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.832 0.358 0.896 0.402 ;
        RECT 0.83 0.158 0.898 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.138 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.138 0.022 ;
        RECT 3.854 -0.022 3.922 0.112 ;
        RECT 3.638 -0.022 3.706 0.112 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 3.424 0.048 3.488 0.092 ;
        RECT 3.64 0.048 3.704 0.092 ;
        RECT 3.856 0.048 3.92 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.154 0.428 2.558 0.472 ;
      RECT 2.646 0.068 3.206 0.112 ;
    LAYER v0 ;
      RECT 3.962 0.158 4.03 0.202 ;
      RECT 3.962 0.518 4.03 0.562 ;
      RECT 3.856 0.358 3.92 0.402 ;
      RECT 3.746 0.158 3.814 0.202 ;
      RECT 3.746 0.518 3.814 0.562 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.53 0.158 3.598 0.202 ;
      RECT 3.53 0.518 3.598 0.562 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.314 0.518 3.382 0.562 ;
      RECT 3.206 0.248 3.274 0.292 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 3.098 0.518 3.166 0.562 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.882 0.518 2.95 0.562 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
    LAYER m1 ;
      RECT 0.486 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.158 3.098 0.202 ;
      RECT 3.098 0.158 3.166 0.292 ;
      RECT 2.754 0.428 3.314 0.472 ;
      RECT 3.166 0.248 3.314 0.292 ;
      RECT 3.314 0.248 3.382 0.472 ;
      RECT 3.382 0.428 3.854 0.472 ;
      RECT 3.854 0.338 3.922 0.472 ;
      RECT 2.558 0.428 2.626 0.562 ;
      RECT 2.626 0.518 4.05 0.562 ;
      RECT 3.206 0.068 3.274 0.202 ;
      RECT 3.274 0.158 4.05 0.202 ;
  END
END b15ao0022as1n32x5

MACRO b15aoai13as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoai13as1n02x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.594 0.112 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.4335 0.466 0.4775 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
END b15aoai13as1n02x3

MACRO b15aoai13as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoai13as1n02x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.702 0.202 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.388 0.574 0.432 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.3835 0.25 0.4275 ;
        RECT 0.614 0.538 0.682 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.202 ;
      RECT 0.25 0.158 0.398 0.202 ;
      RECT 0.398 0.068 0.466 0.202 ;
      RECT 0.466 0.068 0.594 0.112 ;
  END
END b15aoai13as1n02x5

MACRO b15aoai13as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoai13as1n03x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.3605 0.898 0.4045 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.3605 0.574 0.4045 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.45666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.473 0.466 0.517 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.248 0.574 0.292 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.79 0.382 ;
        RECT 0.722 0.068 0.79 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.473 0.682 0.517 ;
        RECT 0.722 0.1365 0.79 0.1805 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
        RECT 0.722 0.473 0.79 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.114 0.142 0.158 ;
        RECT 0.506 0.048 0.574 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.202 ;
    LAYER v0 ;
      RECT 0.616 0.228 0.68 0.272 ;
      RECT 0.29 0.473 0.358 0.517 ;
      RECT 0.292 0.088 0.356 0.132 ;
      RECT 0.074 0.473 0.142 0.517 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.142 0.338 0.29 0.382 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.358 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.292 ;
  END
END b15aoai13as1n03x5

MACRO b15aoai13as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoai13as1n04x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.31901225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.31901225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4128395 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
        RECT 0.378 0.338 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 1.026 0.112 ;
        RECT 0.83 0.068 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.4535 0.898 0.4975 ;
        RECT 0.938 0.068 1.006 0.112 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.472 0.25 0.516 ;
        RECT 0.398 0.472 0.466 0.516 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.682 0.202 ;
    LAYER v0 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
  END
END b15aoai13as1n04x5

MACRO b15aoai13as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoai13as1n06x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.158 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.355873 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38324775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.289 0.79 0.333 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03978 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 3.20285725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.428 1.33 0.472 ;
        RECT 1.046 0.248 1.222 0.292 ;
        RECT 1.154 0.158 1.222 0.292 ;
        RECT 0.83 0.518 1.114 0.562 ;
        RECT 1.046 0.248 1.114 0.562 ;
        RECT 0.83 0.338 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.383 0.898 0.427 ;
        RECT 1.156 0.178 1.22 0.222 ;
        RECT 1.154 0.428 1.222 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 1.264 0.538 1.328 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.83 0.112 ;
      RECT 0.074 0.158 0.79 0.202 ;
    LAYER v0 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.184 0.408 0.248 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.472 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.158 1.046 0.202 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.114 0.068 1.35 0.112 ;
  END
END b15aoai13as1n06x5

MACRO b15aoai13as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoai13as1n08x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.158 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.293 1.438 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.436875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.436875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.178 0.898 0.222 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 0.79 0.472 ;
        RECT 0.486 0.338 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 0.66617275 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 1.458 0.472 ;
        RECT 1.262 0.158 1.33 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.262 0.178 1.33 0.222 ;
        RECT 1.37 0.428 1.438 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.046 0.178 1.114 0.222 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 0.614 0.472 ;
      RECT 0.486 0.068 0.938 0.112 ;
    LAYER v0 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.1355 0.25 0.1795 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.25 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.682 0.518 1.134 0.562 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.006 0.338 1.154 0.382 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.222 0.068 1.458 0.112 ;
  END
END b15aoai13as1n08x5

MACRO b15aob012as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aob012as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.594 0.112 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.4505 0.466 0.4945 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4505 0.142 0.4945 ;
        RECT 0.29 0.4505 0.358 0.4945 ;
        RECT 0.506 0.4505 0.574 0.4945 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.4505 0.25 0.4945 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15aob012as1n02x5

MACRO b15aob012as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aob012as1n03x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.574 0.202 ;
        RECT 0.506 0.068 0.574 0.202 ;
        RECT 0.398 0.158 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.508 0.088 0.572 0.132 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15aob012as1n03x5

MACRO b15aob012as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aob012as1n04x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.574 0.202 ;
        RECT 0.506 0.068 0.574 0.202 ;
        RECT 0.398 0.158 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.508 0.088 0.572 0.132 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.076 0.088 0.14 0.132 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.202 ;
      RECT 0.142 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
  END
END b15aob012as1n04x5

MACRO b15aob012as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aob012as1n06x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 0.614 0.448 0.682 0.492 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.722 0.048 0.79 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.076 0.088 0.14 0.132 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.202 ;
      RECT 0.142 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
  END
END b15aob012as1n06x5

MACRO b15aob012as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aob012as1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.4505 0.466 0.4945 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 0.614 0.4505 0.682 0.4945 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.4505 0.358 0.4945 ;
        RECT 0.506 0.4505 0.574 0.4945 ;
        RECT 0.722 0.4505 0.79 0.4945 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.722 0.158 0.79 0.202 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.4505 0.25 0.4945 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15aob012as1n08x5

MACRO b15aob012as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aob012as1n12x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.158 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.293 1.438 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.594 0.382 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.472 ;
        RECT 1.262 0.158 1.33 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.262 0.178 1.33 0.222 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.478 0.178 1.546 0.222 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.046 0.538 1.114 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.182 0.472 ;
      RECT 0.938 0.158 1.006 0.382 ;
    LAYER v0 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.428 0.722 0.472 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 1.006 0.338 1.154 0.382 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.222 0.068 1.546 0.112 ;
  END
END b15aob012as1n12x5

MACRO b15aob012as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aob012as1n16x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.158 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.293 1.978 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.07416675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.555625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.158 0.79 0.202 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.562 ;
        RECT 1.046 0.338 1.87 0.382 ;
        RECT 1.586 0.158 1.654 0.562 ;
        RECT 1.262 0.338 1.33 0.562 ;
        RECT 1.046 0.338 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.4485 1.114 0.4925 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.586 0.4465 1.654 0.4905 ;
        RECT 1.586 0.178 1.654 0.222 ;
        RECT 1.802 0.4405 1.87 0.4845 ;
        RECT 1.802 0.1785 1.87 0.2225 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.938 0.068 1.006 0.292 ;
    LAYER v0 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.372 0.178 1.436 0.222 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.25 0.338 0.506 0.382 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.574 0.338 0.83 0.382 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.438 0.068 1.998 0.112 ;
  END
END b15aob012as1n16x5

MACRO b15aob012as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aob012as1n24x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5831945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.293 1.654 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.472 ;
        RECT 1.694 0.158 1.762 0.472 ;
        RECT 1.478 0.158 1.546 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.478 0.178 1.546 0.222 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.694 0.1785 1.762 0.2225 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.91 0.1785 1.978 0.2225 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.938 0.068 1.006 0.382 ;
    LAYER v0 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.37 0.178 1.438 0.222 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.1785 0.466 0.2225 ;
      RECT 0.29 0.1785 0.358 0.2225 ;
      RECT 0.182 0.068 0.25 0.112 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.1785 0.142 0.2225 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.068 0.682 0.382 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.358 0.428 0.83 0.472 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.006 0.338 1.154 0.382 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.068 1.438 0.382 ;
      RECT 1.438 0.068 1.978 0.112 ;
  END
END b15aob012as1n24x5

MACRO b15aobi12as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aobi12as1n02x3 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.6075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.6075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.4595 0.358 0.5035 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.398 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.574 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.4595 0.466 0.5035 ;
        RECT 0.506 0.205 0.574 0.249 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.614 0.4685 0.682 0.5125 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.209 0.142 0.253 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.722 0.048 0.79 0.092 ;
    END
  END vssx
END b15aobi12as1n02x3

MACRO b15aobi12as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aobi12as1n02x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.6075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.6075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.4595 0.358 0.5035 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.398 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.574 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.4595 0.466 0.5035 ;
        RECT 0.506 0.205 0.574 0.249 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.614 0.4685 0.682 0.5125 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.209 0.142 0.253 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.722 0.048 0.79 0.092 ;
    END
  END vssx
END b15aobi12as1n02x5

MACRO b15aobi12as1n02x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aobi12as1n02x7 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.4555 0.466 0.4995 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.186 0.358 0.23 ;
        RECT 0.83 0.048 0.898 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
    LAYER v0 ;
      RECT 0.83 0.436 0.898 0.48 ;
      RECT 0.506 0.4555 0.574 0.4995 ;
      RECT 0.182 0.186 0.25 0.23 ;
      RECT 0.182 0.4055 0.25 0.4495 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.83 0.202 ;
      RECT 0.83 0.158 0.898 0.562 ;
  END
END b15aobi12as1n02x7

MACRO b15aobi12as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aobi12as1n04x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.506 0.068 0.898 0.112 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.1855 0.574 0.2295 ;
        RECT 0.83 0.153 0.898 0.197 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.046 0.338 1.114 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.83 0.4555 0.898 0.4995 ;
        RECT 1.046 0.4005 1.114 0.4445 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.073 0.142 0.117 ;
        RECT 0.398 0.1855 0.466 0.2295 ;
        RECT 1.046 0.198 1.114 0.242 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
    LAYER v0 ;
      RECT 0.614 0.42 0.682 0.464 ;
      RECT 0.398 0.4505 0.466 0.4945 ;
      RECT 0.182 0.203 0.25 0.247 ;
      RECT 0.182 0.3905 0.25 0.4345 ;
    LAYER m1 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
  END
END b15aobi12as1n04x5

MACRO b15aobi12as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aobi12as1n06x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.248 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.37 0.293 1.438 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.83 0.068 1.114 0.112 ;
        RECT 0.506 0.248 0.898 0.292 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.508 0.176 0.572 0.22 ;
        RECT 0.83 0.153 0.898 0.197 ;
        RECT 1.046 0.153 1.114 0.197 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 1.262 0.338 1.33 0.652 ;
        RECT 1.046 0.338 1.114 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.3905 0.142 0.4345 ;
        RECT 0.83 0.4005 0.898 0.4445 ;
        RECT 1.046 0.4555 1.114 0.4995 ;
        RECT 1.262 0.4005 1.33 0.4445 ;
        RECT 1.478 0.4005 1.546 0.4445 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 1.262 -0.022 1.33 0.292 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.073 0.142 0.117 ;
        RECT 0.398 0.077 0.466 0.121 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 1.262 0.198 1.33 0.242 ;
        RECT 1.478 0.198 1.546 0.242 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
    LAYER v0 ;
      RECT 0.614 0.42 0.682 0.464 ;
      RECT 0.398 0.4505 0.466 0.4945 ;
      RECT 0.182 0.203 0.25 0.247 ;
      RECT 0.182 0.3905 0.25 0.4345 ;
    LAYER m1 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
  END
END b15aobi12as1n06x5

MACRO b15aobi12as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aobi12as1n08x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5875925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5875925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.158 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.293 1.762 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06732 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.292 ;
        RECT 0.83 0.068 1.33 0.112 ;
        RECT 0.83 0.068 0.898 0.472 ;
        RECT 0.614 0.248 0.898 0.292 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.616 0.178 0.68 0.222 ;
        RECT 0.614 0.3665 0.682 0.4105 ;
        RECT 0.832 0.178 0.896 0.222 ;
        RECT 0.83 0.3665 0.898 0.4105 ;
        RECT 1.046 0.068 1.114 0.112 ;
        RECT 1.262 0.178 1.33 0.222 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.49 0.358 0.534 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.096 0.142 0.14 ;
        RECT 0.29 0.096 0.358 0.14 ;
        RECT 0.506 0.096 0.574 0.14 ;
        RECT 0.722 0.096 0.79 0.14 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.154 0.158 1.222 0.382 ;
      RECT 0.506 0.428 0.574 0.562 ;
    LAYER v0 ;
      RECT 1.586 0.178 1.654 0.222 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.178 1.438 0.222 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.724 0.448 0.788 0.492 ;
      RECT 0.508 0.448 0.572 0.492 ;
      RECT 0.398 0.268 0.466 0.312 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.184 0.408 0.248 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.248 0.466 0.382 ;
      RECT 1.222 0.338 1.37 0.382 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 0.574 0.518 0.722 0.562 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.79 0.518 0.938 0.562 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 1.006 0.428 1.762 0.472 ;
  END
END b15aobi12as1n08x5

MACRO b15aobi12as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aobi12as1n12x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.998 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.586 0.338 1.654 0.382 ;
        RECT 1.91 0.338 1.978 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.35 0.248 2.086 0.292 ;
        RECT 2.018 0.158 2.086 0.292 ;
      LAYER v0 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.10098 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 2.106 0.112 ;
        RECT 1.262 0.158 1.978 0.202 ;
        RECT 1.91 0.068 1.978 0.202 ;
        RECT 1.262 0.068 1.33 0.202 ;
        RECT 0.938 0.068 1.33 0.112 ;
        RECT 0.938 0.068 1.006 0.472 ;
        RECT 0.506 0.248 1.006 0.292 ;
        RECT 0.722 0.158 0.79 0.472 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.508 0.178 0.572 0.222 ;
        RECT 0.506 0.3665 0.574 0.4105 ;
        RECT 0.724 0.178 0.788 0.222 ;
        RECT 0.722 0.3665 0.79 0.4105 ;
        RECT 0.94 0.178 1.004 0.222 ;
        RECT 0.938 0.3665 1.006 0.4105 ;
        RECT 1.154 0.068 1.222 0.112 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.018 0.068 2.086 0.112 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.614 0.0945 0.682 0.1385 ;
        RECT 0.83 0.0945 0.898 0.1385 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.428 0.682 0.562 ;
    LAYER v0 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 0.832 0.448 0.896 0.492 ;
      RECT 0.616 0.448 0.68 0.492 ;
      RECT 0.398 0.268 0.466 0.312 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.184 0.408 0.248 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.248 0.466 0.382 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.898 0.518 1.046 0.562 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.114 0.428 2.086 0.472 ;
  END
END b15aobi12as1n12x5

MACRO b15aobi12as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aobi12as1n16x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 2.538 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
        RECT 1.694 0.338 1.762 0.382 ;
        RECT 2.126 0.338 2.194 0.382 ;
        RECT 2.45 0.338 2.518 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.35 0.248 2.626 0.292 ;
        RECT 2.558 0.158 2.626 0.292 ;
      LAYER v0 ;
        RECT 1.478 0.248 1.546 0.292 ;
        RECT 1.91 0.248 1.978 0.292 ;
        RECT 2.342 0.248 2.41 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14076 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.646 0.112 ;
        RECT 1.37 0.158 2.518 0.202 ;
        RECT 2.45 0.068 2.518 0.202 ;
        RECT 1.37 0.068 1.438 0.202 ;
        RECT 1.046 0.068 1.438 0.112 ;
        RECT 1.046 0.068 1.114 0.472 ;
        RECT 0.614 0.248 1.114 0.292 ;
        RECT 0.83 0.068 0.898 0.472 ;
        RECT 0.614 0.068 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.3995 0.682 0.4435 ;
        RECT 0.614 0.15 0.682 0.194 ;
        RECT 0.83 0.3995 0.898 0.4435 ;
        RECT 0.83 0.15 0.898 0.194 ;
        RECT 1.046 0.3995 1.114 0.4435 ;
        RECT 1.046 0.15 1.114 0.194 ;
        RECT 1.262 0.068 1.33 0.112 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.558 0.068 2.626 0.112 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.594 0.518 1.154 0.562 ;
    LAYER v0 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.2575 0.574 0.3015 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.4535 0.466 0.4975 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.4535 0.25 0.4975 ;
    LAYER m1 ;
      RECT 0.358 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.506 0.382 ;
      RECT 0.358 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.25 0.338 0.29 0.382 ;
      RECT 0.074 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.382 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.222 0.428 2.626 0.472 ;
  END
END b15aobi12as1n16x5

MACRO b15aoi012as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi012as1n02x3 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.518 0.486 0.562 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.1285 0.358 0.1725 ;
        RECT 0.398 0.518 0.466 0.562 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.398 0.048 0.466 0.092 ;
    END
  END vssx
END b15aoi012as1n02x3

MACRO b15aoi012as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi012as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.518 0.486 0.562 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.1285 0.358 0.1725 ;
        RECT 0.398 0.518 0.466 0.562 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
    END
  END vssx
END b15aoi012as1n02x5

MACRO b15aoi012as1n02x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi012as1n02x7 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.15333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.182 0.2 0.25 0.244 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.182 0.518 0.25 0.562 ;
    LAYER m1 ;
      RECT 0.162 0.518 0.29 0.562 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.594 0.472 ;
  END
END b15aoi012as1n02x7

MACRO b15aoi012as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi012as1n04x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.472 ;
        RECT 0.398 0.068 0.79 0.112 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.166 0.466 0.21 ;
        RECT 0.722 0.388 0.79 0.432 ;
        RECT 0.722 0.171 0.79 0.215 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4105 0.25 0.4545 ;
        RECT 0.398 0.448 0.466 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.166 0.25 0.21 ;
        RECT 0.83 0.0905 0.898 0.1345 ;
    END
  END vssx
END b15aoi012as1n04x5

MACRO b15aoi012as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi012as1n06x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.702 0.382 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.81 0.338 1.006 0.382 ;
        RECT 0.938 0.248 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04284 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.79 0.112 ;
        RECT 0.074 0.428 0.358 0.472 ;
        RECT 0.29 0.068 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.183 0.142 0.227 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.29 0.183 0.358 0.227 ;
        RECT 0.614 0.068 0.682 0.112 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
      LAYER v0 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.292 ;
    LAYER v0 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.508 0.228 0.572 0.272 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.398 0.562 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.428 1.026 0.472 ;
      RECT 0.574 0.158 1.026 0.202 ;
  END
END b15aoi012as1n06x5

MACRO b15aoi012as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi012as1n08x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.3155 0.25 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.81 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.338 1.222 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.898 0.112 ;
        RECT 0.074 0.158 0.466 0.202 ;
        RECT 0.398 0.068 0.466 0.202 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.408 0.142 0.452 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.29 0.408 0.358 0.452 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 0.722 0.068 0.79 0.112 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
      LAYER v0 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.518 0.398 0.562 ;
    LAYER v0 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.048 0.228 1.112 0.272 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.616 0.228 0.68 0.272 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.182 0.518 0.25 0.562 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.428 1.242 0.472 ;
  END
END b15aoi012as1n08x5

MACRO b15aoi012as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi012as1n12x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 1.026 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.134 0.338 1.546 0.382 ;
        RECT 1.478 0.248 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 1.114 0.112 ;
        RECT 0.398 0.068 0.466 0.472 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.182 0.136 0.25 0.18 ;
        RECT 0.398 0.408 0.466 0.452 ;
        RECT 0.398 0.162 0.466 0.206 ;
        RECT 0.722 0.068 0.79 0.112 ;
        RECT 0.938 0.068 1.006 0.112 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
      LAYER v0 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.292 ;
    LAYER v0 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.616 0.228 0.68 0.272 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.614 0.562 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.682 0.428 1.566 0.472 ;
      RECT 0.682 0.158 1.566 0.202 ;
  END
END b15aoi012as1n12x5

MACRO b15aoi012as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi012as1n16x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63973075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.293 1.654 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.473923 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.473923 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11934 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.428 1.89 0.472 ;
        RECT 1.694 0.158 1.762 0.472 ;
        RECT 1.478 0.158 1.546 0.472 ;
        RECT 1.262 0.068 1.33 0.472 ;
        RECT 0.614 0.068 1.33 0.112 ;
      LAYER v0 ;
        RECT 0.722 0.068 0.79 0.112 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 1.154 0.068 1.222 0.112 ;
        RECT 1.262 0.203 1.33 0.247 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.478 0.203 1.546 0.247 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.694 0.203 1.762 0.247 ;
        RECT 1.802 0.428 1.87 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 1.37 0.203 1.438 0.247 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 1.802 0.203 1.87 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 1.154 0.472 ;
    LAYER v0 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.048 0.178 1.112 0.222 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.832 0.178 0.896 0.222 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.158 0.898 0.292 ;
      RECT 0.898 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.222 0.518 1.89 0.562 ;
  END
END b15aoi012as1n16x5

MACRO b15aoi012as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi012as1n24x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.50276925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68083325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
        RECT 0.27 0.248 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.543611 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.543611 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.782 0.382 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.694 0.338 1.762 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.543611 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.543611 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.89 0.338 2.734 0.382 ;
        RECT 2.666 0.248 2.734 0.382 ;
      LAYER v0 ;
        RECT 1.91 0.338 1.978 0.382 ;
        RECT 2.126 0.338 2.194 0.382 ;
        RECT 2.342 0.338 2.41 0.382 ;
        RECT 2.558 0.338 2.626 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14382 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 1.782 0.112 ;
        RECT 0.074 0.158 0.898 0.202 ;
        RECT 0.83 0.068 0.898 0.202 ;
        RECT 0.722 0.158 0.79 0.472 ;
        RECT 0.506 0.338 0.574 0.472 ;
        RECT 0.074 0.338 0.574 0.382 ;
        RECT 0.29 0.338 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.076 0.408 0.14 0.452 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.292 0.408 0.356 0.452 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.508 0.408 0.572 0.452 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.724 0.408 0.788 0.452 ;
        RECT 1.046 0.068 1.114 0.112 ;
        RECT 1.262 0.068 1.33 0.112 ;
        RECT 1.478 0.068 1.546 0.112 ;
        RECT 1.694 0.068 1.762 0.112 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
      LAYER v0 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.292 ;
    LAYER v0 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.94 0.228 1.004 0.272 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.182 0.518 0.25 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.938 0.562 ;
      RECT 0.938 0.428 1.006 0.562 ;
      RECT 1.006 0.428 2.754 0.472 ;
      RECT 1.006 0.158 2.754 0.202 ;
  END
END b15aoi012as1n24x5

MACRO b15aoi012as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi012as1n32x5 0 0 ;
  SIZE 3.996 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.47793825 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.724375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.682 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5524075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5524075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 2.538 0.292 ;
        RECT 1.154 0.248 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.586 0.248 1.654 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.018 0.248 2.086 0.292 ;
        RECT 2.234 0.248 2.302 0.292 ;
        RECT 2.45 0.248 2.518 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5524075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5524075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.248 3.922 0.382 ;
        RECT 2.646 0.248 3.922 0.292 ;
      LAYER v0 ;
        RECT 2.666 0.248 2.734 0.292 ;
        RECT 2.882 0.248 2.95 0.292 ;
        RECT 3.098 0.248 3.166 0.292 ;
        RECT 3.314 0.248 3.382 0.292 ;
        RECT 3.53 0.248 3.598 0.292 ;
        RECT 3.746 0.248 3.814 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.19584 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 2.626 0.112 ;
        RECT 1.046 0.068 1.114 0.472 ;
        RECT 0.054 0.158 1.114 0.202 ;
        RECT 0.182 0.428 1.006 0.472 ;
        RECT 0.722 0.158 0.79 0.472 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.184 0.358 0.248 0.402 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.408 1.114 0.452 ;
        RECT 1.37 0.068 1.438 0.112 ;
        RECT 1.586 0.068 1.654 0.112 ;
        RECT 1.802 0.068 1.87 0.112 ;
        RECT 2.018 0.068 2.086 0.112 ;
        RECT 2.234 0.068 2.302 0.112 ;
        RECT 2.45 0.068 2.518 0.112 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
      LAYER v0 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
        RECT 3.748 0.538 3.812 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.03 0.022 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.316 0.048 3.38 0.092 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.748 0.048 3.812 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.154 0.158 3.942 0.202 ;
    LAYER v0 ;
      RECT 3.854 0.158 3.922 0.202 ;
      RECT 3.854 0.428 3.922 0.472 ;
      RECT 3.638 0.158 3.706 0.202 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 1.262 0.562 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.33 0.428 3.942 0.472 ;
  END
END b15aoi012as1n32x5

MACRO b15aoi013as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi013as1n02x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 0.594 0.562 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.506 0.518 0.574 0.562 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
    END
  END vssx
END b15aoi013as1n02x3

MACRO b15aoi013as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi013as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 0.594 0.562 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.136 0.466 0.18 ;
        RECT 0.506 0.518 0.574 0.562 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
    END
  END vssx
END b15aoi013as1n02x5

MACRO b15aoi013as1n02x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi013as1n02x7 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.2705 0.682 0.3145 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.2705 0.466 0.3145 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.2705 0.358 0.3145 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.518 0.702 0.562 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.1575 0.574 0.2015 ;
        RECT 0.614 0.518 0.682 0.562 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.398 0.448 0.466 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
    END
  END vssx
END b15aoi013as1n02x7

MACRO b15aoi013as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi013as1n03x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.760139 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.173426 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.403 0.574 0.447 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.330139 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.553426 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.403 0.682 0.447 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.594 0.202 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.158 0.574 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 1.046 0.138 1.114 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.248 0.358 0.472 ;
    LAYER v0 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.29 0.408 0.358 0.452 ;
    LAYER m1 ;
      RECT 0.378 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.79 0.158 0.918 0.202 ;
      RECT 0.358 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.472 ;
  END
END b15aoi013as1n03x5

MACRO b15aoi013as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi013as1n04x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.3155 0.682 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.222 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.574 0.292 ;
        RECT 0.506 0.158 0.574 0.292 ;
        RECT 0.29 0.158 0.358 0.292 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.292 0.178 0.356 0.222 ;
        RECT 0.508 0.178 0.572 0.222 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.518 0.398 0.562 ;
    LAYER v0 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.94 0.088 1.004 0.132 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.158 0.938 0.202 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.428 1.242 0.472 ;
  END
END b15aoi013as1n04x5

MACRO b15aoi013as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi013as1n06x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.134 0.382 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.242 0.338 1.546 0.382 ;
        RECT 1.478 0.158 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05814 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.292 ;
        RECT 0.398 0.158 0.79 0.202 ;
        RECT 0.054 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.472 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.724 0.228 0.788 0.272 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
      LAYER v0 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.046 0.538 1.114 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 1.478 0.048 1.546 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.594 0.068 1.134 0.112 ;
      RECT 0.162 0.518 0.506 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.372 0.228 1.436 0.272 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.94 0.228 1.004 0.272 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.182 0.518 0.25 0.562 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.37 0.202 ;
      RECT 1.37 0.158 1.438 0.292 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.428 1.546 0.472 ;
  END
END b15aoi013as1n06x5

MACRO b15aoi013as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi013as1n08x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.28915825 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.28915825 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.134 0.382 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.35267975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.242 0.338 1.546 0.382 ;
        RECT 1.478 0.158 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07038 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.292 ;
        RECT 0.398 0.158 0.79 0.202 ;
        RECT 0.054 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.472 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.724 0.228 0.788 0.272 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
      LAYER v0 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.594 0.068 1.134 0.112 ;
      RECT 0.162 0.518 0.506 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.372 0.228 1.436 0.272 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.94 0.228 1.004 0.272 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.182 0.518 0.25 0.562 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.37 0.202 ;
      RECT 1.37 0.158 1.438 0.292 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.428 1.546 0.472 ;
  END
END b15aoi013as1n08x5

MACRO b15aoi022as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi022as1n02x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.398 0.428 0.466 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
END b15aoi022as1n02x3

MACRO b15aoi022as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi022as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.203 0.574 0.247 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
        RECT 0.182 0.068 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.398 0.318 0.466 0.362 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.398 0.472 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.518 0.594 0.562 ;
  END
END b15aoi022as1n02x5

MACRO b15aoi022as1n04x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi022as1n04x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.562 ;
        RECT 0.29 0.158 0.466 0.202 ;
        RECT 0.29 0.068 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.292 0.088 0.356 0.132 ;
        RECT 0.398 0.433 0.466 0.477 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
END b15aoi022as1n04x3

MACRO b15aoi022as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi022as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
        RECT 0.398 0.158 0.574 0.202 ;
        RECT 0.398 0.068 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.4 0.088 0.464 0.132 ;
        RECT 0.506 0.408 0.574 0.452 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.518 0.702 0.562 ;
  END
END b15aoi022as1n04x5

MACRO b15aoi022as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi022as1n06x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.562 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.518 1.114 0.562 ;
        RECT 1.046 0.338 1.114 0.562 ;
        RECT 0.83 0.158 0.898 0.562 ;
        RECT 0.614 0.158 0.682 0.562 ;
        RECT 0.378 0.158 0.682 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.83 0.408 0.898 0.452 ;
        RECT 0.83 0.178 0.898 0.222 ;
        RECT 1.046 0.408 1.114 0.452 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 1.046 0.158 1.114 0.202 ;
    END
  END vssx
END b15aoi022as1n06x5

MACRO b15aoi022as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi022as1n08x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 0.66617275 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.81 0.428 1.35 0.472 ;
        RECT 0.938 0.068 1.006 0.472 ;
        RECT 0.506 0.068 1.006 0.112 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.508 0.138 0.572 0.182 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.938 0.1805 1.006 0.2245 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.262 0.428 1.33 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 0.074 0.428 0.702 0.472 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.614 0.428 0.682 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 1.154 -0.022 1.222 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.29 0.1795 0.358 0.2235 ;
        RECT 1.154 0.1805 1.222 0.2245 ;
        RECT 1.37 0.158 1.438 0.202 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.27 0.518 1.458 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.29 0.518 0.358 0.562 ;
  END
END b15aoi022as1n08x5

MACRO b15aoi022as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi022as1n12x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.158 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.158 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.293 1.762 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.428 1.762 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.614 0.338 1.006 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.178 0.682 0.222 ;
        RECT 0.938 0.178 1.006 0.222 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.154 0.178 1.222 0.222 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.586 0.428 1.654 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.938 0.068 1.37 0.112 ;
      RECT 0.054 0.428 0.83 0.472 ;
    LAYER v0 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.178 1.654 0.222 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.382 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.466 0.068 0.81 0.112 ;
      RECT 1.37 0.068 1.438 0.382 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.898 0.518 1.782 0.562 ;
  END
END b15aoi022as1n12x5

MACRO b15aoi022as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi022as1n16x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 1.006 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 1.006 0.292 ;
        RECT 0.938 0.158 1.006 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.978 0.292 ;
        RECT 1.91 0.068 1.978 0.292 ;
      LAYER v0 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 2.086 0.382 ;
        RECT 2.018 0.158 2.086 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.586 0.338 1.654 0.382 ;
        RECT 1.91 0.338 1.978 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11016 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.87 0.202 ;
        RECT 1.802 0.068 1.87 0.202 ;
        RECT 0.074 0.428 1.114 0.472 ;
        RECT 1.046 0.068 1.114 0.472 ;
        RECT 0.83 0.068 1.114 0.112 ;
        RECT 0.182 0.158 0.898 0.202 ;
        RECT 0.83 0.068 0.898 0.202 ;
        RECT 0.182 0.068 0.25 0.202 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.804 0.088 1.868 0.132 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
      LAYER v0 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 1.154 0.562 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.222 0.428 2.106 0.472 ;
  END
END b15aoi022as1n16x5

MACRO b15aoi022as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi022as1n24x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAGATEAREA 0.0441 LAYER m2 ;
      ANTENNAMAXAREACAR 0.48081625 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68743775 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.1955555 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAGATEAREA 0.0441 LAYER m2 ;
      ANTENNAMAXAREACAR 0.48081625 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68743775 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.1955555 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.87 0.382 ;
        RECT 1.586 0.248 1.654 0.382 ;
      LAYER m2 ;
        RECT 1.568 0.338 2.012 0.382 ;
      LAYER v1 ;
        RECT 1.59 0.338 1.65 0.382 ;
        RECT 1.806 0.338 1.866 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.293 1.654 0.337 ;
        RECT 1.802 0.293 1.87 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAGATEAREA 0.0441 LAYER m2 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63746025 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.1955555 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAGATEAREA 0.0441 LAYER m2 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63746025 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.1955555 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.248 2.518 0.382 ;
        RECT 2.126 0.248 2.194 0.382 ;
      LAYER m2 ;
        RECT 2.092 0.338 2.552 0.382 ;
      LAYER v1 ;
        RECT 2.13 0.338 2.19 0.382 ;
        RECT 2.454 0.338 2.514 0.382 ;
      LAYER v0 ;
        RECT 2.126 0.293 2.194 0.337 ;
        RECT 2.45 0.293 2.518 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAGATEAREA 0.0441 LAYER m2 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63746025 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.26340125 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAGATEAREA 0.0441 LAYER m2 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63746025 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.26340125 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.382 ;
        RECT 0.938 0.248 1.006 0.382 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER m2 ;
        RECT 0.688 0.338 1.24 0.382 ;
      LAYER v1 ;
        RECT 0.726 0.338 0.786 0.382 ;
        RECT 0.942 0.338 1.002 0.382 ;
        RECT 1.158 0.338 1.218 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
        RECT 0.938 0.293 1.006 0.337 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAGATEAREA 0.0441 LAYER m2 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63746025 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.26340125 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAGATEAREA 0.0441 LAYER m2 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63746025 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.26340125 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.382 ;
        RECT 0.29 0.248 0.358 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER m2 ;
        RECT 0.04 0.338 0.608 0.382 ;
      LAYER v1 ;
        RECT 0.078 0.338 0.138 0.382 ;
        RECT 0.294 0.338 0.354 0.382 ;
        RECT 0.51 0.338 0.57 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.17748 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.432 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.428 2.518 0.472 ;
        RECT 1.694 0.158 1.762 0.472 ;
        RECT 1.478 0.158 1.546 0.472 ;
        RECT 1.262 0.068 1.33 0.472 ;
        RECT 0.702 0.068 1.33 0.112 ;
      LAYER v0 ;
        RECT 0.722 0.068 0.79 0.112 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 1.262 0.178 1.33 0.222 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.478 0.178 1.546 0.222 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.694 0.178 1.762 0.222 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.342 0.428 2.41 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.382 ;
      RECT 0.29 0.248 0.358 0.382 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.722 0.248 0.79 0.382 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 0.074 0.158 1.222 0.202 ;
      RECT 1.586 0.248 1.654 0.382 ;
      RECT 1.802 0.248 1.87 0.382 ;
      RECT 2.126 0.248 2.194 0.382 ;
      RECT 2.45 0.248 2.518 0.382 ;
      RECT 0.054 0.428 1.154 0.472 ;
    LAYER v0 ;
      RECT 2.45 0.518 2.518 0.562 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.37 0.178 1.438 0.222 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.438 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.202 ;
      RECT 1.978 0.158 2.518 0.202 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.222 0.518 2.538 0.562 ;
  END
END b15aoi022as1n24x5

MACRO b15aoi022as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi022as1n32x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAGATEAREA 0.0585 LAYER m2 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62085475 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.14741875 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAGATEAREA 0.0585 LAYER m2 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62085475 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.14741875 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.382 ;
        RECT 2.018 0.248 2.086 0.382 ;
      LAYER m2 ;
        RECT 2 0.338 2.428 0.382 ;
      LAYER v1 ;
        RECT 2.022 0.338 2.082 0.382 ;
        RECT 2.238 0.338 2.298 0.382 ;
      LAYER v0 ;
        RECT 2.018 0.293 2.086 0.337 ;
        RECT 2.234 0.293 2.302 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAGATEAREA 0.0585 LAYER m2 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62085475 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.14741875 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAGATEAREA 0.0585 LAYER m2 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62085475 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.14741875 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.248 3.274 0.382 ;
        RECT 2.99 0.248 3.058 0.382 ;
      LAYER m2 ;
        RECT 2.864 0.338 3.308 0.382 ;
      LAYER v1 ;
        RECT 2.994 0.338 3.054 0.382 ;
        RECT 3.21 0.338 3.27 0.382 ;
      LAYER v0 ;
        RECT 2.99 0.293 3.058 0.337 ;
        RECT 3.206 0.293 3.274 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAGATEAREA 0.0585 LAYER m2 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62085475 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.2497095 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAGATEAREA 0.0585 LAYER m2 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62085475 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.2497095 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.248 1.654 0.382 ;
        RECT 1.37 0.248 1.438 0.382 ;
        RECT 1.154 0.248 1.222 0.382 ;
        RECT 0.938 0.248 1.006 0.382 ;
      LAYER m2 ;
        RECT 0.904 0.338 1.672 0.382 ;
      LAYER v1 ;
        RECT 0.942 0.338 1.002 0.382 ;
        RECT 1.158 0.338 1.218 0.382 ;
        RECT 1.374 0.338 1.434 0.382 ;
        RECT 1.59 0.338 1.65 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
        RECT 1.154 0.293 1.222 0.337 ;
        RECT 1.37 0.293 1.438 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAGATEAREA 0.0585 LAYER m2 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62085475 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.2497095 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAGATEAREA 0.0585 LAYER m2 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62085475 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.2497095 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
        RECT 0.29 0.248 0.358 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER m2 ;
        RECT 0.04 0.338 0.824 0.382 ;
      LAYER v1 ;
        RECT 0.078 0.338 0.138 0.382 ;
        RECT 0.294 0.338 0.354 0.382 ;
        RECT 0.51 0.338 0.57 0.382 ;
        RECT 0.726 0.338 0.786 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2142 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.432 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.428 3.294 0.472 ;
        RECT 2.342 0.158 2.41 0.472 ;
        RECT 2.126 0.158 2.194 0.472 ;
        RECT 1.91 0.158 1.978 0.472 ;
        RECT 1.694 0.068 1.762 0.472 ;
        RECT 0.918 0.068 1.762 0.112 ;
      LAYER v0 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 1.154 0.068 1.222 0.112 ;
        RECT 1.37 0.068 1.438 0.112 ;
        RECT 1.694 0.178 1.762 0.222 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.91 0.178 1.978 0.222 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.126 0.178 2.194 0.222 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.342 0.178 2.41 0.222 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 3.098 0.428 3.166 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 3.206 -0.022 3.274 0.112 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
        RECT 3.208 0.048 3.272 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.382 ;
      RECT 0.29 0.248 0.358 0.382 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.722 0.248 0.79 0.382 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.37 0.248 1.438 0.382 ;
      RECT 1.586 0.248 1.654 0.382 ;
      RECT 0.074 0.158 1.654 0.202 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 2.234 0.248 2.302 0.382 ;
      RECT 2.99 0.248 3.058 0.382 ;
      RECT 3.206 0.248 3.274 0.382 ;
      RECT 0.054 0.428 1.586 0.472 ;
    LAYER v0 ;
      RECT 3.206 0.518 3.274 0.562 ;
      RECT 3.098 0.158 3.166 0.202 ;
      RECT 2.99 0.518 3.058 0.562 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.774 0.518 2.842 0.562 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.558 0.518 2.626 0.562 ;
      RECT 2.45 0.178 2.518 0.222 ;
      RECT 2.342 0.518 2.41 0.562 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.126 0.518 2.194 0.562 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.87 0.068 2.45 0.112 ;
      RECT 2.45 0.068 2.518 0.382 ;
      RECT 2.518 0.338 2.774 0.382 ;
      RECT 2.558 0.158 2.774 0.202 ;
      RECT 2.774 0.158 2.842 0.382 ;
      RECT 2.842 0.158 3.274 0.202 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.654 0.518 3.294 0.562 ;
  END
END b15aoi022as1n32x5

MACRO b15aoi022as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi022as1n48x5 0 0 ;
  SIZE 4.86 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAGATEAREA 0.0873 LAYER m2 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5570675 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.1330585 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAGATEAREA 0.0873 LAYER m2 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5570675 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.1330585 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 3.422 0.248 3.49 0.382 ;
        RECT 3.206 0.248 3.274 0.382 ;
        RECT 2.99 0.248 3.058 0.382 ;
      LAYER m2 ;
        RECT 2.972 0.338 3.508 0.382 ;
      LAYER v1 ;
        RECT 2.994 0.338 3.054 0.382 ;
        RECT 3.21 0.338 3.27 0.382 ;
        RECT 3.426 0.338 3.486 0.382 ;
      LAYER v0 ;
        RECT 2.99 0.293 3.058 0.337 ;
        RECT 3.206 0.293 3.274 0.337 ;
        RECT 3.422 0.293 3.49 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAGATEAREA 0.0873 LAYER m2 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5570675 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.167331 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAGATEAREA 0.0873 LAYER m2 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5570675 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.167331 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.718 0.248 4.786 0.382 ;
        RECT 4.502 0.248 4.57 0.382 ;
        RECT 4.286 0.248 4.354 0.382 ;
        RECT 4.07 0.248 4.138 0.382 ;
      LAYER m2 ;
        RECT 4.052 0.338 4.82 0.382 ;
      LAYER v1 ;
        RECT 4.074 0.338 4.134 0.382 ;
        RECT 4.29 0.338 4.35 0.382 ;
        RECT 4.506 0.338 4.566 0.382 ;
        RECT 4.722 0.338 4.782 0.382 ;
      LAYER v0 ;
        RECT 4.07 0.293 4.138 0.337 ;
        RECT 4.286 0.293 4.354 0.337 ;
        RECT 4.502 0.293 4.57 0.337 ;
        RECT 4.718 0.293 4.786 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAGATEAREA 0.0873 LAYER m2 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5570675 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.20160375 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAGATEAREA 0.0873 LAYER m2 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5570675 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.20160375 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.382 ;
        RECT 2.018 0.248 2.086 0.382 ;
        RECT 1.802 0.248 1.87 0.382 ;
        RECT 1.586 0.248 1.654 0.382 ;
        RECT 1.37 0.248 1.438 0.382 ;
      LAYER m2 ;
        RECT 1.352 0.338 2.32 0.382 ;
      LAYER v1 ;
        RECT 1.374 0.338 1.434 0.382 ;
        RECT 1.59 0.338 1.65 0.382 ;
        RECT 1.806 0.338 1.866 0.382 ;
        RECT 2.022 0.338 2.082 0.382 ;
        RECT 2.238 0.338 2.298 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.293 1.438 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
        RECT 1.802 0.293 1.87 0.337 ;
        RECT 2.018 0.293 2.086 0.337 ;
        RECT 2.234 0.293 2.302 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAGATEAREA 0.0873 LAYER m2 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5570675 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.20160375 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAGATEAREA 0.0873 LAYER m2 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5570675 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.20160375 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.382 ;
        RECT 0.722 0.248 0.79 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
        RECT 0.29 0.248 0.358 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER m2 ;
        RECT 0.04 0.338 1.024 0.382 ;
      LAYER v1 ;
        RECT 0.078 0.338 0.138 0.382 ;
        RECT 0.294 0.338 0.354 0.382 ;
        RECT 0.51 0.338 0.57 0.382 ;
        RECT 0.726 0.338 0.786 0.382 ;
        RECT 0.942 0.338 1.002 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.31212 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.428 4.806 0.472 ;
        RECT 3.53 0.158 3.598 0.472 ;
        RECT 3.314 0.158 3.382 0.472 ;
        RECT 3.098 0.158 3.166 0.472 ;
        RECT 2.882 0.158 2.95 0.472 ;
        RECT 2.666 0.158 2.734 0.472 ;
        RECT 2.45 0.068 2.518 0.472 ;
        RECT 1.242 0.068 2.518 0.112 ;
      LAYER v0 ;
        RECT 1.262 0.068 1.33 0.112 ;
        RECT 1.478 0.068 1.546 0.112 ;
        RECT 1.694 0.068 1.762 0.112 ;
        RECT 1.91 0.068 1.978 0.112 ;
        RECT 2.126 0.068 2.194 0.112 ;
        RECT 2.558 0.428 2.626 0.472 ;
        RECT 2.666 0.178 2.734 0.222 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.882 0.178 2.95 0.222 ;
        RECT 2.99 0.428 3.058 0.472 ;
        RECT 3.098 0.178 3.166 0.222 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.314 0.178 3.382 0.222 ;
        RECT 3.422 0.428 3.49 0.472 ;
        RECT 3.53 0.178 3.598 0.222 ;
        RECT 3.638 0.428 3.706 0.472 ;
        RECT 3.854 0.428 3.922 0.472 ;
        RECT 4.07 0.428 4.138 0.472 ;
        RECT 4.286 0.428 4.354 0.472 ;
        RECT 4.502 0.428 4.57 0.472 ;
        RECT 4.718 0.428 4.786 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.894 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.894 0.022 ;
        RECT 4.61 -0.022 4.678 0.112 ;
        RECT 4.394 -0.022 4.462 0.112 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 3.748 0.048 3.812 0.092 ;
        RECT 3.964 0.048 4.028 0.092 ;
        RECT 4.18 0.048 4.244 0.092 ;
        RECT 4.396 0.048 4.46 0.092 ;
        RECT 4.612 0.048 4.676 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.382 ;
      RECT 0.29 0.248 0.358 0.382 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.722 0.248 0.79 0.382 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.37 0.248 1.438 0.382 ;
      RECT 1.586 0.248 1.654 0.382 ;
      RECT 1.802 0.248 1.87 0.382 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 2.234 0.248 2.302 0.382 ;
      RECT 0.054 0.158 2.322 0.202 ;
      RECT 2.99 0.248 3.058 0.382 ;
      RECT 3.206 0.248 3.274 0.382 ;
      RECT 3.422 0.248 3.49 0.382 ;
      RECT 4.07 0.248 4.138 0.382 ;
      RECT 4.286 0.248 4.354 0.382 ;
      RECT 4.502 0.248 4.57 0.382 ;
      RECT 2.558 0.068 2.626 0.292 ;
      RECT 4.718 0.248 4.786 0.382 ;
    LAYER v0 ;
      RECT 4.718 0.158 4.786 0.202 ;
      RECT 4.61 0.518 4.678 0.562 ;
      RECT 4.502 0.158 4.57 0.202 ;
      RECT 4.394 0.518 4.462 0.562 ;
      RECT 4.286 0.158 4.354 0.202 ;
      RECT 4.178 0.518 4.246 0.562 ;
      RECT 4.07 0.158 4.138 0.202 ;
      RECT 3.962 0.518 4.03 0.562 ;
      RECT 3.854 0.158 3.922 0.202 ;
      RECT 3.746 0.518 3.814 0.562 ;
      RECT 3.638 0.178 3.706 0.222 ;
      RECT 3.53 0.518 3.598 0.562 ;
      RECT 3.422 0.068 3.49 0.112 ;
      RECT 3.314 0.518 3.382 0.562 ;
      RECT 3.206 0.068 3.274 0.112 ;
      RECT 3.098 0.518 3.166 0.562 ;
      RECT 2.99 0.068 3.058 0.112 ;
      RECT 2.882 0.518 2.95 0.562 ;
      RECT 2.774 0.068 2.842 0.112 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.558 0.178 2.626 0.222 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.428 2.342 0.472 ;
      RECT 2.342 0.428 2.41 0.562 ;
      RECT 2.41 0.518 4.698 0.562 ;
      RECT 2.626 0.068 3.638 0.112 ;
      RECT 3.638 0.068 3.706 0.382 ;
      RECT 3.706 0.338 3.962 0.382 ;
      RECT 3.746 0.158 3.962 0.202 ;
      RECT 3.962 0.158 4.03 0.382 ;
      RECT 4.03 0.158 4.806 0.202 ;
  END
END b15aoi022as1n48x5

MACRO b15aoi112as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi112as1n02x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.518 0.358 0.562 ;
        RECT 0.29 0.068 0.358 0.562 ;
        RECT 0.054 0.068 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.518 0.142 0.562 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.29 0.158 0.358 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.4505 0.466 0.4945 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.048 0.574 0.092 ;
    END
  END vssx
END b15aoi112as1n02x3

MACRO b15aoi112as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi112as1n02x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.48622225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.702 0.382 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.4955 0.142 0.5395 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.614 0.1355 0.682 0.1795 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.428 0.702 0.472 ;
    LAYER v0 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.428 0.466 0.472 ;
  END
END b15aoi112as1n02x5

MACRO b15aoi112as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi112as1n03x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68158725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.59037025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03978 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 2.66 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.81 0.112 ;
        RECT 0.398 0.158 0.682 0.202 ;
        RECT 0.614 0.068 0.682 0.202 ;
        RECT 0.398 0.068 0.466 0.202 ;
        RECT 0.182 0.068 0.466 0.112 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.182 0.148 0.25 0.192 ;
        RECT 0.722 0.068 0.79 0.112 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
      LAYER v0 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.938 0.406 1.006 0.45 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.29 0.408 0.358 0.452 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.29 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.358 0.518 0.506 0.562 ;
      RECT 0.506 0.338 0.574 0.562 ;
  END
END b15aoi112as1n03x5

MACRO b15aoi112as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi112as1n04x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.518 0.358 0.562 ;
        RECT 0.29 0.338 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.518 0.25 0.562 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.060247 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.84941175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.20333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 1.026 0.202 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.076 0.228 0.14 0.272 ;
        RECT 0.074 0.384 0.142 0.428 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.938 0.158 1.006 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 1.046 0.338 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
      LAYER v0 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 1.046 0.383 1.114 0.427 ;
        RECT 1.37 0.406 1.438 0.45 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 1.478 0.048 1.546 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.81 0.068 1.154 0.112 ;
    LAYER v0 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.614 0.4055 0.682 0.4495 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.384 0.25 0.428 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.248 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 1.154 0.068 1.222 0.202 ;
      RECT 1.222 0.158 1.546 0.202 ;
  END
END b15aoi112as1n04x5

MACRO b15aoi112as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi112as1n06x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.37925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7775925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.55518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.158 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.068 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.293 1.762 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 1.438 0.292 ;
        RECT 0.83 0.068 1.438 0.112 ;
        RECT 1.154 0.068 1.222 0.292 ;
        RECT 0.182 0.248 0.898 0.292 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.398 0.248 0.466 0.472 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.408 0.466 0.452 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.154 0.1605 1.222 0.2045 ;
        RECT 1.37 0.18 1.438 0.224 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
      LAYER v0 ;
        RECT 1.154 0.538 1.222 0.582 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.538 1.654 0.582 ;
        RECT 1.802 0.538 1.87 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.586 0.1805 1.654 0.2245 ;
        RECT 1.802 0.1805 1.87 0.2245 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.614 0.408 0.682 0.452 ;
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.518 1.046 0.562 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.114 0.428 1.87 0.472 ;
  END
END b15aoi112as1n06x5

MACRO b15aoi112as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi112as1n08x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63973075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.3194445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.70370375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.451389 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5875925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.158 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.382 ;
      LAYER v0 ;
        RECT 1.91 0.293 1.978 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.068 1.654 0.292 ;
        RECT 1.046 0.068 1.654 0.112 ;
        RECT 1.37 0.068 1.438 0.292 ;
        RECT 0.506 0.158 1.114 0.202 ;
        RECT 1.046 0.068 1.114 0.202 ;
        RECT 0.506 0.068 0.574 0.472 ;
        RECT 0.29 0.068 0.574 0.112 ;
        RECT 0.29 0.068 0.358 0.472 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.408 0.142 0.452 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.408 0.358 0.452 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.408 0.574 0.452 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.37 0.178 1.438 0.222 ;
        RECT 1.586 0.178 1.654 0.222 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
      LAYER v0 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.538 1.654 0.582 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.018 0.538 2.086 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 0.338 2.214 0.382 ;
        RECT 2.018 -0.022 2.086 0.382 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.802 0.178 1.87 0.222 ;
        RECT 2.018 0.158 2.086 0.202 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.518 1.134 0.562 ;
      RECT 0.702 0.428 2.214 0.472 ;
    LAYER v0 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.182 0.518 0.25 0.562 ;
  END
END b15aoi112as1n08x5

MACRO b15aoi122as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi122as1n02x3 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.113 0.898 0.157 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.113 0.682 0.157 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END e
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.42 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 0.898 0.562 ;
        RECT 0.506 0.338 0.898 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.203 0.574 0.247 ;
        RECT 0.83 0.423 0.898 0.467 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.2035 0.142 0.2475 ;
        RECT 0.722 0.2035 0.79 0.2475 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 0.702 0.472 ;
    LAYER v0 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.182 0.428 0.25 0.472 ;
  END
END b15aoi122as1n02x3

MACRO b15aoi122as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi122as1n02x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.760139 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.34685175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.203 0.79 0.247 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.466 0.112 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
    END
  END e
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.472 ;
        RECT 0.398 0.338 0.898 0.382 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.203 0.466 0.247 ;
        RECT 0.832 0.408 0.896 0.452 ;
        RECT 0.83 0.203 0.898 0.247 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.614 0.203 0.682 0.247 ;
        RECT 0.938 0.048 1.006 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.702 0.472 ;
      RECT 0.486 0.518 1.026 0.562 ;
    LAYER v0 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
  END
END b15aoi122as1n02x5

MACRO b15aoi122as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi122as1n04x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.914375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.6255555 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.088 0.79 0.132 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 1.546 0.472 ;
        RECT 0.938 0.338 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.6625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.04615375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.202 ;
      LAYER v0 ;
        RECT 1.478 0.138 1.546 0.182 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.769375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.35916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.088 0.682 0.132 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END e
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 1.33 0.292 ;
        RECT 0.29 0.338 0.79 0.382 ;
        RECT 0.722 0.248 0.79 0.382 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.1855 0.358 0.2295 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.154 0.248 1.222 0.292 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.506 0.1685 0.574 0.2125 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.37 0.138 1.438 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 1.438 0.472 ;
      RECT 0.702 0.518 1.546 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.428 0.25 0.472 ;
  END
END b15aoi122as1n04x5

MACRO b15aoi122as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi122as1n06x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.41708325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.83416675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.382 ;
      LAYER v0 ;
        RECT 1.91 0.138 1.978 0.182 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.458 0.382 ;
        RECT 1.046 0.158 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.97359475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.318 0.898 0.362 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.338 0.25 0.382 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.594 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END e
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07038 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.674 0.428 1.998 0.472 ;
        RECT 1.802 0.248 1.87 0.472 ;
        RECT 1.154 0.248 1.87 0.292 ;
        RECT 1.694 0.068 1.762 0.292 ;
        RECT 1.154 0.068 1.222 0.292 ;
        RECT 0.506 0.068 1.222 0.112 ;
        RECT 0.938 0.068 1.006 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.18 0.574 0.224 ;
        RECT 0.722 0.18 0.79 0.224 ;
        RECT 0.938 0.18 1.006 0.224 ;
        RECT 1.156 0.178 1.22 0.222 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 1.91 0.428 1.978 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.18 0.142 0.224 ;
        RECT 0.29 0.18 0.358 0.224 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 1.802 0.138 1.87 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 1.566 0.472 ;
      RECT 0.918 0.518 1.998 0.562 ;
    LAYER v0 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.428 0.25 0.472 ;
  END
END b15aoi122as1n06x5

MACRO b15aoi122as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi122as1n08x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 1.484375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.484375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.322 0.338 2.518 0.382 ;
        RECT 2.45 0.068 2.518 0.382 ;
      LAYER v0 ;
        RECT 2.342 0.338 2.41 0.382 ;
        RECT 2.45 0.088 2.518 0.132 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63658125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.338 1.89 0.382 ;
        RECT 1.37 0.158 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 1.33 0.382 ;
        RECT 0.938 0.158 1.006 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.378 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.898 0.382 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END e
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07956 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.428 2.518 0.472 ;
        RECT 2.126 0.068 2.194 0.472 ;
        RECT 1.478 0.248 2.194 0.292 ;
        RECT 1.478 0.068 1.546 0.292 ;
        RECT 0.614 0.068 1.546 0.112 ;
        RECT 1.262 0.068 1.33 0.292 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.614 0.068 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.18 0.682 0.224 ;
        RECT 0.83 0.18 0.898 0.224 ;
        RECT 1.262 0.166 1.33 0.21 ;
        RECT 1.478 0.166 1.546 0.21 ;
        RECT 2.126 0.346 2.194 0.39 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.342 0.428 2.41 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 1.91 0.138 1.978 0.182 ;
        RECT 2.234 0.138 2.302 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 1.998 0.472 ;
      RECT 1.134 0.518 2.538 0.562 ;
    LAYER v0 ;
      RECT 2.45 0.518 2.518 0.562 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.428 0.25 0.472 ;
  END
END b15aoi122as1n08x5

MACRO b15aoi222as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi222as1n02x3 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 1.026 0.202 ;
        RECT 0.83 0.158 0.898 0.472 ;
        RECT 0.614 0.068 0.682 0.202 ;
        RECT 0.182 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.83 0.408 0.898 0.452 ;
        RECT 0.938 0.158 1.006 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.682 0.472 ;
      RECT 0.29 0.518 1.026 0.562 ;
    LAYER v0 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
  END
END b15aoi222as1n02x3

MACRO b15aoi222as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi222as1n02x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 1.026 0.202 ;
        RECT 0.83 0.158 0.898 0.472 ;
        RECT 0.614 0.068 0.682 0.202 ;
        RECT 0.182 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.83 0.408 0.898 0.452 ;
        RECT 0.938 0.158 1.006 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.682 0.472 ;
      RECT 0.29 0.518 1.026 0.562 ;
    LAYER v0 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
  END
END b15aoi222as1n02x5

MACRO b15aoi222as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi222as1n04x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.338 1.458 0.382 ;
        RECT 1.262 0.158 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.23925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.162 0.338 0.358 0.382 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.23925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 2.491111 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.428 1.458 0.472 ;
        RECT 1.046 0.068 1.458 0.112 ;
        RECT 0.83 0.248 1.114 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.938 0.248 1.006 0.472 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.506 0.068 0.898 0.112 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.15 0.574 0.194 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.068 1.438 0.112 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.594 0.518 1.458 0.562 ;
    LAYER v0 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.358 0.898 0.402 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.83 0.472 ;
      RECT 0.83 0.338 0.898 0.472 ;
  END
END b15aoi222as1n04x5

MACRO b15aoi222as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi222as1n06x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.802 0.3155 1.87 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.1056945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.47425925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.158 1.33 0.292 ;
      LAYER v0 ;
        RECT 1.262 0.228 1.33 0.272 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.338 1.33 0.472 ;
        RECT 1.026 0.338 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 0.918 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.378 0.338 0.574 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.158 1.762 0.472 ;
        RECT 1.37 0.248 1.762 0.292 ;
        RECT 1.478 0.248 1.546 0.472 ;
        RECT 1.37 0.068 1.438 0.292 ;
        RECT 1.154 0.068 1.438 0.112 ;
        RECT 0.83 0.248 1.222 0.292 ;
        RECT 1.154 0.068 1.222 0.292 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.398 0.068 0.898 0.112 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.1805 0.466 0.2245 ;
        RECT 0.832 0.1685 0.896 0.2125 ;
        RECT 1.478 0.408 1.546 0.452 ;
        RECT 1.696 0.178 1.76 0.222 ;
        RECT 1.694 0.408 1.762 0.452 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 1.134 0.472 ;
      RECT 0.702 0.518 1.89 0.562 ;
    LAYER v0 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
  END
END b15aoi222as1n06x5

MACRO b15aoi222as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi222as1n08x5 0 0 ;
  SIZE 2.376 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.158 2.194 0.472 ;
      LAYER v0 ;
        RECT 2.126 0.3155 2.194 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88754625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2530065 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.478 0.273 1.546 0.317 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.134 0.338 1.438 0.382 ;
        RECT 1.37 0.248 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.026 0.382 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.486 0.338 0.682 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.068 2.302 0.472 ;
        RECT 2.018 0.068 2.302 0.112 ;
        RECT 2.018 0.068 2.086 0.472 ;
        RECT 1.586 0.248 2.086 0.292 ;
        RECT 1.802 0.248 1.87 0.472 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.262 0.158 1.654 0.202 ;
        RECT 0.938 0.248 1.33 0.292 ;
        RECT 1.262 0.158 1.33 0.292 ;
        RECT 0.938 0.068 1.006 0.292 ;
        RECT 0.506 0.068 1.006 0.112 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.191 0.574 0.235 ;
        RECT 0.722 0.191 0.79 0.235 ;
        RECT 0.94 0.1685 1.004 0.2125 ;
        RECT 1.586 0.408 1.654 0.452 ;
        RECT 1.802 0.408 1.87 0.452 ;
        RECT 2.018 0.408 2.086 0.452 ;
        RECT 2.018 0.1575 2.086 0.2015 ;
        RECT 2.234 0.408 2.302 0.452 ;
        RECT 2.234 0.203 2.302 0.247 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.41 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.41 0.022 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.802 0.138 1.87 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 1.546 0.472 ;
      RECT 0.81 0.518 2.302 0.562 ;
    LAYER v0 ;
      RECT 2.126 0.518 2.194 0.562 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
  END
END b15aoi222as1n08x5

MACRO b15aoi222as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15aoi222as1n12x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.54239325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.538 0.338 2.734 0.382 ;
        RECT 2.666 0.158 2.734 0.382 ;
      LAYER v0 ;
        RECT 2.558 0.338 2.626 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.54239325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.338 2.43 0.382 ;
        RECT 2.234 0.158 2.302 0.382 ;
      LAYER v0 ;
        RECT 2.342 0.338 2.41 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.54239325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.566 0.338 1.978 0.382 ;
        RECT 1.91 0.158 1.978 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.54239325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.35 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.54239325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.378 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.54239325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.594 0.338 0.79 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.428 2.95 0.472 ;
        RECT 2.882 0.248 2.95 0.472 ;
        RECT 2.774 0.248 2.95 0.292 ;
        RECT 2.774 0.068 2.842 0.292 ;
        RECT 2.558 0.068 2.842 0.112 ;
        RECT 2.558 0.068 2.626 0.202 ;
        RECT 2.018 0.068 2.086 0.472 ;
        RECT 1.802 0.068 2.086 0.112 ;
        RECT 1.262 0.248 1.87 0.292 ;
        RECT 1.802 0.068 1.87 0.292 ;
        RECT 1.262 0.068 1.33 0.292 ;
        RECT 0.614 0.068 1.33 0.112 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.614 0.068 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.191 0.682 0.235 ;
        RECT 0.83 0.191 0.898 0.235 ;
        RECT 1.046 0.191 1.114 0.235 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.56 0.138 2.624 0.182 ;
        RECT 2.558 0.428 2.626 0.472 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.774 0.1575 2.842 0.2015 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.342 0.138 2.41 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 1.89 0.472 ;
      RECT 1.026 0.518 2.97 0.562 ;
    LAYER v0 ;
      RECT 2.882 0.518 2.95 0.562 ;
      RECT 2.666 0.518 2.734 0.562 ;
      RECT 2.45 0.518 2.518 0.562 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
  END
END b15aoi222as1n12x5

MACRO b15bfm201as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfm201as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.383 0.466 0.427 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.383 0.358 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.383 0.142 0.427 ;
  END
END b15bfm201as1n02x5

MACRO b15bfm201as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfm201as1n04x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.988 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.988 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.428 0.358 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.158 0.358 0.202 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
    LAYER v0 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.383 0.142 0.427 ;
  END
END b15bfm201as1n04x5

MACRO b15bfm201as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfm201as1n08x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49822225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49822225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.432 0.466 0.476 ;
        RECT 0.398 0.163 0.466 0.207 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.432 0.358 0.476 ;
        RECT 0.506 0.432 0.574 0.476 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.163 0.358 0.207 ;
        RECT 0.506 0.163 0.574 0.207 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
    LAYER v0 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.386 0.142 0.43 ;
  END
END b15bfm201as1n08x5

MACRO b15bfm201as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfm201as1n16x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.398 0.338 0.682 0.382 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.113 0.466 0.157 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.614 0.113 0.682 0.157 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.113 0.358 0.157 ;
        RECT 0.506 0.113 0.574 0.157 ;
        RECT 0.722 0.113 0.79 0.157 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.074 0.113 0.142 0.157 ;
      RECT 0.076 0.498 0.14 0.542 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.248 0.358 0.472 ;
  END
END b15bfm201as1n16x5

MACRO b15bfm402as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfm402as1n02x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.383 1.006 0.427 ;
        RECT 0.938 0.203 1.006 0.247 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 0.83 0.383 0.898 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.2025 0.25 0.2465 ;
        RECT 0.83 0.203 0.898 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.614 0.158 0.682 0.472 ;
    LAYER v0 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.2025 0.682 0.2465 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.398 0.2025 0.466 0.2465 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.074 0.2025 0.142 0.2465 ;
      RECT 0.074 0.383 0.142 0.427 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.518 0.722 0.562 ;
      RECT 0.722 0.248 0.79 0.562 ;
  END
END b15bfm402as1n02x5

MACRO b15bfm402as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfm402as1n04x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.383 1.006 0.427 ;
        RECT 0.938 0.203 1.006 0.247 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 0.83 0.4725 0.898 0.5165 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.2025 0.25 0.2465 ;
        RECT 0.83 0.114 0.898 0.158 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.614 0.158 0.682 0.472 ;
    LAYER v0 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.2025 0.682 0.2465 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.398 0.2025 0.466 0.2465 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.074 0.2025 0.142 0.2465 ;
      RECT 0.074 0.383 0.142 0.427 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.518 0.722 0.562 ;
      RECT 0.722 0.248 0.79 0.562 ;
  END
END b15bfm402as1n04x5

MACRO b15bfm402as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfm402as1n08x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.383 1.006 0.427 ;
        RECT 0.938 0.203 1.006 0.247 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 0.83 0.4725 0.898 0.5165 ;
        RECT 1.046 0.4725 1.114 0.5165 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.2025 0.25 0.2465 ;
        RECT 0.83 0.114 0.898 0.158 ;
        RECT 1.046 0.114 1.114 0.158 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.614 0.158 0.682 0.472 ;
    LAYER v0 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.614 0.2025 0.682 0.2465 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.398 0.2025 0.466 0.2465 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.074 0.2025 0.142 0.2465 ;
      RECT 0.074 0.383 0.142 0.427 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.518 0.722 0.562 ;
      RECT 0.722 0.248 0.79 0.562 ;
  END
END b15bfm402as1n08x5

MACRO b15bfm402as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfm402as1n16x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.088 0.358 0.132 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.472 ;
        RECT 0.938 0.248 1.222 0.292 ;
        RECT 0.938 0.068 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.383 1.006 0.427 ;
        RECT 0.938 0.1285 1.006 0.1725 ;
        RECT 1.154 0.383 1.222 0.427 ;
        RECT 1.154 0.1285 1.222 0.1725 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.046 0.4725 1.114 0.5165 ;
        RECT 1.262 0.4725 1.33 0.5165 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.2025 0.25 0.2465 ;
        RECT 0.83 0.1285 0.898 0.1725 ;
        RECT 1.046 0.1285 1.114 0.1725 ;
        RECT 1.262 0.1285 1.33 0.1725 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.398 0.158 0.466 0.472 ;
    LAYER v0 ;
      RECT 0.83 0.293 0.898 0.337 ;
      RECT 0.614 0.186 0.682 0.23 ;
      RECT 0.614 0.3435 0.682 0.3875 ;
      RECT 0.398 0.2025 0.466 0.2465 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.074 0.2025 0.142 0.2465 ;
      RECT 0.074 0.383 0.142 0.427 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.428 0.83 0.472 ;
      RECT 0.83 0.248 0.898 0.472 ;
  END
END b15bfm402as1n16x5

MACRO b15bfn000as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n02x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.408 0.358 0.452 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
    LAYER v0 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.408 0.142 0.452 ;
  END
END b15bfn000as1n02x5

MACRO b15bfn000as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n03x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.383 0.358 0.427 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
    LAYER v0 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.383 0.142 0.427 ;
  END
END b15bfn000as1n03x5

MACRO b15bfn000as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n04x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.3155 0.25 0.3595 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.423 0.466 0.467 ;
        RECT 0.398 0.1305 0.466 0.1745 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.523 0.358 0.567 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.2305 0.358 0.2745 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
    LAYER v0 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.408 0.142 0.452 ;
  END
END b15bfn000as1n04x5

MACRO b15bfn000as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n06x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.383 0.358 0.427 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.383 0.466 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.1225 0.25 0.1665 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
    LAYER v0 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.383 0.142 0.427 ;
  END
END b15bfn000as1n06x5

MACRO b15bfn000as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n08x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.506 0.428 0.574 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.158 0.574 0.202 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
    LAYER v0 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.383 0.142 0.427 ;
  END
END b15bfn000as1n08x5

MACRO b15bfn000as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n12x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.398 0.338 0.682 0.382 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.4405 0.466 0.4845 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.4405 0.682 0.4845 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.074 0.1695 0.142 0.2135 ;
      RECT 0.076 0.498 0.14 0.542 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.248 0.358 0.472 ;
  END
END b15bfn000as1n12x5

MACRO b15bfn000as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n16x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.428 0.79 0.472 ;
        RECT 0.722 0.158 0.79 0.472 ;
        RECT 0.29 0.158 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.29 0.248 0.358 0.292 ;
      RECT 0.074 0.068 0.142 0.112 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.248 0.594 0.292 ;
  END
END b15bfn000as1n16x5

MACRO b15bfn000as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n24x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
        RECT 0.398 0.338 0.898 0.382 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.455 0.466 0.499 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.455 0.682 0.499 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 0.83 0.455 0.898 0.499 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.455 0.358 0.499 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.938 0.455 1.006 0.499 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.455 0.25 0.499 ;
  END
END b15bfn000as1n24x5

MACRO b15bfn000as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n32x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.29 0.158 1.222 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
        RECT 1.154 0.538 1.222 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.182 0.1365 0.25 0.1805 ;
      RECT 0.182 0.4385 0.25 0.4825 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.248 1.006 0.292 ;
  END
END b15bfn000as1n32x5

MACRO b15bfn000as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n48x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14688 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.472 ;
        RECT 0.398 0.158 1.762 0.202 ;
        RECT 1.478 0.158 1.546 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 1.478 0.048 1.546 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.292 0.228 0.356 0.272 ;
      RECT 0.074 0.428 0.142 0.472 ;
      RECT 0.076 0.228 0.14 0.272 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.358 0.338 1.438 0.382 ;
  END
END b15bfn000as1n48x5

MACRO b15bfn000as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n64x5 0 0 ;
  SIZE 2.376 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.19584 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.472 ;
        RECT 0.506 0.158 2.302 0.202 ;
        RECT 2.018 0.158 2.086 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.158 2.194 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.41 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.41 0.022 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.234 0.048 2.302 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.466 0.338 1.654 0.382 ;
  END
END b15bfn000as1n64x5

MACRO b15bfn000as1n80x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn000as1n80x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.52777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.52777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.428 2.842 0.472 ;
        RECT 2.774 0.158 2.842 0.472 ;
        RECT 0.614 0.158 2.842 0.202 ;
        RECT 2.558 0.158 2.626 0.472 ;
        RECT 2.342 0.158 2.41 0.472 ;
        RECT 2.126 0.158 2.194 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.158 2.734 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.776 0.538 2.84 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 1.478 0.048 1.546 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 1.91 0.048 1.978 0.092 ;
        RECT 2.126 0.048 2.194 0.092 ;
        RECT 2.342 0.048 2.41 0.092 ;
        RECT 2.558 0.048 2.626 0.092 ;
        RECT 2.774 0.048 2.842 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.508 0.228 0.572 0.272 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.292 0.228 0.356 0.272 ;
      RECT 0.074 0.428 0.142 0.472 ;
      RECT 0.076 0.228 0.14 0.272 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.358 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.338 2.086 0.382 ;
  END
END b15bfn000as1n80x5

MACRO b15bfn001as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn001as1n06x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.3155 0.25 0.3595 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.455 0.358 0.499 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.455 0.466 0.499 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.455 0.142 0.499 ;
  END
END b15bfn001as1n06x5

MACRO b15bfn001as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn001as1n08x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.473 0.466 0.517 ;
        RECT 0.398 0.153 0.466 0.197 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.506 0.473 0.574 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.153 0.574 0.197 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.074 0.24 0.142 0.284 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.472 ;
  END
END b15bfn001as1n08x5

MACRO b15bfn001as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn001as1n12x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.398 0.338 0.682 0.382 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.4485 0.682 0.4925 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.448 0.25 0.492 ;
  END
END b15bfn001as1n12x5

MACRO b15bfn001as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn001as1n16x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.398 0.338 0.682 0.382 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.429 0.466 0.473 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.429 0.682 0.473 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.428 0.824 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.722 0.248 0.79 0.472 ;
    LAYER v1 ;
      RECT 0.726 0.428 0.786 0.472 ;
      RECT 0.186 0.428 0.246 0.472 ;
    LAYER v0 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.429 0.25 0.473 ;
  END
END b15bfn001as1n16x5

MACRO b15bfn001as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn001as1n24x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.79 0.472 ;
        RECT 0.074 0.248 0.682 0.292 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.398 0.068 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.046 0.44 1.114 0.484 ;
      RECT 1.048 0.228 1.112 0.272 ;
      RECT 0.83 0.44 0.898 0.484 ;
      RECT 0.832 0.228 0.896 0.272 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.29 0.338 0.358 0.382 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.83 0.382 ;
      RECT 0.83 0.158 0.898 0.562 ;
      RECT 0.898 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.562 ;
  END
END b15bfn001as1n24x5

MACRO b15bfn001as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn001as1n32x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 0.506 0.158 1.438 0.202 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.398 0.452 0.466 0.496 ;
      RECT 0.4 0.228 0.464 0.272 ;
      RECT 0.182 0.452 0.25 0.496 ;
      RECT 0.184 0.228 0.248 0.272 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.338 1.33 0.382 ;
  END
END b15bfn001as1n32x5

MACRO b15bfn001as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn001as1n48x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.574 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14688 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.472 ;
        RECT 0.722 0.158 2.086 0.202 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 0.83 0.338 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.832 0.358 0.896 0.402 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.074 0.428 0.722 0.472 ;
      RECT 0.682 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 0.79 0.248 1.762 0.292 ;
  END
END b15bfn001as1n48x5

MACRO b15bfn001as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn001as1n64x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.898 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.19584 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.428 2.734 0.472 ;
        RECT 2.666 0.158 2.734 0.472 ;
        RECT 0.938 0.158 2.734 0.202 ;
        RECT 2.45 0.158 2.518 0.472 ;
        RECT 2.234 0.158 2.302 0.472 ;
        RECT 1.046 0.338 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.048 0.358 1.112 0.402 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.428 2.626 0.472 ;
        RECT 2.558 0.158 2.626 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.832 0.178 0.896 0.222 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.158 0.898 0.292 ;
      RECT 0.074 0.428 0.938 0.472 ;
      RECT 0.898 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.006 0.248 2.194 0.292 ;
  END
END b15bfn001as1n64x5

MACRO b15bfn001as1n80x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15bfn001as1n80x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5795 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5795 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 1.006 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 0.614 0.338 0.682 0.382 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.428 3.382 0.472 ;
        RECT 3.314 0.158 3.382 0.472 ;
        RECT 1.154 0.158 3.382 0.202 ;
        RECT 3.098 0.158 3.166 0.472 ;
        RECT 2.882 0.158 2.95 0.472 ;
        RECT 2.666 0.158 2.734 0.472 ;
        RECT 1.262 0.338 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.264 0.358 1.328 0.402 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.428 2.626 0.472 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.774 0.158 2.842 0.202 ;
        RECT 2.99 0.428 3.058 0.472 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.206 0.158 3.274 0.202 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.316 0.538 3.38 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.316 0.048 3.38 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 1.048 0.178 1.112 0.222 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.832 0.178 0.896 0.222 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.158 0.898 0.292 ;
      RECT 0.898 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 0.074 0.428 1.154 0.472 ;
      RECT 1.114 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.222 0.248 2.626 0.292 ;
  END
END b15bfn001as1n80x5

MACRO b15cand02as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cand02as1n02x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2455555 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.83037025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.616 0.113 0.68 0.157 ;
        RECT 0.614 0.473 0.682 0.517 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.398 0.473 0.466 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.398 0.048 0.466 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.29 0.473 0.358 0.517 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.358 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.472 ;
  END
END b15cand02as1n02x5

MACRO b15cand02as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cand02as1n03x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2455555 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.83037025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.616 0.113 0.68 0.157 ;
        RECT 0.614 0.473 0.682 0.517 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.398 0.473 0.466 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.4 0.048 0.464 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.29 0.473 0.358 0.517 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.358 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.472 ;
  END
END b15cand02as1n03x5

MACRO b15cand02as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cand02as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.408 0.574 0.452 ;
        RECT 0.506 0.113 0.574 0.157 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4735 0.142 0.5175 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.113 0.466 0.157 ;
        RECT 0.614 0.113 0.682 0.157 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.398 0.3155 0.466 0.3595 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.113 0.25 0.157 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.428 0.398 0.472 ;
      RECT 0.398 0.248 0.466 0.472 ;
  END
END b15cand02as1n04x5

MACRO b15cand02as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cand02as1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.64666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03366 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.562 ;
        RECT 0.506 0.248 0.79 0.292 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.4505 0.574 0.4945 ;
        RECT 0.506 0.09 0.574 0.134 ;
        RECT 0.722 0.4505 0.79 0.4945 ;
        RECT 0.722 0.09 0.79 0.134 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4735 0.142 0.5175 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.614 0.4505 0.682 0.4945 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.09 0.466 0.134 ;
        RECT 0.614 0.09 0.682 0.134 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.398 0.3155 0.466 0.3595 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.113 0.25 0.157 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.428 0.398 0.472 ;
      RECT 0.398 0.248 0.466 0.472 ;
  END
END b15cand02as1n08x5

MACRO b15cand02as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cand02as1n12x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.34685175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.173426 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.383 0.466 0.427 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
        RECT 0.614 0.338 0.898 0.382 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.473 0.682 0.517 ;
        RECT 0.614 0.113 0.682 0.157 ;
        RECT 0.83 0.473 0.898 0.517 ;
        RECT 0.83 0.113 0.898 0.157 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.506 0.473 0.574 0.517 ;
        RECT 0.722 0.473 0.79 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.113 0.574 0.157 ;
        RECT 0.722 0.113 0.79 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 0.466 0.112 ;
    LAYER v0 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.29 0.473 0.358 0.517 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.358 0.248 0.574 0.292 ;
  END
END b15cand02as1n12x5

MACRO b15cand02as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cand02as1n16x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.2705 0.466 0.3145 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06426 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
        RECT 0.614 0.248 1.114 0.292 ;
        RECT 0.83 0.068 0.898 0.562 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.473 0.682 0.517 ;
        RECT 0.614 0.113 0.682 0.157 ;
        RECT 0.83 0.473 0.898 0.517 ;
        RECT 0.83 0.113 0.898 0.157 ;
        RECT 1.046 0.473 1.114 0.517 ;
        RECT 1.046 0.113 1.114 0.157 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.722 0.473 0.79 0.517 ;
        RECT 0.938 0.473 1.006 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.113 0.574 0.157 ;
        RECT 0.722 0.113 0.79 0.157 ;
        RECT 0.938 0.113 1.006 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 0.466 0.112 ;
    LAYER v0 ;
      RECT 0.506 0.2705 0.574 0.3145 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.428 0.506 0.472 ;
      RECT 0.506 0.248 0.574 0.472 ;
  END
END b15cand02as1n16x5

MACRO b15cand02as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cand02as1n24x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 1.79931625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 1.79931625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.158 0.79 0.202 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09486 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.428 1.458 0.472 ;
        RECT 1.262 0.068 1.33 0.472 ;
        RECT 0.83 0.248 1.33 0.292 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.506 -0.022 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 0.29 0.472 ;
      RECT 1.37 0.158 1.438 0.382 ;
    LAYER v0 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.508 0.408 0.572 0.452 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.054 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.574 0.338 1.222 0.382 ;
  END
END b15cand02as1n24x5

MACRO b15cand02as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cand02as1n32x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.881389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0189 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6715345 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9963195 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9963195 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.428 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.4505 0.682 0.4945 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11628 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.428 1.998 0.472 ;
        RECT 0.938 0.158 1.998 0.202 ;
        RECT 1.802 0.158 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.428 0.506 0.472 ;
      RECT 1.91 0.248 1.978 0.382 ;
    LAYER v0 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 0.83 0.1575 0.898 0.2015 ;
      RECT 0.83 0.45 0.898 0.494 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 0.074 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.338 0.938 0.382 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.006 0.248 1.762 0.292 ;
  END
END b15cand02as1n32x5

MACRO b15cand02as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cand02as1n64x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41377775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.574 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41477125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.898 0.382 ;
        RECT 0.83 0.248 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.21726 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.428 2.97 0.472 ;
        RECT 1.262 0.158 2.97 0.202 ;
        RECT 2.774 0.158 2.842 0.472 ;
        RECT 2.558 0.158 2.626 0.472 ;
        RECT 2.342 0.158 2.41 0.472 ;
        RECT 2.126 0.158 2.194 0.472 ;
        RECT 1.91 0.158 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 2.882 0.158 2.95 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.776 0.538 2.84 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.472 ;
      RECT 2.882 0.248 2.95 0.382 ;
    LAYER v0 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.158 1.006 0.202 ;
      RECT 0.142 0.248 0.182 0.292 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.142 0.428 0.938 0.472 ;
      RECT 0.938 0.338 1.006 0.472 ;
      RECT 1.006 0.338 1.87 0.382 ;
  END
END b15cand02as1n64x5

MACRO b15cbf000as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.383 0.466 0.427 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.383 0.358 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.074 0.216 0.142 0.26 ;
      RECT 0.074 0.3925 0.142 0.4365 ;
  END
END b15cbf000as1n02x5

MACRO b15cbf000as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n03x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.394 0.466 0.438 ;
        RECT 0.398 0.1965 0.466 0.2405 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.113 0.358 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
    LAYER v0 ;
      RECT 0.182 0.1935 0.25 0.2375 ;
      RECT 0.182 0.3875 0.25 0.4315 ;
  END
END b15cbf000as1n03x5

MACRO b15cbf000as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n04x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.4565 0.574 0.5005 ;
        RECT 0.506 0.1585 0.574 0.2025 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.473 0.358 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.398 0.293 0.466 0.337 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.162 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.382 ;
  END
END b15cbf000as1n04x5

MACRO b15cbf000as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n06x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.4225 0.466 0.4665 ;
        RECT 0.398 0.1935 0.466 0.2375 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.4225 0.574 0.4665 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.113 0.358 0.157 ;
        RECT 0.506 0.1935 0.574 0.2375 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
    LAYER v0 ;
      RECT 0.182 0.1945 0.25 0.2385 ;
      RECT 0.182 0.3845 0.25 0.4285 ;
  END
END b15cbf000as1n06x5

MACRO b15cbf000as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.408 0.574 0.452 ;
        RECT 0.506 0.184 0.574 0.228 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.398 0.293 0.466 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.398 0.472 ;
      RECT 0.398 0.158 0.466 0.472 ;
  END
END b15cbf000as1n08x5

MACRO b15cbf000as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n12x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.562 ;
        RECT 0.506 0.248 0.79 0.292 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.4505 0.574 0.4945 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.4505 0.79 0.4945 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.614 0.338 0.682 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.493 0.358 0.537 ;
        RECT 0.614 0.4505 0.682 0.4945 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.398 0.293 0.466 0.337 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.562 ;
  END
END b15cbf000as1n12x5

MACRO b15cbf000as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n16x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05814 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.562 ;
        RECT 0.506 0.248 0.79 0.292 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.83 0.448 0.898 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.398 0.293 0.466 0.337 ;
      RECT 0.182 0.423 0.25 0.467 ;
      RECT 0.184 0.088 0.248 0.132 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.382 ;
  END
END b15cbf000as1n16x5

MACRO b15cbf000as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n24x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.428 1.134 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.29 0.158 1.006 0.202 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.046 0.248 1.114 0.382 ;
    LAYER v0 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.682 0.382 ;
  END
END b15cbf000as1n24x5

MACRO b15cbf000as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n32x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1071 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.29 0.158 1.222 0.202 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.29 0.248 0.358 0.292 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.248 0.898 0.292 ;
  END
END b15cbf000as1n32x5

MACRO b15cbf000as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n48x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16524 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 1.998 0.472 ;
        RECT 0.506 0.158 1.998 0.202 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.91 0.248 1.978 0.382 ;
    LAYER v0 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.134 0.466 0.178 ;
      RECT 0.398 0.43 0.466 0.474 ;
      RECT 0.074 0.248 0.142 0.292 ;
    LAYER m1 ;
      RECT 0.054 0.248 0.398 0.292 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.466 0.248 1.114 0.292 ;
  END
END b15cbf000as1n48x5

MACRO b15cbf000as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n64x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 2.43 0.472 ;
        RECT 0.506 0.158 2.43 0.202 ;
        RECT 2.234 0.158 2.302 0.472 ;
        RECT 2.018 0.158 2.086 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 1.586 0.158 1.654 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.342 0.158 2.41 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 2.342 0.248 2.41 0.382 ;
    LAYER v0 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.466 0.248 1.046 0.292 ;
      RECT 1.046 0.248 1.114 0.382 ;
      RECT 1.114 0.338 1.458 0.382 ;
  END
END b15cbf000as1n64x5

MACRO b15cbf000as1n80x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf000as1n80x5 0 0 ;
  SIZE 3.132 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.589 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.589 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.486 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.26928 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.135 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.428 3.058 0.472 ;
        RECT 2.99 0.158 3.058 0.472 ;
        RECT 1.046 0.158 3.058 0.202 ;
        RECT 2.342 0.158 2.41 0.472 ;
        RECT 2.126 0.158 2.194 0.472 ;
        RECT 1.046 0.158 1.114 0.472 ;
        RECT 0.83 0.248 1.114 0.292 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 2.882 0.158 2.95 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.166 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.776 0.538 2.84 0.582 ;
        RECT 2.992 0.538 3.056 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.166 0.022 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.154 0.338 1.586 0.382 ;
      RECT 2.45 0.248 2.862 0.292 ;
    LAYER v0 ;
      RECT 2.774 0.248 2.842 0.292 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.398 0.472 ;
      RECT 0.398 0.338 0.466 0.472 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.054 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 0.682 0.338 1.006 0.382 ;
      RECT 1.586 0.248 1.654 0.382 ;
      RECT 1.654 0.248 2.086 0.292 ;
  END
END b15cbf000as1n80x5

MACRO b15cbf034as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf034as1n02x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.2705 0.25 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 1.91 0.113 1.978 0.157 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.33 0.472 ;
        RECT 0.29 0.428 0.574 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.694 0.383 1.762 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 0.614 0.518 1.114 0.562 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.614 -0.022 0.682 0.562 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.113 0.466 0.157 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.938 0.518 1.006 0.562 ;
        RECT 1.046 0.168 1.114 0.212 ;
        RECT 1.694 0.113 1.762 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 1.478 0.068 1.546 0.472 ;
    LAYER v0 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.1475 1.546 0.1915 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.79 0.338 1.37 0.382 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.546 0.248 1.87 0.292 ;
  END
END b15cbf034as1n02x5

MACRO b15cbf034as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf034as1n03x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.2705 0.25 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 1.91 0.113 1.978 0.157 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.33 0.472 ;
        RECT 0.29 0.428 0.574 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.694 0.383 1.762 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 0.614 0.518 1.114 0.562 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.614 -0.022 0.682 0.562 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.113 0.466 0.157 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.938 0.518 1.006 0.562 ;
        RECT 1.046 0.168 1.114 0.212 ;
        RECT 1.694 0.113 1.762 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 1.478 0.068 1.546 0.472 ;
    LAYER v0 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.1475 1.546 0.1915 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.79 0.338 1.37 0.382 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.546 0.248 1.87 0.292 ;
  END
END b15cbf034as1n03x5

MACRO b15cbf034as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf034as1n04x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.2705 0.25 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 1.91 0.113 1.978 0.157 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.33 0.472 ;
        RECT 0.29 0.428 0.574 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.694 0.383 1.762 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 0.614 0.518 1.114 0.562 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.614 -0.022 0.682 0.562 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.113 0.466 0.157 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.938 0.518 1.006 0.562 ;
        RECT 1.046 0.168 1.114 0.212 ;
        RECT 1.694 0.113 1.762 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 1.478 0.068 1.546 0.472 ;
    LAYER v0 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.478 0.1475 1.546 0.1915 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.79 0.338 1.37 0.382 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.546 0.248 1.762 0.292 ;
  END
END b15cbf034as1n04x5

MACRO b15cbf034as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf034as1n08x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.2705 0.25 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.113 1.978 0.157 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.33 0.472 ;
        RECT 0.29 0.428 0.574 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.694 0.383 1.762 0.427 ;
        RECT 2.018 0.428 2.086 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 0.614 0.518 1.114 0.562 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.614 -0.022 0.682 0.562 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.113 0.466 0.157 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.938 0.518 1.006 0.562 ;
        RECT 1.046 0.168 1.114 0.212 ;
        RECT 1.694 0.113 1.762 0.157 ;
        RECT 2.018 0.113 2.086 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 1.478 0.068 1.546 0.472 ;
    LAYER v0 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.478 0.1475 1.546 0.1915 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.79 0.338 1.37 0.382 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.546 0.248 1.762 0.292 ;
  END
END b15cbf034as1n08x5

MACRO b15cbf034as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf034as1n12x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.2705 0.25 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.562 ;
        RECT 1.91 0.248 2.194 0.292 ;
        RECT 1.91 0.068 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.113 1.978 0.157 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.113 2.194 0.157 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.33 0.472 ;
        RECT 0.29 0.428 0.574 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 2.018 0.428 2.086 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 0.614 0.518 1.114 0.562 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.614 -0.022 0.682 0.562 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.113 0.466 0.157 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.938 0.518 1.006 0.562 ;
        RECT 1.046 0.168 1.114 0.212 ;
        RECT 1.694 0.113 1.762 0.157 ;
        RECT 2.018 0.113 2.086 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 1.478 0.068 1.546 0.472 ;
    LAYER v0 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.478 0.1475 1.546 0.1915 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.79 0.338 1.37 0.382 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.546 0.248 1.762 0.292 ;
  END
END b15cbf034as1n12x5

MACRO b15cbf034as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf034as1n16x5 0 0 ;
  SIZE 2.376 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.2705 0.25 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06426 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.562 ;
        RECT 1.694 0.248 2.194 0.292 ;
        RECT 1.91 0.068 1.978 0.562 ;
        RECT 1.694 0.068 1.762 0.562 ;
      LAYER v0 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.113 1.762 0.157 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.113 1.978 0.157 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.113 2.194 0.157 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.41 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 2.018 0.338 2.086 0.652 ;
        RECT 1.802 0.338 1.87 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.33 0.472 ;
        RECT 0.29 0.428 0.574 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.234 0.428 2.302 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.41 0.022 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 0.614 0.518 1.114 0.562 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.614 -0.022 0.682 0.562 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.113 0.466 0.157 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.938 0.518 1.006 0.562 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.802 0.113 1.87 0.157 ;
        RECT 2.018 0.113 2.086 0.157 ;
        RECT 2.234 0.113 2.302 0.157 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 0.83 0.158 1.33 0.202 ;
      RECT 1.478 0.068 1.546 0.472 ;
    LAYER v0 ;
      RECT 1.478 0.1475 1.546 0.1915 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.79 0.338 1.37 0.382 ;
      RECT 1.37 0.158 1.438 0.382 ;
  END
END b15cbf034as1n16x5

MACRO b15cbf034as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf034as1n24x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.2705 0.25 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07956 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.338 2.626 0.382 ;
        RECT 2.558 0.158 2.626 0.382 ;
        RECT 1.91 0.158 2.626 0.202 ;
        RECT 2.45 0.338 2.518 0.562 ;
        RECT 2.342 0.158 2.41 0.382 ;
        RECT 2.234 0.338 2.302 0.562 ;
        RECT 2.126 0.158 2.194 0.382 ;
        RECT 2.018 0.338 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.45 0.158 2.518 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.29 0.428 0.574 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 0.398 0.518 1.114 0.562 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.614 -0.022 0.682 0.562 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.113 0.466 0.157 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 0.938 0.518 1.006 0.562 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.262 0.428 1.586 0.472 ;
    LAYER v0 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.156 0.158 1.22 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.79 0.338 1.262 0.382 ;
      RECT 1.262 0.248 1.33 0.382 ;
      RECT 1.33 0.248 1.546 0.292 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.068 1.654 0.112 ;
      RECT 1.262 0.158 1.586 0.202 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.654 0.248 2.086 0.292 ;
  END
END b15cbf034as1n24x5

MACRO b15cbf034as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf034as1n32x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.2705 0.25 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.10404 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.338 2.842 0.382 ;
        RECT 2.774 0.158 2.842 0.382 ;
        RECT 1.91 0.158 2.842 0.202 ;
        RECT 2.666 0.338 2.734 0.562 ;
        RECT 2.558 0.158 2.626 0.382 ;
        RECT 2.45 0.338 2.518 0.562 ;
        RECT 2.342 0.158 2.41 0.382 ;
        RECT 2.234 0.338 2.302 0.562 ;
        RECT 2.126 0.158 2.194 0.382 ;
        RECT 2.018 0.338 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.666 0.158 2.734 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.338 1.978 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.29 0.428 0.574 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 0.398 0.518 1.114 0.562 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.614 -0.022 0.682 0.562 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.113 0.466 0.157 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 0.938 0.518 1.006 0.562 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.262 0.428 1.586 0.472 ;
    LAYER v0 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.156 0.158 1.22 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.79 0.338 1.262 0.382 ;
      RECT 1.262 0.248 1.33 0.382 ;
      RECT 1.33 0.248 1.546 0.292 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.068 1.654 0.112 ;
      RECT 1.262 0.158 1.586 0.202 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.654 0.248 2.086 0.292 ;
  END
END b15cbf034as1n32x5

MACRO b15cbf034as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cbf034as1n64x5 0 0 ;
  SIZE 4.536 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.2705 0.25 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.428 4.482 0.472 ;
        RECT 2.558 0.158 4.482 0.202 ;
        RECT 4.286 0.158 4.354 0.472 ;
        RECT 4.07 0.158 4.138 0.472 ;
        RECT 3.854 0.158 3.922 0.472 ;
        RECT 3.638 0.158 3.706 0.472 ;
        RECT 3.422 0.158 3.49 0.472 ;
        RECT 3.206 0.158 3.274 0.472 ;
      LAYER v0 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 2.882 0.158 2.95 0.202 ;
        RECT 3.098 0.428 3.166 0.472 ;
        RECT 3.098 0.158 3.166 0.202 ;
        RECT 3.314 0.428 3.382 0.472 ;
        RECT 3.314 0.158 3.382 0.202 ;
        RECT 3.53 0.428 3.598 0.472 ;
        RECT 3.53 0.158 3.598 0.202 ;
        RECT 3.746 0.428 3.814 0.472 ;
        RECT 3.746 0.158 3.814 0.202 ;
        RECT 3.962 0.428 4.03 0.472 ;
        RECT 3.962 0.158 4.03 0.202 ;
        RECT 4.178 0.428 4.246 0.472 ;
        RECT 4.178 0.158 4.246 0.202 ;
        RECT 4.394 0.428 4.462 0.472 ;
        RECT 4.394 0.158 4.462 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.57 0.652 ;
        RECT 4.286 0.518 4.354 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.854 0.518 3.922 0.652 ;
        RECT 3.638 0.518 3.706 0.652 ;
        RECT 3.422 0.518 3.49 0.652 ;
        RECT 3.206 0.518 3.274 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.29 0.428 0.574 0.472 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.776 0.538 2.84 0.582 ;
        RECT 2.992 0.538 3.056 0.582 ;
        RECT 3.208 0.538 3.272 0.582 ;
        RECT 3.424 0.538 3.488 0.582 ;
        RECT 3.64 0.538 3.704 0.582 ;
        RECT 3.856 0.538 3.92 0.582 ;
        RECT 4.072 0.538 4.136 0.582 ;
        RECT 4.288 0.538 4.352 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.57 0.022 ;
        RECT 4.286 -0.022 4.354 0.112 ;
        RECT 4.07 -0.022 4.138 0.112 ;
        RECT 3.854 -0.022 3.922 0.112 ;
        RECT 3.638 -0.022 3.706 0.112 ;
        RECT 3.422 -0.022 3.49 0.112 ;
        RECT 3.206 -0.022 3.274 0.112 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.486 0.518 1.33 0.562 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.83 -0.022 0.898 0.562 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.113 0.466 0.157 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 0.83 0.113 0.898 0.157 ;
        RECT 1.046 0.518 1.114 0.562 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
        RECT 3.208 0.048 3.272 0.092 ;
        RECT 3.424 0.048 3.488 0.092 ;
        RECT 3.64 0.048 3.704 0.092 ;
        RECT 3.856 0.048 3.92 0.092 ;
        RECT 4.072 0.048 4.136 0.092 ;
        RECT 4.286 0.048 4.354 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 0.938 0.158 2.41 0.202 ;
      RECT 4.394 0.248 4.462 0.382 ;
    LAYER v0 ;
      RECT 2.99 0.338 3.058 0.382 ;
      RECT 2.774 0.338 2.842 0.382 ;
      RECT 2.558 0.338 2.626 0.382 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.694 0.42 1.762 0.464 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.402 1.006 0.446 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.402 0.682 0.446 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 1.006 0.248 2.302 0.292 ;
      RECT 1.762 0.338 2.45 0.382 ;
      RECT 1.586 0.068 2.45 0.112 ;
      RECT 2.45 0.068 2.518 0.382 ;
      RECT 2.518 0.338 3.166 0.382 ;
  END
END b15cbf034as1n64x5

MACRO b15cinv00as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.383 0.358 0.427 ;
        RECT 0.29 0.178 0.358 0.222 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.178 0.25 0.222 ;
    END
  END vssx
END b15cinv00as1n02x5

MACRO b15cinv00as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n03x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.64666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.64666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3995 0.358 0.4435 ;
        RECT 0.29 0.1285 0.358 0.1725 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.3995 0.25 0.4435 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.1285 0.25 0.1725 ;
    END
  END vssx
END b15cinv00as1n03x5

MACRO b15cinv00as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n04x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.29 0.113 0.358 0.157 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
    END
  END vssx
END b15cinv00as1n04x5

MACRO b15cinv00as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n06x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.20333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.20333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.408 0.358 0.452 ;
        RECT 0.29 0.178 0.358 0.222 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.398 0.408 0.466 0.452 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.095 0.25 0.139 ;
        RECT 0.398 0.095 0.466 0.139 ;
    END
  END vssx
END b15cinv00as1n06x5

MACRO b15cinv00as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n08x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.9025 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.9025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.29 0.113 0.358 0.157 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.398 0.113 0.466 0.157 ;
    END
  END vssx
END b15cinv00as1n08x5

MACRO b15cinv00as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n12x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
        RECT 0.29 0.248 0.574 0.292 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.292 0.178 0.356 0.222 ;
        RECT 0.29 0.384 0.358 0.428 ;
        RECT 0.508 0.178 0.572 0.222 ;
        RECT 0.506 0.384 0.574 0.428 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4755 0.25 0.5195 ;
        RECT 0.398 0.4755 0.466 0.5195 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
    END
  END vssx
END b15cinv00as1n12x5

MACRO b15cinv00as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n16x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0333 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63675675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.73625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05814 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.702 0.472 ;
        RECT 0.506 0.158 0.574 0.472 ;
        RECT 0.074 0.158 0.574 0.202 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.382 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.616 0.113 0.68 0.157 ;
    END
  END vssx
END b15cinv00as1n16x5

MACRO b15cinv00as1n20x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n20x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.48081625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.589 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07956 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
        RECT 0.182 0.338 0.682 0.382 ;
        RECT 0.054 0.158 0.682 0.202 ;
        RECT 0.398 0.158 0.466 0.472 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.184 0.408 0.248 0.452 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.4 0.408 0.464 0.452 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.616 0.408 0.68 0.452 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
    END
  END vssx
END b15cinv00as1n20x5

MACRO b15cinv00as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n24x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0513 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.486 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07956 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.79 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
        RECT 0.074 0.158 0.79 0.202 ;
        RECT 0.614 0.338 0.682 0.562 ;
        RECT 0.398 0.338 0.466 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
END b15cinv00as1n24x5

MACRO b15cinv00as1n28x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n28x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.50276925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0504 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5835715 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.486 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.10404 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.472 ;
        RECT 0.182 0.338 0.898 0.382 ;
        RECT 0.054 0.158 0.898 0.202 ;
        RECT 0.614 0.158 0.682 0.472 ;
        RECT 0.398 0.338 0.466 0.472 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.184 0.408 0.248 0.452 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.4 0.408 0.464 0.452 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.616 0.408 0.68 0.452 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.832 0.408 0.896 0.452 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
    END
  END vssx
END b15cinv00as1n28x5

MACRO b15cinv00as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n32x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0657 LAYER m1 ;
      ANTENNAMAXAREACAR 0.510137 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.682 0.292 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.10404 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.006 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.074 0.158 1.006 0.202 ;
        RECT 0.722 0.158 0.79 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
END b15cinv00as1n32x5

MACRO b15cinv00as1n40x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n40x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0801 LAYER m1 ;
      ANTENNAMAXAREACAR 0.520899 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5795 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.594 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.12852 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 1.222 0.382 ;
        RECT 1.154 0.158 1.222 0.382 ;
        RECT 0.074 0.158 1.222 0.202 ;
        RECT 1.046 0.338 1.114 0.472 ;
        RECT 0.938 0.158 1.006 0.382 ;
        RECT 0.83 0.338 0.898 0.472 ;
        RECT 0.722 0.158 0.79 0.382 ;
        RECT 0.614 0.338 0.682 0.472 ;
        RECT 0.398 0.338 0.466 0.472 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.184 0.408 0.248 0.452 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.4 0.408 0.464 0.452 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.616 0.408 0.68 0.452 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.832 0.408 0.896 0.452 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.048 0.408 1.112 0.452 ;
        RECT 1.046 0.158 1.114 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
END b15cinv00as1n40x5

MACRO b15cinv00as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n48x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0945 LAYER m1 ;
      ANTENNAMAXAREACAR 0.528381 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57791675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.81 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 0.074 0.158 1.438 0.202 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.184 0.358 0.248 0.402 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
END b15cinv00as1n48x5

MACRO b15cinv00as1n56x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n56x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57633325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.1008 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 1.33 0.382 ;
        RECT 0.83 0.248 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.782 0.472 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 0.074 0.158 1.654 0.202 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.382 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.696 0.132 1.76 0.176 ;
    END
  END vssx
END b15cinv00as1n56x5

MACRO b15cinv00as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n64x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.1224 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57558825 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.1152 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6115625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 1.546 0.382 ;
        RECT 1.046 0.248 1.114 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.20808 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.998 0.472 ;
        RECT 1.802 0.068 1.87 0.472 ;
        RECT 1.586 0.248 1.87 0.292 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 0.074 0.158 1.654 0.202 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.802 0.113 1.87 0.157 ;
        RECT 1.91 0.428 1.978 0.472 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.91 -0.022 1.978 0.382 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.694 0.113 1.762 0.157 ;
        RECT 1.91 0.113 1.978 0.157 ;
    END
  END vssx
END b15cinv00as1n64x5

MACRO b15cinv00as1n80x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cinv00as1n80x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.1584 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57431825 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.1449 LAYER m1 ;
      ANTENNAMAXAREACAR 0.627826 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 1.762 0.292 ;
        RECT 1.262 0.248 1.33 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.586 0.248 1.654 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.25704 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 2.518 0.472 ;
        RECT 2.45 0.158 2.518 0.472 ;
        RECT 0.074 0.158 2.518 0.202 ;
        RECT 2.234 0.158 2.302 0.472 ;
        RECT 2.018 0.158 2.086 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 0.506 0.158 0.574 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.342 0.158 2.41 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
    END
  END vssx
END b15cinv00as1n80x5

MACRO b15clb0a2as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n02x3 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.383 0.682 0.427 ;
        RECT 0.614 0.203 0.682 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.113 0.358 0.157 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.203 0.142 0.247 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.142 0.428 0.506 0.472 ;
      RECT 0.506 0.248 0.574 0.472 ;
  END
END b15clb0a2as1n02x3

MACRO b15clb0a2as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n02x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.478 0.682 0.522 ;
        RECT 0.614 0.203 0.682 0.247 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.398 0.048 0.466 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.29 0.453 0.358 0.497 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.358 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.472 ;
  END
END b15clb0a2as1n02x5

MACRO b15clb0a2as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n03x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.491 0.682 0.535 ;
        RECT 0.614 0.1805 0.682 0.2245 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.398 0.048 0.466 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.29 0.453 0.358 0.497 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.358 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.472 ;
  END
END b15clb0a2as1n03x5

MACRO b15clb0a2as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.473 0.682 0.517 ;
        RECT 0.614 0.118 0.682 0.162 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.4 0.538 0.464 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.4 0.048 0.464 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.118 0.25 0.162 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
  END
END b15clb0a2as1n04x5

MACRO b15clb0a2as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n06x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.498 0.682 0.542 ;
        RECT 0.614 0.1645 0.682 0.2085 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.506 0.498 0.574 0.542 ;
        RECT 0.722 0.498 0.79 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.722 0.1645 0.79 0.2085 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.473 0.358 0.517 ;
      RECT 0.182 0.068 0.25 0.112 ;
      RECT 0.074 0.203 0.142 0.247 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.142 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.562 ;
  END
END b15clb0a2as1n06x5

MACRO b15clb0a2as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.473 0.682 0.517 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.3155 0.466 0.3595 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.722 0.473 0.79 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.3155 0.574 0.3595 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.203 0.25 0.247 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.428 0.506 0.472 ;
      RECT 0.506 0.248 0.574 0.472 ;
  END
END b15clb0a2as1n08x5

MACRO b15clb0a2as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n12x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.562 ;
        RECT 0.722 0.248 1.006 0.292 ;
        RECT 0.722 0.068 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.23925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.4795 0.358 0.5235 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.83 0.448 0.898 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.398 0.4795 0.466 0.5235 ;
      RECT 0.29 0.158 0.358 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
  END
END b15clb0a2as1n12x5

MACRO b15clb0a2as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n16x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.23925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.562 ;
        RECT 0.722 0.248 1.006 0.292 ;
        RECT 0.722 0.068 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.23925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.29 0.158 0.358 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.382 ;
  END
END b15clb0a2as1n16x5

MACRO b15clb0a2as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n24x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08262 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 0.722 0.158 1.438 0.202 ;
        RECT 0.83 0.338 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.832 0.358 0.896 0.402 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.199111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5450505 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.682 0.382 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
    LAYER v0 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.616 0.228 0.68 0.272 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.202 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.074 0.428 0.29 0.472 ;
      RECT 0.25 0.248 0.29 0.292 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.358 0.428 0.722 0.472 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 0.79 0.248 1.242 0.292 ;
  END
END b15clb0a2as1n24x5

MACRO b15clb0a2as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n32x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.84941175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5553845 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.10404 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.472 ;
        RECT 0.83 0.158 1.762 0.202 ;
        RECT 0.938 0.338 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.94 0.358 1.004 0.402 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.0314285 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.424706 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
    LAYER v0 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.724 0.228 0.788 0.272 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.182 0.068 0.25 0.112 ;
      RECT 0.182 0.441 0.25 0.485 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.162 0.068 0.506 0.112 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.292 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.428 0.83 0.472 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 0.898 0.248 1.654 0.292 ;
  END
END b15clb0a2as1n32x5

MACRO b15clb0a2as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n48x5 0 0 ;
  SIZE 2.376 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1683 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 2.322 0.472 ;
        RECT 1.154 0.158 2.322 0.202 ;
        RECT 2.126 0.158 2.194 0.472 ;
        RECT 1.91 0.158 1.978 0.472 ;
        RECT 1.694 0.158 1.762 0.472 ;
        RECT 1.154 0.158 1.222 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.156 0.228 1.22 0.272 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.4725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.589 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 1.114 0.292 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.41 0.022 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 2.234 0.248 2.302 0.382 ;
    LAYER v0 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.202 ;
      RECT 0.466 0.158 1.114 0.202 ;
      RECT 0.074 0.428 0.506 0.472 ;
      RECT 0.25 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.574 0.428 0.722 0.472 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.338 1.654 0.382 ;
  END
END b15clb0a2as1n48x5

MACRO b15clb0a2as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n64x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0387 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3849095 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.486 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.20808 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 2.754 0.472 ;
        RECT 2.558 0.068 2.626 0.472 ;
        RECT 1.478 0.248 2.626 0.292 ;
        RECT 2.342 0.068 2.41 0.472 ;
        RECT 2.126 0.068 2.194 0.472 ;
        RECT 1.91 0.068 1.978 0.472 ;
        RECT 1.694 0.068 1.762 0.292 ;
        RECT 1.478 0.068 1.546 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.478 0.1275 1.546 0.1715 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.694 0.1275 1.762 0.1715 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.91 0.1275 1.978 0.1715 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.126 0.1275 2.194 0.1715 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.342 0.1275 2.41 0.1715 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.558 0.1275 2.626 0.1715 ;
        RECT 2.666 0.428 2.734 0.472 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.25962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0504 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53984125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 1.438 0.292 ;
        RECT 1.37 0.158 1.438 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.262 0.248 1.33 0.292 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.666 -0.022 2.734 0.382 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.666 0.1275 2.734 0.1715 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
    LAYER v0 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.202 ;
      RECT 0.466 0.158 1.242 0.202 ;
      RECT 0.054 0.428 0.614 0.472 ;
      RECT 0.25 0.248 0.614 0.292 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.682 0.338 1.87 0.382 ;
  END
END b15clb0a2as1n64x5

MACRO b15clb0a2as1n80x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0a2as1n80x5 0 0 ;
  SIZE 4.104 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.703 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0513 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.682 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.25704 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.428 4.03 0.472 ;
        RECT 3.962 0.158 4.03 0.472 ;
        RECT 1.586 0.158 4.03 0.202 ;
        RECT 3.746 0.158 3.814 0.472 ;
        RECT 3.53 0.158 3.598 0.472 ;
        RECT 3.314 0.158 3.382 0.472 ;
        RECT 3.098 0.158 3.166 0.472 ;
        RECT 2.882 0.158 2.95 0.472 ;
        RECT 1.694 0.338 1.762 0.472 ;
      LAYER v0 ;
        RECT 1.696 0.358 1.76 0.402 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.428 2.626 0.472 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.774 0.158 2.842 0.202 ;
        RECT 2.99 0.428 3.058 0.472 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.206 0.158 3.274 0.202 ;
        RECT 3.422 0.428 3.49 0.472 ;
        RECT 3.422 0.158 3.49 0.202 ;
        RECT 3.638 0.428 3.706 0.472 ;
        RECT 3.638 0.158 3.706 0.202 ;
        RECT 3.854 0.428 3.922 0.472 ;
        RECT 3.854 0.158 3.922 0.202 ;
    END
  END clkout
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.91609425 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0675 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4030815 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.438 0.382 ;
        RECT 0.83 0.248 0.898 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END en
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.138 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 3.964 0.538 4.028 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.138 0.022 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
      LAYER v0 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.316 0.048 3.38 0.092 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.748 0.048 3.812 0.092 ;
        RECT 3.964 0.048 4.028 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
    LAYER v0 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.158 1.154 0.202 ;
      RECT 1.154 0.158 1.222 0.292 ;
      RECT 1.222 0.248 1.478 0.292 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 0.25 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.074 0.428 0.722 0.472 ;
      RECT 0.682 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 0.79 0.428 1.586 0.472 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.654 0.248 2.842 0.292 ;
  END
END b15clb0a2as1n80x5

MACRO b15clb0o2as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0o2as1n02x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.383 0.574 0.427 ;
        RECT 0.506 0.212 0.574 0.256 ;
    END
  END clkout
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END enb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.398 0.1315 0.466 0.1755 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.1315 0.358 0.1755 ;
      RECT 0.074 0.383 0.142 0.427 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.142 0.518 0.29 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
  END
END b15clb0o2as1n02x5

MACRO b15clb0o2as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0o2as1n03x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.408 0.574 0.452 ;
        RECT 0.506 0.212 0.574 0.256 ;
    END
  END clkout
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END enb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.212 0.142 0.256 ;
        RECT 0.398 0.1305 0.466 0.1745 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.1305 0.358 0.1745 ;
      RECT 0.074 0.387 0.142 0.431 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.142 0.518 0.29 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
  END
END b15clb0o2as1n03x5

MACRO b15clb0o2as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0o2as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.408 0.574 0.452 ;
        RECT 0.506 0.209 0.574 0.253 ;
    END
  END clkout
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END enb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.398 0.127 0.466 0.171 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.127 0.358 0.171 ;
      RECT 0.182 0.518 0.25 0.562 ;
    LAYER m1 ;
      RECT 0.162 0.518 0.29 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
  END
END b15clb0o2as1n04x5

MACRO b15clb0o2as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0o2as1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END clkout
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END enb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.338 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.182 0.518 0.25 0.562 ;
    LAYER m1 ;
      RECT 0.162 0.518 0.29 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
  END
END b15clb0o2as1n08x5

MACRO b15clb0o2as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0o2as1n12x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
        RECT 0.614 0.248 0.898 0.292 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.473 0.682 0.517 ;
        RECT 0.614 0.1375 0.682 0.1815 ;
        RECT 0.83 0.473 0.898 0.517 ;
        RECT 0.83 0.1375 0.898 0.1815 ;
    END
  END clkout
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END enb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.506 0.473 0.574 0.517 ;
        RECT 0.722 0.473 0.79 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.722 0.1375 0.79 0.1815 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.382 ;
  END
END b15clb0o2as1n12x5

MACRO b15clb0o2as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0o2as1n16x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.825679 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.472 ;
        RECT 0.83 0.248 1.114 0.292 ;
        RECT 0.83 0.068 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.3905 0.898 0.4345 ;
        RECT 0.83 0.1375 0.898 0.1815 ;
        RECT 1.046 0.3905 1.114 0.4345 ;
        RECT 1.046 0.1375 1.114 0.1815 ;
    END
  END clkout
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0171 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.40666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.682 0.382 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END enb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.938 0.485 1.006 0.529 ;
        RECT 1.154 0.485 1.222 0.529 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.938 0.1375 1.006 0.1815 ;
        RECT 1.154 0.1375 1.222 0.1815 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
    LAYER v0 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.182 0.408 0.25 0.452 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.398 0.562 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.428 0.79 0.472 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.382 ;
  END
END b15clb0o2as1n16x5

MACRO b15clb0o2as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0o2as1n24x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07956 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.438 0.382 ;
        RECT 1.37 0.158 1.438 0.382 ;
        RECT 0.722 0.158 1.438 0.202 ;
        RECT 1.262 0.338 1.33 0.562 ;
        RECT 1.046 0.338 1.114 0.562 ;
        RECT 0.83 0.338 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.262 0.158 1.33 0.202 ;
    END
  END clkout
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 0.65636375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 1.31272725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.702 0.382 ;
        RECT 0.29 0.338 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END enb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
    LAYER v0 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.614 0.133 0.682 0.177 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.182 0.133 0.25 0.177 ;
      RECT 0.182 0.408 0.25 0.452 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.398 0.562 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.428 0.79 0.472 ;
      RECT 0.25 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.248 1.242 0.292 ;
  END
END b15clb0o2as1n24x5

MACRO b15clb0o2as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0o2as1n32x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.2255 0.25 0.2695 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.10404 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 1.762 0.382 ;
        RECT 1.694 0.158 1.762 0.382 ;
        RECT 0.83 0.158 1.762 0.202 ;
        RECT 1.586 0.338 1.654 0.562 ;
        RECT 1.478 0.158 1.546 0.382 ;
        RECT 1.37 0.338 1.438 0.562 ;
        RECT 1.154 0.338 1.222 0.562 ;
        RECT 0.938 0.338 1.006 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.586 0.158 1.654 0.202 ;
    END
  END clkout
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.92239325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.594 0.292 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END enb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
      LAYER v0 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
    LAYER v0 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.722 0.133 0.79 0.177 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.133 0.358 0.177 ;
      RECT 0.292 0.408 0.356 0.452 ;
      RECT 0.182 0.518 0.25 0.562 ;
      RECT 0.074 0.133 0.142 0.177 ;
      RECT 0.076 0.408 0.14 0.452 ;
    LAYER m1 ;
      RECT 0.074 0.518 0.398 0.562 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.428 0.898 0.472 ;
      RECT 0.142 0.338 0.29 0.382 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.358 0.338 0.722 0.382 ;
      RECT 0.722 0.068 0.79 0.382 ;
      RECT 0.79 0.248 1.35 0.292 ;
  END
END b15clb0o2as1n32x5

MACRO b15clb0o2as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15clb0o2as1n64x5 0 0 ;
  SIZE 3.24 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41377775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END clk
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.428 3.186 0.472 ;
        RECT 1.262 0.158 3.186 0.202 ;
        RECT 2.99 0.158 3.058 0.472 ;
        RECT 2.774 0.158 2.842 0.472 ;
        RECT 2.558 0.158 2.626 0.472 ;
        RECT 2.342 0.158 2.41 0.472 ;
        RECT 1.37 0.338 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.372 0.358 1.436 0.402 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 2.882 0.158 2.95 0.202 ;
        RECT 3.098 0.428 3.166 0.472 ;
        RECT 3.098 0.158 3.166 0.202 ;
    END
  END clkout
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0513 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.33 0.382 ;
        RECT 1.046 0.248 1.114 0.382 ;
        RECT 0.614 0.248 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END enb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.274 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
      LAYER v0 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.776 0.538 2.84 0.582 ;
        RECT 2.992 0.538 3.056 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.274 0.022 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.472 ;
      RECT 3.098 0.248 3.166 0.382 ;
    LAYER v0 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.694 0.248 1.762 0.292 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.338 0.466 0.382 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.184 0.408 0.248 0.452 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.398 0.562 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.428 1.33 0.472 ;
      RECT 0.25 0.338 0.506 0.382 ;
      RECT 0.074 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.574 0.158 1.154 0.202 ;
      RECT 1.154 0.158 1.222 0.292 ;
      RECT 1.222 0.248 2.302 0.292 ;
  END
END b15clb0o2as1n64x5

MACRO b15cmbn22as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cmbn22as1n02x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.006 0.382 ;
        RECT 0.722 0.338 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
        RECT 0.182 0.158 0.358 0.202 ;
        RECT 0.182 0.068 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.178 0.142 0.222 ;
    END
  END clkout
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.248889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.248889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END s
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.248 0.608 0.292 ;
      RECT 0.688 0.248 1.256 0.292 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 1.154 0.248 1.222 0.472 ;
    LAYER v1 ;
      RECT 1.158 0.248 1.218 0.292 ;
      RECT 0.726 0.248 0.786 0.292 ;
      RECT 0.51 0.248 0.57 0.292 ;
      RECT 0.186 0.248 0.246 0.292 ;
    LAYER v0 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.338 0.25 0.382 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.702 0.202 ;
      RECT 0.682 0.248 0.81 0.292 ;
  END
END b15cmbn22as1n02x5

MACRO b15cmbn22as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cmbn22as1n03x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.006 0.382 ;
        RECT 0.722 0.338 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
        RECT 0.182 0.158 0.358 0.202 ;
        RECT 0.182 0.068 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.78666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.178 0.142 0.222 ;
    END
  END clkout
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.248889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.248889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END s
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.248 0.608 0.292 ;
      RECT 0.688 0.248 1.256 0.292 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 1.154 0.248 1.222 0.472 ;
    LAYER v1 ;
      RECT 1.158 0.248 1.218 0.292 ;
      RECT 0.726 0.248 0.786 0.292 ;
      RECT 0.51 0.248 0.57 0.292 ;
      RECT 0.186 0.248 0.246 0.292 ;
    LAYER v0 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.338 0.25 0.382 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.702 0.202 ;
      RECT 0.682 0.248 0.81 0.292 ;
  END
END b15cmbn22as1n03x5

MACRO b15cmbn22as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cmbn22as1n04x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.006 0.382 ;
        RECT 0.722 0.338 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
        RECT 0.182 0.158 0.358 0.202 ;
        RECT 0.182 0.068 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.178 0.142 0.222 ;
    END
  END clkout
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.248889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 6.248889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END s
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.248 0.608 0.292 ;
      RECT 0.688 0.248 1.256 0.292 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 1.154 0.248 1.222 0.472 ;
    LAYER v1 ;
      RECT 1.158 0.248 1.218 0.292 ;
      RECT 0.726 0.248 0.786 0.292 ;
      RECT 0.51 0.248 0.57 0.292 ;
      RECT 0.186 0.248 0.246 0.292 ;
    LAYER v0 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.338 0.25 0.382 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.702 0.202 ;
      RECT 0.682 0.248 0.81 0.292 ;
  END
END b15cmbn22as1n04x5

MACRO b15cmbn22as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cmbn22as1n08x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.3155 0.25 0.3595 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.562 ;
      LAYER v0 ;
        RECT 1.802 0.3155 1.87 0.3595 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.068 1.654 0.562 ;
      LAYER v0 ;
        RECT 1.586 0.498 1.654 0.542 ;
        RECT 1.586 0.138 1.654 0.182 ;
    END
  END clkout
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 2.48507925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 5.7985185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.3115 0.682 0.3555 ;
    END
  END s
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 1.478 0.498 1.546 0.542 ;
        RECT 1.694 0.498 1.762 0.542 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.694 0.138 1.762 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.338 0.932 0.382 ;
      RECT 1.012 0.338 2.012 0.382 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 1.91 0.068 1.978 0.562 ;
    LAYER v1 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.834 0.338 0.894 0.382 ;
      RECT 0.078 0.338 0.138 0.382 ;
    LAYER v0 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.498 1.978 0.542 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.408 0.79 0.452 ;
      RECT 0.506 0.152 0.574 0.196 ;
      RECT 0.506 0.429 0.574 0.473 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.562 ;
      RECT 0.79 0.518 0.938 0.562 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.006 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 0.574 0.068 1.33 0.112 ;
  END
END b15cmbn22as1n08x5

MACRO b15cmbn22as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cmbn22as1n12x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.3155 0.25 0.3595 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.472 ;
      LAYER v0 ;
        RECT 2.018 0.3155 2.086 0.3595 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.068 1.762 0.562 ;
        RECT 1.478 0.338 1.762 0.382 ;
        RECT 1.478 0.068 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 1.694 0.138 1.762 0.182 ;
    END
  END clkout
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 2.046536 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 6.95822225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.3155 0.79 0.3595 ;
    END
  END s
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.018 0.538 2.086 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.338 1.04 0.382 ;
      RECT 1.12 0.338 2.12 0.382 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 1.91 0.068 1.978 0.562 ;
    LAYER v1 ;
      RECT 1.914 0.338 1.974 0.382 ;
      RECT 1.158 0.338 1.218 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.294 0.338 0.354 0.382 ;
    LAYER v0 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.223 1.33 0.267 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.154 0.223 1.222 0.267 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 1.046 0.223 1.114 0.267 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.938 0.223 1.006 0.267 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.83 0.223 0.898 0.267 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.614 0.408 0.682 0.452 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.29 0.448 0.358 0.492 ;
    LAYER m1 ;
      RECT 0.83 0.158 0.898 0.562 ;
      RECT 0.898 0.518 1.046 0.562 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 0.682 0.068 1.35 0.112 ;
  END
END b15cmbn22as1n12x5

MACRO b15cmbn22as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cmbn22as1n16x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.43712425 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.248 2.41 0.292 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.428 2.194 0.472 ;
        RECT 2.126 0.158 2.194 0.472 ;
        RECT 1.694 0.158 2.194 0.202 ;
      LAYER v0 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.202 ;
    END
  END clkout
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 1.16686875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 1.16686875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.898 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END s
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.428 2.32 0.472 ;
    LAYER m1 ;
      RECT 0.83 0.428 1.114 0.472 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 1.154 0.158 1.478 0.202 ;
      RECT 0.722 0.518 1.586 0.562 ;
      RECT 2.234 0.068 2.302 0.472 ;
    LAYER v1 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 0.942 0.428 1.002 0.472 ;
    LAYER v0 ;
      RECT 2.234 0.149 2.302 0.193 ;
      RECT 2.234 0.408 2.302 0.452 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.574 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.382 ;
      RECT 1.006 0.338 1.33 0.382 ;
      RECT 0.142 0.428 0.466 0.472 ;
      RECT 0.142 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 1.154 0.428 1.37 0.472 ;
      RECT 1.114 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 0.722 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 1.654 0.248 1.978 0.292 ;
  END
END b15cmbn22as1n16x5

MACRO b15cmbn22as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cmbn22as1n24x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0189 LAYER m1 ;
      ANTENNAMAXAREACAR 0.687619 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0189 LAYER m1 ;
      ANTENNAMAXAREACAR 0.687619 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.158 2.842 0.472 ;
      LAYER v0 ;
        RECT 2.774 0.338 2.842 0.382 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07956 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.428 2.626 0.472 ;
        RECT 2.558 0.158 2.626 0.472 ;
        RECT 1.91 0.158 2.626 0.202 ;
      LAYER v0 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.45 0.158 2.518 0.202 ;
    END
  END clkout
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0279 LAYER m1 ;
      ANTENNAMAXAREACAR 1.0541935 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0279 LAYER m1 ;
      ANTENNAMAXAREACAR 1.0541935 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.898 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END s
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.776 0.538 2.84 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.92 0.338 2.984 0.382 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.054 0.428 0.398 0.472 ;
      RECT 1.262 0.158 1.694 0.202 ;
      RECT 0.83 0.518 1.802 0.562 ;
      RECT 2.666 0.068 2.734 0.562 ;
      RECT 2.882 0.068 2.95 0.562 ;
    LAYER v1 ;
      RECT 2.886 0.338 2.946 0.382 ;
      RECT 2.67 0.338 2.73 0.382 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
    LAYER v0 ;
      RECT 2.882 0.156 2.95 0.2 ;
      RECT 2.882 0.4405 2.95 0.4845 ;
      RECT 2.666 0.156 2.734 0.2 ;
      RECT 2.666 0.4405 2.734 0.4845 ;
      RECT 2.342 0.248 2.41 0.292 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 1.91 0.248 1.978 0.292 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.506 0.4505 0.574 0.4945 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.722 0.428 0.938 0.472 ;
      RECT 0.938 0.338 1.006 0.472 ;
      RECT 1.006 0.428 1.222 0.472 ;
      RECT 0.574 0.248 1.046 0.292 ;
      RECT 1.046 0.248 1.114 0.382 ;
      RECT 1.114 0.338 1.438 0.382 ;
      RECT 0.054 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.158 1.154 0.202 ;
      RECT 1.154 0.158 1.222 0.292 ;
      RECT 1.262 0.428 1.478 0.472 ;
      RECT 1.222 0.248 1.478 0.292 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 1.546 0.428 1.762 0.472 ;
      RECT 1.694 0.158 1.762 0.382 ;
      RECT 0.83 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.562 ;
      RECT 1.87 0.248 2.518 0.292 ;
  END
END b15cmbn22as1n24x5

MACRO b15cmbn22as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cmbn22as1n32x5 0 0 ;
  SIZE 3.672 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
        RECT 0.182 0.248 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.158 3.598 0.472 ;
      LAYER v0 ;
        RECT 3.53 0.338 3.598 0.382 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.10404 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.428 3.166 0.472 ;
        RECT 3.098 0.158 3.166 0.472 ;
        RECT 2.234 0.158 3.166 0.202 ;
      LAYER v0 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.428 2.626 0.472 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.774 0.158 2.842 0.202 ;
        RECT 2.99 0.428 3.058 0.472 ;
        RECT 2.99 0.158 3.058 0.202 ;
    END
  END clkout
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.931 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.931 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.222 0.382 ;
        RECT 0.722 0.338 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END s
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.706 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.706 0.022 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
        RECT 3.316 0.048 3.38 0.092 ;
        RECT 3.532 0.048 3.596 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.028 0.428 3.508 0.472 ;
    LAYER m1 ;
      RECT 0.938 0.428 1.438 0.472 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 1.478 0.158 2.018 0.202 ;
      RECT 0.83 0.518 2.126 0.562 ;
      RECT 3.206 0.068 3.274 0.562 ;
      RECT 3.422 0.068 3.49 0.562 ;
    LAYER v1 ;
      RECT 3.426 0.428 3.486 0.472 ;
      RECT 3.21 0.428 3.27 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.266 0.428 1.326 0.472 ;
      RECT 1.05 0.428 1.11 0.472 ;
    LAYER v0 ;
      RECT 3.422 0.152 3.49 0.196 ;
      RECT 3.422 0.435 3.49 0.479 ;
      RECT 3.206 0.152 3.274 0.196 ;
      RECT 3.206 0.435 3.274 0.479 ;
      RECT 2.882 0.248 2.95 0.292 ;
      RECT 2.666 0.248 2.734 0.292 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.4505 0.682 0.4945 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.4 0.358 0.464 0.402 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 0.682 0.248 1.262 0.292 ;
      RECT 1.262 0.248 1.33 0.382 ;
      RECT 1.33 0.338 1.87 0.382 ;
      RECT 0.142 0.428 0.398 0.472 ;
      RECT 0.398 0.338 0.466 0.472 ;
      RECT 0.142 0.158 1.37 0.202 ;
      RECT 1.37 0.158 1.438 0.292 ;
      RECT 1.478 0.428 1.91 0.472 ;
      RECT 1.438 0.248 1.91 0.292 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 0.83 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.562 ;
      RECT 2.194 0.248 3.058 0.292 ;
  END
END b15cmbn22as1n32x5

MACRO b15cmbn22as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15cmbn22as1n64x5 0 0 ;
  SIZE 6.48 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.072 LAYER m1 ;
      ANTENNAGATEAREA 0.072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.6935 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2820555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.16133325 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.072 LAYER m1 ;
      ANTENNAGATEAREA 0.072 LAYER m2 ;
      ANTENNAMAXAREACAR 0.6935 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2820555 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.16133325 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.338 2.086 0.382 ;
        RECT 1.262 0.338 1.33 0.472 ;
      LAYER m2 ;
        RECT 0.92 0.428 1.472 0.472 ;
      LAYER v1 ;
        RECT 1.266 0.428 1.326 0.472 ;
      LAYER v0 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.694 0.338 1.762 0.382 ;
        RECT 1.91 0.338 1.978 0.382 ;
    END
  END s
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.543611 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.543611 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.898 0.292 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 6.338 0.248 6.406 0.472 ;
        RECT 5.582 0.248 6.406 0.292 ;
      LAYER v0 ;
        RECT 5.69 0.248 5.758 0.292 ;
        RECT 5.906 0.248 5.974 0.292 ;
        RECT 6.122 0.248 6.19 0.292 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.20808 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.428 5.434 0.472 ;
        RECT 5.366 0.158 5.434 0.472 ;
        RECT 3.53 0.158 5.434 0.202 ;
        RECT 3.53 0.338 3.598 0.472 ;
      LAYER v0 ;
        RECT 3.532 0.358 3.596 0.402 ;
        RECT 3.638 0.158 3.706 0.202 ;
        RECT 3.746 0.428 3.814 0.472 ;
        RECT 3.854 0.158 3.922 0.202 ;
        RECT 3.962 0.428 4.03 0.472 ;
        RECT 4.07 0.158 4.138 0.202 ;
        RECT 4.178 0.428 4.246 0.472 ;
        RECT 4.286 0.158 4.354 0.202 ;
        RECT 4.394 0.428 4.462 0.472 ;
        RECT 4.502 0.158 4.57 0.202 ;
        RECT 4.61 0.428 4.678 0.472 ;
        RECT 4.718 0.158 4.786 0.202 ;
        RECT 4.826 0.428 4.894 0.472 ;
        RECT 4.934 0.158 5.002 0.202 ;
        RECT 5.042 0.428 5.11 0.472 ;
        RECT 5.15 0.158 5.218 0.202 ;
        RECT 5.258 0.428 5.326 0.472 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.514 0.652 ;
        RECT 6.338 0.518 6.406 0.652 ;
        RECT 6.122 0.518 6.19 0.652 ;
        RECT 5.906 0.518 5.974 0.652 ;
        RECT 5.69 0.518 5.758 0.652 ;
        RECT 5.474 0.518 5.542 0.652 ;
        RECT 5.15 0.518 5.218 0.652 ;
        RECT 4.934 0.518 5.002 0.652 ;
        RECT 4.718 0.518 4.786 0.652 ;
        RECT 4.502 0.518 4.57 0.652 ;
        RECT 4.286 0.518 4.354 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.854 0.518 3.922 0.652 ;
        RECT 3.638 0.518 3.706 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 3.64 0.538 3.704 0.582 ;
        RECT 3.856 0.538 3.92 0.582 ;
        RECT 4.072 0.538 4.136 0.582 ;
        RECT 4.288 0.538 4.352 0.582 ;
        RECT 4.504 0.538 4.568 0.582 ;
        RECT 4.72 0.538 4.784 0.582 ;
        RECT 4.936 0.538 5 0.582 ;
        RECT 5.152 0.538 5.216 0.582 ;
        RECT 5.476 0.538 5.54 0.582 ;
        RECT 5.692 0.538 5.756 0.582 ;
        RECT 5.908 0.538 5.972 0.582 ;
        RECT 6.124 0.538 6.188 0.582 ;
        RECT 6.34 0.538 6.404 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.514 0.022 ;
        RECT 6.338 -0.022 6.406 0.112 ;
        RECT 6.122 -0.022 6.19 0.112 ;
        RECT 5.906 -0.022 5.974 0.112 ;
        RECT 5.69 -0.022 5.758 0.112 ;
        RECT 5.474 -0.022 5.542 0.112 ;
        RECT 5.258 -0.022 5.326 0.112 ;
        RECT 5.042 -0.022 5.11 0.112 ;
        RECT 4.826 -0.022 4.894 0.112 ;
        RECT 4.61 -0.022 4.678 0.112 ;
        RECT 4.394 -0.022 4.462 0.112 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.748 0.048 3.812 0.092 ;
        RECT 3.964 0.048 4.028 0.092 ;
        RECT 4.18 0.048 4.244 0.092 ;
        RECT 4.396 0.048 4.46 0.092 ;
        RECT 4.612 0.048 4.676 0.092 ;
        RECT 4.828 0.048 4.892 0.092 ;
        RECT 5.044 0.048 5.108 0.092 ;
        RECT 5.26 0.048 5.324 0.092 ;
        RECT 5.476 0.048 5.54 0.092 ;
        RECT 5.692 0.048 5.756 0.092 ;
        RECT 5.908 0.048 5.972 0.092 ;
        RECT 6.124 0.048 6.188 0.092 ;
        RECT 6.34 0.048 6.404 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.552 0.428 6.316 0.472 ;
    LAYER m1 ;
      RECT 0.938 0.428 1.154 0.472 ;
      RECT 1.37 0.428 2.302 0.472 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 2.342 0.158 3.314 0.202 ;
      RECT 1.262 0.518 3.422 0.562 ;
      RECT 5.474 0.158 5.542 0.472 ;
    LAYER v1 ;
      RECT 6.234 0.428 6.294 0.472 ;
      RECT 6.018 0.428 6.078 0.472 ;
      RECT 5.802 0.428 5.862 0.472 ;
      RECT 5.586 0.428 5.646 0.472 ;
      RECT 3.318 0.428 3.378 0.472 ;
      RECT 2.238 0.428 2.298 0.472 ;
      RECT 2.022 0.428 2.082 0.472 ;
      RECT 1.806 0.428 1.866 0.472 ;
      RECT 1.59 0.428 1.65 0.472 ;
    LAYER v0 ;
      RECT 6.23 0.158 6.298 0.202 ;
      RECT 6.232 0.358 6.296 0.402 ;
      RECT 6.014 0.158 6.082 0.202 ;
      RECT 6.014 0.428 6.082 0.472 ;
      RECT 5.798 0.158 5.866 0.202 ;
      RECT 5.798 0.428 5.866 0.472 ;
      RECT 5.582 0.158 5.65 0.202 ;
      RECT 5.582 0.428 5.65 0.472 ;
      RECT 5.15 0.338 5.218 0.382 ;
      RECT 4.934 0.338 5.002 0.382 ;
      RECT 4.718 0.338 4.786 0.382 ;
      RECT 4.502 0.338 4.57 0.382 ;
      RECT 4.286 0.248 4.354 0.292 ;
      RECT 4.07 0.248 4.138 0.292 ;
      RECT 3.854 0.248 3.922 0.292 ;
      RECT 3.638 0.248 3.706 0.292 ;
      RECT 3.206 0.068 3.274 0.112 ;
      RECT 3.206 0.518 3.274 0.562 ;
      RECT 3.098 0.158 3.166 0.202 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.99 0.068 3.058 0.112 ;
      RECT 2.99 0.338 3.058 0.382 ;
      RECT 2.99 0.518 3.058 0.562 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.882 0.428 2.95 0.472 ;
      RECT 2.774 0.068 2.842 0.112 ;
      RECT 2.774 0.338 2.842 0.382 ;
      RECT 2.774 0.518 2.842 0.562 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.558 0.338 2.626 0.382 ;
      RECT 2.558 0.518 2.626 0.562 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.832 0.358 0.896 0.402 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.33 0.338 2.086 0.382 ;
      RECT 0.938 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.222 0.248 2.126 0.292 ;
      RECT 2.126 0.248 2.194 0.382 ;
      RECT 2.194 0.338 3.166 0.382 ;
      RECT 0.142 0.428 0.83 0.472 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.142 0.158 2.234 0.202 ;
      RECT 2.234 0.158 2.302 0.292 ;
      RECT 2.342 0.428 3.206 0.472 ;
      RECT 2.302 0.248 3.206 0.292 ;
      RECT 3.206 0.248 3.274 0.472 ;
      RECT 3.314 0.158 3.382 0.472 ;
      RECT 1.262 0.068 3.422 0.112 ;
      RECT 3.422 0.068 3.49 0.562 ;
      RECT 3.49 0.248 4.394 0.292 ;
      RECT 4.394 0.248 4.462 0.382 ;
      RECT 4.462 0.338 5.326 0.382 ;
      RECT 5.542 0.428 6.23 0.472 ;
      RECT 6.23 0.338 6.298 0.472 ;
      RECT 5.542 0.158 6.406 0.202 ;
  END
END b15cmbn22as1n64x5

MACRO b15corn02as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15corn02as1n02x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.383 0.574 0.427 ;
        RECT 0.506 0.212 0.574 0.256 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.398 0.13 0.466 0.174 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.13 0.358 0.174 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.162 0.428 0.29 0.472 ;
      RECT 0.29 0.068 0.358 0.472 ;
  END
END b15corn02as1n02x5

MACRO b15corn02as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15corn02as1n03x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.388 0.574 0.432 ;
        RECT 0.506 0.211 0.574 0.255 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.398 0.13 0.466 0.174 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.13 0.358 0.174 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.162 0.428 0.29 0.472 ;
      RECT 0.29 0.068 0.358 0.472 ;
  END
END b15corn02as1n03x5

MACRO b15corn02as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15corn02as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.506 0.136 0.574 0.18 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.398 0.136 0.466 0.18 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.136 0.358 0.18 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.162 0.428 0.29 0.472 ;
      RECT 0.29 0.068 0.358 0.472 ;
  END
END b15corn02as1n04x5

MACRO b15corn02as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15corn02as1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.451 0.574 0.495 ;
        RECT 0.506 0.13 0.574 0.174 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.614 0.451 0.682 0.495 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.398 0.13 0.466 0.174 ;
        RECT 0.614 0.13 0.682 0.174 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.13 0.358 0.174 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.162 0.428 0.29 0.472 ;
      RECT 0.29 0.068 0.358 0.472 ;
  END
END b15corn02as1n08x5

MACRO b15corn02as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15corn02as1n12x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.562 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.456 0.574 0.5 ;
        RECT 0.506 0.13 0.574 0.174 ;
        RECT 0.722 0.456 0.79 0.5 ;
        RECT 0.722 0.13 0.79 0.174 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.614 0.456 0.682 0.5 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.398 0.13 0.466 0.174 ;
        RECT 0.614 0.13 0.682 0.174 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.13 0.358 0.174 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.162 0.428 0.29 0.472 ;
      RECT 0.29 0.068 0.358 0.472 ;
  END
END b15corn02as1n12x5

MACRO b15corn02as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15corn02as1n16x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 1.4114285 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0135 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7994075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.682 0.382 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06426 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.562 ;
        RECT 0.83 0.248 1.33 0.292 ;
        RECT 1.046 0.068 1.114 0.562 ;
        RECT 0.83 0.068 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.457 0.898 0.501 ;
        RECT 0.83 0.1045 0.898 0.1485 ;
        RECT 1.046 0.457 1.114 0.501 ;
        RECT 1.046 0.1045 1.114 0.1485 ;
        RECT 1.262 0.457 1.33 0.501 ;
        RECT 1.262 0.1045 1.33 0.1485 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.938 0.457 1.006 0.501 ;
        RECT 1.154 0.457 1.222 0.501 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.938 0.1045 1.006 0.1485 ;
        RECT 1.154 0.1045 1.222 0.1485 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
    LAYER v0 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.182 0.408 0.25 0.452 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.398 0.562 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.428 0.79 0.472 ;
      RECT 0.25 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.382 ;
  END
END b15corn02as1n16x5

MACRO b15corn02as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15corn02as1n24x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.825679 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 0.65636375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 1.11076925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.702 0.382 ;
        RECT 0.29 0.338 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.428 1.566 0.472 ;
        RECT 0.722 0.158 1.566 0.202 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 0.938 0.338 1.006 0.472 ;
        RECT 0.81 0.338 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.13 0.142 0.174 ;
        RECT 0.398 0.13 0.466 0.174 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 1.478 0.248 1.546 0.382 ;
    LAYER v0 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.614 0.133 0.682 0.177 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.182 0.13 0.25 0.174 ;
      RECT 0.182 0.408 0.25 0.452 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.398 0.562 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.428 0.898 0.472 ;
      RECT 0.25 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.248 1.242 0.292 ;
  END
END b15corn02as1n24x5

MACRO b15corn02as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15corn02as1n32x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.20333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.9025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11628 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.428 1.89 0.472 ;
        RECT 0.83 0.158 1.89 0.202 ;
        RECT 1.694 0.158 1.762 0.472 ;
        RECT 1.046 0.338 1.114 0.472 ;
        RECT 0.83 0.338 1.114 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
      LAYER v0 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 1.802 0.248 1.87 0.382 ;
    LAYER v0 ;
      RECT 1.478 0.248 1.546 0.292 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.518 0.25 0.562 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.518 0.506 0.562 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.428 0.898 0.472 ;
      RECT 0.054 0.428 0.182 0.472 ;
      RECT 0.142 0.248 0.182 0.292 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.25 0.428 0.398 0.472 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.292 ;
      RECT 0.79 0.248 1.566 0.292 ;
  END
END b15corn02as1n32x5

MACRO b15corn02as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15corn02as1n64x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.52777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.81196575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.486 0.292 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60462225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0324 LAYER m1 ;
      ANTENNAMAXAREACAR 0.839753 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.35 0.382 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END clk2
  PIN clkout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.428 3.294 0.472 ;
        RECT 1.37 0.158 3.294 0.202 ;
        RECT 3.098 0.158 3.166 0.472 ;
        RECT 2.882 0.158 2.95 0.472 ;
        RECT 2.666 0.158 2.734 0.472 ;
        RECT 2.45 0.158 2.518 0.472 ;
        RECT 2.234 0.158 2.302 0.472 ;
        RECT 1.586 0.338 1.654 0.472 ;
        RECT 1.458 0.338 1.654 0.382 ;
      LAYER v0 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.428 2.626 0.472 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.774 0.158 2.842 0.202 ;
        RECT 2.99 0.428 3.058 0.472 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.206 0.158 3.274 0.202 ;
    END
  END clkout
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
      LAYER v0 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.472 ;
      RECT 3.206 0.248 3.274 0.382 ;
    LAYER v0 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.292 0.408 0.356 0.452 ;
      RECT 0.182 0.518 0.25 0.562 ;
      RECT 0.076 0.408 0.14 0.452 ;
    LAYER m1 ;
      RECT 0.074 0.518 0.506 0.562 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.428 1.546 0.472 ;
      RECT 0.142 0.338 0.29 0.382 ;
      RECT 0.29 0.338 0.358 0.472 ;
      RECT 0.358 0.338 0.614 0.382 ;
      RECT 0.182 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 0.682 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.33 0.248 2.194 0.292 ;
  END
END b15corn02as1n64x5

MACRO b15inv000as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n02x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
    END
  END vssx
END b15inv000as1n02x5

MACRO b15inv000as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n03x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
    END
  END vssx
END b15inv000as1n03x5

MACRO b15inv000as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n04x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
    END
  END vssx
END b15inv000as1n04x5

MACRO b15inv000as1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n05x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
    END
  END vssx
END b15inv000as1n05x5

MACRO b15inv000as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n06x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
END b15inv000as1n06x5

MACRO b15inv000as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n08x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
    END
  END vssx
END b15inv000as1n08x5

MACRO b15inv000as1n10x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n10x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 0.494 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 0.494 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
    END
  END vssx
END b15inv000as1n10x5

MACRO b15inv000as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n12x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
END b15inv000as1n12x5

MACRO b15inv000as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n16x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.158 0.466 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.158 0.574 0.202 ;
    END
  END vssx
END b15inv000as1n16x5

MACRO b15inv000as1n20x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n20x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.589 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.589 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.182 0.338 0.682 0.382 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.158 0.574 0.202 ;
    END
  END vssx
END b15inv000as1n20x5

MACRO b15inv000as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n24x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.378 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.79 0.472 ;
        RECT 0.722 0.248 0.79 0.472 ;
        RECT 0.182 0.248 0.79 0.292 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.506 0.248 0.574 0.472 ;
        RECT 0.398 0.068 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.1275 0.25 0.1715 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.1275 0.466 0.1715 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.1275 0.682 0.1715 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
END b15inv000as1n24x5

MACRO b15inv000as1n28x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n28x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0504 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5835715 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0504 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5835715 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.486 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.472 ;
        RECT 0.054 0.158 0.898 0.202 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.722 0.158 0.79 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
    END
  END vssx
END b15inv000as1n28x5

MACRO b15inv000as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n32x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.682 0.382 ;
        RECT 0.614 0.248 0.682 0.382 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.006 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.074 0.158 1.006 0.202 ;
        RECT 0.722 0.158 0.79 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
END b15inv000as1n32x5

MACRO b15inv000as1n40x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n40x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5795 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5795 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.898 0.382 ;
        RECT 0.83 0.248 0.898 0.382 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.074 0.158 1.222 0.202 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
END b15inv000as1n40x5

MACRO b15inv000as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n48x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57791675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57791675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.898 0.382 ;
        RECT 0.83 0.248 0.898 0.382 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14688 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 0.074 0.158 1.438 0.202 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
END b15inv000as1n48x5

MACRO b15inv000as1n56x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n56x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.1008 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57678575 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.1008 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57678575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.114 0.382 ;
        RECT 1.046 0.248 1.114 0.382 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.17136 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 0.074 0.158 1.654 0.202 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.506 0.158 0.574 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
    END
  END vssx
END b15inv000as1n56x5

MACRO b15inv000as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n64x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.1152 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5759375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.1152 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5759375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.33 0.382 ;
        RECT 1.262 0.248 1.33 0.382 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.19584 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 0.074 0.158 1.87 0.202 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 0.506 0.158 0.574 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
    END
  END vssx
END b15inv000as1n64x5

MACRO b15inv000as1n80x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv000as1n80x5 0 0 ;
  SIZE 2.376 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 1.762 0.382 ;
        RECT 0.83 0.248 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.472 ;
        RECT 0.074 0.158 2.302 0.202 ;
        RECT 2.018 0.158 2.086 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.158 2.194 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.41 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.41 0.022 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
    END
  END vssx
END b15inv000as1n80x5

MACRO b15inv020as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n03x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.1105 0.25 0.1545 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.1105 0.142 0.1545 ;
    END
  END vssx
END b15inv020as1n03x5

MACRO b15inv020as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n04x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.452 0.25 0.496 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
    END
  END vssx
END b15inv020as1n04x5

MACRO b15inv020as1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n05x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.4775 0.25 0.5215 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4775 0.142 0.5215 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
    END
  END vssx
END b15inv020as1n05x5

MACRO b15inv020as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n06x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.158 0.358 0.202 ;
    END
  END vssx
END b15inv020as1n06x5

MACRO b15inv020as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n08x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.455 0.25 0.499 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.455 0.358 0.499 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
END b15inv020as1n08x5

MACRO b15inv020as1n10x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n10x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 0.494 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.4755 0.25 0.5195 ;
        RECT 0.182 0.1115 0.25 0.1555 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4755 0.142 0.5195 ;
        RECT 0.29 0.4755 0.358 0.5195 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.1115 0.142 0.1555 ;
        RECT 0.29 0.1115 0.358 0.1555 ;
    END
  END vssx
END b15inv020as1n10x5

MACRO b15inv020as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n12x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.84941175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03978 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.476 0.25 0.52 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.476 0.466 0.52 ;
        RECT 0.398 0.158 0.466 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.476 0.142 0.52 ;
        RECT 0.29 0.476 0.358 0.52 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.158 0.358 0.202 ;
    END
  END vssx
END b15inv020as1n12x5

MACRO b15inv020as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n16x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04284 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.4765 0.25 0.5205 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.4765 0.466 0.5205 ;
        RECT 0.398 0.158 0.466 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4765 0.142 0.5205 ;
        RECT 0.29 0.4765 0.358 0.5205 ;
        RECT 0.506 0.4765 0.574 0.5205 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.158 0.574 0.202 ;
    END
  END vssx
END b15inv020as1n16x5

MACRO b15inv020as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n24x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7139395 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.48081625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.182 0.248 0.682 0.292 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.518 0.358 0.562 ;
        RECT 0.506 0.518 0.574 0.562 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END vssx
END b15inv020as1n24x5

MACRO b15inv020as1n28x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n28x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0369 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68585375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0513 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.182 0.338 0.682 0.382 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.518 0.358 0.562 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 0.722 0.518 0.79 0.562 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.068 0.358 0.112 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 0.722 0.068 0.79 0.112 ;
    END
  END vssx
END b15inv020as1n28x5

MACRO b15inv020as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n32x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0594 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4260605 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08874 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.562 ;
        RECT 0.182 0.338 0.682 0.382 ;
        RECT 0.182 0.158 0.682 0.202 ;
        RECT 0.398 0.338 0.466 0.562 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.184 0.23 0.248 0.274 ;
        RECT 0.182 0.4535 0.25 0.4975 ;
        RECT 0.398 0.4535 0.466 0.4975 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.616 0.23 0.68 0.274 ;
        RECT 0.614 0.4535 0.682 0.4975 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
END b15inv020as1n32x5

MACRO b15inv020as1n40x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n40x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0504 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5835715 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0738 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3985365 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.574 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11934 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 0.898 0.472 ;
        RECT 0.83 0.068 0.898 0.472 ;
        RECT 0.182 0.248 0.898 0.292 ;
        RECT 0.614 0.068 0.682 0.472 ;
        RECT 0.398 0.068 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
END b15inv020as1n40x5

MACRO b15inv020as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n48x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0648 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5805555 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0882 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4265305 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 1.006 0.382 ;
        RECT 0.938 0.248 1.006 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14382 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.472 ;
        RECT 0.054 0.158 1.114 0.202 ;
        RECT 0.398 0.158 0.466 0.472 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 0.938 0.158 1.006 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.382 ;
  END
END b15inv020as1n48x5

MACRO b15inv020as1n56x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n56x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5795 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.1026 LAYER m1 ;
      ANTENNAMAXAREACAR 0.40666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.898 0.382 ;
        RECT 0.83 0.248 0.898 0.382 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14994 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.074 0.158 1.222 0.202 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
END b15inv020as1n56x5

MACRO b15inv020as1n64x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n64x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57791675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.42676925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.898 0.382 ;
        RECT 0.83 0.248 0.898 0.382 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.17442 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 0.074 0.158 1.438 0.202 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
END b15inv020as1n64x5

MACRO b15inv020as1n80x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv020as1n80x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57633325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.1458 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4269135 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 1.222 0.382 ;
        RECT 1.154 0.248 1.222 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2295 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.472 ;
        RECT 0.054 0.158 1.762 0.202 ;
        RECT 1.478 0.158 1.546 0.472 ;
        RECT 1.262 0.158 1.33 0.472 ;
        RECT 0.398 0.158 0.466 0.472 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.382 ;
  END
END b15inv020as1n80x5

MACRO b15inv040as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n02x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.3835 0.25 0.4275 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4645 0.142 0.5085 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
    END
  END vssx
END b15inv040as1n02x5

MACRO b15inv040as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n03x5 0 0 ;
  SIZE 0.324 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.3885 0.25 0.4325 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.488 0.142 0.532 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.358 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
    END
  END vssx
END b15inv040as1n03x5

MACRO b15inv040as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.363 0.25 0.407 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
END b15inv040as1n04x5

MACRO b15inv040as1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n05x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 0.89818175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.182 0.196 0.25 0.24 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4925 0.142 0.5365 ;
        RECT 0.29 0.493 0.358 0.537 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.196 0.358 0.24 ;
    END
  END vssx
END b15inv040as1n05x5

MACRO b15inv040as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n06x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.3925 0.25 0.4365 ;
        RECT 0.182 0.158 0.25 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.29 0.473 0.358 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.158 0.358 0.202 ;
    END
  END vssx
END b15inv040as1n06x5

MACRO b15inv040as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n08x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.84941175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04284 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.452 0.25 0.496 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.452 0.466 0.496 ;
        RECT 0.398 0.158 0.466 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.452 0.142 0.496 ;
        RECT 0.29 0.452 0.358 0.496 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.158 0.358 0.202 ;
    END
  END vssx
END b15inv040as1n08x5

MACRO b15inv040as1n10x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n10x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0261 LAYER m1 ;
      ANTENNAMAXAREACAR 0.497931 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0189 LAYER m1 ;
      ANTENNAMAXAREACAR 0.687619 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.446 0.25 0.49 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.446 0.466 0.49 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.446 0.358 0.49 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
END b15inv040as1n10x5

MACRO b15inv040as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n12x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04284 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.3935 0.25 0.4375 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.3935 0.466 0.4375 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.477 0.142 0.521 ;
        RECT 0.29 0.477 0.358 0.521 ;
        RECT 0.506 0.477 0.574 0.521 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END vssx
END b15inv040as1n12x5

MACRO b15inv040as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n16x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.48081625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7139395 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.182 0.338 0.682 0.382 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.423 0.25 0.467 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.431 0.466 0.475 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.425 0.682 0.469 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END vssx
END b15inv040as1n16x5

MACRO b15inv040as1n20x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n20x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0513 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0369 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68585375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.182 0.338 0.682 0.382 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.722 0.428 0.79 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
END b15inv040as1n20x5

MACRO b15inv040as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n24x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0657 LAYER m1 ;
      ANTENNAMAXAREACAR 0.510137 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.77583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
        RECT 0.182 0.338 0.898 0.382 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
END b15inv040as1n24x5

MACRO b15inv040as1n28x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n28x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4655 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0513 LAYER m1 ;
      ANTENNAMAXAREACAR 0.65333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.10404 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
        RECT 0.182 0.338 0.898 0.382 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.4435 0.25 0.4875 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.4435 0.466 0.4875 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.4435 0.682 0.4875 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 0.83 0.4435 0.898 0.4875 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
END b15inv040as1n28x5

MACRO b15inv040as1n36x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n36x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.47793825 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0657 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6350685 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.382 ;
        RECT 0.398 0.248 0.898 0.292 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.12852 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.074 0.158 1.222 0.202 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.154 0.538 1.222 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.154 0.048 1.222 0.092 ;
    END
  END vssx
END b15inv040as1n36x5

MACRO b15inv040as1n40x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n40x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.1017 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4909735 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0729 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68493825 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.382 ;
        RECT 0.398 0.248 0.898 0.292 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14688 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 0.074 0.158 1.438 0.202 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.154 0.538 1.222 0.582 ;
        RECT 1.37 0.538 1.438 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
    END
  END vssx
END b15inv040as1n40x5

MACRO b15inv040as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n48x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.1161 LAYER m1 ;
      ANTENNAMAXAREACAR 0.46542625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.618969 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.382 ;
        RECT 0.398 0.248 0.898 0.292 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.566 0.472 ;
        RECT 0.074 0.158 1.566 0.202 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.478 0.248 1.546 0.382 ;
  END
END b15inv040as1n48x5

MACRO b15inv040as1n60x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15inv040as1n60x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.46075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.1089 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60925625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.382 ;
        RECT 0.074 0.248 0.574 0.292 ;
        RECT 0.29 0.248 0.358 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END a
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 0.074 0.158 1.87 0.202 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.158 1.762 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 1.802 0.048 1.87 0.092 ;
    END
  END vssx
END b15inv040as1n60x5

MACRO b15mbn022as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mbn022as1n02x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.383 1.222 0.427 ;
        RECT 1.154 0.158 1.222 0.202 ;
    END
  END o
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.5625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.5625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.403 0.898 0.447 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.046 0.467 1.114 0.511 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
    LAYER v0 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.403 0.79 0.447 ;
      RECT 0.614 0.403 0.682 0.447 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.287 0.466 0.331 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.006 0.338 1.046 0.382 ;
      RECT 1.046 0.158 1.114 0.382 ;
  END
END b15mbn022as1n02x5

MACRO b15mbn022as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mbn022as1n03x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.383 1.222 0.427 ;
        RECT 1.154 0.158 1.222 0.202 ;
    END
  END o
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.16666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.16666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.403 0.898 0.447 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.046 0.467 1.114 0.511 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
    LAYER v0 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.403 0.79 0.447 ;
      RECT 0.614 0.403 0.682 0.447 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.287 0.466 0.331 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.006 0.338 1.046 0.382 ;
      RECT 1.046 0.158 1.114 0.382 ;
  END
END b15mbn022as1n03x5

MACRO b15mbn022as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mbn022as1n04x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.383 1.222 0.427 ;
        RECT 1.154 0.158 1.222 0.202 ;
    END
  END o
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.85 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.85 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.403 0.898 0.447 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.046 0.467 1.114 0.511 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
    LAYER v0 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.403 0.79 0.447 ;
      RECT 0.614 0.403 0.682 0.447 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.287 0.466 0.331 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.006 0.338 1.046 0.382 ;
      RECT 1.046 0.158 1.114 0.382 ;
  END
END b15mbn022as1n04x5

MACRO b15mbn022as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mbn022as1n06x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.383 1.222 0.427 ;
        RECT 1.154 0.158 1.222 0.202 ;
    END
  END o
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.16666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.16666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.403 0.898 0.447 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.046 0.467 1.114 0.511 ;
        RECT 1.262 0.538 1.33 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
    LAYER v0 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.403 0.79 0.447 ;
      RECT 0.614 0.403 0.682 0.447 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.287 0.466 0.331 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.428 0.506 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.006 0.338 1.046 0.382 ;
      RECT 1.046 0.158 1.114 0.382 ;
  END
END b15mbn022as1n06x5

MACRO b15mbn022as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mbn022as1n08x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.448 1.114 0.492 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 1.438 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.37 0.1355 1.438 0.1795 ;
    END
  END o
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.831 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.831 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.088 0.574 0.132 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.478 0.448 1.546 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.1805 0.358 0.2245 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.478 0.1355 1.546 0.1795 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.614 0.158 1.262 0.202 ;
    LAYER v0 ;
      RECT 1.262 0.2705 1.33 0.3145 ;
      RECT 1.154 0.363 1.222 0.407 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.832 0.408 0.896 0.452 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.616 0.268 0.68 0.312 ;
      RECT 0.182 0.1805 0.25 0.2245 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.338 0.614 0.382 ;
      RECT 0.614 0.248 0.682 0.382 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.722 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.562 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.262 0.158 1.33 0.382 ;
  END
END b15mbn022as1n08x5

MACRO b15mbn022as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mbn022as1n12x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 1.6953845 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 1.6953845 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.448 1.114 0.492 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.068 1.762 0.562 ;
        RECT 1.478 0.248 1.762 0.292 ;
        RECT 1.478 0.068 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.478 0.1315 1.546 0.1755 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 1.694 0.1315 1.762 0.1755 ;
    END
  END o
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.158 0.574 0.202 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.586 0.448 1.654 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.178 0.358 0.222 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.586 0.1315 1.654 0.1755 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.614 0.158 1.37 0.202 ;
    LAYER v0 ;
      RECT 1.37 0.2705 1.438 0.3145 ;
      RECT 1.262 0.363 1.33 0.407 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.832 0.408 0.896 0.452 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.616 0.268 0.68 0.312 ;
      RECT 0.616 0.448 0.68 0.492 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.445 0.25 0.489 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.338 0.614 0.382 ;
      RECT 0.614 0.248 0.682 0.382 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.722 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.562 ;
      RECT 1.006 0.248 1.262 0.292 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.37 0.158 1.438 0.382 ;
  END
END b15mbn022as1n12x5

MACRO b15mbn022as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mbn022as1n16x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.3775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.3775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.448 1.114 0.492 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.068 1.762 0.562 ;
        RECT 1.478 0.248 1.762 0.292 ;
        RECT 1.478 0.068 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.478 0.132 1.546 0.176 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 1.694 0.132 1.762 0.176 ;
    END
  END o
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 2.2935715 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 2.2935715 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.158 0.574 0.202 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.178 0.358 0.222 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.586 0.132 1.654 0.176 ;
        RECT 1.802 0.132 1.87 0.176 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.614 0.158 1.37 0.202 ;
    LAYER v0 ;
      RECT 1.37 0.2705 1.438 0.3145 ;
      RECT 1.262 0.363 1.33 0.407 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.832 0.408 0.896 0.452 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.616 0.268 0.68 0.312 ;
      RECT 0.616 0.448 0.68 0.492 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.445 0.25 0.489 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.338 0.614 0.382 ;
      RECT 0.614 0.248 0.682 0.382 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.722 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.562 ;
      RECT 1.006 0.248 1.262 0.292 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.37 0.158 1.438 0.382 ;
  END
END b15mbn022as1n16x5

MACRO b15mbn022as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mbn022as1n24x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.14791675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.14791675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.158 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.408 1.33 0.452 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5553845 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.158 2.302 0.472 ;
        RECT 1.802 0.248 2.302 0.292 ;
        RECT 2.018 0.158 2.086 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.804 0.178 1.868 0.222 ;
        RECT 1.802 0.363 1.87 0.407 ;
        RECT 2.02 0.178 2.084 0.222 ;
        RECT 2.018 0.363 2.086 0.407 ;
        RECT 2.236 0.178 2.3 0.222 ;
        RECT 2.234 0.363 2.302 0.407 ;
    END
  END o
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.71791675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 1.6492 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.694 0.4635 1.762 0.5075 ;
        RECT 1.91 0.4635 1.978 0.5075 ;
        RECT 2.126 0.4635 2.194 0.5075 ;
        RECT 2.342 0.4635 2.41 0.5075 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.722 0.068 0.79 0.292 ;
    LAYER v0 ;
      RECT 1.694 0.2705 1.762 0.3145 ;
      RECT 1.586 0.363 1.654 0.407 ;
      RECT 1.37 0.322 1.438 0.366 ;
      RECT 1.156 0.138 1.22 0.182 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.048 0.408 1.112 0.452 ;
      RECT 0.94 0.138 1.004 0.182 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.832 0.448 0.896 0.492 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.29 0.248 0.358 0.292 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.506 0.472 ;
      RECT 0.182 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.574 0.518 0.722 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.338 0.83 0.382 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.472 ;
      RECT 0.898 0.518 1.154 0.562 ;
      RECT 0.938 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 1.222 0.518 1.37 0.562 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.438 0.248 1.586 0.292 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.006 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.202 ;
      RECT 1.222 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.438 0.158 1.694 0.202 ;
      RECT 1.694 0.158 1.762 0.382 ;
  END
END b15mbn022as1n24x5

MACRO b15mdn022as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mdn022as1n02x3 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.3155 0.898 0.3595 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.562 ;
        RECT 0.398 0.158 0.682 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.614 0.448 0.682 0.492 ;
    END
  END o1
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.8425 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.8425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.448 0.466 0.492 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.83 0.538 0.898 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.83 0.048 0.898 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.722 0.158 0.79 0.562 ;
    LAYER v0 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.29 0.448 0.358 0.492 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.562 ;
  END
END b15mdn022as1n02x3

MACRO b15mdn022as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mdn022as1n02x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 3.35666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 3.35666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.088 0.79 0.132 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.408 0.574 0.452 ;
        RECT 0.506 0.178 0.574 0.222 ;
    END
  END o1
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.86333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 6.954 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.178 0.358 0.222 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.938 0.448 1.006 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.938 0.1355 1.006 0.1795 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.562 ;
    LAYER v0 ;
      RECT 1.046 0.217 1.114 0.261 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.614 0.408 0.682 0.452 ;
      RECT 0.398 0.178 0.466 0.222 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.158 1.114 0.562 ;
  END
END b15mdn022as1n02x5

MACRO b15mdn022as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mdn022as1n03x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.5175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.088 0.79 0.132 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.408 0.574 0.452 ;
        RECT 0.506 0.178 0.574 0.222 ;
    END
  END o1
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.6746155 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 5.795 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.178 0.358 0.222 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.938 0.448 1.006 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.938 0.1355 1.006 0.1795 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.562 ;
    LAYER v0 ;
      RECT 1.046 0.217 1.114 0.261 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.614 0.408 0.682 0.452 ;
      RECT 0.398 0.178 0.466 0.222 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.158 1.114 0.562 ;
  END
END b15mdn022as1n03x5

MACRO b15mdn022as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mdn022as1n04x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.2035 0.682 0.2475 ;
    END
  END o1
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.55769225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.55769225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.318 0.898 0.362 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.262 0.538 1.33 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.181 0.358 0.225 ;
        RECT 1.046 0.178 1.114 0.222 ;
        RECT 1.262 0.048 1.33 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.292 ;
    LAYER v0 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.448 1.222 0.492 ;
      RECT 0.722 0.2035 0.79 0.2475 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.2035 0.574 0.2475 ;
      RECT 0.508 0.408 0.572 0.452 ;
      RECT 0.182 0.181 0.25 0.225 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.506 0.382 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 0.702 0.428 0.938 0.472 ;
      RECT 0.574 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.472 ;
      RECT 1.006 0.338 1.154 0.382 ;
      RECT 1.154 0.158 1.222 0.562 ;
  END
END b15mdn022as1n04x5

MACRO b15mdn022as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mdn022as1n06x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.158 1.546 0.472 ;
      LAYER v0 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.518 1.114 0.562 ;
        RECT 1.046 0.338 1.114 0.562 ;
        RECT 0.83 0.338 0.898 0.562 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.4 0.682 0.444 ;
        RECT 0.83 0.4 0.898 0.444 ;
        RECT 1.046 0.4 1.114 0.444 ;
    END
  END o1
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0171 LAYER m1 ;
      ANTENNAMAXAREACAR 2.17 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0171 LAYER m1 ;
      ANTENNAMAXAREACAR 2.17 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.178 0.574 0.222 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.493 0.358 0.537 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.202 ;
    LAYER v0 ;
      RECT 1.37 0.408 1.438 0.452 ;
      RECT 1.372 0.178 1.436 0.222 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.4 1.006 0.444 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.4 0.79 0.444 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.184 0.408 0.248 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.466 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.472 ;
      RECT 0.79 0.248 0.83 0.292 ;
      RECT 0.83 0.158 0.898 0.292 ;
      RECT 0.898 0.158 1.114 0.202 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 0.79 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.158 1.438 0.472 ;
  END
END b15mdn022as1n06x5

MACRO b15mdn022as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mdn022as1n08x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.248 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.293 1.762 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.292 ;
        RECT 0.614 0.068 1.114 0.112 ;
        RECT 0.83 0.068 0.898 0.382 ;
        RECT 0.614 0.068 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.194 0.682 0.238 ;
        RECT 0.83 0.194 0.898 0.238 ;
        RECT 1.046 0.194 1.114 0.238 ;
    END
  END o1
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.59916675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.59916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.33 0.382 ;
        RECT 1.154 0.248 1.33 0.292 ;
        RECT 1.154 0.068 1.222 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.091 1.222 0.135 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.586 0.538 1.654 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.093 0.358 0.137 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.048 1.654 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.382 ;
    LAYER v0 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 0.938 0.194 1.006 0.238 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.722 0.194 0.79 0.238 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.398 0.178 0.466 0.222 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.338 0.722 0.382 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.79 0.428 1.026 0.472 ;
      RECT 0.702 0.518 1.154 0.562 ;
      RECT 1.006 0.338 1.154 0.382 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.222 0.428 1.37 0.472 ;
      RECT 1.37 0.248 1.438 0.472 ;
      RECT 1.438 0.248 1.478 0.292 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 1.438 0.428 1.586 0.472 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.654 0.428 1.782 0.472 ;
      RECT 1.654 0.158 1.782 0.202 ;
  END
END b15mdn022as1n08x5

MACRO b15mdn022as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mdn022as1n12x5 0 0 ;
  SIZE 2.376 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.382 ;
      LAYER v0 ;
        RECT 2.234 0.293 2.302 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.546 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END o1
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0342 LAYER m1 ;
      ANTENNAMAXAREACAR 2.3614285 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0342 LAYER m1 ;
      ANTENNAMAXAREACAR 2.3614285 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.702 0.518 1.762 0.562 ;
        RECT 1.694 0.338 1.762 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 1.586 0.518 1.654 0.562 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.41 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.538 2.302 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.41 0.022 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.234 0.048 2.302 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.83 0.158 0.898 0.292 ;
    LAYER v0 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.448 2.194 0.492 ;
      RECT 1.91 0.138 1.978 0.182 ;
      RECT 1.91 0.448 1.978 0.492 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.48 0.138 1.544 0.182 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.264 0.138 1.328 0.182 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 1.048 0.178 1.112 0.222 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.832 0.178 0.896 0.222 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 0.682 0.428 1.134 0.472 ;
      RECT 0.682 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.068 1.478 0.112 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 0.898 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 1.242 0.428 1.586 0.472 ;
      RECT 1.114 0.248 1.586 0.292 ;
      RECT 1.586 0.248 1.654 0.472 ;
      RECT 1.654 0.248 1.91 0.292 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 1.978 0.248 2.126 0.292 ;
      RECT 2.126 0.068 2.194 0.562 ;
  END
END b15mdn022as1n12x5

MACRO b15mdn022as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15mdn022as1n16x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.248 2.95 0.382 ;
      LAYER v0 ;
        RECT 2.882 0.293 2.95 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.12546 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.026 0.338 1.978 0.382 ;
        RECT 1.91 0.158 1.978 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.694 0.338 1.762 0.382 ;
        RECT 1.912 0.2645 1.976 0.3085 ;
    END
  END o1
  PIN sa
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 1.82875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 1.82875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.518 2.194 0.562 ;
        RECT 2.126 0.338 2.194 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.518 1.006 0.562 ;
        RECT 2.018 0.518 2.086 0.562 ;
    END
  END sa
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.882 0.538 2.95 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 2.666 0.138 2.734 0.182 ;
        RECT 2.882 0.048 2.95 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.154 0.068 1.222 0.202 ;
    LAYER v0 ;
      RECT 2.774 0.138 2.842 0.182 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.558 0.138 2.626 0.182 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.804 0.178 1.868 0.222 ;
      RECT 1.586 0.248 1.654 0.292 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.372 0.138 1.436 0.182 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.156 0.138 1.22 0.182 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 0.898 0.428 1.458 0.472 ;
      RECT 0.898 0.248 1.802 0.292 ;
      RECT 1.802 0.158 1.87 0.292 ;
      RECT 1.222 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.566 0.428 2.018 0.472 ;
      RECT 1.438 0.068 2.018 0.112 ;
      RECT 2.018 0.068 2.086 0.472 ;
      RECT 2.086 0.248 2.342 0.292 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.41 0.248 2.558 0.292 ;
      RECT 2.558 0.068 2.626 0.562 ;
      RECT 2.626 0.248 2.774 0.292 ;
      RECT 2.774 0.068 2.842 0.562 ;
  END
END b15mdn022as1n16x5

MACRO b15nanb02as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb02as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.113 0.358 0.157 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.466 0.382 ;
        RECT 0.398 0.158 0.466 0.382 ;
        RECT 0.29 0.338 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.468 0.358 0.512 ;
        RECT 0.398 0.253 0.466 0.297 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.468 0.25 0.512 ;
        RECT 0.398 0.468 0.466 0.512 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.182 -0.022 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.253 0.25 0.297 ;
    END
  END vssx
END b15nanb02as1n02x5

MACRO b15nanb02as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb02as1n03x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.574 0.382 ;
        RECT 0.506 0.068 0.574 0.382 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.473 0.466 0.517 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
        RECT 0.506 0.473 0.574 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
END b15nanb02as1n03x5

MACRO b15nanb02as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb02as1n04x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.574 0.382 ;
        RECT 0.506 0.068 0.574 0.382 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.473 0.466 0.517 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
        RECT 0.506 0.473 0.574 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
END b15nanb02as1n04x5

MACRO b15nanb02as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb02as1n06x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.76277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.0073015 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.486 0.068 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.682 0.562 ;
        RECT 0.398 0.338 0.682 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.614 0.448 0.682 0.492 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.184 0.358 0.228 ;
        RECT 0.722 0.184 0.79 0.228 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.074 0.188 0.142 0.232 ;
      RECT 0.074 0.448 0.142 0.492 ;
  END
END b15nanb02as1n06x5

MACRO b15nanb02as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb02as1n08x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.562 ;
        RECT 0.398 0.248 0.79 0.292 ;
        RECT 0.398 0.428 0.682 0.472 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.724 0.428 0.788 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.453 0.25 0.497 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.506 0.112 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.574 0.158 0.918 0.202 ;
  END
END b15nanb02as1n08x5

MACRO b15nanb02as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb02as1n12x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.382 ;
        RECT 0.938 0.248 1.222 0.292 ;
      LAYER v0 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 1.222 0.472 ;
        RECT 0.83 0.248 0.898 0.472 ;
        RECT 0.486 0.248 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.046 0.428 1.114 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.594 0.068 0.722 0.112 ;
    LAYER v0 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.453 0.25 0.497 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.594 0.382 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.79 0.158 1.222 0.202 ;
  END
END b15nanb02as1n12x5

MACRO b15nanb02as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb02as1n16x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.248 1.438 0.472 ;
        RECT 1.134 0.248 1.438 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 1.33 0.472 ;
        RECT 1.262 0.338 1.33 0.472 ;
        RECT 0.938 0.248 1.006 0.472 ;
        RECT 0.486 0.248 1.006 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.264 0.358 1.328 0.402 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.486 0.068 0.83 0.112 ;
    LAYER v0 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.453 0.25 0.497 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.81 0.382 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.158 1.458 0.202 ;
  END
END b15nanb02as1n16x5

MACRO b15nanb02as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb02as1n24x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.87875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.87 0.472 ;
        RECT 1.458 0.248 1.87 0.292 ;
      LAYER v0 ;
        RECT 1.586 0.248 1.654 0.292 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 1.762 0.472 ;
        RECT 1.694 0.338 1.762 0.472 ;
        RECT 1.154 0.248 1.222 0.472 ;
        RECT 0.486 0.248 1.222 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.696 0.358 1.76 0.402 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.486 0.158 1.89 0.202 ;
    LAYER v0 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.453 0.25 0.497 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 1.026 0.382 ;
  END
END b15nanb02as1n24x5

MACRO b15nanb03as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb03as1n02x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.398 0.068 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.562 ;
        RECT 0.398 0.248 0.682 0.292 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.616 0.178 0.68 0.222 ;
        RECT 0.614 0.428 0.682 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.506 0.428 0.574 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.204 0.25 0.248 ;
    END
  END vssx
END b15nanb03as1n02x5

MACRO b15nanb03as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb03as1n03x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.398 0.068 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.562 ;
        RECT 0.398 0.248 0.682 0.292 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.616 0.178 0.68 0.222 ;
        RECT 0.614 0.428 0.682 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.506 0.428 0.574 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
    END
  END vssx
END b15nanb03as1n03x5

MACRO b15nanb03as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb03as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.472 ;
        RECT 0.398 0.068 0.682 0.112 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.3835 0.466 0.4275 ;
        RECT 0.614 0.3835 0.682 0.4275 ;
        RECT 0.614 0.181 0.682 0.225 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 0.506 0.468 0.574 0.512 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
    END
  END vssx
END b15nanb03as1n04x5

MACRO b15nanb03as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb03as1n06x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
        RECT 0.506 0.158 0.79 0.202 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.472 ;
        RECT 0.29 0.068 0.898 0.112 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.83 0.383 0.898 0.427 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03366 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.428 0.682 0.472 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.4505 0.142 0.4945 ;
  END
END b15nanb03as1n06x5

MACRO b15nanb03as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb03as1n08x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 1.006 0.292 ;
        RECT 0.29 0.338 0.466 0.382 ;
        RECT 0.398 0.248 0.466 0.382 ;
        RECT 0.29 0.338 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.382 ;
        RECT 0.938 0.158 1.114 0.202 ;
        RECT 0.938 0.068 1.006 0.202 ;
        RECT 0.506 0.068 1.006 0.112 ;
        RECT 0.29 0.158 0.574 0.202 ;
        RECT 0.506 0.068 0.574 0.202 ;
        RECT 0.29 0.158 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.292 0.228 0.356 0.272 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03978 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 1.006 0.562 ;
        RECT 0.506 0.338 1.006 0.382 ;
        RECT 0.722 0.338 0.79 0.562 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.518 0.142 0.562 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 1.046 0.538 1.114 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
    LAYER v0 ;
      RECT 0.182 0.1475 0.25 0.1915 ;
      RECT 0.182 0.3985 0.25 0.4425 ;
  END
END b15nanb03as1n08x5

MACRO b15nanb03as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb03as1n12x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.596389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.134 0.292 ;
        RECT 0.938 0.248 1.006 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 1.546 0.472 ;
        RECT 1.242 0.248 1.546 0.292 ;
      LAYER v0 ;
        RECT 1.262 0.248 1.33 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.428 1.438 0.472 ;
        RECT 1.37 0.338 1.438 0.472 ;
        RECT 0.486 0.158 0.81 0.202 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.372 0.358 1.436 0.402 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
        RECT 1.154 0.538 1.222 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.486 0.068 1.134 0.112 ;
      RECT 0.918 0.158 1.546 0.202 ;
    LAYER v0 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.182 0.1355 0.25 0.1795 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.248 0.574 0.292 ;
  END
END b15nanb03as1n12x5

MACRO b15nanb03as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nanb03as1n16x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7775925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.548889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.458 0.292 ;
        RECT 1.046 0.248 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.248 1.978 0.472 ;
        RECT 1.566 0.248 1.978 0.292 ;
      LAYER v0 ;
        RECT 1.694 0.248 1.762 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07956 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 1.87 0.472 ;
        RECT 1.802 0.338 1.87 0.472 ;
        RECT 0.486 0.158 0.918 0.202 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.804 0.358 1.868 0.402 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.046 0.538 1.114 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
        RECT 1.694 0.538 1.762 0.582 ;
        RECT 1.91 0.538 1.978 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.486 0.068 1.458 0.112 ;
      RECT 1.026 0.158 1.998 0.202 ;
    LAYER v0 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.136 0.25 0.18 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.248 0.594 0.292 ;
  END
END b15nanb03as1n16x5

MACRO b15nand02as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand02as1n02x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.182 0.4285 0.25 0.4725 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
    END
  END vssx
END b15nand02as1n02x5

MACRO b15nand02as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand02as1n03x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.182 0.428 0.25 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
    END
  END vssx
END b15nand02as1n03x5

MACRO b15nand02as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand02as1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 0.378 0.472 ;
        RECT 0.182 0.068 0.25 0.472 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.29 0.428 0.358 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
    END
  END vssx
END b15nand02as1n04x5

MACRO b15nand02as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand02as1n06x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.448 0.466 0.492 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END vssx
END b15nand02as1n06x5

MACRO b15nand02as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand02as1n08x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3605 0.142 0.4045 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.3605 0.574 0.4045 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.453 0.25 0.497 ;
        RECT 0.182 0.228 0.25 0.272 ;
        RECT 0.398 0.453 0.466 0.497 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.398 0.048 0.466 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.292 0.138 0.356 0.182 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.292 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
  END
END b15nand02as1n08x5

MACRO b15nand02as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand02as1n12x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.79 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.178 0.142 0.222 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.29 0.178 0.358 0.222 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.614 0.428 0.682 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.136 0.682 0.18 ;
      RECT 0.398 0.178 0.466 0.222 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.068 0.682 0.382 ;
  END
END b15nand02as1n12x5

MACRO b15nand02as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand02as1n16x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 1.114 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07956 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.78666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 1.134 0.472 ;
        RECT 0.398 0.158 0.466 0.472 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.182 0.178 0.25 0.222 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.398 0.178 0.466 0.222 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.046 0.428 1.114 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.046 0.136 1.114 0.18 ;
      RECT 0.83 0.136 0.898 0.18 ;
      RECT 0.616 0.138 0.68 0.182 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 0.898 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
  END
END b15nand02as1n16x5

MACRO b15nand02as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand02as1n24x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63973075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.222 0.472 ;
        RECT 0.506 0.158 0.574 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.178 0.142 0.222 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.29 0.178 0.358 0.222 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.506 0.178 0.574 0.222 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.046 0.428 1.114 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.046 0.136 1.114 0.18 ;
      RECT 0.83 0.136 0.898 0.18 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.382 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.068 1.114 0.382 ;
  END
END b15nand02as1n24x5

MACRO b15nand02as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand02as1n32x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6169615 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.338 1.546 0.382 ;
        RECT 1.262 0.248 1.33 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6169615 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.81 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.12852 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.654 0.472 ;
        RECT 1.586 0.068 1.654 0.472 ;
        RECT 0.918 0.068 1.654 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.938 0.068 1.006 0.112 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.154 0.068 1.222 0.112 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.37 0.068 1.438 0.112 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.588 0.138 1.652 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.538 1.654 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.48 0.228 1.544 0.272 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.184 0.228 0.248 0.272 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.292 ;
  END
END b15nand02as1n32x5

MACRO b15nand02as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand02as1n48x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60540175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4056815 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.338 1.978 0.382 ;
        RECT 1.91 0.248 1.978 0.382 ;
        RECT 1.262 0.248 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60540175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4056815 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.79 0.382 ;
        RECT 0.722 0.248 0.79 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.472 ;
        RECT 1.154 0.158 2.086 0.202 ;
        RECT 1.154 0.158 1.222 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.154 0.2455 1.222 0.2895 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.018 0.2455 2.086 0.2895 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
        RECT 1.154 0.538 1.222 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.046 0.2455 1.114 0.2895 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.184 0.228 0.248 0.272 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.158 1.046 0.202 ;
      RECT 1.046 0.068 1.114 0.382 ;
      RECT 1.114 0.068 2.086 0.112 ;
  END
END b15nand02as1n48x5

MACRO b15nand03as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand03as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
        RECT 0.074 0.068 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.068 0.25 0.112 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.466 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.198 0.142 0.242 ;
        RECT 0.29 0.428 0.358 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.398 0.048 0.466 0.092 ;
    END
  END vssx
END b15nand03as1n02x5

MACRO b15nand03as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand03as1n03x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
        RECT 0.074 0.068 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.068 0.25 0.112 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.466 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.198 0.142 0.242 ;
        RECT 0.29 0.428 0.358 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.398 0.048 0.466 0.092 ;
    END
  END vssx
END b15nand03as1n03x5

MACRO b15nand03as1n04x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand03as1n04x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 0.574 0.472 ;
        RECT 0.182 0.068 0.25 0.472 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.398 0.428 0.466 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
END b15nand03as1n04x3

MACRO b15nand03as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand03as1n04x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 0.574 0.472 ;
        RECT 0.182 0.068 0.25 0.472 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.398 0.428 0.466 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
END b15nand03as1n04x5

MACRO b15nand03as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand03as1n06x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.466 0.472 ;
        RECT 0.398 0.248 0.466 0.472 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.158 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.184 0.178 0.248 0.222 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
      LAYER v0 ;
        RECT 0.83 0.048 0.898 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 0.702 0.112 ;
      RECT 0.398 0.158 1.026 0.202 ;
    LAYER v0 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
  END
END b15nand03as1n06x5

MACRO b15nand03as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand03as1n08x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.553426 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.1650695 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.2455 0.466 0.2895 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.006 0.382 ;
        RECT 0.938 0.248 1.006 0.382 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03978 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 1.006 0.472 ;
        RECT 0.182 0.518 0.466 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.184 0.448 0.248 0.492 ;
        RECT 0.182 0.198 0.25 0.242 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
      LAYER v0 ;
        RECT 0.83 0.048 0.898 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 0.702 0.112 ;
    LAYER v0 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.506 0.2455 0.574 0.2895 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.574 0.158 1.026 0.202 ;
  END
END b15nand03as1n08x5

MACRO b15nand03as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand03as1n12x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3670085 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3670085 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.338 1.114 0.382 ;
        RECT 1.046 0.158 1.114 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06426 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 1.114 0.472 ;
        RECT 0.398 0.158 0.466 0.472 ;
        RECT 0.182 0.158 0.466 0.202 ;
        RECT 0.182 0.068 0.25 0.202 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.938 0.428 1.006 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.046 0.538 1.114 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
      LAYER v0 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.938 0.138 1.006 0.182 ;
      RECT 0.724 0.138 0.788 0.182 ;
      RECT 0.508 0.138 0.572 0.182 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
  END
END b15nand03as1n12x5

MACRO b15nand03as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand03as1n16x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.338 0.25 0.382 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.2806535 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.594 0.382 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.28915825 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.81 0.338 1.114 0.382 ;
        RECT 1.046 0.158 1.114 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09486 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.134 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.054 0.158 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.29 0.243 0.358 0.287 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.046 0.428 1.114 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.202 ;
      LAYER v0 ;
        RECT 0.83 0.06 0.898 0.104 ;
        RECT 1.048 0.048 1.112 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.702 0.112 ;
    LAYER v0 ;
      RECT 0.938 0.153 1.006 0.197 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.508 0.178 0.572 0.222 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.292 ;
      RECT 0.574 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
  END
END b15nand03as1n16x5

MACRO b15nand03as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand03as1n24x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.134 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.242 0.338 1.762 0.382 ;
        RECT 1.694 0.158 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.478 0.338 1.546 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.12546 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 1.762 0.472 ;
        RECT 0.182 0.248 0.574 0.292 ;
        RECT 0.506 0.158 0.574 0.292 ;
        RECT 0.398 0.248 0.466 0.472 ;
        RECT 0.182 0.158 0.25 0.292 ;
        RECT 0.054 0.158 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.508 0.178 0.572 0.222 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.586 0.428 1.654 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
        RECT 1.694 0.538 1.762 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
      LAYER v0 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 1.134 0.112 ;
    LAYER v0 ;
      RECT 1.588 0.228 1.652 0.272 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.724 0.228 0.788 0.272 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.292 ;
      RECT 0.79 0.158 1.586 0.202 ;
      RECT 1.586 0.158 1.654 0.292 ;
  END
END b15nand03as1n24x5

MACRO b15nand04as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand04as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.203 0.574 0.247 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.574 0.472 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.048 0.574 0.092 ;
    END
  END vssx
END b15nand04as1n02x5

MACRO b15nand04as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand04as1n03x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.574 0.472 ;
        RECT 0.506 0.068 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.506 0.203 0.574 0.247 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
    END
  END vssx
END b15nand04as1n03x5

MACRO b15nand04as1n04x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand04as1n04x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.118 0.142 0.162 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
END b15nand04as1n04x3

MACRO b15nand04as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand04as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 0.702 0.472 ;
        RECT 0.182 0.068 0.25 0.472 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.614 0.428 0.682 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.614 0.048 0.682 0.092 ;
    END
  END vssx
END b15nand04as1n04x5

MACRO b15nand04as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand04as1n06x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.398 0.158 0.466 0.292 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.23925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.378 0.338 0.574 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.81 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.382 ;
        RECT 0.81 0.248 1.006 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.026 0.472 ;
        RECT 0.074 0.158 0.27 0.202 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.938 0.428 1.006 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
      LAYER v0 ;
        RECT 0.832 0.048 0.896 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 0.466 0.112 ;
    LAYER v0 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.79 0.158 1.026 0.202 ;
  END
END b15nand04as1n06x5

MACRO b15nand04as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand04as1n08x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.43712425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.43712425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.293072 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.918 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.43712425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.026 0.338 1.222 0.382 ;
        RECT 1.154 0.248 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.428 1.222 0.472 ;
        RECT 0.398 0.518 0.682 0.562 ;
        RECT 0.614 0.428 0.682 0.562 ;
        RECT 0.398 0.338 0.466 0.562 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.4535 0.25 0.4975 ;
        RECT 0.182 0.223 0.25 0.267 ;
        RECT 0.4 0.44 0.464 0.484 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.046 0.428 1.114 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
        RECT 1.154 0.538 1.222 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
      LAYER v0 ;
        RECT 1.046 0.048 1.114 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.292 ;
    LAYER v0 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.94 0.138 1.004 0.182 ;
      RECT 0.724 0.138 0.788 0.182 ;
      RECT 0.508 0.138 0.572 0.182 ;
      RECT 0.292 0.138 0.356 0.182 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.358 0.068 0.506 0.112 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 0.79 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 1.114 0.158 1.242 0.202 ;
  END
END b15nand04as1n08x5

MACRO b15nand04as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand04as1n12x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4796445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.381689 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.702 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.381689 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.81 0.338 1.006 0.382 ;
        RECT 0.938 0.158 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4796445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.242 0.338 1.438 0.382 ;
        RECT 1.37 0.158 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08874 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 1.458 0.472 ;
        RECT 0.398 0.248 0.466 0.472 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.158 0.25 0.292 ;
        RECT 0.054 0.158 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.37 0.428 1.438 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.046 0.538 1.114 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
      LAYER v0 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.83 0.068 0.898 0.202 ;
    LAYER v0 ;
      RECT 1.262 0.139 1.33 0.183 ;
      RECT 1.048 0.138 1.112 0.182 ;
      RECT 0.832 0.138 0.896 0.182 ;
      RECT 0.616 0.138 0.68 0.182 ;
      RECT 0.4 0.138 0.464 0.182 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.202 ;
      RECT 0.466 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.898 0.068 1.046 0.112 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.248 1.262 0.292 ;
      RECT 1.262 0.068 1.33 0.292 ;
  END
END b15nand04as1n12x5

MACRO b15nand04as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nand04as1n16x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.378 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4867975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.006 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4867975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.338 1.566 0.382 ;
        RECT 1.262 0.158 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.478 0.338 1.546 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.782 0.338 2.086 0.382 ;
        RECT 2.018 0.248 2.086 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 2.086 0.472 ;
        RECT 0.506 0.158 0.574 0.472 ;
        RECT 0.182 0.158 0.574 0.202 ;
        RECT 0.182 0.158 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.184 0.228 0.248 0.272 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.91 0.428 1.978 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
        RECT 1.154 0.538 1.222 0.582 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.538 1.654 0.582 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.018 0.538 2.086 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
      LAYER v0 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 1.91 0.048 1.978 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.154 0.068 1.222 0.292 ;
    LAYER v0 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.372 0.228 1.436 0.272 ;
      RECT 1.154 0.228 1.222 0.272 ;
      RECT 0.938 0.228 1.006 0.272 ;
      RECT 0.722 0.228 0.79 0.272 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.222 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.438 0.158 2.106 0.202 ;
  END
END b15nand04as1n16x5

MACRO b15nandp2as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp2as1n02x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
        RECT 0.054 0.158 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.182 0.395 0.25 0.439 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
END b15nandp2as1n02x5

MACRO b15nandp2as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp2as1n03x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
        RECT 0.054 0.158 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.182 0.428 0.25 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
END b15nandp2as1n03x5

MACRO b15nandp2as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp2as1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.182 0.428 0.25 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
    END
  END vssx
END b15nandp2as1n04x5

MACRO b15nandp2as1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp2as1n05x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.182 0.428 0.25 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
    END
  END vssx
END b15nandp2as1n05x5

MACRO b15nandp2as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp2as1n08x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.682 0.292 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.574 0.382 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.428 0.79 0.472 ;
        RECT 0.722 0.158 0.79 0.472 ;
        RECT 0.182 0.158 0.79 0.202 ;
        RECT 0.614 0.068 0.682 0.202 ;
        RECT 0.182 0.068 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.184 0.088 0.248 0.132 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.616 0.088 0.68 0.132 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.4 0.048 0.464 0.092 ;
    END
  END vssx
END b15nandp2as1n08x5

MACRO b15nandp2as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp2as1n12x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.79 0.472 ;
        RECT 0.722 0.158 0.79 0.472 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.506 0.178 0.574 0.222 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.722 0.178 0.79 0.222 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.398 0.178 0.466 0.222 ;
      RECT 0.182 0.178 0.25 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.466 0.068 0.79 0.112 ;
  END
END b15nandp2as1n12x5

MACRO b15nandp2as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp2as1n16x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 0.898 0.562 ;
        RECT 0.182 0.338 0.898 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
        RECT 0.398 0.158 0.466 0.562 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.435 0.25 0.479 ;
        RECT 0.182 0.201 0.25 0.245 ;
        RECT 0.398 0.435 0.466 0.479 ;
        RECT 0.398 0.2175 0.466 0.2615 ;
        RECT 0.614 0.435 0.682 0.479 ;
        RECT 0.83 0.435 0.898 0.479 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
      LAYER v0 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.508 0.138 0.572 0.182 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.506 0.112 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.574 0.248 0.83 0.292 ;
      RECT 0.83 0.158 0.898 0.292 ;
      RECT 0.898 0.158 1.026 0.202 ;
  END
END b15nandp2as1n16x5

MACRO b15nandp2as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp2as1n24x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11934 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.222 0.472 ;
        RECT 0.506 0.158 0.574 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.178 0.142 0.222 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.29 0.178 0.358 0.222 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.506 0.178 0.574 0.222 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.046 0.428 1.114 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.382 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.158 1.114 0.382 ;
  END
END b15nandp2as1n24x5

MACRO b15nandp2as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp2as1n32x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.15606 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.938 0.178 1.006 0.222 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.154 0.1785 1.222 0.2225 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.37 0.1785 1.438 0.2225 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.586 0.1785 1.654 0.2225 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.068 0.466 0.382 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.068 0.682 0.382 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.068 0.898 0.382 ;
      RECT 0.898 0.068 1.654 0.112 ;
  END
END b15nandp2as1n32x5

MACRO b15nandp2as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp2as1n48x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.382 ;
      LAYER v0 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49970225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49970225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.23562 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 2.43 0.472 ;
        RECT 2.234 0.158 2.302 0.472 ;
        RECT 2.018 0.158 2.086 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.37 0.178 1.438 0.222 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.586 0.178 1.654 0.222 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.802 0.178 1.87 0.222 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.018 0.178 2.086 0.222 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.234 0.178 2.302 0.222 ;
        RECT 2.342 0.428 2.41 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 2.342 0.068 2.41 0.112 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.398 0.178 0.466 0.222 ;
      RECT 0.182 0.178 0.25 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.382 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.158 0.466 0.382 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.158 1.114 0.382 ;
      RECT 1.114 0.338 1.262 0.382 ;
      RECT 1.262 0.068 1.33 0.382 ;
      RECT 1.33 0.068 2.43 0.112 ;
  END
END b15nandp2as1n48x5

MACRO b15nandp3as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp3as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.466 0.472 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.346 0.142 0.39 ;
        RECT 0.074 0.115 0.142 0.159 ;
        RECT 0.29 0.428 0.358 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.398 0.048 0.466 0.092 ;
    END
  END vssx
END b15nandp3as1n02x5

MACRO b15nandp3as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp3as1n03x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.2255 0.25 0.2695 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.2255 0.466 0.2695 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 0.486 0.472 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.115 0.142 0.159 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.4 0.048 0.464 0.092 ;
    END
  END vssx
END b15nandp3as1n03x5

MACRO b15nandp3as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp3as1n04x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.466 0.112 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.4505 0.25 0.4945 ;
        RECT 0.182 0.15 0.25 0.194 ;
        RECT 0.398 0.4555 0.466 0.4995 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
END b15nandp3as1n04x5

MACRO b15nandp3as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp3as1n08x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.702 0.292 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.382 ;
        RECT 0.81 0.248 1.006 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.428 1.006 0.472 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.182 0.178 0.25 0.222 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
      LAYER v0 ;
        RECT 0.832 0.048 0.896 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 0.702 0.112 ;
      RECT 0.486 0.158 1.026 0.202 ;
    LAYER v0 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
  END
END b15nandp3as1n08x5

MACRO b15nandp3as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp3as1n12x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    ANTENNADIFFAREA 0.08568 LAYER m2 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 1.006 0.562 ;
        RECT 0.722 0.338 0.79 0.562 ;
        RECT 0.506 0.338 0.574 0.562 ;
        RECT 0.29 0.158 0.358 0.562 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER m2 ;
        RECT 0.04 0.428 1.024 0.472 ;
      LAYER v1 ;
        RECT 0.078 0.428 0.138 0.472 ;
        RECT 0.294 0.428 0.354 0.472 ;
        RECT 0.51 0.428 0.57 0.472 ;
        RECT 0.726 0.428 0.786 0.472 ;
        RECT 0.942 0.428 1.002 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.428 0.142 0.472 ;
        RECT 0.074 0.201 0.142 0.245 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.29 0.201 0.358 0.245 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.938 0.428 1.006 0.472 ;
    END
  END o1
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END c
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
      LAYER v0 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.074 0.068 0.702 0.112 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
    LAYER v0 ;
      RECT 0.94 0.228 1.004 0.272 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.938 0.202 ;
      RECT 0.938 0.158 1.006 0.292 ;
  END
END b15nandp3as1n12x5

MACRO b15nandp3as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp3as1n16x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41477125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.574 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41477125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.81 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.50154875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.026 0.338 1.438 0.382 ;
        RECT 1.37 0.158 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1071 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.428 1.438 0.472 ;
        RECT 0.074 0.248 0.378 0.292 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.076 0.178 0.14 0.222 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.262 0.428 1.33 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
      LAYER v0 ;
        RECT 1.046 0.0905 1.114 0.1345 ;
        RECT 1.262 0.0905 1.33 0.1345 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.918 0.112 ;
    LAYER v0 ;
      RECT 1.154 0.0905 1.222 0.1345 ;
      RECT 0.938 0.248 1.006 0.292 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.724 0.178 0.788 0.222 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.292 ;
      RECT 0.79 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.292 ;
  END
END b15nandp3as1n16x5

MACRO b15nandp3as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nandp3as1n24x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.293 1.87 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.17442 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.428 1.89 0.472 ;
        RECT 0.614 0.158 0.682 0.472 ;
        RECT 0.054 0.158 0.682 0.202 ;
        RECT 0.398 0.158 0.466 0.562 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.802 0.428 1.87 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.112 ;
      LAYER v0 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 1.804 0.048 1.868 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.162 0.068 1.33 0.112 ;
    LAYER v0 ;
      RECT 1.694 0.138 1.762 0.182 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.264 0.178 1.328 0.222 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.048 0.178 1.112 0.222 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.832 0.178 0.896 0.222 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.182 0.068 0.25 0.112 ;
    LAYER m1 ;
      RECT 0.83 0.158 0.898 0.292 ;
      RECT 0.898 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.292 ;
      RECT 1.114 0.248 1.262 0.292 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.33 0.248 1.478 0.292 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 1.546 0.248 1.694 0.292 ;
      RECT 1.694 0.068 1.762 0.292 ;
  END
END b15nandp3as1n24x5

MACRO b15nano22as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano22as1n02x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.383 0.358 0.427 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.518 0.702 0.562 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.614 0.518 0.682 0.562 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.4 0.538 0.464 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.498 0.25 0.542 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15nano22as1n02x5

MACRO b15nano22as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano22as1n03x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.383 0.358 0.427 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.518 0.702 0.562 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.614 0.518 0.682 0.562 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.4 0.538 0.464 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.498 0.25 0.542 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15nano22as1n03x5

MACRO b15nano22as1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano22as1n05x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.068 0.142 0.112 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.532 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.432 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.562 ;
        RECT 0.506 0.158 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.722 0.465 0.79 0.509 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.223 0.142 0.267 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.142 0.428 0.614 0.472 ;
      RECT 0.614 0.248 0.682 0.472 ;
  END
END b15nano22as1n05x5

MACRO b15nano22as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano22as1n06x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.383 0.358 0.427 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.603125 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83214275 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.133 0.466 0.177 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 0.898 0.472 ;
        RECT 0.83 0.248 0.898 0.472 ;
        RECT 0.506 0.248 0.898 0.292 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.133 0.574 0.177 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.498 0.142 0.542 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.133 0.358 0.177 ;
        RECT 0.614 0.133 0.682 0.177 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.182 0.498 0.25 0.542 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.248 0.466 0.382 ;
      RECT 0.466 0.338 0.79 0.382 ;
  END
END b15nano22as1n06x5

MACRO b15nano22as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano22as1n08x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.96875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.97916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.498 0.574 0.542 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.114 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.428 1.33 0.562 ;
        RECT 0.722 0.428 1.33 0.472 ;
        RECT 1.154 0.068 1.222 0.472 ;
        RECT 0.722 0.248 1.222 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.264 0.498 1.328 0.542 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.383 0.142 0.427 ;
        RECT 0.29 0.4705 0.358 0.5145 ;
        RECT 0.614 0.498 0.682 0.542 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.1715 0.142 0.2155 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.383 0.25 0.427 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.472 ;
  END
END b15nano22as1n08x5

MACRO b15nano22as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano22as1n12x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.574 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.338 1.762 0.382 ;
        RECT 1.694 0.248 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 1.654 0.292 ;
        RECT 1.586 0.068 1.654 0.292 ;
        RECT 1.37 0.068 1.438 0.292 ;
        RECT 1.046 0.068 1.114 0.472 ;
        RECT 0.83 0.068 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.408 0.898 0.452 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.046 0.408 1.114 0.452 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.694 0.138 1.762 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.518 1.262 0.562 ;
    LAYER v0 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.3155 0.682 0.3595 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.292 0.088 0.356 0.132 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.074 0.428 0.614 0.472 ;
      RECT 0.358 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.33 0.428 1.782 0.472 ;
  END
END b15nano22as1n12x5

MACRO b15nano22as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano22as1n16x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.48081625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7139395 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.248 2.194 0.472 ;
        RECT 1.694 0.248 2.194 0.292 ;
      LAYER v0 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.018 0.248 2.086 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1071 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 2.214 0.202 ;
        RECT 0.938 0.248 1.654 0.292 ;
        RECT 1.586 0.158 1.654 0.292 ;
        RECT 1.37 0.068 1.438 0.472 ;
        RECT 1.154 0.068 1.222 0.472 ;
        RECT 0.938 0.068 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.154 0.408 1.222 0.452 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.158 2.194 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 0.83 0.472 ;
      RECT 0.938 0.518 1.586 0.562 ;
    LAYER v0 ;
      RECT 2.018 0.427 2.086 0.471 ;
      RECT 1.802 0.427 1.87 0.471 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.398 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.562 ;
  END
END b15nano22as1n16x5

MACRO b15nano22as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano22as1n24x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.50276925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.66693875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.248 2.626 0.472 ;
        RECT 1.91 0.248 2.626 0.292 ;
      LAYER v0 ;
        RECT 2.018 0.248 2.086 0.292 ;
        RECT 2.234 0.248 2.302 0.292 ;
        RECT 2.45 0.248 2.518 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14382 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 2.646 0.202 ;
        RECT 1.586 0.248 1.87 0.292 ;
        RECT 1.802 0.158 1.87 0.292 ;
        RECT 1.586 0.068 1.654 0.472 ;
        RECT 0.938 0.338 1.654 0.382 ;
        RECT 1.37 0.068 1.438 0.472 ;
        RECT 1.154 0.068 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.94 0.408 1.004 0.452 ;
        RECT 0.938 0.223 1.006 0.267 ;
        RECT 1.156 0.408 1.22 0.452 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.372 0.408 1.436 0.452 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.588 0.408 1.652 0.452 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.158 2.626 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.91 0.538 1.978 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 0.83 0.472 ;
      RECT 0.938 0.518 1.802 0.562 ;
    LAYER v0 ;
      RECT 2.45 0.429 2.518 0.473 ;
      RECT 2.234 0.429 2.302 0.473 ;
      RECT 2.018 0.429 2.086 0.473 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.398 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.086 0.338 2.234 0.382 ;
      RECT 2.234 0.338 2.302 0.562 ;
      RECT 2.302 0.338 2.45 0.382 ;
      RECT 2.45 0.338 2.518 0.562 ;
  END
END b15nano22as1n24x5

MACRO b15nano23as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano23as1n02x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.518 0.79 0.562 ;
        RECT 0.722 0.068 0.79 0.562 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.724 0.448 0.788 0.492 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.453 0.142 0.497 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.453 0.25 0.497 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15nano23as1n02x5

MACRO b15nano23as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano23as1n03x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.518 0.79 0.562 ;
        RECT 0.722 0.068 0.79 0.562 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.724 0.448 0.788 0.492 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
  END
END b15nano23as1n03x5

MACRO b15nano23as1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano23as1n05x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.292 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.068 0.142 0.112 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
        RECT 0.398 0.158 0.898 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.832 0.088 0.896 0.132 ;
        RECT 0.83 0.464 0.898 0.508 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
      LAYER v0 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.2025 0.142 0.2465 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.142 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.518 0.722 0.562 ;
      RECT 0.722 0.248 0.79 0.562 ;
  END
END b15nano23as1n05x5

MACRO b15nano23as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano23as1n06x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.472 ;
        RECT 0.722 0.248 1.222 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.114 0.382 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03978 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 1.222 0.202 ;
        RECT 0.506 0.428 0.79 0.472 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.158 1.114 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.518 0.83 0.562 ;
    LAYER v0 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.182 0.448 0.25 0.492 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.182 0.112 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.382 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.898 0.428 1.046 0.472 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.114 0.518 1.242 0.562 ;
  END
END b15nano23as1n06x5

MACRO b15nano23as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano23as1n08x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.53875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.35916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.498 0.682 0.542 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.654 0.292 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.478 0.248 1.546 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.89818175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.762 0.382 ;
        RECT 1.694 0.248 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06732 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 1.782 0.202 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.158 1.762 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.383 0.142 0.427 ;
        RECT 0.29 0.4675 0.358 0.5115 ;
        RECT 0.506 0.383 0.574 0.427 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.694 0.478 1.762 0.522 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.162 0.142 0.206 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.518 1.154 0.562 ;
    LAYER v0 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.616 0.228 0.68 0.272 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.383 0.25 0.427 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.222 0.428 1.37 0.472 ;
      RECT 1.37 0.428 1.438 0.562 ;
      RECT 1.438 0.518 1.654 0.562 ;
  END
END b15nano23as1n08x5

MACRO b15nano23as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano23as1n12x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.574 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.248 2.086 0.472 ;
        RECT 1.154 0.248 2.086 0.292 ;
      LAYER v0 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.586 0.248 1.654 0.292 ;
        RECT 1.91 0.248 1.978 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.978 0.382 ;
        RECT 1.046 0.248 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07956 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 2.086 0.202 ;
        RECT 0.722 0.428 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.158 1.978 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.518 1.262 0.562 ;
    LAYER v0 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.292 0.088 0.356 0.132 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.074 0.428 0.614 0.472 ;
      RECT 0.358 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 1.262 0.428 1.33 0.562 ;
      RECT 1.33 0.428 1.91 0.472 ;
      RECT 1.91 0.428 1.978 0.562 ;
      RECT 1.978 0.518 2.106 0.562 ;
  END
END b15nano23as1n12x5

MACRO b15nano23as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano23as1n16x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 1.978 0.292 ;
        RECT 1.478 0.248 1.546 0.472 ;
      LAYER v0 ;
        RECT 1.586 0.248 1.654 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63973075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.248 2.626 0.472 ;
        RECT 2.126 0.248 2.626 0.292 ;
      LAYER v0 ;
        RECT 2.234 0.248 2.302 0.292 ;
        RECT 2.45 0.248 2.518 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.12852 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 2.646 0.202 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.154 0.408 1.222 0.452 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.158 2.626 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.45 0.048 2.518 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 0.83 0.472 ;
      RECT 1.586 0.338 1.654 0.472 ;
      RECT 0.938 0.518 2.086 0.562 ;
    LAYER v0 ;
      RECT 2.452 0.408 2.516 0.452 ;
      RECT 2.236 0.408 2.3 0.452 ;
      RECT 2.02 0.408 2.084 0.452 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.804 0.408 1.868 0.452 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.588 0.408 1.652 0.452 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.398 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.472 ;
      RECT 1.87 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.472 ;
      RECT 2.086 0.338 2.234 0.382 ;
      RECT 2.234 0.338 2.302 0.472 ;
      RECT 2.302 0.338 2.45 0.382 ;
      RECT 2.45 0.338 2.518 0.472 ;
  END
END b15nano23as1n16x5

MACRO b15nano23as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nano23as1n24x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6169615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 2.518 0.292 ;
        RECT 1.802 0.248 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.248 1.978 0.292 ;
        RECT 2.126 0.248 2.194 0.292 ;
        RECT 2.342 0.248 2.41 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6169615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.248 3.382 0.472 ;
        RECT 2.666 0.248 3.382 0.292 ;
      LAYER v0 ;
        RECT 2.774 0.248 2.842 0.292 ;
        RECT 2.99 0.248 3.058 0.292 ;
        RECT 3.206 0.248 3.274 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.17442 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 3.382 0.202 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 0.938 0.338 1.654 0.382 ;
        RECT 1.37 0.068 1.438 0.472 ;
        RECT 1.154 0.068 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.94 0.408 1.004 0.452 ;
        RECT 0.938 0.223 1.006 0.267 ;
        RECT 1.156 0.408 1.22 0.452 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.372 0.408 1.436 0.452 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.588 0.408 1.652 0.452 ;
        RECT 1.588 0.228 1.652 0.272 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 2.774 0.158 2.842 0.202 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.206 0.158 3.274 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.314 0.538 3.382 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.098 0.048 3.166 0.092 ;
        RECT 3.314 0.048 3.382 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 0.83 0.472 ;
      RECT 1.91 0.338 1.978 0.472 ;
      RECT 0.938 0.518 2.626 0.562 ;
    LAYER v0 ;
      RECT 3.208 0.408 3.272 0.452 ;
      RECT 2.992 0.408 3.056 0.452 ;
      RECT 2.776 0.408 2.84 0.452 ;
      RECT 2.56 0.408 2.624 0.452 ;
      RECT 2.45 0.518 2.518 0.562 ;
      RECT 2.344 0.408 2.408 0.452 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.128 0.408 2.192 0.452 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.912 0.408 1.976 0.452 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.4 0.178 0.464 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.398 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 1.978 0.338 2.126 0.382 ;
      RECT 2.126 0.338 2.194 0.472 ;
      RECT 2.194 0.338 2.342 0.382 ;
      RECT 2.342 0.338 2.41 0.472 ;
      RECT 2.41 0.338 2.558 0.382 ;
      RECT 2.558 0.338 2.626 0.472 ;
      RECT 2.626 0.338 2.774 0.382 ;
      RECT 2.774 0.338 2.842 0.472 ;
      RECT 2.842 0.338 2.99 0.382 ;
      RECT 2.99 0.338 3.058 0.472 ;
      RECT 3.058 0.338 3.206 0.382 ;
      RECT 3.206 0.338 3.274 0.472 ;
  END
END b15nano23as1n24x5

MACRO b15nona22as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona22as1n02x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3605 0.142 0.4045 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.3605 0.358 0.4045 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.702 0.202 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.473 0.574 0.517 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.614 0.248 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.473 0.466 0.517 ;
        RECT 0.614 0.473 0.682 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15nona22as1n02x5

MACRO b15nona22as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona22as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.591111 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.702 0.202 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.453 0.574 0.497 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.614 0.248 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.614 0.453 0.682 0.497 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15nona22as1n04x5

MACRO b15nona22as1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona22as1n05x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.432 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.3995 0.574 0.4435 ;
        RECT 0.722 0.184 0.79 0.228 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.722 0.462 0.79 0.506 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.4 0.048 0.464 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.428 0.398 0.472 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
  END
END b15nona22as1n05x5

MACRO b15nona22as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona22as1n08x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
        RECT 0.722 0.248 0.898 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.398 0.068 0.79 0.112 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 0.79 0.562 ;
        RECT 0.506 0.338 0.79 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.614 0.178 0.682 0.222 ;
        RECT 0.722 0.448 0.79 0.492 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.83 0.538 0.898 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.83 0.1105 0.898 0.1545 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15nona22as1n08x5

MACRO b15nona22as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona22as1n12x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.91583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.87375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5301235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3670085 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.33 0.382 ;
        RECT 1.262 0.158 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.702 0.428 1.33 0.472 ;
        RECT 0.83 0.158 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.83 0.228 0.898 0.272 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.594 0.472 ;
      RECT 0.722 0.068 0.79 0.292 ;
    LAYER v0 ;
      RECT 1.154 0.138 1.222 0.182 ;
      RECT 0.94 0.138 1.004 0.182 ;
      RECT 0.722 0.228 0.79 0.272 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.25 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.574 0.338 0.79 0.382 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.068 1.222 0.292 ;
  END
END b15nona22as1n12x5

MACRO b15nona22as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona22as1n16x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.436875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.91583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.202 ;
      LAYER v0 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.378 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.134 0.338 1.438 0.382 ;
        RECT 1.37 0.158 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07038 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.428 1.438 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.228 0.79 0.272 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.938 0.228 1.006 0.272 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.262 0.428 1.33 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.722 0.068 1.046 0.112 ;
    LAYER v0 ;
      RECT 1.262 0.1355 1.33 0.1795 ;
      RECT 1.048 0.138 1.112 0.182 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.508 0.498 0.572 0.542 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.25 0.248 0.614 0.292 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.248 1.262 0.292 ;
      RECT 1.262 0.068 1.33 0.292 ;
  END
END b15nona22as1n16x5

MACRO b15nona22as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona22as1n24x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
        RECT 0.506 0.248 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3732445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.674 0.338 1.978 0.382 ;
        RECT 1.91 0.158 1.978 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.338 1.762 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.428 1.998 0.472 ;
        RECT 1.37 0.248 1.438 0.472 ;
        RECT 0.938 0.248 1.438 0.292 ;
        RECT 1.154 0.248 1.222 0.472 ;
        RECT 0.938 0.248 1.006 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.91 0.428 1.978 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.802 0.538 1.87 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 1.91 0.048 1.978 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.518 0.83 0.562 ;
      RECT 0.83 0.068 1.262 0.112 ;
    LAYER v0 ;
      RECT 1.804 0.228 1.868 0.272 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.616 0.408 0.68 0.452 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.4 0.408 0.464 0.452 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.184 0.408 0.248 0.452 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.472 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.472 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.472 ;
      RECT 0.054 0.158 0.83 0.202 ;
      RECT 0.83 0.158 0.898 0.562 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.158 1.802 0.202 ;
      RECT 1.802 0.158 1.87 0.292 ;
  END
END b15nona22as1n24x5

MACRO b15nona22as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona22as1n32x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
        RECT 0.614 0.248 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.378 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53481475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.39494025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.338 2.518 0.382 ;
        RECT 2.45 0.248 2.518 0.382 ;
      LAYER v0 ;
        RECT 2.126 0.338 2.194 0.382 ;
        RECT 2.342 0.338 2.41 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.428 2.538 0.472 ;
        RECT 1.802 0.248 1.87 0.472 ;
        RECT 1.154 0.248 1.87 0.292 ;
        RECT 1.586 0.248 1.654 0.472 ;
        RECT 1.37 0.248 1.438 0.472 ;
        RECT 1.154 0.248 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.248 1.546 0.292 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.694 0.248 1.762 0.292 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.342 0.428 2.41 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 1.046 0.068 1.694 0.112 ;
    LAYER v0 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.184 0.228 0.248 0.272 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.614 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.682 0.518 1.114 0.562 ;
      RECT 0.25 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.428 1.006 0.472 ;
      RECT 0.574 0.158 1.222 0.202 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 1.762 0.158 2.538 0.202 ;
  END
END b15nona22as1n32x5

MACRO b15nona23as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona23as1n02x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.562 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.722 0.151 0.79 0.195 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.614 0.448 0.682 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15nona23as1n02x5

MACRO b15nona23as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona23as1n04x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.31901225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.562 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.722 0.151 0.79 0.195 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.614 0.538 0.682 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15nona23as1n04x5

MACRO b15nona23as1n05x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona23as1n05x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 0.287111 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.472 ;
        RECT 0.506 0.068 0.898 0.112 ;
        RECT 0.506 0.068 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.408 0.574 0.452 ;
        RECT 0.83 0.408 0.898 0.452 ;
        RECT 0.83 0.154 0.898 0.198 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.722 0.293 0.79 0.337 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.428 0.398 0.472 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.682 0.428 0.722 0.472 ;
      RECT 0.722 0.158 0.79 0.472 ;
  END
END b15nona23as1n05x5

MACRO b15nona23as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona23as1n08x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.242 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.248 1.222 0.292 ;
        RECT 1.154 0.158 1.222 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.486 0.428 1.242 0.472 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.178 0.682 0.222 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.493 0.14 0.537 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.046 0.538 1.114 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.382 ;
    LAYER v0 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.138 0.25 0.182 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.428 0.378 0.472 ;
      RECT 0.574 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.158 1.046 0.202 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.114 0.068 1.242 0.112 ;
  END
END b15nona23as1n08x5

MACRO b15nona23as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona23as1n12x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.91583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.87375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5301235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3670085 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 1.242 0.382 ;
        RECT 0.938 0.248 1.006 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.35 0.338 1.654 0.382 ;
        RECT 1.586 0.158 1.654 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07038 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.702 0.428 1.674 0.472 ;
        RECT 0.83 0.158 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.83 0.228 0.898 0.272 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.586 0.428 1.654 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.588 0.048 1.652 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.594 0.472 ;
      RECT 0.722 0.068 0.79 0.292 ;
      RECT 0.938 0.158 1.154 0.202 ;
    LAYER v0 ;
      RECT 1.478 0.138 1.546 0.182 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.722 0.228 0.79 0.272 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.25 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.574 0.338 0.79 0.382 ;
      RECT 0.79 0.068 1.33 0.112 ;
      RECT 1.154 0.158 1.222 0.292 ;
      RECT 1.222 0.248 1.478 0.292 ;
      RECT 1.478 0.068 1.546 0.292 ;
  END
END b15nona23as1n12x5

MACRO b15nona23as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona23as1n16x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.436875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.91583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.202 ;
      LAYER v0 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.28915825 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.35 0.382 ;
        RECT 1.046 0.158 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.458 0.338 1.762 0.382 ;
        RECT 1.694 0.158 1.762 0.382 ;
      LAYER v0 ;
        RECT 1.478 0.338 1.546 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09486 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.428 1.782 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.228 0.79 0.272 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.938 0.228 1.006 0.272 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.694 0.428 1.762 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 1.154 0.158 1.222 0.292 ;
    LAYER v0 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.156 0.178 1.22 0.222 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.83 0.228 0.898 0.272 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.508 0.498 0.572 0.542 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.25 0.248 0.614 0.292 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.898 0.068 1.35 0.112 ;
      RECT 1.222 0.248 1.586 0.292 ;
      RECT 1.586 0.068 1.654 0.292 ;
  END
END b15nona23as1n16x5

MACRO b15nona23as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona23as1n24x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.14791675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 1.62058825 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.84941175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3732445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.338 1.89 0.382 ;
        RECT 1.37 0.158 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.338 1.654 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63973075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.998 0.338 2.518 0.382 ;
        RECT 2.45 0.158 2.518 0.382 ;
      LAYER v0 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.234 0.338 2.302 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 2.538 0.472 ;
        RECT 1.262 0.158 1.33 0.472 ;
        RECT 1.046 0.158 1.114 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.046 0.228 1.114 0.272 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.262 0.228 1.33 0.272 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.45 0.428 2.518 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.694 0.538 1.762 0.582 ;
        RECT 1.91 0.538 1.978 0.582 ;
        RECT 2.126 0.538 2.194 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.478 0.158 1.546 0.292 ;
    LAYER v0 ;
      RECT 2.344 0.228 2.408 0.272 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.48 0.228 1.544 0.272 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.154 0.228 1.222 0.272 ;
      RECT 0.938 0.228 1.006 0.272 ;
      RECT 0.722 0.408 0.79 0.452 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.616 0.498 0.68 0.542 ;
      RECT 0.506 0.318 0.574 0.362 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.614 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.466 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.574 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.562 ;
      RECT 1.006 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.068 1.89 0.112 ;
      RECT 1.546 0.158 2.342 0.202 ;
      RECT 2.342 0.158 2.41 0.292 ;
  END
END b15nona23as1n24x5

MACRO b15nona23as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nona23as1n32x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.574 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.222 0.382 ;
        RECT 1.046 0.158 1.114 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5556445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0603 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41466 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.338 2.538 0.382 ;
        RECT 1.802 0.158 1.87 0.382 ;
      LAYER v0 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.234 0.338 2.302 0.382 ;
        RECT 2.45 0.338 2.518 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53481475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.39494025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.646 0.338 3.274 0.382 ;
        RECT 3.206 0.248 3.274 0.382 ;
      LAYER v0 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 2.882 0.338 2.95 0.382 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.16524 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.134 0.428 3.274 0.472 ;
        RECT 1.694 0.158 1.762 0.472 ;
        RECT 1.478 0.158 1.546 0.472 ;
        RECT 1.262 0.158 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.262 0.228 1.33 0.272 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.478 0.228 1.546 0.272 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.694 0.228 1.762 0.272 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 3.098 0.428 3.166 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 3.206 0.518 3.274 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
      LAYER v0 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.342 0.538 2.41 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.776 0.538 2.84 0.582 ;
        RECT 2.992 0.538 3.056 0.582 ;
        RECT 3.208 0.538 3.272 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.518 0.398 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.91 0.158 1.978 0.292 ;
    LAYER v0 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 1.912 0.228 1.976 0.272 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.37 0.228 1.438 0.272 ;
      RECT 1.154 0.228 1.222 0.272 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.94 0.228 1.004 0.272 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.338 0.466 0.382 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.184 0.408 0.248 0.452 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.472 ;
      RECT 0.25 0.338 0.614 0.382 ;
      RECT 0.054 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 0.682 0.158 0.938 0.202 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.428 1.026 0.472 ;
      RECT 1.222 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.438 0.068 2.538 0.112 ;
      RECT 1.978 0.158 3.294 0.202 ;
  END
END b15nona23as1n32x5

MACRO b15nonb02as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb02as1n02x3 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.473 0.358 0.517 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
        RECT 0.29 0.248 0.466 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.398 0.372 0.466 0.416 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.372 0.25 0.416 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END vssx
END b15nonb02as1n02x3

MACRO b15nonb02as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb02as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
        RECT 0.398 0.338 0.574 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.506 0.4385 0.574 0.4825 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.074 0.1535 0.142 0.1975 ;
      RECT 0.074 0.448 0.142 0.492 ;
  END
END b15nonb02as1n02x5

MACRO b15nonb02as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb02as1n03x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
        RECT 0.398 0.338 0.574 0.382 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.506 0.4395 0.574 0.4835 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.448 0.142 0.492 ;
  END
END b15nonb02as1n03x5

MACRO b15nonb02as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb02as1n04x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.382 ;
        RECT 0.29 0.248 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.472 ;
        RECT 0.29 0.158 0.898 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.074 0.1245 0.142 0.1685 ;
      RECT 0.076 0.498 0.14 0.542 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.338 0.358 0.472 ;
      RECT 0.358 0.338 0.682 0.382 ;
  END
END b15nonb02as1n04x5

MACRO b15nonb02as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb02as1n06x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.382 ;
        RECT 0.29 0.248 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.472 ;
        RECT 0.29 0.158 0.898 0.202 ;
        RECT 0.506 0.428 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.508 0.498 0.572 0.542 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.074 0.1245 0.142 0.1685 ;
      RECT 0.076 0.498 0.14 0.542 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.338 0.358 0.472 ;
      RECT 0.358 0.338 0.682 0.382 ;
  END
END b15nonb02as1n06x5

MACRO b15nonb02as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb02as1n08x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.898 0.382 ;
        RECT 0.29 0.338 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.562 ;
        RECT 0.506 0.428 1.006 0.472 ;
        RECT 0.29 0.158 1.006 0.202 ;
        RECT 0.506 0.428 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.508 0.498 0.572 0.542 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.94 0.498 1.004 0.542 ;
        RECT 0.94 0.088 1.004 0.132 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.248 0.898 0.292 ;
  END
END b15nonb02as1n08x5

MACRO b15nonb02as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb02as1n12x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.382 ;
        RECT 0.29 0.248 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06732 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 1.222 0.472 ;
        RECT 1.154 0.068 1.222 0.472 ;
        RECT 0.29 0.158 1.222 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.156 0.088 1.22 0.132 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.435 0.25 0.479 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 1.006 0.382 ;
  END
END b15nonb02as1n12x5

MACRO b15nonb02as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb02as1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0315 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 1.546 0.382 ;
        RECT 0.29 0.248 1.546 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09486 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 0.29 0.158 1.654 0.202 ;
      LAYER v0 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.454 0.25 0.498 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 1.438 0.382 ;
  END
END b15nonb02as1n16x5

MACRO b15nonb03as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb03as1n02x3 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.473 0.466 0.517 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.398 0.248 0.682 0.292 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.383 0.682 0.427 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.204 0.25 0.248 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END vssx
END b15nonb03as1n02x3

MACRO b15nonb03as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb03as1n02x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.518 0.25 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.518 0.142 0.562 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 0.594 0.562 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.518 0.574 0.562 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 0.682 0.472 ;
        RECT 0.614 0.068 0.682 0.472 ;
        RECT 0.398 0.248 0.682 0.292 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.616 0.358 0.68 0.402 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END vssx
END b15nonb03as1n02x5

MACRO b15nonb03as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb03as1n03x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 0.682 0.562 ;
        RECT 0.614 0.068 0.682 0.562 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END vssx
END b15nonb03as1n03x5

MACRO b15nonb03as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb03as1n04x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.81 0.382 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 1.006 0.472 ;
        RECT 0.938 0.248 1.006 0.472 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.898 0.292 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.614 0.068 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.938 0.538 1.006 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.1305 0.25 0.1745 ;
        RECT 0.398 0.1355 0.466 0.1795 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.074 0.2305 0.142 0.2745 ;
      RECT 0.074 0.448 0.142 0.492 ;
  END
END b15nonb03as1n04x5

MACRO b15nonb03as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb03as1n06x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.918 0.382 ;
        RECT 0.506 0.338 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.83037025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.428 1.114 0.472 ;
        RECT 1.046 0.248 1.114 0.472 ;
        RECT 0.398 0.518 0.682 0.562 ;
        RECT 0.614 0.428 0.682 0.562 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03978 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 1.006 0.292 ;
        RECT 0.938 0.068 1.006 0.292 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.4505 0.358 0.4945 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.4505 0.25 0.4945 ;
  END
END b15nonb03as1n06x5

MACRO b15nonb03as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb03as1n08x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.596389 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 1.134 0.382 ;
        RECT 0.938 0.248 1.006 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.242 0.338 1.546 0.382 ;
        RECT 1.478 0.068 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.158 1.438 0.292 ;
        RECT 0.614 0.158 1.438 0.202 ;
        RECT 0.486 0.428 0.81 0.472 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.262 0.158 1.33 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.135 0.142 0.179 ;
        RECT 0.29 0.135 0.358 0.179 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.594 0.518 1.134 0.562 ;
      RECT 0.918 0.428 1.546 0.472 ;
    LAYER v0 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.338 0.466 0.382 ;
      RECT 0.182 0.135 0.25 0.179 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.574 0.382 ;
  END
END b15nonb03as1n08x5

MACRO b15nonb03as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nonb03as1n12x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.566 0.382 ;
        RECT 1.154 0.248 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.478 0.338 1.546 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.674 0.338 2.086 0.382 ;
        RECT 2.018 0.158 2.086 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.338 1.762 0.382 ;
        RECT 1.91 0.338 1.978 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 1.978 0.202 ;
        RECT 0.486 0.428 1.006 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.802 0.158 1.87 0.202 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.135 0.142 0.179 ;
        RECT 0.29 0.135 0.358 0.179 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 1.91 0.048 1.978 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.486 0.518 1.566 0.562 ;
      RECT 1.134 0.428 2.106 0.472 ;
    LAYER v0 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.182 0.135 0.25 0.179 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.81 0.382 ;
  END
END b15nonb03as1n12x5

MACRO b15nor002as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor002as1n02x3 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.428 0.378 0.472 ;
        RECT 0.054 0.158 0.378 0.202 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.29 0.158 0.358 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
    END
  END vssx
END b15nor002as1n02x3

MACRO b15nor002as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor002as1n02x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.428 0.378 0.472 ;
        RECT 0.054 0.158 0.378 0.202 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.29 0.158 0.358 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
    END
  END vssx
END b15nor002as1n02x5

MACRO b15nor002as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor002as1n03x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.428 0.358 0.562 ;
        RECT 0.182 0.428 0.358 0.472 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.292 0.498 0.356 0.542 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
END b15nor002as1n03x5

MACRO b15nor002as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor002as1n04x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END vssx
END b15nor002as1n04x5

MACRO b15nor002as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor002as1n06x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2255 0.142 0.2695 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.2255 0.574 0.2695 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.466 0.292 ;
        RECT 0.398 0.068 0.466 0.292 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.363 0.25 0.407 ;
        RECT 0.182 0.133 0.25 0.177 ;
        RECT 0.398 0.133 0.466 0.177 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.133 0.358 0.177 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.292 0.448 0.356 0.492 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.29 0.562 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.338 0.574 0.562 ;
  END
END b15nor002as1n06x5

MACRO b15nor002as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor002as1n08x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.79 0.382 ;
        RECT 0.722 0.248 0.79 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.682 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.428 0.898 0.472 ;
        RECT 0.83 0.158 0.898 0.472 ;
        RECT 0.074 0.158 0.898 0.202 ;
        RECT 0.29 0.428 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.292 0.498 0.356 0.542 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.722 0.428 0.79 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
    END
  END vssx
END b15nor002as1n08x5

MACRO b15nor002as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor002as1n12x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 1.006 0.562 ;
        RECT 0.378 0.338 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
        RECT 0.27 0.248 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 1.114 0.202 ;
        RECT 0.83 0.428 0.898 0.562 ;
        RECT 0.074 0.428 0.898 0.472 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.832 0.498 0.896 0.542 ;
        RECT 0.938 0.158 1.006 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
    END
  END vssx
END b15nor002as1n12x5

MACRO b15nor002as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor002as1n16x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.382 ;
        RECT 0.614 0.248 1.006 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.466 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.518 1.222 0.562 ;
        RECT 1.154 0.158 1.222 0.562 ;
        RECT 0.074 0.158 1.222 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.518 1.006 0.562 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.154 0.428 1.222 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.722 0.382 ;
      RECT 0.722 0.338 0.79 0.472 ;
      RECT 0.79 0.428 1.046 0.472 ;
      RECT 1.046 0.248 1.114 0.472 ;
  END
END b15nor002as1n16x5

MACRO b15nor002as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor002as1n24x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.42741875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56698425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.33 0.382 ;
        RECT 0.83 0.248 1.33 0.292 ;
        RECT 0.83 0.248 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.154 0.248 1.222 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0594 LAYER m1 ;
      ANTENNAMAXAREACAR 0.42094275 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56698425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.382 ;
        RECT 0.074 0.248 0.682 0.292 ;
        RECT 0.398 0.248 0.466 0.382 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.13158 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.518 1.654 0.562 ;
        RECT 1.586 0.158 1.654 0.562 ;
        RECT 0.074 0.158 1.654 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.518 1.006 0.562 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.154 0.518 1.222 0.562 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.37 0.518 1.438 0.562 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.588 0.428 1.652 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.478 0.3405 1.546 0.3845 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.184 0.358 0.248 0.402 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.472 ;
      RECT 0.25 0.428 1.478 0.472 ;
      RECT 1.478 0.248 1.546 0.472 ;
  END
END b15nor002as1n24x5

MACRO b15nor002as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor002as1n32x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.474456 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.70803425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.382 ;
        RECT 1.37 0.248 2.302 0.292 ;
        RECT 2.018 0.248 2.086 0.382 ;
        RECT 1.802 0.248 1.87 0.382 ;
        RECT 1.586 0.248 1.654 0.382 ;
        RECT 1.37 0.248 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.478 0.248 1.546 0.292 ;
        RECT 1.694 0.248 1.762 0.292 ;
        RECT 1.91 0.248 1.978 0.292 ;
        RECT 2.126 0.248 2.194 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4274455 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63788025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.382 ;
        RECT 0.074 0.248 1.222 0.292 ;
        RECT 0.938 0.248 1.006 0.382 ;
        RECT 0.722 0.248 0.79 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.18972 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.518 2.518 0.562 ;
        RECT 2.45 0.158 2.518 0.562 ;
        RECT 0.162 0.158 2.518 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.37 0.518 1.438 0.562 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.586 0.518 1.654 0.562 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.802 0.518 1.87 0.562 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.018 0.518 2.086 0.562 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.234 0.518 2.302 0.562 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.45 0.338 2.518 0.382 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
        RECT 2.234 0.048 2.302 0.092 ;
        RECT 2.45 0.048 2.518 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 2.342 0.338 2.41 0.382 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.184 0.358 0.248 0.402 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.472 ;
      RECT 0.25 0.428 2.342 0.472 ;
      RECT 2.342 0.248 2.41 0.472 ;
  END
END b15nor002as1n32x5

MACRO b15nor003as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor003as1n02x3 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.473 0.466 0.517 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.486 0.202 ;
        RECT 0.074 0.158 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.363 0.142 0.407 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
END b15nor003as1n02x3

MACRO b15nor003as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor003as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.383 0.358 0.427 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.383 0.142 0.427 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.562 ;
        RECT 0.074 0.158 0.466 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.479 0.466 0.523 ;
        RECT 0.398 0.2455 0.466 0.2895 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
END b15nor003as1n02x5

MACRO b15nor003as1n02x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor003as1n02x7 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.484 0.466 0.528 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
END b15nor003as1n02x7

MACRO b15nor003as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor003as1n03x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.64666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.574 0.562 ;
        RECT 0.506 0.068 0.574 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.113 0.25 0.157 ;
        RECT 0.506 0.434 0.574 0.478 ;
        RECT 0.506 0.113 0.574 0.157 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.113 0.142 0.157 ;
        RECT 0.398 0.113 0.466 0.157 ;
    END
  END vssx
END b15nor003as1n03x5

MACRO b15nor003as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor003as1n04x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68158725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.19277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03978 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.4675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.158 0.918 0.202 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.399 0.79 0.443 ;
        RECT 0.83 0.158 0.898 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.406 0.25 0.45 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.4 0.448 0.464 0.492 ;
    LAYER m1 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.518 0.918 0.562 ;
  END
END b15nor003as1n04x5

MACRO b15nor003as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor003as1n06x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 0.477111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0126 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68158725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.472 ;
        RECT 0.506 0.248 0.79 0.292 ;
        RECT 0.506 0.068 0.574 0.292 ;
        RECT 0.074 0.068 0.574 0.112 ;
        RECT 0.29 0.068 0.358 0.382 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.1785 0.142 0.2225 ;
        RECT 0.29 0.176 0.358 0.22 ;
        RECT 0.508 0.1735 0.572 0.2175 ;
        RECT 0.724 0.173 0.788 0.217 ;
        RECT 0.722 0.408 0.79 0.452 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
      LAYER v0 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.682 0.472 ;
      RECT 0.29 0.518 0.918 0.562 ;
    LAYER v0 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
  END
END b15nor003as1n06x5

MACRO b15nor003as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor003as1n08x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.84941175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06426 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 1.242 0.472 ;
        RECT 0.074 0.158 1.242 0.202 ;
        RECT 1.046 0.158 1.114 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.518 1.222 0.562 ;
    LAYER v0 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.616 0.408 0.68 0.452 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.4 0.408 0.464 0.452 ;
      RECT 0.184 0.408 0.248 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.472 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.472 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.472 ;
  END
END b15nor003as1n08x5

MACRO b15nor003as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor003as1n12x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 1.546 0.472 ;
      LAYER v0 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0324 LAYER m1 ;
      ANTENNAMAXAREACAR 0.518395 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 1.566 0.202 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.182 0.338 0.574 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.181 0.25 0.225 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.154 0.408 1.222 0.452 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 1.114 0.472 ;
      RECT 0.506 0.518 1.566 0.562 ;
    LAYER v0 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
  END
END b15nor003as1n12x5

MACRO b15nor003as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor003as1n16x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63973075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.87 0.562 ;
        RECT 1.566 0.248 1.87 0.292 ;
      LAYER v0 ;
        RECT 1.586 0.248 1.654 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 1.026 0.292 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63973075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.12546 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 1.782 0.202 ;
        RECT 1.242 0.428 1.762 0.472 ;
        RECT 1.694 0.338 1.762 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 0.182 0.338 0.574 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.1565 0.25 0.2005 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.696 0.358 1.76 0.402 ;
        RECT 1.694 0.158 1.762 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 1.134 0.472 ;
      RECT 0.614 0.518 1.762 0.562 ;
    LAYER v0 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.428 0.25 0.472 ;
  END
END b15nor003as1n16x5

MACRO b15nor004as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor004as1n02x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.4505 0.574 0.4945 ;
        RECT 0.506 0.1355 0.574 0.1795 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.118 0.25 0.162 ;
        RECT 0.398 0.1355 0.466 0.1795 ;
    END
  END vssx
END b15nor004as1n02x3

MACRO b15nor004as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor004as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.436 0.574 0.48 ;
        RECT 0.506 0.118 0.574 0.162 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.1305 0.25 0.1745 ;
        RECT 0.398 0.118 0.466 0.162 ;
    END
  END vssx
END b15nor004as1n02x5

MACRO b15nor004as1n02x7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor004as1n02x7 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.4955 0.574 0.5395 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.118 0.25 0.162 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END vssx
END b15nor004as1n02x7

MACRO b15nor004as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor004as1n03x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03978 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.682 0.562 ;
        RECT 0.614 0.428 0.682 0.562 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.1355 0.25 0.1795 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.616 0.448 0.68 0.492 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
    END
  END vssx
END b15nor004as1n03x5

MACRO b15nor004as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor004as1n04x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03366 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
      LAYER v0 ;
        RECT 1.046 0.448 1.114 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.832 0.448 0.896 0.492 ;
      RECT 0.4 0.448 0.464 0.492 ;
    LAYER m1 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.518 0.83 0.562 ;
      RECT 0.83 0.428 0.898 0.562 ;
  END
END b15nor004as1n04x5

MACRO b15nor004as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor004as1n06x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.222 0.562 ;
        RECT 1.026 0.338 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.486 0.382 ;
        RECT 0.29 0.338 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.33 0.562 ;
        RECT 0.29 0.248 1.33 0.292 ;
        RECT 0.938 0.068 1.006 0.292 ;
        RECT 0.83 0.248 0.898 0.382 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.83 0.318 0.898 0.362 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.262 0.4555 1.33 0.4995 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.048 0.498 1.112 0.542 ;
      RECT 0.4 0.498 0.464 0.542 ;
    LAYER m1 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.428 1.046 0.472 ;
      RECT 1.046 0.428 1.114 0.562 ;
  END
END b15nor004as1n06x5

MACRO b15nor004as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor004as1n08x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.97359475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.702 0.292 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.472 ;
        RECT 0.938 0.248 1.222 0.292 ;
      LAYER v0 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.84941175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.248 1.654 0.472 ;
        RECT 1.35 0.248 1.654 0.292 ;
      LAYER v0 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08874 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.78666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 1.654 0.202 ;
        RECT 0.398 0.158 0.466 0.472 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.398 0.408 0.466 0.452 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
      LAYER v0 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.538 1.654 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.518 0.81 0.562 ;
      RECT 0.918 0.518 1.262 0.562 ;
    LAYER v0 ;
      RECT 1.48 0.408 1.544 0.452 ;
      RECT 1.264 0.408 1.328 0.452 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.048 0.408 1.112 0.452 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.616 0.408 0.68 0.452 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.29 0.518 0.358 0.562 ;
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.472 ;
      RECT 0.682 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.472 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 1.33 0.338 1.478 0.382 ;
      RECT 1.478 0.338 1.546 0.472 ;
  END
END b15nor004as1n08x5

MACRO b15nor004as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15nor004as1n12x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.918 0.292 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.248 1.654 0.472 ;
        RECT 1.134 0.248 1.654 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.248 2.194 0.382 ;
        RECT 1.802 0.248 2.194 0.292 ;
      LAYER v0 ;
        RECT 1.91 0.248 1.978 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1071 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.158 2.194 0.202 ;
        RECT 0.398 0.158 0.466 0.472 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.338 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.184 0.408 0.248 0.452 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.4 0.408 0.464 0.452 ;
        RECT 0.506 0.158 0.574 0.202 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.018 0.158 2.086 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
      LAYER v0 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.018 0.538 2.086 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 1.91 0.048 1.978 0.092 ;
        RECT 2.126 0.048 2.194 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.518 1.026 0.562 ;
      RECT 1.134 0.518 1.694 0.562 ;
    LAYER v0 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.48 0.408 1.544 0.452 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.264 0.408 1.328 0.452 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.832 0.408 0.896 0.452 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.616 0.408 0.68 0.452 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.614 0.338 0.682 0.472 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.338 1.262 0.382 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.33 0.338 1.478 0.382 ;
      RECT 1.478 0.338 1.546 0.472 ;
      RECT 1.694 0.428 1.762 0.562 ;
      RECT 1.762 0.428 2.214 0.472 ;
  END
END b15nor004as1n12x5

MACRO b15norp02as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp02as1n02x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.157 0.25 0.201 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
END b15norp02as1n02x5

MACRO b15norp02as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp02as1n03x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3605 0.358 0.4045 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.157 0.25 0.201 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
END b15norp02as1n03x5

MACRO b15norp02as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp02as1n04x5 0 0 ;
  SIZE 0.432 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.157 0.25 0.201 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.466 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
    END
  END vssx
END b15norp02as1n04x5

MACRO b15norp02as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp02as1n08x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.596389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.596389 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 0.682 0.472 ;
        RECT 0.614 0.248 0.682 0.472 ;
        RECT 0.182 0.518 0.574 0.562 ;
        RECT 0.506 0.428 0.574 0.562 ;
        RECT 0.182 0.428 0.25 0.562 ;
        RECT 0.074 0.428 0.25 0.472 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.682 0.202 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.408 0.466 0.452 ;
        RECT 0.506 0.158 0.574 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
    END
  END vssx
END b15norp02as1n08x5

MACRO b15norp02as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp02as1n12x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.472 ;
        RECT 0.074 0.158 0.79 0.202 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.506 0.408 0.574 0.452 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.722 0.408 0.79 0.452 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.248 0.466 0.562 ;
      RECT 0.466 0.518 0.79 0.562 ;
  END
END b15norp02as1n12x5

MACRO b15norp02as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp02as1n16x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.898 0.292 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.614 0.068 0.682 0.292 ;
        RECT 0.398 0.068 0.466 0.472 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.385 0.25 0.429 ;
        RECT 0.182 0.151 0.25 0.195 ;
        RECT 0.398 0.3685 0.466 0.4125 ;
        RECT 0.398 0.151 0.466 0.195 ;
        RECT 0.614 0.151 0.682 0.195 ;
        RECT 0.83 0.151 0.898 0.195 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
      LAYER v0 ;
        RECT 0.614 0.538 0.682 0.582 ;
        RECT 0.83 0.538 0.898 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.508 0.448 0.572 0.492 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.506 0.562 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.574 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.428 1.026 0.472 ;
  END
END b15norp02as1n16x5

MACRO b15norp02as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp02as1n24x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11934 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.074 0.158 1.222 0.202 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.722 0.158 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.154 0.408 1.222 0.452 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.614 0.408 0.682 0.452 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 0.682 0.518 1.222 0.562 ;
  END
END b15norp02as1n24x5

MACRO b15norp02as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp02as1n32x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.15606 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 0.074 0.158 1.654 0.202 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.938 0.158 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.154 0.408 1.222 0.452 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.586 0.408 1.654 0.452 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.722 0.408 0.79 0.452 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.614 0.408 0.682 0.452 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 0.898 0.518 1.654 0.562 ;
  END
END b15norp02as1n32x5

MACRO b15norp02as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp02as1n48x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.45269175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.248 2.41 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49970225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0873 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49970225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.23562 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.158 2.43 0.202 ;
        RECT 2.234 0.158 2.302 0.472 ;
        RECT 2.018 0.158 2.086 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.37 0.158 1.438 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.586 0.408 1.654 0.452 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.802 0.408 1.87 0.452 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.018 0.408 2.086 0.452 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.234 0.408 2.302 0.452 ;
        RECT 2.342 0.158 2.41 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 2.342 0.518 2.41 0.562 ;
      RECT 2.126 0.518 2.194 0.562 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.614 0.408 0.682 0.452 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 0.898 0.248 1.046 0.292 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 1.114 0.248 1.262 0.292 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.33 0.518 2.43 0.562 ;
  END
END b15norp02as1n48x5

MACRO b15norp03as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp03as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.383 0.358 0.427 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.383 0.142 0.427 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
        RECT 0.29 0.248 0.466 0.292 ;
        RECT 0.29 0.068 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.398 0.498 0.466 0.542 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.4 0.048 0.464 0.092 ;
    END
  END vssx
END b15norp03as1n02x5

MACRO b15norp03as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp03as1n03x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.486 0.562 ;
        RECT 0.182 0.428 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.518 0.466 0.562 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.383 0.466 0.427 ;
        RECT 0.398 0.1355 0.466 0.1795 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.1355 0.358 0.1795 ;
    END
  END vssx
END b15norp03as1n03x5

MACRO b15norp03as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp03as1n04x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.466 0.562 ;
        RECT 0.398 0.068 0.466 0.562 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.436 0.25 0.48 ;
        RECT 0.182 0.1305 0.25 0.1745 ;
        RECT 0.398 0.15 0.466 0.194 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
END b15norp03as1n04x5

MACRO b15norp03as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp03as1n08x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 1.006 0.202 ;
        RECT 0.83 0.338 0.898 0.472 ;
        RECT 0.722 0.338 0.898 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.832 0.408 0.896 0.452 ;
        RECT 0.83 0.158 0.898 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.518 1.026 0.562 ;
    LAYER v0 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.408 0.574 0.452 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.182 0.472 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.25 0.428 0.466 0.472 ;
      RECT 0.25 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.472 ;
  END
END b15norp03as1n08x5

MACRO b15norp03as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp03as1n12x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.29 0.158 1.222 0.202 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.182 0.338 0.574 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
        RECT 0.182 0.068 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.154 0.408 1.222 0.452 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.428 0.81 0.472 ;
      RECT 0.506 0.518 1.222 0.562 ;
    LAYER v0 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.428 0.358 0.472 ;
  END
END b15norp03as1n12x5

MACRO b15norp03as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp03as1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.382 ;
        RECT 0.83 0.248 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.248 1.654 0.472 ;
        RECT 1.262 0.248 1.654 0.292 ;
      LAYER v0 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 1.654 0.202 ;
        RECT 0.182 0.338 0.79 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
        RECT 0.398 0.068 0.466 0.472 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.184 0.408 0.248 0.452 ;
        RECT 0.182 0.1285 0.25 0.1725 ;
        RECT 0.4 0.408 0.464 0.452 ;
        RECT 0.398 0.1285 0.466 0.1725 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
      LAYER v0 ;
        RECT 1.154 0.538 1.222 0.582 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.538 1.654 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.518 1.026 0.562 ;
    LAYER v0 ;
      RECT 1.48 0.358 1.544 0.402 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.506 0.428 1.478 0.472 ;
      RECT 1.478 0.338 1.546 0.472 ;
  END
END b15norp03as1n16x5

MACRO b15norp03as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15norp03as1n24x5 0 0 ;
  SIZE 2.376 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53481475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53481475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53481475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53481475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 1.546 0.382 ;
        RECT 1.046 0.248 1.546 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.382 ;
        RECT 1.694 0.248 2.302 0.292 ;
      LAYER v0 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.018 0.248 2.086 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14688 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 2.302 0.202 ;
        RECT 0.182 0.338 1.006 0.382 ;
        RECT 0.938 0.158 1.006 0.382 ;
        RECT 0.614 0.068 0.682 0.472 ;
        RECT 0.398 0.068 0.466 0.472 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.184 0.408 0.248 0.452 ;
        RECT 0.182 0.1285 0.25 0.1725 ;
        RECT 0.4 0.408 0.464 0.452 ;
        RECT 0.398 0.1285 0.466 0.1725 ;
        RECT 0.616 0.408 0.68 0.452 ;
        RECT 0.614 0.1285 0.682 0.1725 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.158 2.194 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.41 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
      LAYER v0 ;
        RECT 1.586 0.538 1.654 0.582 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.018 0.538 2.086 0.582 ;
        RECT 2.234 0.538 2.302 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.41 0.022 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.518 1.458 0.562 ;
    LAYER v0 ;
      RECT 2.128 0.358 2.192 0.402 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.37 0.518 1.438 0.562 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.722 0.428 2.126 0.472 ;
      RECT 2.126 0.338 2.194 0.472 ;
  END
END b15norp03as1n24x5

MACRO b15oa0012as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0012as1n02x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0018 LAYER m1 ;
      ANTENNAMAXAREACAR 6.46 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.408 0.466 0.452 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.614 0.448 0.682 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
    LAYER m1 ;
      RECT 0.27 0.518 0.506 0.562 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.562 ;
  END
END b15oa0012as1n02x5

MACRO b15oa0012as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0012as1n03x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0027 LAYER m1 ;
      ANTENNAMAXAREACAR 4.94 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.408 0.466 0.452 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.614 0.448 0.682 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
    LAYER m1 ;
      RECT 0.27 0.518 0.506 0.562 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.158 0.722 0.202 ;
      RECT 0.722 0.158 0.79 0.562 ;
  END
END b15oa0012as1n03x5

MACRO b15oa0012as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0012as1n04x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.436 0.79 0.48 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.378 0.202 ;
    LAYER v0 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.382 ;
  END
END b15oa0012as1n04x5

MACRO b15oa0012as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0012as1n06x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9985185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
        RECT 0.054 0.248 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.4495 0.898 0.4935 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.518 0.142 0.562 ;
        RECT 0.614 0.4505 0.682 0.4945 ;
        RECT 0.938 0.4495 1.006 0.4935 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.338 0.466 0.562 ;
    LAYER v0 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.4 0.228 0.464 0.272 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.398 0.202 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.382 ;
  END
END b15oa0012as1n06x5

MACRO b15oa0012as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0012as1n08x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.25076925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.25076925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.088 0.466 0.132 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.4265 1.114 0.4705 ;
        RECT 1.046 0.138 1.114 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.938 0.4265 1.006 0.4705 ;
        RECT 1.154 0.4265 1.222 0.4705 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.221 0.574 0.265 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 0.29 0.112 ;
    LAYER v0 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.29 0.178 0.358 0.222 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.428 0.378 0.472 ;
      RECT 0.29 0.068 0.358 0.382 ;
      RECT 0.358 0.338 0.614 0.382 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.068 0.898 0.562 ;
  END
END b15oa0012as1n08x5

MACRO b15oa0012as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0012as1n12x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.068 1.654 0.562 ;
        RECT 1.37 0.338 1.654 0.382 ;
        RECT 1.37 0.068 1.438 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.436 1.438 0.48 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.436 1.654 0.48 ;
        RECT 1.586 0.138 1.654 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.046 0.538 1.114 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.722 0.202 ;
      RECT 0.506 0.338 0.574 0.472 ;
    LAYER v0 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.94 0.408 1.004 0.452 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.508 0.408 0.572 0.452 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.518 0.702 0.562 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.79 0.068 1.134 0.112 ;
      RECT 0.574 0.338 0.83 0.382 ;
      RECT 0.83 0.158 0.898 0.382 ;
      RECT 0.898 0.338 0.938 0.382 ;
      RECT 0.938 0.338 1.006 0.472 ;
      RECT 0.898 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.382 ;
  END
END b15oa0012as1n12x5

MACRO b15oa0012as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0012as1n16x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.97359475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.562 ;
        RECT 1.586 0.338 1.87 0.382 ;
        RECT 1.586 0.068 1.654 0.562 ;
      LAYER v0 ;
        RECT 1.586 0.436 1.654 0.48 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 1.802 0.436 1.87 0.48 ;
        RECT 1.802 0.138 1.87 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 1.046 0.538 1.114 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
        RECT 1.694 0.538 1.762 0.582 ;
        RECT 1.91 0.538 1.978 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.83 0.202 ;
      RECT 0.614 0.338 0.682 0.472 ;
    LAYER v0 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.156 0.408 1.22 0.452 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.832 0.408 0.896 0.452 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.616 0.408 0.68 0.452 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.184 0.408 0.248 0.452 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.918 0.562 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.242 0.112 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.472 ;
      RECT 0.898 0.338 0.938 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.006 0.338 1.154 0.382 ;
      RECT 1.154 0.338 1.222 0.472 ;
      RECT 1.006 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
  END
END b15oa0012as1n16x5

MACRO b15oa0012as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0012as1n24x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.87962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.65972225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.248 1.762 0.472 ;
      LAYER v0 ;
        RECT 1.694 0.293 1.762 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.65972225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.65972225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.518 0.562 ;
        RECT 2.018 0.338 2.518 0.382 ;
        RECT 2.234 0.068 2.302 0.562 ;
        RECT 2.018 0.068 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.436 2.086 0.48 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.234 0.436 2.302 0.48 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.45 0.436 2.518 0.48 ;
        RECT 2.45 0.138 2.518 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
        RECT 1.694 0.538 1.762 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 1.154 0.202 ;
      RECT 0.722 0.338 0.79 0.472 ;
    LAYER v0 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.588 0.408 1.652 0.452 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.372 0.408 1.436 0.452 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.94 0.408 1.004 0.452 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.724 0.408 0.788 0.452 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.518 1.134 0.562 ;
      RECT 1.154 0.068 1.222 0.202 ;
      RECT 1.222 0.068 1.782 0.112 ;
      RECT 0.79 0.338 0.938 0.382 ;
      RECT 0.938 0.338 1.006 0.472 ;
      RECT 1.006 0.338 1.262 0.382 ;
      RECT 1.262 0.158 1.33 0.382 ;
      RECT 1.33 0.338 1.37 0.382 ;
      RECT 1.37 0.338 1.438 0.472 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.338 1.654 0.472 ;
      RECT 1.33 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.382 ;
  END
END b15oa0012as1n24x5

MACRO b15oa0012as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0012as1n32x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7139395 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.48081625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.248 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.293 1.978 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.52390025 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.52390025 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11016 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.068 2.842 0.562 ;
        RECT 2.126 0.338 2.842 0.382 ;
        RECT 2.558 0.068 2.626 0.562 ;
        RECT 2.342 0.068 2.41 0.562 ;
        RECT 2.126 0.068 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.436 2.194 0.48 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.342 0.436 2.41 0.48 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.436 2.626 0.48 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.774 0.436 2.842 0.48 ;
        RECT 2.774 0.138 2.842 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 1.262 0.202 ;
      RECT 0.83 0.338 0.898 0.472 ;
    LAYER v0 ;
      RECT 2.018 0.293 2.086 0.337 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.804 0.408 1.868 0.452 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.588 0.408 1.652 0.452 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.264 0.408 1.328 0.452 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.048 0.408 1.112 0.452 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.832 0.408 0.896 0.452 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.4 0.408 0.464 0.452 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.184 0.408 0.248 0.452 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 1.35 0.562 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.068 1.89 0.112 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.472 ;
      RECT 1.114 0.338 1.262 0.382 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.33 0.338 1.37 0.382 ;
      RECT 1.37 0.158 1.438 0.382 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.338 1.654 0.472 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.472 ;
      RECT 1.438 0.158 2.018 0.202 ;
      RECT 2.018 0.158 2.086 0.382 ;
  END
END b15oa0012as1n32x5

MACRO b15oa0022as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0022as1n02x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 0.83 0.178 0.898 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.722 0.448 0.79 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.29 0.178 0.358 0.222 ;
      RECT 0.29 0.408 0.358 0.452 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.25 0.518 0.614 0.562 ;
      RECT 0.614 0.158 0.682 0.562 ;
  END
END b15oa0022as1n02x5

MACRO b15oa0022as1n03x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0022as1n03x3 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 0.83 0.178 0.898 0.222 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.722 0.448 0.79 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.29 0.178 0.358 0.222 ;
      RECT 0.29 0.408 0.358 0.452 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.25 0.518 0.614 0.562 ;
      RECT 0.614 0.158 0.682 0.562 ;
  END
END b15oa0022as1n03x3

MACRO b15oa0022as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0022as1n03x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.4055 0.898 0.4495 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.29 0.178 0.358 0.222 ;
      RECT 0.29 0.408 0.358 0.452 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.25 0.518 0.614 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
  END
END b15oa0022as1n03x5

MACRO b15oa0022as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0022as1n04x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.4055 0.898 0.4495 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.29 0.178 0.358 0.222 ;
      RECT 0.29 0.408 0.358 0.452 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.29 0.112 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.25 0.518 0.614 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
  END
END b15oa0022as1n04x5

MACRO b15oa0022as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0022as1n06x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.451 0.898 0.495 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.938 0.451 1.006 0.495 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.398 0.338 0.466 0.382 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.398 0.112 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 0.25 0.518 0.614 0.562 ;
      RECT 0.614 0.068 0.682 0.562 ;
  END
END b15oa0022as1n06x5

MACRO b15oa0022as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0022as1n08x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.158 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.382 ;
        RECT 0.506 0.248 1.006 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.81 0.382 ;
        RECT 0.614 0.338 0.682 0.472 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.473 0.25 0.517 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.37 0.448 1.438 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.614 0.048 0.682 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.158 0.938 0.202 ;
    LAYER v0 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.372 0.178 1.436 0.222 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.156 0.178 1.22 0.222 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.293 0.358 0.337 ;
    LAYER m1 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.428 0.574 0.562 ;
      RECT 0.574 0.518 0.722 0.562 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 1.154 0.158 1.222 0.292 ;
      RECT 0.79 0.428 1.262 0.472 ;
      RECT 1.222 0.248 1.262 0.292 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.33 0.248 1.37 0.292 ;
      RECT 1.37 0.158 1.438 0.292 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.006 0.068 1.566 0.112 ;
  END
END b15oa0022as1n08x5

MACRO b15oa0022as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0022as1n12x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.486 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.114 0.472 ;
        RECT 0.83 0.338 1.114 0.382 ;
        RECT 0.83 0.338 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 1.134 0.292 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.068 1.654 0.562 ;
        RECT 1.37 0.338 1.654 0.382 ;
        RECT 1.37 0.068 1.438 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.586 0.138 1.654 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
      LAYER v0 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 0.722 0.112 ;
    LAYER v0 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.292 0.498 0.356 0.542 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.614 0.472 ;
      RECT 0.074 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.518 1.154 0.562 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 1.222 0.428 1.262 0.472 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.79 0.158 1.33 0.202 ;
  END
END b15oa0022as1n12x5

MACRO b15oa0022as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0022as1n16x5 0 0 ;
  SIZE 2.376 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.248 1.762 0.562 ;
      LAYER v0 ;
        RECT 1.694 0.293 1.762 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.562 ;
        RECT 1.91 0.248 2.194 0.292 ;
        RECT 1.91 0.068 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.4555 1.978 0.4995 ;
        RECT 1.91 0.138 1.978 0.182 ;
        RECT 2.126 0.4555 2.194 0.4995 ;
        RECT 2.126 0.138 2.194 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.41 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.538 1.654 0.582 ;
        RECT 1.802 0.4555 1.87 0.4995 ;
        RECT 2.018 0.4555 2.086 0.4995 ;
        RECT 2.234 0.4555 2.302 0.4995 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.41 0.022 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.234 0.138 2.302 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.046 0.248 1.114 0.472 ;
      RECT 0.054 0.158 0.83 0.202 ;
      RECT 0.398 0.518 0.938 0.562 ;
    LAYER v0 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.408 1.546 0.452 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.408 0.682 0.452 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.408 0.25 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.248 0.466 0.472 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.248 0.682 0.472 ;
      RECT 1.114 0.248 1.262 0.292 ;
      RECT 1.262 0.248 1.33 0.472 ;
      RECT 1.33 0.248 1.478 0.292 ;
      RECT 1.478 0.248 1.546 0.472 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.674 0.112 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.006 0.518 1.33 0.562 ;
      RECT 1.006 0.158 1.802 0.202 ;
      RECT 1.802 0.158 1.87 0.382 ;
  END
END b15oa0022as1n16x5

MACRO b15oa0022as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0022as1n24x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.89722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.89722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.222 0.562 ;
      LAYER v0 ;
        RECT 1.154 0.408 1.222 0.452 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.65972225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.65972225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.293 2.302 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.89722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.89722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.408 1.114 0.452 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.562 ;
        RECT 2.45 0.248 2.95 0.292 ;
        RECT 2.666 0.068 2.734 0.562 ;
        RECT 2.45 0.068 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.4555 2.518 0.4995 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 2.666 0.4555 2.734 0.4995 ;
        RECT 2.666 0.138 2.734 0.182 ;
        RECT 2.882 0.4555 2.95 0.4995 ;
        RECT 2.882 0.138 2.95 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.018 0.538 2.086 0.582 ;
        RECT 2.342 0.4555 2.41 0.4995 ;
        RECT 2.558 0.4555 2.626 0.4995 ;
        RECT 2.774 0.4555 2.842 0.4995 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 1.046 0.202 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 0.614 0.248 0.682 0.472 ;
    LAYER v0 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.408 1.762 0.452 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.408 1.546 0.452 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.37 0.408 1.438 0.452 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.722 0.408 0.79 0.452 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.408 0.682 0.452 ;
      RECT 0.506 0.408 0.574 0.452 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.182 0.472 ;
      RECT 0.182 0.248 0.25 0.472 ;
      RECT 0.25 0.428 0.466 0.472 ;
      RECT 0.25 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.574 0.518 0.722 0.562 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.114 0.068 2.106 0.112 ;
      RECT 1.33 0.518 1.478 0.562 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.546 0.518 1.694 0.562 ;
      RECT 1.694 0.248 1.762 0.562 ;
      RECT 1.762 0.248 1.91 0.292 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 1.978 0.248 2.126 0.292 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 0.898 0.248 1.154 0.292 ;
      RECT 1.154 0.158 1.222 0.292 ;
      RECT 1.222 0.158 1.37 0.202 ;
      RECT 1.37 0.158 1.438 0.472 ;
      RECT 1.438 0.158 1.586 0.202 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.654 0.158 2.342 0.202 ;
      RECT 2.342 0.158 2.41 0.382 ;
  END
END b15oa0022as1n24x5

MACRO b15oa0022as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oa0022as1n32x5 0 0 ;
  SIZE 3.672 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.67900225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.67900225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.338 1.438 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.408 1.438 0.452 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6596145 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6596145 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.248 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.374 2.734 0.418 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.67900225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.67900225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.338 1.33 0.562 ;
      LAYER v0 ;
        RECT 1.262 0.408 1.33 0.452 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11628 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.598 0.562 ;
        RECT 2.882 0.248 3.598 0.292 ;
        RECT 3.314 0.068 3.382 0.562 ;
        RECT 3.098 0.068 3.166 0.562 ;
        RECT 2.882 0.068 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.4555 2.95 0.4995 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.098 0.4555 3.166 0.4995 ;
        RECT 3.098 0.138 3.166 0.182 ;
        RECT 3.314 0.4555 3.382 0.4995 ;
        RECT 3.314 0.138 3.382 0.182 ;
        RECT 3.53 0.4555 3.598 0.4995 ;
        RECT 3.53 0.138 3.598 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.706 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.774 0.4555 2.842 0.4995 ;
        RECT 2.99 0.4555 3.058 0.4995 ;
        RECT 3.206 0.4555 3.274 0.4995 ;
        RECT 3.422 0.4555 3.49 0.4995 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.706 0.022 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
        RECT 3.206 0.138 3.274 0.182 ;
        RECT 3.422 0.138 3.49 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.586 0.338 1.654 0.562 ;
      RECT 0.074 0.158 1.262 0.202 ;
      RECT 0.722 0.248 0.79 0.472 ;
    LAYER v0 ;
      RECT 2.774 0.293 2.842 0.337 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.342 0.068 2.41 0.112 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.408 1.87 0.452 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.694 0.408 1.762 0.452 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.478 0.408 1.546 0.452 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.722 0.408 0.79 0.452 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.408 0.682 0.452 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.29 0.472 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.358 0.428 0.574 0.472 ;
      RECT 0.358 0.248 0.614 0.292 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.518 1.046 0.562 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 1.654 0.518 1.802 0.562 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 2.018 0.562 ;
      RECT 2.018 0.248 2.086 0.562 ;
      RECT 2.126 0.428 2.342 0.472 ;
      RECT 2.086 0.248 2.342 0.292 ;
      RECT 2.342 0.248 2.41 0.472 ;
      RECT 2.41 0.428 2.626 0.472 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.068 2.646 0.112 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.222 0.248 1.478 0.292 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.546 0.158 1.694 0.202 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.762 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.472 ;
      RECT 1.978 0.158 2.774 0.202 ;
      RECT 2.774 0.158 2.842 0.382 ;
  END
END b15oa0022as1n32x5

MACRO b15oab012as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oab012as1n02x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.3155 0.574 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 0.594 0.562 ;
        RECT 0.398 0.158 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.1985 0.466 0.2425 ;
        RECT 0.506 0.518 0.574 0.562 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.118 0.358 0.162 ;
        RECT 0.506 0.048 0.574 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.1985 0.25 0.2425 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.158 0.25 0.562 ;
  END
END b15oab012as1n02x3

MACRO b15oab012as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oab012as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.3155 0.574 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 0.594 0.562 ;
        RECT 0.398 0.158 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.1985 0.466 0.2425 ;
        RECT 0.506 0.518 0.574 0.562 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.118 0.358 0.162 ;
        RECT 0.506 0.048 0.574 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.1985 0.25 0.2425 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.158 0.25 0.562 ;
  END
END b15oab012as1n02x5

MACRO b15oab012as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oab012as1n03x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.3155 0.574 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 0.594 0.562 ;
        RECT 0.398 0.158 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.1985 0.466 0.2425 ;
        RECT 0.506 0.518 0.574 0.562 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.118 0.358 0.162 ;
        RECT 0.506 0.048 0.574 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.1985 0.25 0.2425 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.158 0.25 0.562 ;
  END
END b15oab012as1n03x5

MACRO b15oab012as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oab012as1n04x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.3155 0.574 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.518 0.682 0.562 ;
        RECT 0.614 0.158 0.682 0.562 ;
        RECT 0.398 0.158 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.1985 0.466 0.2425 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 0.614 0.1985 0.682 0.2425 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.118 0.358 0.162 ;
        RECT 0.506 0.118 0.574 0.162 ;
        RECT 0.722 0.118 0.79 0.162 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.1985 0.25 0.2425 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.158 0.25 0.562 ;
  END
END b15oab012as1n04x5

MACRO b15oab012as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oab012as1n06x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.3155 0.574 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.472 ;
        RECT 0.506 0.428 0.574 0.562 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.1985 0.466 0.2425 ;
        RECT 0.508 0.498 0.572 0.542 ;
        RECT 0.614 0.1985 0.682 0.2425 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.118 0.358 0.162 ;
        RECT 0.506 0.118 0.574 0.162 ;
        RECT 0.722 0.118 0.79 0.162 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.1985 0.25 0.2425 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.158 0.25 0.562 ;
  END
END b15oab012as1n06x5

MACRO b15oab012as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oab012as1n08x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0117 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 3.29925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0081 LAYER m2 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
      ANTENNAMAXAREACAR 4.948889 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER m2 ;
        RECT 0.04 0.428 0.592 0.472 ;
      LAYER v1 ;
        RECT 0.078 0.428 0.138 0.472 ;
        RECT 0.51 0.428 0.57 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
        RECT 0.506 0.3155 0.574 0.3595 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.222 0.472 ;
        RECT 0.81 0.338 1.222 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.4675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.33 0.562 ;
        RECT 0.614 0.248 1.33 0.292 ;
        RECT 0.83 0.068 0.898 0.292 ;
        RECT 0.614 0.518 0.81 0.562 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.1285 0.682 0.1725 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.83 0.1285 0.898 0.1725 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.262 0.458 1.33 0.502 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.128 0.358 0.172 ;
        RECT 0.506 0.1285 0.574 0.1725 ;
        RECT 0.722 0.1285 0.79 0.1725 ;
        RECT 0.938 0.1285 1.006 0.1725 ;
        RECT 1.262 0.048 1.33 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.472 ;
      RECT 0.506 0.248 0.574 0.472 ;
    LAYER v0 ;
      RECT 0.398 0.209 0.466 0.253 ;
      RECT 0.29 0.518 0.358 0.562 ;
    LAYER m1 ;
      RECT 0.27 0.518 0.398 0.562 ;
      RECT 0.398 0.158 0.466 0.562 ;
  END
END b15oab012as1n08x5

MACRO b15oab012as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oab012as1n12x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0144 LAYER m2 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
      ANTENNAMAXAREACAR 2.4744445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
      ANTENNAMAXAREACAR 3.29925925 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.042963 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER m2 ;
        RECT 0.04 0.428 0.592 0.472 ;
      LAYER v1 ;
        RECT 0.078 0.428 0.138 0.472 ;
        RECT 0.51 0.428 0.57 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
        RECT 0.506 0.3155 0.574 0.3595 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.81 0.338 1.242 0.382 ;
        RECT 0.938 0.338 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07038 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.78666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.242 0.518 1.438 0.562 ;
        RECT 1.37 0.068 1.438 0.562 ;
        RECT 0.614 0.248 1.438 0.292 ;
        RECT 1.154 0.068 1.222 0.292 ;
        RECT 0.938 0.068 1.006 0.292 ;
        RECT 0.614 0.518 0.81 0.562 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.262 0.518 1.33 0.562 ;
        RECT 1.37 0.138 1.438 0.182 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.472 ;
      RECT 0.506 0.248 0.574 0.472 ;
    LAYER v0 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.29 0.518 0.358 0.562 ;
    LAYER m1 ;
      RECT 0.27 0.518 0.398 0.562 ;
      RECT 0.398 0.068 0.466 0.562 ;
  END
END b15oab012as1n12x5

MACRO b15oab012as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oab012as1n16x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.63973075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.382 ;
      LAYER v0 ;
        RECT 2.018 0.248 2.086 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.89818175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.682 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.27 0.338 0.79 0.382 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.428 2.106 0.472 ;
        RECT 1.91 0.068 1.978 0.472 ;
        RECT 1.046 0.338 1.978 0.382 ;
        RECT 1.694 0.068 1.762 0.382 ;
        RECT 1.478 0.068 1.546 0.382 ;
        RECT 1.262 0.068 1.33 0.382 ;
        RECT 1.046 0.068 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.586 0.338 1.654 0.382 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 1.802 0.338 1.87 0.382 ;
        RECT 1.91 0.138 1.978 0.182 ;
        RECT 2.018 0.428 2.086 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.018 0.048 2.086 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.938 0.428 1.586 0.472 ;
    LAYER v0 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.428 0.25 0.562 ;
      RECT 0.25 0.428 0.83 0.472 ;
      RECT 0.074 0.158 0.83 0.202 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.654 0.518 1.998 0.562 ;
  END
END b15oab012as1n16x5

MACRO b15oabi12as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oabi12as1n02x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0018 LAYER m1 ;
      ANTENNAMAXAREACAR 5.51 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.498 0.358 0.542 ;
        RECT 0.29 0.1355 0.358 0.1795 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.398 0.386 0.466 0.43 ;
        RECT 0.722 0.538 0.79 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.614 0.048 0.682 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.486 0.158 0.81 0.202 ;
    LAYER v0 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.182 0.1355 0.25 0.1795 ;
      RECT 0.182 0.387 0.25 0.431 ;
  END
END b15oabi12as1n02x5

MACRO b15oabi12as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oabi12as1n03x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.383 0.574 0.427 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 2.204 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.473 0.466 0.517 ;
        RECT 0.398 0.153 0.466 0.197 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.473 0.358 0.517 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.614 0.1855 0.682 0.2295 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.29 0.293 0.358 0.337 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.478 0.142 0.522 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.382 ;
  END
END b15oabi12as1n03x5

MACRO b15oabi12as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oabi12as1n04x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.3155 0.25 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.81 0.382 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.52 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.518 0.574 0.562 ;
        RECT 0.506 0.338 0.574 0.562 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.1355 0.358 0.1795 ;
        RECT 0.506 0.433 0.574 0.477 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4505 0.25 0.4945 ;
        RECT 0.722 0.523 0.79 0.567 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.1355 0.25 0.1795 ;
        RECT 0.614 0.048 0.682 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.722 0.153 0.79 0.197 ;
      RECT 0.506 0.1405 0.574 0.1845 ;
      RECT 0.074 0.2205 0.142 0.2645 ;
      RECT 0.074 0.4505 0.142 0.4945 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.574 0.248 0.722 0.292 ;
      RECT 0.722 0.068 0.79 0.292 ;
  END
END b15oabi12as1n04x5

MACRO b15oabi12as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oabi12as1n06x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.594 0.562 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
        RECT 0.506 0.518 0.574 0.562 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.562 ;
        RECT 0.722 0.068 1.006 0.112 ;
        RECT 0.398 0.248 0.79 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.388 0.466 0.432 ;
        RECT 0.722 0.166 0.79 0.21 ;
        RECT 0.938 0.4505 1.006 0.4945 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4055 0.142 0.4495 ;
        RECT 0.722 0.4055 0.79 0.4495 ;
        RECT 1.046 0.538 1.114 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.292 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.118 0.358 0.162 ;
        RECT 0.506 0.118 0.574 0.162 ;
        RECT 1.262 0.1805 1.33 0.2245 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.1805 1.114 0.2245 ;
    LAYER m1 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.114 0.428 1.242 0.472 ;
  END
END b15oabi12as1n06x5

MACRO b15oabi12as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oabi12as1n08x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 1.006 0.562 ;
        RECT 0.81 0.338 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
        RECT 0.702 0.248 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03366 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 0.898 0.562 ;
        RECT 0.29 0.428 0.898 0.472 ;
        RECT 0.29 0.068 0.594 0.112 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 0.832 0.498 0.896 0.542 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
    LAYER v0 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.4 0.228 0.464 0.272 ;
      RECT 0.182 0.141 0.25 0.185 ;
      RECT 0.182 0.4365 0.25 0.4805 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.158 1.134 0.202 ;
  END
END b15oabi12as1n08x5

MACRO b15oabi12as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oabi12as1n12x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 1.546 0.472 ;
        RECT 0.938 0.338 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 1.35 0.292 ;
        RECT 0.83 0.248 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.154 0.248 1.222 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.518 1.566 0.562 ;
        RECT 1.37 0.428 1.438 0.562 ;
        RECT 0.506 0.428 1.438 0.472 ;
        RECT 1.046 0.428 1.114 0.562 ;
        RECT 0.506 0.068 0.81 0.112 ;
        RECT 0.506 0.068 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.508 0.138 0.572 0.182 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.722 0.068 0.79 0.112 ;
        RECT 1.048 0.498 1.112 0.542 ;
        RECT 1.478 0.518 1.546 0.562 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.292 ;
    LAYER v0 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.616 0.228 0.68 0.272 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.141 0.25 0.185 ;
      RECT 0.182 0.437 0.25 0.481 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.466 0.382 ;
      RECT 0.682 0.158 1.566 0.202 ;
  END
END b15oabi12as1n12x5

MACRO b15oabi12as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oabi12as1n16x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.674 0.382 ;
        RECT 0.83 0.248 0.898 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.478 0.338 1.546 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.87 0.472 ;
        RECT 1.026 0.248 1.87 0.292 ;
      LAYER v0 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.694 0.248 1.762 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 1.674 0.472 ;
        RECT 1.154 0.428 1.222 0.562 ;
        RECT 0.398 0.068 0.918 0.112 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.068 0.898 0.112 ;
        RECT 1.156 0.498 1.22 0.542 ;
        RECT 1.586 0.428 1.654 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.158 0.574 0.292 ;
    LAYER v0 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.508 0.228 0.572 0.272 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.182 0.141 0.25 0.185 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.182 0.472 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.428 0.29 0.472 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.518 0.574 0.562 ;
      RECT 0.574 0.158 1.89 0.202 ;
  END
END b15oabi12as1n16x5

MACRO b15oabi12as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oabi12as1n24x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 2.322 0.382 ;
        RECT 1.046 0.248 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
        RECT 2.234 0.338 2.302 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.248 2.518 0.472 ;
        RECT 1.242 0.248 2.518 0.292 ;
      LAYER v0 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.478 0.248 1.546 0.292 ;
        RECT 1.91 0.248 1.978 0.292 ;
        RECT 2.342 0.248 2.41 0.292 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11016 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.428 2.302 0.562 ;
        RECT 0.614 0.428 2.302 0.472 ;
        RECT 1.802 0.428 1.87 0.562 ;
        RECT 1.37 0.428 1.438 0.562 ;
        RECT 0.614 0.068 1.134 0.112 ;
        RECT 0.614 0.068 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.616 0.1395 0.68 0.1835 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.83 0.068 0.898 0.112 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.068 1.114 0.112 ;
        RECT 1.372 0.498 1.436 0.542 ;
        RECT 1.804 0.498 1.868 0.542 ;
        RECT 2.236 0.498 2.3 0.542 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.292 ;
    LAYER v0 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.724 0.228 0.788 0.272 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.29 0.141 0.358 0.185 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.141 0.142 0.185 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.142 0.428 0.29 0.472 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 0.358 0.428 0.506 0.472 ;
      RECT 0.506 0.248 0.574 0.472 ;
      RECT 0.79 0.158 2.538 0.202 ;
  END
END b15oabi12as1n24x5

MACRO b15oai012as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai012as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.4505 0.466 0.4945 ;
        RECT 0.398 0.153 0.466 0.197 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.4505 0.358 0.4945 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END vssx
END b15oai012as1n02x5

MACRO b15oai012as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai012as1n03x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.383 0.142 0.427 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.466 0.202 ;
        RECT 0.398 0.068 0.466 0.202 ;
        RECT 0.29 0.158 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.4505 0.358 0.4945 ;
        RECT 0.4 0.088 0.464 0.132 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.1305 0.25 0.1745 ;
    END
  END vssx
END b15oai012as1n03x5

MACRO b15oai012as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai012as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.378 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.15333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.486 0.428 0.682 0.472 ;
        RECT 0.614 0.068 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.108 0.682 0.152 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4505 0.142 0.4945 ;
        RECT 0.614 0.538 0.682 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.063 0.358 0.107 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.182 0.15 0.25 0.194 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.068 0.466 0.292 ;
  END
END b15oai012as1n04x5

MACRO b15oai012as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai012as1n06x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.594 0.562 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
        RECT 0.506 0.518 0.574 0.562 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.472 ;
        RECT 0.398 0.248 0.898 0.292 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.408 0.466 0.452 ;
        RECT 0.83 0.4055 0.898 0.4495 ;
        RECT 0.83 0.163 0.898 0.207 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4055 0.142 0.4495 ;
        RECT 0.722 0.4055 0.79 0.4495 ;
        RECT 0.938 0.538 1.006 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.118 0.574 0.162 ;
    END
  END vssx
END b15oai012as1n06x5

MACRO b15oai012as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai012as1n08x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.682 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.358 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04284 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.562 ;
        RECT 0.722 0.158 1.006 0.202 ;
        RECT 0.378 0.518 0.79 0.562 ;
        RECT 0.722 0.158 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.518 0.466 0.562 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.938 0.448 1.006 0.492 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.682 0.472 ;
    LAYER v0 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.506 0.202 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.574 0.068 1.026 0.112 ;
  END
END b15oai012as1n08x5

MACRO b15oai012as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai012as1n12x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 0.79401225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59550925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.291 1.006 0.335 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.382 ;
        RECT 0.182 0.248 0.79 0.292 ;
        RECT 0.182 0.158 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.594 0.382 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05814 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.428 1.114 0.472 ;
        RECT 1.046 0.068 1.114 0.472 ;
        RECT 0.83 0.068 0.898 0.472 ;
        RECT 0.29 0.428 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.292 0.498 0.356 0.542 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.046 0.138 1.114 0.182 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.068 1.024 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.202 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.938 0.068 1.006 0.202 ;
    LAYER v1 ;
      RECT 0.942 0.068 1.002 0.112 ;
      RECT 0.726 0.068 0.786 0.112 ;
      RECT 0.51 0.068 0.57 0.112 ;
      RECT 0.294 0.068 0.354 0.112 ;
      RECT 0.078 0.068 0.138 0.112 ;
    LAYER v0 ;
      RECT 0.938 0.138 1.006 0.182 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.074 0.138 0.142 0.182 ;
  END
END b15oai012as1n12x5

MACRO b15oai012as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai012as1n16x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.158 1.546 0.472 ;
      LAYER v0 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
        RECT 0.594 0.248 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.486 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.158 1.438 0.562 ;
        RECT 1.154 0.338 1.438 0.382 ;
        RECT 0.594 0.518 1.222 0.562 ;
        RECT 1.154 0.158 1.222 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.518 0.682 0.562 ;
        RECT 0.83 0.518 0.898 0.562 ;
        RECT 1.156 0.178 1.22 0.222 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.178 1.438 0.222 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 1.046 0.202 ;
    LAYER v0 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.94 0.358 1.004 0.402 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.938 0.472 ;
      RECT 0.938 0.338 1.006 0.472 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.114 0.068 1.566 0.112 ;
  END
END b15oai012as1n16x5

MACRO b15oai012as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai012as1n24x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.87875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.158 2.194 0.472 ;
      LAYER v0 ;
        RECT 2.126 0.2705 2.194 0.3145 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53481475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53481475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 1.546 0.382 ;
        RECT 1.478 0.158 1.546 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.79 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11016 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.562 ;
        RECT 1.586 0.338 2.086 0.382 ;
        RECT 1.802 0.158 1.87 0.562 ;
        RECT 0.81 0.518 1.654 0.562 ;
        RECT 1.586 0.158 1.654 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.518 0.898 0.562 ;
        RECT 1.046 0.518 1.114 0.562 ;
        RECT 1.262 0.518 1.33 0.562 ;
        RECT 1.478 0.518 1.546 0.562 ;
        RECT 1.586 0.178 1.654 0.222 ;
        RECT 1.802 0.4545 1.87 0.4985 ;
        RECT 1.802 0.178 1.87 0.222 ;
        RECT 2.018 0.4545 2.086 0.4985 ;
        RECT 2.018 0.178 2.086 0.222 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 1.458 0.472 ;
    LAYER v0 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.158 1.37 0.202 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.438 0.068 2.214 0.112 ;
  END
END b15oai012as1n24x5

MACRO b15oai012as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai012as1n32x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.338 2.842 0.382 ;
        RECT 2.774 0.158 2.842 0.382 ;
      LAYER v0 ;
        RECT 2.342 0.338 2.41 0.382 ;
        RECT 2.558 0.338 2.626 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.543611 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.543611 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.026 0.338 1.978 0.382 ;
        RECT 1.91 0.158 1.978 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.694 0.338 1.762 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.918 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14076 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0027 LAYER m1 ;
      ANTENNAMAXAREACAR 3.99 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.428 2.842 0.472 ;
        RECT 2.666 0.158 2.734 0.292 ;
        RECT 2.018 0.158 2.734 0.202 ;
        RECT 1.026 0.518 2.086 0.562 ;
        RECT 2.018 0.158 2.086 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.518 1.114 0.562 ;
        RECT 1.262 0.518 1.33 0.562 ;
        RECT 1.478 0.518 1.546 0.562 ;
        RECT 1.694 0.518 1.762 0.562 ;
        RECT 1.91 0.518 1.978 0.562 ;
        RECT 2.018 0.245 2.086 0.289 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.668 0.228 2.732 0.272 ;
        RECT 2.666 0.428 2.734 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
        RECT 2.776 0.538 2.84 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 1.89 0.472 ;
    LAYER v0 ;
      RECT 2.774 0.068 2.842 0.112 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.342 0.068 2.41 0.112 ;
      RECT 2.126 0.068 2.194 0.112 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.158 1.802 0.202 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 1.87 0.068 2.862 0.112 ;
  END
END b15oai012as1n32x5

MACRO b15oai012as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai012as1n48x5 0 0 ;
  SIZE 4.212 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.8535385 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57791675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.248 4.138 0.472 ;
        RECT 3.422 0.248 4.138 0.292 ;
      LAYER v0 ;
        RECT 3.53 0.248 3.598 0.292 ;
        RECT 3.746 0.248 3.814 0.292 ;
        RECT 3.962 0.248 4.03 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57791675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57791675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.248 2.95 0.472 ;
        RECT 1.478 0.248 2.95 0.292 ;
      LAYER v0 ;
        RECT 1.586 0.248 1.654 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.018 0.248 2.086 0.292 ;
        RECT 2.234 0.248 2.302 0.292 ;
        RECT 2.45 0.248 2.518 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57791675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57791675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 1.33 0.382 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END c
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.20196 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.158 4.138 0.202 ;
        RECT 3.854 0.338 3.922 0.562 ;
        RECT 2.99 0.338 3.922 0.382 ;
        RECT 3.638 0.338 3.706 0.562 ;
        RECT 3.422 0.338 3.49 0.562 ;
        RECT 3.206 0.158 3.274 0.562 ;
        RECT 1.458 0.518 3.058 0.562 ;
        RECT 2.99 0.158 3.058 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.518 1.546 0.562 ;
        RECT 1.694 0.518 1.762 0.562 ;
        RECT 1.91 0.518 1.978 0.562 ;
        RECT 2.126 0.518 2.194 0.562 ;
        RECT 2.342 0.518 2.41 0.562 ;
        RECT 2.558 0.518 2.626 0.562 ;
        RECT 2.882 0.158 2.95 0.202 ;
        RECT 2.99 0.4295 3.058 0.4735 ;
        RECT 3.098 0.158 3.166 0.202 ;
        RECT 3.206 0.4295 3.274 0.4735 ;
        RECT 3.314 0.158 3.382 0.202 ;
        RECT 3.422 0.4295 3.49 0.4735 ;
        RECT 3.53 0.158 3.598 0.202 ;
        RECT 3.638 0.4295 3.706 0.4735 ;
        RECT 3.746 0.158 3.814 0.202 ;
        RECT 3.854 0.4295 3.922 0.4735 ;
        RECT 3.962 0.158 4.03 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.246 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 3.964 0.538 4.028 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.246 0.022 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 2.842 0.472 ;
    LAYER v0 ;
      RECT 4.07 0.068 4.138 0.112 ;
      RECT 3.854 0.068 3.922 0.112 ;
      RECT 3.638 0.068 3.706 0.112 ;
      RECT 3.422 0.068 3.49 0.112 ;
      RECT 3.206 0.068 3.274 0.112 ;
      RECT 2.99 0.068 3.058 0.112 ;
      RECT 2.774 0.068 2.842 0.112 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.158 2.666 0.202 ;
      RECT 2.666 0.068 2.734 0.202 ;
      RECT 2.734 0.068 4.158 0.112 ;
  END
END b15oai012as1n48x5

MACRO b15oai013as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai013as1n02x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.506 0.118 0.574 0.162 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.448 0.466 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
END b15oai013as1n02x3

MACRO b15oai013as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai013as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.574 0.202 ;
        RECT 0.506 0.068 0.574 0.202 ;
        RECT 0.398 0.158 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.4505 0.466 0.4945 ;
        RECT 0.508 0.088 0.572 0.132 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.1355 0.358 0.1795 ;
    END
  END vssx
END b15oai013as1n02x5

MACRO b15oai013as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai013as1n03x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
        RECT 0.074 0.248 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.25 0.562 ;
        RECT 0.054 0.338 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.682 0.382 ;
        RECT 0.614 0.068 0.682 0.382 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.468 0.574 0.512 ;
        RECT 0.614 0.0905 0.682 0.1345 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.526 0.142 0.57 ;
        RECT 0.614 0.468 0.682 0.512 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.108 0.142 0.152 ;
        RECT 0.398 0.048 0.466 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.508 0.228 0.572 0.272 ;
      RECT 0.29 0.158 0.358 0.202 ;
    LAYER m1 ;
      RECT 0.27 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.292 ;
  END
END b15oai013as1n03x5

MACRO b15oai013as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai013as1n04x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.134 0.202 ;
        RECT 0.938 0.158 1.006 0.472 ;
        RECT 0.722 0.248 1.006 0.292 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 1.046 0.158 1.114 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 1.046 0.538 1.114 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.83 0.202 ;
    LAYER v0 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.4 0.448 0.464 0.492 ;
      RECT 0.29 0.158 0.358 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.518 0.83 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.026 0.112 ;
  END
END b15oai013as1n04x5

MACRO b15oai013as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai013as1n06x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.881389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.17518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0459 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.472 ;
        RECT 0.722 0.248 1.114 0.292 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 1.048 0.178 1.112 0.222 ;
        RECT 1.046 0.408 1.114 0.452 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.1805 0.142 0.2245 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.682 0.472 ;
      RECT 0.378 0.518 1.006 0.562 ;
    LAYER v0 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.428 0.142 0.472 ;
  END
END b15oai013as1n06x5

MACRO b15oai013as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai013as1n08x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.158 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.293 1.438 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.596389 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 1.84571425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.81 0.428 1.458 0.472 ;
        RECT 1.262 0.158 1.33 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.262 0.178 1.33 0.222 ;
        RECT 1.37 0.428 1.438 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 0.702 0.472 ;
      RECT 0.486 0.518 1.026 0.562 ;
    LAYER v0 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 0.938 0.15 1.006 0.194 ;
      RECT 0.938 0.518 1.006 0.562 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.184 0.178 0.248 0.222 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.292 ;
      RECT 0.466 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.382 ;
      RECT 0.682 0.158 0.898 0.202 ;
      RECT 0.682 0.338 0.938 0.382 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.006 0.068 1.458 0.112 ;
  END
END b15oai013as1n08x5

MACRO b15oai013as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai013as1n12x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.293 1.87 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.83784725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.11712975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.292 ;
      LAYER v0 ;
        RECT 1.046 0.228 1.114 0.272 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.69534725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.92712975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.228 1.006 0.272 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.158 1.978 0.562 ;
        RECT 1.134 0.428 1.978 0.472 ;
        RECT 1.694 0.158 1.762 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.694 0.178 1.762 0.222 ;
        RECT 1.912 0.498 1.976 0.542 ;
        RECT 1.91 0.178 1.978 0.222 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 1.026 0.472 ;
      RECT 0.594 0.518 1.566 0.562 ;
    LAYER v0 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.382 ;
      RECT 0.25 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.574 0.338 0.722 0.382 ;
      RECT 0.722 0.158 0.79 0.382 ;
      RECT 0.79 0.338 1.262 0.382 ;
      RECT 1.262 0.158 1.33 0.382 ;
      RECT 1.33 0.338 1.478 0.382 ;
      RECT 1.478 0.068 1.546 0.382 ;
      RECT 1.546 0.068 1.978 0.112 ;
  END
END b15oai013as1n12x5

MACRO b15oai022as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai022as1n02x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 0.574 0.562 ;
        RECT 0.398 0.428 0.574 0.472 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.118 0.466 0.162 ;
        RECT 0.508 0.498 0.572 0.542 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.468 0.358 0.512 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END vssx
END b15oai022as1n02x3

MACRO b15oai022as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai022as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.428 0.466 0.472 ;
        RECT 0.398 0.068 0.466 0.472 ;
        RECT 0.29 0.428 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.292 0.498 0.356 0.542 ;
        RECT 0.398 0.153 0.466 0.197 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
    END
  END vssx
END b15oai022as1n02x5

MACRO b15oai022as1n04x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai022as1n04x3 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.518 0.79 0.562 ;
        RECT 0.722 0.158 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.518 0.682 0.562 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.3155 0.898 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.682 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
        RECT 0.506 0.338 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.508 0.408 0.572 0.452 ;
        RECT 0.614 0.2205 0.682 0.2645 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.518 0.142 0.562 ;
        RECT 0.83 0.518 0.898 0.562 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.068 0.358 0.112 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.508 0.138 0.572 0.182 ;
      RECT 0.182 0.163 0.25 0.207 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.25 0.248 0.506 0.292 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.574 0.068 0.898 0.112 ;
  END
END b15oai022as1n04x3

MACRO b15oai022as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai022as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.27 0.518 0.574 0.562 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
        RECT 0.506 0.178 0.574 0.222 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.358 0.068 0.702 0.112 ;
  END
END b15oai022as1n04x5

MACRO b15oai022as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai022as1n06x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.562 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.382 ;
        RECT 0.83 0.068 1.114 0.112 ;
        RECT 0.398 0.518 0.898 0.562 ;
        RECT 0.83 0.068 0.898 0.562 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.42 0.466 0.464 ;
        RECT 0.83 0.4125 0.898 0.4565 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.153 1.114 0.197 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 1.046 0.468 1.114 0.512 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.118 0.358 0.162 ;
        RECT 0.506 0.118 0.574 0.162 ;
    END
  END vssx
END b15oai022as1n06x5

MACRO b15oai022as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai022as1n08x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.114 0.562 ;
        RECT 0.83 0.338 1.114 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.472 ;
        RECT 0.722 0.248 1.222 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.574 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 1.222 0.202 ;
        RECT 0.938 0.428 1.006 0.562 ;
        RECT 0.29 0.428 1.006 0.472 ;
        RECT 0.614 0.158 0.682 0.472 ;
        RECT 0.29 0.428 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.292 0.498 0.356 0.542 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 0.94 0.498 1.004 0.542 ;
        RECT 1.046 0.158 1.114 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.506 0.202 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.574 0.068 1.242 0.112 ;
  END
END b15oai022as1n08x5

MACRO b15oai022as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai022as1n12x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.338 1.546 0.562 ;
        RECT 1.026 0.338 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.248 1.654 0.472 ;
        RECT 1.046 0.248 1.654 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.478 0.248 1.546 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.702 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.682 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 1.566 0.202 ;
        RECT 1.37 0.428 1.438 0.562 ;
        RECT 0.29 0.428 1.438 0.472 ;
        RECT 0.83 0.158 0.898 0.472 ;
        RECT 0.29 0.428 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.292 0.498 0.356 0.542 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.372 0.498 1.436 0.542 ;
        RECT 1.478 0.158 1.546 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.722 0.202 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.79 0.068 1.674 0.112 ;
  END
END b15oai022as1n12x5

MACRO b15oai022as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai022as1n16x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.338 1.978 0.562 ;
        RECT 1.262 0.338 1.978 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.248 2.086 0.472 ;
        RECT 1.154 0.248 2.086 0.292 ;
      LAYER v0 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.586 0.248 1.654 0.292 ;
        RECT 1.91 0.248 1.978 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.898 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 1.006 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.998 0.202 ;
        RECT 1.802 0.428 1.87 0.562 ;
        RECT 0.29 0.428 1.87 0.472 ;
        RECT 1.37 0.428 1.438 0.562 ;
        RECT 1.046 0.158 1.114 0.472 ;
        RECT 0.722 0.428 0.79 0.562 ;
        RECT 0.29 0.428 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.292 0.498 0.356 0.542 ;
        RECT 0.724 0.498 0.788 0.542 ;
        RECT 1.262 0.158 1.33 0.202 ;
        RECT 1.372 0.498 1.436 0.542 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.804 0.498 1.868 0.542 ;
        RECT 1.91 0.158 1.978 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.938 0.202 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.006 0.068 2.106 0.112 ;
  END
END b15oai022as1n16x5

MACRO b15oai022as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai022as1n24x5 0 0 ;
  SIZE 3.024 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.338 2.842 0.562 ;
        RECT 1.694 0.338 2.842 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.338 1.87 0.382 ;
        RECT 2.234 0.338 2.302 0.382 ;
        RECT 2.666 0.338 2.734 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.248 2.95 0.472 ;
        RECT 1.586 0.248 2.95 0.292 ;
      LAYER v0 ;
        RECT 1.694 0.248 1.762 0.292 ;
        RECT 2.018 0.248 2.086 0.292 ;
        RECT 2.45 0.248 2.518 0.292 ;
        RECT 2.774 0.248 2.842 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 1.33 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 1.438 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.262 0.248 1.33 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14688 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.158 2.862 0.202 ;
        RECT 2.666 0.428 2.734 0.562 ;
        RECT 0.29 0.428 2.734 0.472 ;
        RECT 2.234 0.428 2.302 0.562 ;
        RECT 1.802 0.428 1.87 0.562 ;
        RECT 1.478 0.158 1.546 0.472 ;
        RECT 1.154 0.428 1.222 0.562 ;
        RECT 0.722 0.428 0.79 0.562 ;
        RECT 0.29 0.428 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.292 0.498 0.356 0.542 ;
        RECT 0.724 0.498 0.788 0.542 ;
        RECT 1.156 0.498 1.22 0.542 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 1.804 0.498 1.868 0.542 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.236 0.498 2.3 0.542 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 2.668 0.498 2.732 0.542 ;
        RECT 2.774 0.158 2.842 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.058 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.058 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 1.37 0.202 ;
      RECT 1.37 0.068 1.438 0.202 ;
      RECT 1.438 0.068 2.97 0.112 ;
  END
END b15oai022as1n24x5

MACRO b15oai022as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai022as1n32x5 0 0 ;
  SIZE 3.888 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.338 3.706 0.562 ;
        RECT 2.126 0.338 3.706 0.382 ;
      LAYER v0 ;
        RECT 2.234 0.338 2.302 0.382 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 3.098 0.338 3.166 0.382 ;
        RECT 3.53 0.338 3.598 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.746 0.248 3.814 0.472 ;
        RECT 2.018 0.248 3.814 0.292 ;
      LAYER v0 ;
        RECT 2.126 0.248 2.194 0.292 ;
        RECT 2.45 0.248 2.518 0.292 ;
        RECT 2.882 0.248 2.95 0.292 ;
        RECT 3.314 0.248 3.382 0.292 ;
        RECT 3.638 0.248 3.706 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 1.762 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 1.87 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.694 0.248 1.762 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.19584 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.158 3.726 0.202 ;
        RECT 3.53 0.428 3.598 0.562 ;
        RECT 0.29 0.428 3.598 0.472 ;
        RECT 3.098 0.428 3.166 0.562 ;
        RECT 2.666 0.428 2.734 0.562 ;
        RECT 2.234 0.428 2.302 0.562 ;
        RECT 1.91 0.158 1.978 0.472 ;
        RECT 1.586 0.428 1.654 0.562 ;
        RECT 1.154 0.428 1.222 0.562 ;
        RECT 0.722 0.428 0.79 0.562 ;
        RECT 0.29 0.428 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.292 0.498 0.356 0.542 ;
        RECT 0.724 0.498 0.788 0.542 ;
        RECT 1.156 0.498 1.22 0.542 ;
        RECT 1.588 0.498 1.652 0.542 ;
        RECT 2.126 0.158 2.194 0.202 ;
        RECT 2.236 0.498 2.3 0.542 ;
        RECT 2.342 0.158 2.41 0.202 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 2.668 0.498 2.732 0.542 ;
        RECT 2.774 0.158 2.842 0.202 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.1 0.498 3.164 0.542 ;
        RECT 3.206 0.158 3.274 0.202 ;
        RECT 3.422 0.158 3.49 0.202 ;
        RECT 3.532 0.498 3.596 0.542 ;
        RECT 3.638 0.158 3.706 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.922 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.748 0.538 3.812 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.922 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 3.746 0.068 3.814 0.112 ;
      RECT 3.53 0.068 3.598 0.112 ;
      RECT 3.314 0.068 3.382 0.112 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 2.882 0.068 2.95 0.112 ;
      RECT 2.666 0.068 2.734 0.112 ;
      RECT 2.45 0.068 2.518 0.112 ;
      RECT 2.234 0.068 2.302 0.112 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 1.802 0.202 ;
      RECT 1.802 0.068 1.87 0.202 ;
      RECT 1.87 0.068 3.834 0.112 ;
  END
END b15oai022as1n32x5

MACRO b15oai022as1n48x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai022as1n48x5 0 0 ;
  SIZE 5.616 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.366 0.338 5.434 0.562 ;
        RECT 2.99 0.338 5.434 0.382 ;
      LAYER v0 ;
        RECT 3.098 0.338 3.166 0.382 ;
        RECT 3.53 0.338 3.598 0.382 ;
        RECT 3.962 0.338 4.03 0.382 ;
        RECT 4.394 0.338 4.462 0.382 ;
        RECT 4.826 0.338 4.894 0.382 ;
        RECT 5.258 0.338 5.326 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.474 0.248 5.542 0.472 ;
        RECT 2.882 0.248 5.542 0.292 ;
      LAYER v0 ;
        RECT 2.99 0.248 3.058 0.292 ;
        RECT 3.314 0.248 3.382 0.292 ;
        RECT 3.746 0.248 3.814 0.292 ;
        RECT 4.178 0.248 4.246 0.292 ;
        RECT 4.61 0.248 4.678 0.292 ;
        RECT 5.042 0.248 5.11 0.292 ;
        RECT 5.366 0.248 5.434 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 2.626 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.586 0.338 1.654 0.382 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.45 0.338 2.518 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 2.734 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.234 0.248 2.302 0.292 ;
        RECT 2.558 0.248 2.626 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.29376 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.158 5.454 0.202 ;
        RECT 5.258 0.428 5.326 0.562 ;
        RECT 0.29 0.428 5.326 0.472 ;
        RECT 4.826 0.428 4.894 0.562 ;
        RECT 4.394 0.428 4.462 0.562 ;
        RECT 3.962 0.428 4.03 0.562 ;
        RECT 3.53 0.428 3.598 0.562 ;
        RECT 3.098 0.428 3.166 0.562 ;
        RECT 2.774 0.158 2.842 0.472 ;
        RECT 2.45 0.428 2.518 0.562 ;
        RECT 2.018 0.428 2.086 0.562 ;
        RECT 1.586 0.428 1.654 0.562 ;
        RECT 1.154 0.428 1.222 0.562 ;
        RECT 0.722 0.428 0.79 0.562 ;
        RECT 0.29 0.428 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.292 0.498 0.356 0.542 ;
        RECT 0.724 0.498 0.788 0.542 ;
        RECT 1.156 0.498 1.22 0.542 ;
        RECT 1.588 0.498 1.652 0.542 ;
        RECT 2.02 0.498 2.084 0.542 ;
        RECT 2.452 0.498 2.516 0.542 ;
        RECT 2.99 0.158 3.058 0.202 ;
        RECT 3.1 0.498 3.164 0.542 ;
        RECT 3.206 0.158 3.274 0.202 ;
        RECT 3.422 0.158 3.49 0.202 ;
        RECT 3.532 0.498 3.596 0.542 ;
        RECT 3.638 0.158 3.706 0.202 ;
        RECT 3.854 0.158 3.922 0.202 ;
        RECT 3.964 0.498 4.028 0.542 ;
        RECT 4.07 0.158 4.138 0.202 ;
        RECT 4.286 0.158 4.354 0.202 ;
        RECT 4.396 0.498 4.46 0.542 ;
        RECT 4.502 0.158 4.57 0.202 ;
        RECT 4.718 0.158 4.786 0.202 ;
        RECT 4.828 0.498 4.892 0.542 ;
        RECT 4.934 0.158 5.002 0.202 ;
        RECT 5.15 0.158 5.218 0.202 ;
        RECT 5.26 0.498 5.324 0.542 ;
        RECT 5.366 0.158 5.434 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.65 0.652 ;
        RECT 5.474 0.518 5.542 0.652 ;
        RECT 5.042 0.518 5.11 0.652 ;
        RECT 4.61 0.518 4.678 0.652 ;
        RECT 4.178 0.518 4.246 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.316 0.538 3.38 0.582 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 4.18 0.538 4.244 0.582 ;
        RECT 4.612 0.538 4.676 0.582 ;
        RECT 5.044 0.538 5.108 0.582 ;
        RECT 5.476 0.538 5.54 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.65 0.022 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 5.474 0.068 5.542 0.112 ;
      RECT 5.258 0.068 5.326 0.112 ;
      RECT 5.042 0.068 5.11 0.112 ;
      RECT 4.826 0.068 4.894 0.112 ;
      RECT 4.61 0.068 4.678 0.112 ;
      RECT 4.394 0.068 4.462 0.112 ;
      RECT 4.178 0.068 4.246 0.112 ;
      RECT 3.962 0.068 4.03 0.112 ;
      RECT 3.746 0.068 3.814 0.112 ;
      RECT 3.53 0.068 3.598 0.112 ;
      RECT 3.314 0.068 3.382 0.112 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 2.774 0.068 2.842 0.112 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 2.666 0.202 ;
      RECT 2.666 0.068 2.734 0.202 ;
      RECT 2.734 0.068 5.562 0.112 ;
  END
END b15oai022as1n48x5

MACRO b15oai112as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai112as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.594 0.112 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.574 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.506 0.2205 0.574 0.2645 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.1355 0.25 0.1795 ;
    END
  END vssx
END b15oai112as1n02x5

MACRO b15oai112as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai112as1n04x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.383 0.466 0.427 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03366 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 2.204 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.562 ;
        RECT 0.506 0.068 0.79 0.112 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.478 0.574 0.522 ;
        RECT 0.722 0.478 0.79 0.522 ;
        RECT 0.722 0.153 0.79 0.197 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.526 0.142 0.57 ;
        RECT 0.614 0.478 0.682 0.522 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.4 0.088 0.464 0.132 ;
      RECT 0.074 0.24 0.142 0.284 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.382 ;
      RECT 0.142 0.158 0.398 0.202 ;
      RECT 0.398 0.068 0.466 0.202 ;
  END
END b15oai112as1n04x5

MACRO b15oai112as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai112as1n06x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.382 ;
        RECT 0.506 0.068 1.006 0.112 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.383 0.574 0.427 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03978 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 9.0725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.428 1.026 0.472 ;
        RECT 0.722 0.158 0.79 0.472 ;
        RECT 0.614 0.428 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.616 0.498 0.68 0.542 ;
        RECT 0.722 0.1835 0.79 0.2275 ;
        RECT 0.938 0.428 1.006 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END vssx
END b15oai112as1n06x5

MACRO b15oai112as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai112as1n08x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.522639 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7613195 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.358 0.79 0.402 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03366 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.562 ;
        RECT 0.614 0.248 1.114 0.292 ;
        RECT 0.83 0.248 0.898 0.562 ;
        RECT 0.398 0.518 0.682 0.562 ;
        RECT 0.614 0.248 0.682 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.4 0.448 0.464 0.492 ;
        RECT 0.83 0.453 0.898 0.497 ;
        RECT 1.048 0.178 1.112 0.222 ;
        RECT 1.046 0.453 1.114 0.497 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.938 0.453 1.006 0.497 ;
        RECT 1.154 0.538 1.222 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 1.006 0.202 ;
      RECT 0.702 0.068 1.242 0.112 ;
    LAYER v0 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.182 0.158 0.25 0.202 ;
  END
END b15oai112as1n08x5

MACRO b15oai112as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai112as1n12x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.20333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.248 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.918 0.292 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5301235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.594 0.292 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.398 0.248 0.466 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0612 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.134 0.158 1.458 0.202 ;
        RECT 1.262 0.158 1.33 0.562 ;
        RECT 1.046 0.338 1.33 0.382 ;
        RECT 0.398 0.428 1.114 0.472 ;
        RECT 1.046 0.338 1.114 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.262 0.453 1.33 0.497 ;
        RECT 1.37 0.158 1.438 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.154 0.453 1.222 0.497 ;
        RECT 1.37 0.538 1.438 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 1.026 0.202 ;
      RECT 0.81 0.068 1.35 0.112 ;
    LAYER v0 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
  END
END b15oai112as1n12x5

MACRO b15oai112as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai112as1n16x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.338 1.674 0.382 ;
        RECT 1.478 0.248 1.546 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.134 0.338 1.33 0.382 ;
        RECT 1.262 0.158 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.204213 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.87579125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.0985 0.898 0.1425 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.363367 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.27 0.382 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 1.674 0.472 ;
        RECT 1.37 0.158 1.674 0.202 ;
        RECT 1.37 0.158 1.438 0.472 ;
        RECT 0.398 0.518 0.898 0.562 ;
        RECT 0.83 0.428 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
        RECT 1.154 0.538 1.222 0.582 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.538 1.654 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.722 0.0985 0.79 0.1425 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 0.79 0.472 ;
      RECT 0.938 0.068 1.674 0.112 ;
    LAYER v0 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.156 0.178 1.22 0.222 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.94 0.178 1.004 0.222 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.136 0.25 0.18 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.25 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.382 ;
      RECT 0.79 0.338 0.938 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.158 1.222 0.292 ;
  END
END b15oai112as1n16x5

MACRO b15oai122as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai122as1n02x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.383 0.574 0.427 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.383 0.79 0.427 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.383 0.142 0.427 ;
    END
  END e
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0018 LAYER m1 ;
      ANTENNAMAXAREACAR 5.035 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.562 ;
        RECT 0.398 0.158 0.682 0.202 ;
        RECT 0.29 0.338 0.466 0.382 ;
        RECT 0.398 0.158 0.466 0.382 ;
        RECT 0.29 0.338 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.433 0.358 0.477 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.614 0.4905 0.682 0.5345 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.398 0.518 0.466 0.562 ;
        RECT 0.83 0.538 0.898 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.163 0.358 0.207 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.506 0.068 0.574 0.112 ;
    LAYER m1 ;
      RECT 0.486 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.292 ;
  END
END b15oai122as1n02x5

MACRO b15oai122as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai122as1n04x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END e
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0027 LAYER m1 ;
      ANTENNAMAXAREACAR 14.88333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.4675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.594 0.292 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.4555 0.466 0.4995 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.51 0.142 0.554 ;
        RECT 0.614 0.468 0.682 0.512 ;
        RECT 1.046 0.538 1.114 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.29 0.048 0.358 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.81 0.068 1.046 0.112 ;
    LAYER v0 ;
      RECT 1.048 0.138 1.112 0.182 ;
      RECT 0.938 0.24 1.006 0.284 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.074 0.243 0.142 0.287 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.382 ;
      RECT 0.142 0.158 0.938 0.202 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.046 0.068 1.114 0.202 ;
  END
END b15oai122as1n04x5

MACRO b15oai122as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai122as1n08x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.158 1.546 0.472 ;
      LAYER v0 ;
        RECT 1.478 0.2705 1.546 0.3145 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.158 1.33 0.382 ;
        RECT 1.026 0.248 1.33 0.292 ;
      LAYER v0 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.918 0.292 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
        RECT 0.378 0.248 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.27 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
    END
  END e
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04284 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.518 1.438 0.562 ;
        RECT 1.37 0.158 1.438 0.562 ;
        RECT 1.046 0.338 1.114 0.562 ;
        RECT 0.722 0.338 1.114 0.382 ;
        RECT 0.398 0.518 0.79 0.562 ;
        RECT 0.722 0.338 0.79 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.4 0.448 0.464 0.492 ;
        RECT 1.048 0.419 1.112 0.463 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.37 0.178 1.438 0.222 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.83 0.448 0.898 0.492 ;
        RECT 1.478 0.538 1.546 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 1.222 0.202 ;
      RECT 0.702 0.068 1.566 0.112 ;
    LAYER v0 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
  END
END b15oai122as1n08x5

MACRO b15oai122as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai122as1n12x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.248 2.194 0.382 ;
      LAYER v0 ;
        RECT 2.126 0.293 2.194 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.158 1.762 0.382 ;
        RECT 1.37 0.248 1.762 0.292 ;
      LAYER v0 ;
        RECT 1.478 0.248 1.546 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 1.222 0.292 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.248 1.114 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.56130725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.682 0.292 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
        RECT 0.054 0.248 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END e
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06732 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.428 2.214 0.472 ;
        RECT 1.802 0.158 2.214 0.202 ;
        RECT 2.018 0.158 2.086 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 1.262 0.338 1.33 0.472 ;
        RECT 0.83 0.338 1.33 0.382 ;
        RECT 0.506 0.518 0.898 0.562 ;
        RECT 0.83 0.338 0.898 0.562 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.406 0.574 0.45 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.158 2.194 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.802 0.538 1.87 0.582 ;
        RECT 2.018 0.538 2.086 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 1.566 0.202 ;
      RECT 0.918 0.068 2.106 0.112 ;
    LAYER v0 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.586 0.068 1.654 0.112 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.182 0.158 0.25 0.202 ;
  END
END b15oai122as1n12x5

MACRO b15oai122as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai122as1n16x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.0344445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.248 2.734 0.382 ;
      LAYER v0 ;
        RECT 2.666 0.293 2.734 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5875925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.998 0.292 ;
        RECT 1.802 0.248 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.248 1.978 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5875925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.458 0.292 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5875925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.898 0.292 ;
        RECT 0.506 0.248 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5875925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.466 0.292 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END e
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.428 2.754 0.472 ;
        RECT 2.214 0.158 2.754 0.202 ;
        RECT 2.558 0.158 2.626 0.472 ;
        RECT 2.342 0.158 2.41 0.472 ;
        RECT 1.694 0.518 2.194 0.562 ;
        RECT 2.126 0.428 2.194 0.562 ;
        RECT 1.91 0.428 1.978 0.562 ;
        RECT 1.694 0.338 1.762 0.562 ;
        RECT 1.154 0.338 1.762 0.382 ;
        RECT 0.614 0.518 1.222 0.562 ;
        RECT 1.154 0.338 1.222 0.562 ;
        RECT 0.83 0.338 0.898 0.562 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.432 0.682 0.476 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.696 0.448 1.76 0.492 ;
        RECT 1.912 0.448 1.976 0.492 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.158 2.734 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 2.342 0.538 2.41 0.582 ;
        RECT 2.558 0.538 2.626 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 2.106 0.202 ;
      RECT 1.242 0.068 2.646 0.112 ;
    LAYER v0 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.342 0.068 2.41 0.112 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
  END
END b15oai122as1n16x5

MACRO b15oai222as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai222as1n02x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.2935 0.682 0.3375 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.158 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.428 0.79 0.562 ;
        RECT 0.398 0.428 0.79 0.472 ;
        RECT 0.182 0.518 0.466 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.178 0.25 0.222 ;
        RECT 0.29 0.518 0.358 0.562 ;
        RECT 0.724 0.498 0.788 0.542 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.508 0.138 0.572 0.182 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
    LAYER m1 ;
      RECT 0.054 0.068 0.506 0.112 ;
      RECT 0.506 0.068 0.574 0.202 ;
  END
END b15oai222as1n02x5

MACRO b15oai222as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai222as1n04x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.383 0.358 0.427 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.383 0.142 0.427 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 3.6575 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.82875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.318 0.682 0.362 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.383 1.006 0.427 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.428 0.79 0.562 ;
        RECT 0.398 0.428 0.79 0.472 ;
        RECT 0.182 0.518 0.466 0.562 ;
        RECT 0.398 0.428 0.466 0.562 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.178 0.25 0.222 ;
        RECT 0.29 0.518 0.358 0.562 ;
        RECT 0.724 0.498 0.788 0.542 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 0.594 0.112 ;
      RECT 0.29 0.158 1.006 0.202 ;
    LAYER v0 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
  END
END b15oai222as1n04x5

MACRO b15oai222as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai222as1n06x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 1.546 0.472 ;
      LAYER v0 ;
        RECT 1.478 0.293 1.546 0.337 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04284 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.518 1.35 0.562 ;
        RECT 0.938 0.428 1.006 0.562 ;
        RECT 0.722 0.428 1.006 0.472 ;
        RECT 0.29 0.518 0.79 0.562 ;
        RECT 0.722 0.428 0.79 0.562 ;
        RECT 0.162 0.158 0.486 0.202 ;
        RECT 0.29 0.158 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.506 0.518 0.574 0.562 ;
        RECT 1.262 0.518 1.33 0.562 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
      LAYER v0 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 1.586 0.048 1.654 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 1.026 0.112 ;
      RECT 0.594 0.158 1.674 0.202 ;
    LAYER v0 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
  END
END b15oai222as1n06x5

MACRO b15oai222as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai222as1n08x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.248 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.37 0.293 1.438 0.337 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.802 0.293 1.87 0.337 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05202 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.518 1.546 0.562 ;
        RECT 1.478 0.338 1.546 0.562 ;
        RECT 1.154 0.248 1.222 0.562 ;
        RECT 0.83 0.248 1.222 0.292 ;
        RECT 0.398 0.518 0.898 0.562 ;
        RECT 0.83 0.248 0.898 0.562 ;
        RECT 0.054 0.158 0.574 0.202 ;
        RECT 0.398 0.338 0.466 0.562 ;
        RECT 0.29 0.338 0.466 0.382 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.478 0.409 1.546 0.453 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
      LAYER v0 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 1.134 0.112 ;
      RECT 0.702 0.158 1.87 0.202 ;
    LAYER v0 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
  END
END b15oai222as1n08x5

MACRO b15oai222as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai222as1n12x5 0 0 ;
  SIZE 2.592 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.248 1.654 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.293 1.654 0.337 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.248 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.293 1.978 0.337 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.248 2.41 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.293 2.41 0.337 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08262 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.518 2.086 0.562 ;
        RECT 2.018 0.338 2.086 0.562 ;
        RECT 1.694 0.428 1.762 0.562 ;
        RECT 1.478 0.428 1.762 0.472 ;
        RECT 1.478 0.248 1.546 0.472 ;
        RECT 1.154 0.248 1.546 0.292 ;
        RECT 0.506 0.518 1.222 0.562 ;
        RECT 1.154 0.248 1.222 0.562 ;
        RECT 0.938 0.428 1.006 0.562 ;
        RECT 0.722 0.428 0.79 0.562 ;
        RECT 0.162 0.158 0.702 0.202 ;
        RECT 0.506 0.158 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.506 0.415 0.574 0.459 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.724 0.448 0.788 0.492 ;
        RECT 0.94 0.448 1.004 0.492 ;
        RECT 1.154 0.4235 1.222 0.4675 ;
        RECT 1.802 0.518 1.87 0.562 ;
        RECT 2.018 0.411 2.086 0.455 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.626 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.626 0.022 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
      LAYER v0 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 1.566 0.112 ;
      RECT 0.918 0.158 2.518 0.202 ;
    LAYER v0 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
  END
END b15oai222as1n12x5

MACRO b15oai222as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oai222as1n16x5 0 0 ;
  SIZE 3.24 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7775925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5831945 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.9675925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7256945 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.248 2.194 0.472 ;
      LAYER v0 ;
        RECT 2.126 0.293 2.194 0.337 ;
    END
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5875925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.248 2.518 0.472 ;
      LAYER v0 ;
        RECT 2.45 0.293 2.518 0.337 ;
    END
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.248 2.95 0.472 ;
      LAYER v0 ;
        RECT 2.882 0.293 2.95 0.337 ;
    END
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.10404 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.518 2.626 0.562 ;
        RECT 2.558 0.338 2.626 0.562 ;
        RECT 2.342 0.338 2.41 0.562 ;
        RECT 2.018 0.248 2.086 0.562 ;
        RECT 1.478 0.248 2.086 0.292 ;
        RECT 0.614 0.518 1.546 0.562 ;
        RECT 1.478 0.248 1.546 0.562 ;
        RECT 1.262 0.338 1.33 0.562 ;
        RECT 0.162 0.158 0.918 0.202 ;
        RECT 0.83 0.338 0.898 0.562 ;
        RECT 0.614 0.338 0.682 0.562 ;
        RECT 0.506 0.338 0.682 0.382 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
        RECT 0.83 0.4075 0.898 0.4515 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.262 0.4075 1.33 0.4515 ;
        RECT 1.478 0.4095 1.546 0.4535 ;
        RECT 2.342 0.4075 2.41 0.4515 ;
        RECT 2.558 0.397 2.626 0.441 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.274 0.022 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
      LAYER v0 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.068 1.998 0.112 ;
      RECT 1.134 0.158 3.186 0.202 ;
    LAYER v0 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.558 0.158 2.626 0.202 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.074 0.068 0.142 0.112 ;
  END
END b15oai222as1n16x5

MACRO b15oaoi13as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oaoi13as1n02x3 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.428 0.594 0.472 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.1445 0.466 0.1885 ;
        RECT 0.506 0.428 0.574 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.506 0.048 0.574 0.092 ;
    END
  END vssx
END b15oaoi13as1n02x3

MACRO b15oaoi13as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oaoi13as1n02x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.428 0.702 0.472 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.1925 0.574 0.2365 ;
        RECT 0.614 0.428 0.682 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.185 0.25 0.229 ;
        RECT 0.614 0.048 0.682 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.398 0.472 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.518 0.594 0.562 ;
  END
END b15oaoi13as1n02x5

MACRO b15oaoi13as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oaoi13as1n03x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.64666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.378 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.486 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.318 0.142 0.362 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.428 0.918 0.472 ;
        RECT 0.722 0.068 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.128 0.79 0.172 ;
        RECT 0.83 0.428 0.898 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.074 0.158 0.486 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.832 0.048 0.896 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.27 0.068 0.682 0.112 ;
    LAYER v0 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.29 0.068 0.358 0.112 ;
      RECT 0.292 0.498 0.356 0.542 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.614 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.682 0.518 0.81 0.562 ;
  END
END b15oaoi13as1n03x5

MACRO b15oaoi13as1n04x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oaoi13as1n04x3 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.378 0.382 ;
        RECT 0.074 0.338 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.486 0.292 ;
        RECT 0.074 0.068 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.428 0.918 0.472 ;
        RECT 0.722 0.068 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.142 0.79 0.186 ;
        RECT 0.83 0.428 0.898 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.114 0.25 0.158 ;
        RECT 0.398 0.114 0.466 0.158 ;
        RECT 0.832 0.048 0.896 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
    LAYER m1 ;
      RECT 0.27 0.428 0.614 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.682 0.518 0.81 0.562 ;
  END
END b15oaoi13as1n04x3

MACRO b15oaoi13as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oaoi13as1n04x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.825679 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.92239325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.293 1.222 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03366 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.158 0.682 0.202 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.158 0.574 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 1.046 0.538 1.114 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.292 ;
        RECT 1.046 -0.022 1.114 0.292 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.046 0.183 1.114 0.227 ;
        RECT 1.262 0.183 1.33 0.227 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.506 0.518 0.918 0.562 ;
      RECT 0.702 0.428 1.33 0.472 ;
    LAYER v0 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.518 0.682 0.562 ;
  END
END b15oaoi13as1n04x5

MACRO b15oaoi13as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15oaoi13as1n08x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.293 0.682 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.8295425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.382 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.97359475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.068 1.654 0.382 ;
      LAYER v0 ;
        RECT 1.586 0.293 1.654 0.337 ;
    END
  END d
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.158 0.682 0.202 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.158 0.142 0.202 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.158 0.574 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 1.262 0.538 1.33 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.518 0.29 0.562 ;
      RECT 0.614 0.428 1.674 0.472 ;
    LAYER v0 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.138 0.79 0.182 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.411 0.574 0.455 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.29 0.408 0.358 0.452 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.378 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.29 0.248 0.358 0.562 ;
      RECT 0.358 0.248 0.506 0.292 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.574 0.518 1.134 0.562 ;
  END
END b15oaoi13as1n08x5

MACRO b15obai22as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15obai22as1n02x3 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.472 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.068 0.142 0.112 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.3155 0.466 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.562 ;
        RECT 0.506 0.248 0.682 0.292 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.614 0.436 0.682 0.48 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.4505 0.358 0.4945 ;
        RECT 0.83 0.538 0.898 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.203 0.358 0.247 ;
        RECT 0.722 0.118 0.79 0.162 ;
    END
  END vssx
END b15obai22as1n02x3

MACRO b15obai22as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15obai22as1n02x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.594 0.382 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.382 ;
        RECT 0.506 0.248 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 0.898 0.562 ;
        RECT 0.29 0.428 0.898 0.472 ;
        RECT 0.506 0.068 0.574 0.202 ;
        RECT 0.29 0.068 0.574 0.112 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.508 0.138 0.572 0.182 ;
        RECT 0.832 0.498 0.896 0.542 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.722 0.118 0.79 0.162 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
    LAYER v0 ;
      RECT 0.182 0.248 0.25 0.292 ;
      RECT 0.182 0.4555 0.25 0.4995 ;
  END
END b15obai22as1n02x5

MACRO b15obai22as1n04x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15obai22as1n04x3 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.114 0.562 ;
        RECT 0.722 0.338 1.114 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.99777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.202 ;
        RECT 0.054 0.068 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.068 0.142 0.112 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 1.026 0.292 ;
        RECT 0.614 0.248 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.4505 0.682 0.4945 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.468 0.358 0.512 ;
        RECT 0.722 0.4505 0.79 0.4945 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.243 0.358 0.287 ;
        RECT 0.506 0.048 0.574 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.832 0.088 0.896 0.132 ;
      RECT 0.398 0.243 0.466 0.287 ;
      RECT 0.074 0.248 0.142 0.292 ;
      RECT 0.074 0.4505 0.142 0.4945 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.382 ;
      RECT 0.466 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
  END
END b15obai22as1n04x3

MACRO b15obai22as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15obai22as1n04x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.113 1.006 0.157 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.486 0.338 0.79 0.382 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.378 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.428 0.898 0.472 ;
        RECT 0.83 0.068 0.898 0.472 ;
        RECT 0.486 0.068 0.898 0.112 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.83 0.2255 0.898 0.2695 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.046 0.468 1.114 0.512 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.382 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.088 0.142 0.132 ;
        RECT 0.29 0.088 0.358 0.132 ;
        RECT 1.046 0.243 1.114 0.287 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.182 0.088 0.25 0.132 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.25 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
  END
END b15obai22as1n04x5

MACRO b15obai22as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15obai22as1n06x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.64666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.702 0.382 ;
        RECT 0.29 0.338 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.338 1.33 0.562 ;
        RECT 1.134 0.338 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.248 1.438 0.472 ;
        RECT 1.026 0.248 1.438 0.292 ;
      LAYER v0 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.262 0.248 1.33 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.428 1.222 0.562 ;
        RECT 0.486 0.428 1.222 0.472 ;
        RECT 0.83 0.248 0.898 0.472 ;
        RECT 0.398 0.248 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.156 0.498 1.22 0.542 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.722 0.538 0.79 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
        RECT 1.37 0.538 1.438 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.378 0.158 1.458 0.202 ;
    LAYER v0 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.4325 0.142 0.4765 ;
  END
END b15obai22as1n06x5

MACRO b15obai22as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15obai22as1n08x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 0.81 0.382 ;
        RECT 0.29 0.338 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.338 1.438 0.562 ;
        RECT 1.242 0.338 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 1.546 0.472 ;
        RECT 1.134 0.248 1.546 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.428 1.33 0.562 ;
        RECT 0.594 0.428 1.33 0.472 ;
        RECT 0.938 0.248 1.006 0.472 ;
        RECT 0.506 0.248 1.006 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.264 0.498 1.328 0.542 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.486 0.158 1.566 0.202 ;
    LAYER v0 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.4325 0.25 0.4765 ;
  END
END b15obai22as1n08x5

MACRO b15obai22as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15obai22as1n12x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 1.026 0.382 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.782 0.292 ;
        RECT 1.262 0.248 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.586 0.248 1.654 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.248 1.978 0.472 ;
        RECT 1.458 0.338 1.978 0.382 ;
      LAYER v0 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.428 1.762 0.562 ;
        RECT 1.37 0.428 1.762 0.472 ;
        RECT 1.154 0.518 1.438 0.562 ;
        RECT 1.37 0.428 1.438 0.562 ;
        RECT 1.154 0.248 1.222 0.562 ;
        RECT 0.702 0.428 1.222 0.472 ;
        RECT 0.486 0.248 1.222 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.262 0.518 1.33 0.562 ;
        RECT 1.696 0.498 1.76 0.542 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.486 0.158 1.998 0.202 ;
    LAYER v0 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.4325 0.25 0.4765 ;
  END
END b15obai22as1n12x5

MACRO b15obai22as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15obai22as1n16x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.338 1.242 0.382 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.248 2.43 0.292 ;
        RECT 1.478 0.248 1.546 0.472 ;
      LAYER v0 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.234 0.248 2.302 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.338 2.41 0.472 ;
        RECT 1.674 0.338 2.41 0.382 ;
      LAYER v0 ;
        RECT 1.694 0.338 1.762 0.382 ;
        RECT 2.126 0.338 2.194 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.518 2.43 0.562 ;
        RECT 2.234 0.428 2.302 0.562 ;
        RECT 1.586 0.428 2.302 0.472 ;
        RECT 1.37 0.518 1.654 0.562 ;
        RECT 1.586 0.428 1.654 0.562 ;
        RECT 1.37 0.248 1.438 0.562 ;
        RECT 0.506 0.428 1.438 0.472 ;
        RECT 0.486 0.248 1.438 0.292 ;
        RECT 0.506 0.428 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.508 0.498 0.572 0.542 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.478 0.518 1.546 0.562 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 2.342 0.518 2.41 0.562 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
        RECT 2.236 0.048 2.3 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.486 0.158 2.43 0.202 ;
    LAYER v0 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.182 0.4325 0.25 0.4765 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.158 0.378 0.202 ;
  END
END b15obai22as1n16x5

MACRO b15obai22as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15obai22as1n24x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 1.782 0.382 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.694 0.338 1.762 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.248 3.402 0.292 ;
        RECT 2.018 0.248 2.086 0.472 ;
      LAYER v0 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.342 0.248 2.41 0.292 ;
        RECT 2.774 0.248 2.842 0.292 ;
        RECT 3.206 0.248 3.274 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.338 3.382 0.472 ;
        RECT 2.214 0.338 3.382 0.382 ;
      LAYER v0 ;
        RECT 2.234 0.338 2.302 0.382 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END d
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.17136 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.615 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.518 3.402 0.562 ;
        RECT 3.206 0.428 3.274 0.562 ;
        RECT 2.126 0.428 3.274 0.472 ;
        RECT 1.91 0.518 2.194 0.562 ;
        RECT 2.126 0.428 2.194 0.562 ;
        RECT 1.91 0.248 1.978 0.562 ;
        RECT 0.614 0.428 1.978 0.472 ;
        RECT 0.594 0.248 1.978 0.292 ;
        RECT 0.614 0.428 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.616 0.498 0.68 0.542 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.586 0.248 1.654 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.018 0.518 2.086 0.562 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 3.314 0.518 3.382 0.562 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.206 -0.022 3.274 0.112 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
        RECT 3.208 0.048 3.272 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.594 0.158 3.402 0.202 ;
    LAYER v0 ;
      RECT 3.314 0.158 3.382 0.202 ;
      RECT 3.098 0.158 3.166 0.202 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.29 0.4325 0.358 0.4765 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.4325 0.142 0.4765 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.358 0.158 0.486 0.202 ;
  END
END b15obai22as1n24x5

MACRO b15orn002as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn002as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.408 0.466 0.452 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15orn002as1n02x5

MACRO b15orn002as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn002as1n03x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.433 0.466 0.477 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15orn002as1n03x5

MACRO b15orn002as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn002as1n04x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
  END
END b15orn002as1n04x5

MACRO b15orn002as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn002as1n08x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.574 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.83 0.448 0.898 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.3155 0.682 0.3595 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.292 0.498 0.356 0.542 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.614 0.472 ;
      RECT 0.074 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
  END
END b15orn002as1n08x5

MACRO b15orn002as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn002as1n12x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.574 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.562 ;
        RECT 0.722 0.338 1.006 0.382 ;
        RECT 0.722 0.068 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.83 0.448 0.898 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.83 0.138 0.898 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.3155 0.682 0.3595 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.292 0.498 0.356 0.542 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.614 0.472 ;
      RECT 0.074 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
  END
END b15orn002as1n12x5

MACRO b15orn002as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn002as1n16x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.682 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.89818175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.79 0.382 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.562 ;
        RECT 0.938 0.338 1.222 0.382 ;
        RECT 0.938 0.068 1.006 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.448 1.006 0.492 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.154 0.138 1.222 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.182 0.428 0.25 0.562 ;
      RECT 0.25 0.428 0.83 0.472 ;
      RECT 0.074 0.158 0.83 0.202 ;
      RECT 0.83 0.158 0.898 0.472 ;
  END
END b15orn002as1n16x5

MACRO b15orn002as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn002as1n24x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.898 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.918 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0918 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.068 1.654 0.562 ;
        RECT 1.154 0.338 1.654 0.382 ;
        RECT 1.37 0.068 1.438 0.562 ;
        RECT 1.154 0.068 1.222 0.562 ;
      LAYER v0 ;
        RECT 1.154 0.4395 1.222 0.4835 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.37 0.4395 1.438 0.4835 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.4395 1.654 0.4835 ;
        RECT 1.586 0.138 1.654 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.292 0.498 0.356 0.542 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 1.046 0.472 ;
      RECT 0.074 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.472 ;
  END
END b15orn002as1n24x5

MACRO b15orn002as1n32x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn002as1n32x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.548889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.574 0.292 ;
        RECT 0.182 0.248 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.38086175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.565522 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.472 ;
        RECT 0.702 0.248 1.222 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END b
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.11322 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.068 2.086 0.562 ;
        RECT 1.37 0.338 2.086 0.382 ;
        RECT 1.802 0.068 1.87 0.562 ;
        RECT 1.586 0.068 1.654 0.562 ;
        RECT 1.37 0.068 1.438 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.018 0.138 2.086 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
      LAYER v0 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 1.912 0.538 1.976 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 1.91 0.138 1.978 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
    LAYER v0 ;
      RECT 1.262 0.293 1.33 0.337 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.448 1.114 0.492 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.616 0.448 0.68 0.492 ;
      RECT 0.508 0.358 0.572 0.402 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.518 0.25 0.562 ;
      RECT 0.076 0.358 0.14 0.402 ;
    LAYER m1 ;
      RECT 0.162 0.518 0.614 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
      RECT 0.142 0.428 0.506 0.472 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 0.142 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.382 ;
  END
END b15orn002as1n32x5

MACRO b15orn003as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn003as1n02x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.473 0.142 0.517 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.473 0.358 0.517 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.381 0.574 0.425 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.381 0.466 0.425 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END vssx
END b15orn003as1n02x5

MACRO b15orn003as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn003as1n03x5 0 0 ;
  SIZE 0.648 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 1.064 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.436 0.574 0.48 ;
        RECT 0.506 0.138 0.574 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
      LAYER v0 ;
        RECT 0.398 0.538 0.466 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.682 0.022 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.202 ;
      LAYER v0 ;
        RECT 0.182 0.138 0.25 0.182 ;
        RECT 0.398 0.138 0.466 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.4405 0.142 0.4845 ;
  END
END b15orn003as1n03x5

MACRO b15orn003as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn003as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.616 0.158 0.68 0.202 ;
        RECT 0.614 0.4225 0.682 0.4665 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
      LAYER v0 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.518 0.182 0.562 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.382 ;
  END
END b15orn003as1n04x5

MACRO b15orn003as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn003as1n08x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.62277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 1.006 0.382 ;
        RECT 0.938 0.248 1.006 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.562 ;
      LAYER v0 ;
        RECT 1.154 0.4725 1.222 0.5165 ;
        RECT 1.154 0.1755 1.222 0.2195 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
      LAYER v0 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.046 0.4725 1.114 0.5165 ;
        RECT 1.262 0.4725 1.33 0.5165 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.518 0.682 0.562 ;
      RECT 0.29 0.428 1.006 0.472 ;
    LAYER v0 ;
      RECT 1.046 0.293 1.114 0.337 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.182 0.408 0.25 0.452 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.158 0.506 0.202 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.574 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 0.79 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.382 ;
  END
END b15orn003as1n08x5

MACRO b15orn003as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn003as1n12x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.293 0.574 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.562 ;
        RECT 0.614 0.248 1.114 0.292 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.562 ;
        RECT 1.262 0.248 1.546 0.292 ;
        RECT 1.262 0.068 1.33 0.562 ;
      LAYER v0 ;
        RECT 1.262 0.439 1.33 0.483 ;
        RECT 1.262 0.132 1.33 0.176 ;
        RECT 1.478 0.42 1.546 0.464 ;
        RECT 1.478 0.1325 1.546 0.1765 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
      LAYER v0 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.518 0.682 0.562 ;
      RECT 0.29 0.428 1.006 0.472 ;
    LAYER v0 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.184 0.408 0.248 0.452 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.518 0.142 0.562 ;
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.158 1.154 0.202 ;
      RECT 1.154 0.158 1.222 0.382 ;
  END
END b15orn003as1n12x5

MACRO b15orn003as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn003as1n16x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.546 0.382 ;
        RECT 1.478 0.248 1.546 0.382 ;
        RECT 1.154 0.248 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.338 1.33 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
        RECT 0.506 0.338 1.006 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.398 0.248 0.466 0.382 ;
        RECT 0.074 0.248 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.562 ;
        RECT 1.694 0.248 1.978 0.292 ;
        RECT 1.694 0.068 1.762 0.562 ;
      LAYER v0 ;
        RECT 1.694 0.4225 1.762 0.4665 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 1.91 0.4225 1.978 0.4665 ;
        RECT 1.91 0.138 1.978 0.182 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.264 0.048 1.328 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.428 0.898 0.472 ;
      RECT 0.506 0.518 1.438 0.562 ;
    LAYER v0 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.518 1.33 0.562 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.114 0.428 1.458 0.472 ;
      RECT 1.114 0.158 1.586 0.202 ;
      RECT 1.586 0.158 1.654 0.472 ;
  END
END b15orn003as1n16x5

MACRO b15orn003as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15orn003as1n24x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.378 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 1.026 0.292 ;
        RECT 0.614 0.248 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.87 0.562 ;
        RECT 1.35 0.248 1.87 0.292 ;
      LAYER v0 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.586 0.248 1.654 0.292 ;
    END
  END c
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.518 0.562 ;
        RECT 2.018 0.248 2.518 0.292 ;
        RECT 2.234 0.068 2.302 0.562 ;
        RECT 2.018 0.068 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.408 2.086 0.452 ;
        RECT 2.018 0.1495 2.086 0.1935 ;
        RECT 2.234 0.408 2.302 0.452 ;
        RECT 2.234 0.1495 2.302 0.1935 ;
        RECT 2.45 0.408 2.518 0.452 ;
        RECT 2.45 0.1495 2.518 0.1935 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.262 0.518 1.33 0.652 ;
      LAYER v0 ;
        RECT 1.264 0.538 1.328 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
      LAYER v0 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 1.478 0.048 1.546 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.518 1.222 0.562 ;
      RECT 0.614 0.428 1.762 0.472 ;
    LAYER v0 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.518 1.114 0.562 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.518 0.898 0.562 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.518 0.682 0.562 ;
      RECT 0.508 0.408 0.572 0.452 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.518 0.466 0.562 ;
      RECT 0.292 0.408 0.356 0.452 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.518 0.25 0.562 ;
    LAYER m1 ;
      RECT 0.29 0.338 0.358 0.472 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.162 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.574 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.472 ;
  END
END b15orn003as1n24x5

MACRO b15ornc04as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ornc04as1n02x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.378 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.518 1.026 0.562 ;
        RECT 0.83 0.338 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.518 1.006 0.562 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0018 LAYER m1 ;
      ANTENNAMAXAREACAR 4.56 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.248 0.682 0.562 ;
        RECT 0.398 0.338 0.682 0.382 ;
        RECT 0.398 0.158 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.203 0.466 0.247 ;
        RECT 0.614 0.42 0.682 0.464 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.4555 0.142 0.4995 ;
        RECT 0.506 0.51 0.574 0.554 ;
        RECT 0.722 0.538 0.79 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.166 0.25 0.21 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.938 0.378 1.006 0.422 ;
      RECT 0.83 0.138 0.898 0.182 ;
    LAYER m1 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 0.898 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.472 ;
  END
END b15ornc04as1n02x5

MACRO b15ornc04as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ornc04as1n03x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.054 0.518 0.25 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.518 0.142 0.562 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0153 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.006 0.382 ;
        RECT 0.938 0.158 1.006 0.382 ;
        RECT 0.83 0.338 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.468 0.898 0.512 ;
        RECT 0.938 0.2305 1.006 0.2745 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.468 0.358 0.512 ;
        RECT 0.722 0.468 0.79 0.512 ;
        RECT 0.938 0.468 1.006 0.512 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.178 0.25 0.222 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
    LAYER v0 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.506 0.448 0.574 0.492 ;
      RECT 0.074 0.178 0.142 0.222 ;
      RECT 0.074 0.343 0.142 0.387 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.574 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
  END
END b15ornc04as1n03x5

MACRO b15ornc04as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ornc04as1n04x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 1.2385185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.518 0.466 0.562 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.518 0.358 0.562 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.006 0.382 ;
        RECT 0.938 0.158 1.006 0.382 ;
        RECT 0.83 0.338 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.468 0.898 0.512 ;
        RECT 0.938 0.24 1.006 0.284 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.468 0.142 0.512 ;
        RECT 0.722 0.468 0.79 0.512 ;
        RECT 0.938 0.468 1.006 0.512 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.198 0.25 0.242 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
    END
  END vssx
  OBS
    LAYER v0 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.506 0.4455 0.574 0.4895 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.574 0.562 ;
      RECT 0.574 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.292 ;
  END
END b15ornc04as1n04x5

MACRO b15ornc04as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ornc04as1n06x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.248 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.293 0.79 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.248 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.293 1.006 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0063 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41015875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.57422225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.3155 0.358 0.3595 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02142 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.574 0.382 ;
        RECT 0.506 0.068 0.574 0.382 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.423 0.466 0.467 ;
        RECT 0.506 0.167 0.574 0.211 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.506 0.523 0.574 0.567 ;
        RECT 0.938 0.538 1.006 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.1285 0.358 0.1725 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.248 0.682 0.562 ;
    LAYER v0 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.293 0.682 0.337 ;
      RECT 0.182 0.2125 0.25 0.2565 ;
      RECT 0.076 0.498 0.14 0.542 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.142 0.428 0.182 0.472 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.068 0.898 0.562 ;
  END
END b15ornc04as1n06x5

MACRO b15ornc04as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ornc04as1n08x5 0 0 ;
  SIZE 1.512 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.158 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.0306 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 0.898 0.562 ;
        RECT 0.614 0.338 0.898 0.382 ;
        RECT 0.614 0.158 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.428 0.898 0.472 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.546 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.938 0.338 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.518 0.142 0.562 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.722 0.518 0.79 0.562 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.37 0.518 1.438 0.562 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.546 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.83 0.158 0.898 0.202 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.046 0.158 1.114 0.562 ;
    LAYER v0 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.398 0.338 0.466 0.382 ;
      RECT 0.29 0.518 0.358 0.562 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.518 0.398 0.562 ;
      RECT 0.398 0.248 0.466 0.562 ;
      RECT 1.114 0.518 1.262 0.562 ;
      RECT 1.262 0.068 1.33 0.562 ;
  END
END b15ornc04as1n08x5

MACRO b15ornc04as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ornc04as1n12x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.158 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.248 1.87 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.562 ;
        RECT 0.722 0.248 1.222 0.292 ;
        RECT 0.938 0.248 1.006 0.562 ;
        RECT 0.722 0.248 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.498 0.79 0.542 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 0.938 0.498 1.006 0.542 ;
        RECT 1.154 0.498 1.222 0.542 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.4705 0.25 0.5145 ;
        RECT 0.83 0.498 0.898 0.542 ;
        RECT 1.046 0.498 1.114 0.542 ;
        RECT 1.694 0.4695 1.762 0.5135 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.158 0.358 0.202 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 1.802 0.048 1.87 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 0.614 0.158 1.33 0.202 ;
    LAYER v0 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.382 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.248 0.682 0.562 ;
      RECT 1.33 0.518 1.478 0.562 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 1.546 0.338 1.694 0.382 ;
      RECT 1.694 0.068 1.762 0.382 ;
  END
END b15ornc04as1n12x5

MACRO b15ornc04as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ornc04as1n16x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.466 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.574 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.338 1.978 0.562 ;
        RECT 1.694 0.338 1.978 0.382 ;
      LAYER v0 ;
        RECT 1.802 0.338 1.87 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.248 2.086 0.472 ;
        RECT 1.586 0.248 2.086 0.292 ;
      LAYER v0 ;
        RECT 1.694 0.248 1.762 0.292 ;
        RECT 1.91 0.248 1.978 0.292 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07038 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.428 1.438 0.472 ;
        RECT 1.154 0.248 1.222 0.472 ;
        RECT 0.722 0.248 1.222 0.292 ;
        RECT 0.722 0.068 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.724 0.178 0.788 0.222 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.262 0.428 1.33 0.472 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 1.262 0.338 1.478 0.382 ;
    LAYER v0 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.804 0.498 1.868 0.542 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.37 0.338 1.438 0.382 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.832 0.088 0.896 0.132 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.292 0.498 0.356 0.542 ;
      RECT 0.182 0.158 0.25 0.202 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.358 0.562 ;
      RECT 0.358 0.428 0.614 0.472 ;
      RECT 0.074 0.158 0.614 0.202 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 1.114 0.382 ;
      RECT 0.898 0.158 1.438 0.202 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.546 0.428 1.802 0.472 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 1.546 0.158 2.086 0.202 ;
  END
END b15ornc04as1n16x5

MACRO b15ornc04as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ornc04as1n24x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.486 0.338 0.682 0.382 ;
        RECT 0.614 0.158 0.682 0.382 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7053595 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.338 0.378 0.382 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.3975925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.596389 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.338 2.41 0.382 ;
        RECT 2.342 0.248 2.41 0.382 ;
        RECT 2.126 0.248 2.194 0.382 ;
      LAYER v0 ;
        RECT 2.234 0.338 2.302 0.382 ;
    END
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.7494445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.338 2.734 0.382 ;
        RECT 2.666 0.158 2.734 0.382 ;
        RECT 2.45 0.248 2.518 0.382 ;
      LAYER v0 ;
        RECT 2.558 0.338 2.626 0.382 ;
    END
  END d
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.428 1.87 0.472 ;
        RECT 1.37 0.248 1.438 0.472 ;
        RECT 0.938 0.248 1.438 0.292 ;
      LAYER v0 ;
        RECT 1.046 0.428 1.114 0.472 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.262 0.428 1.33 0.472 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.694 0.428 1.762 0.472 ;
    END
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.506 -0.022 0.574 0.292 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.178 0.142 0.222 ;
        RECT 0.29 0.178 0.358 0.222 ;
        RECT 0.506 0.178 0.574 0.222 ;
        RECT 0.722 0.178 0.79 0.222 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.428 0.79 0.472 ;
      RECT 0.83 0.068 1.262 0.112 ;
      RECT 1.478 0.338 1.91 0.382 ;
      RECT 2.018 0.428 2.734 0.472 ;
    LAYER v0 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.518 2.302 0.562 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.338 1.87 0.382 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.938 0.338 1.006 0.382 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.518 0.574 0.562 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.398 0.518 0.83 0.562 ;
      RECT 0.83 0.158 0.898 0.562 ;
      RECT 0.898 0.338 1.33 0.382 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.158 1.978 0.202 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.978 0.338 2.018 0.382 ;
      RECT 2.018 0.158 2.086 0.382 ;
      RECT 1.978 0.518 2.322 0.562 ;
      RECT 2.086 0.158 2.626 0.202 ;
  END
END b15ornc04as1n24x5

MACRO b15rm0023as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rm0023as1n02x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 3.7255555 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 3.7255555 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.458 0.068 1.782 0.112 ;
        RECT 0.486 0.068 0.682 0.112 ;
      LAYER m2 ;
        RECT 0.488 0.068 1.564 0.112 ;
      LAYER v1 ;
        RECT 0.51 0.068 0.57 0.112 ;
        RECT 1.482 0.068 1.542 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 1.478 0.068 1.546 0.112 ;
        RECT 1.694 0.068 1.762 0.112 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 1.978 0.292 ;
        RECT 1.91 0.068 1.978 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.338 2.086 0.382 ;
        RECT 2.018 0.158 2.086 0.382 ;
        RECT 1.37 0.518 1.978 0.562 ;
        RECT 1.91 0.338 1.978 0.562 ;
        RECT 1.37 0.338 1.438 0.562 ;
        RECT 0.182 0.338 1.438 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 2.018 0.248 2.086 0.292 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.156 0.142 0.2 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.126 0.138 2.194 0.182 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.473 0.79 0.517 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 2.018 0.048 2.086 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.428 1.564 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.682 0.472 ;
      RECT 0.486 0.068 0.682 0.112 ;
      RECT 0.594 0.158 0.918 0.202 ;
      RECT 1.046 0.158 1.654 0.202 ;
      RECT 1.458 0.068 1.782 0.112 ;
    LAYER v1 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 0.51 0.428 0.57 0.472 ;
    LAYER v0 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 1.478 0.338 1.546 0.472 ;
      RECT 1.546 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.472 ;
  END
END b15rm0023as1n02x5

MACRO b15rm0023as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rm0023as1n04x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 3.7255555 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 3.7255555 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.458 0.068 1.782 0.112 ;
        RECT 0.486 0.068 0.682 0.112 ;
      LAYER m2 ;
        RECT 0.488 0.068 1.564 0.112 ;
      LAYER v1 ;
        RECT 0.51 0.068 0.57 0.112 ;
        RECT 1.482 0.068 1.542 0.112 ;
      LAYER v0 ;
        RECT 0.506 0.068 0.574 0.112 ;
        RECT 1.478 0.068 1.546 0.112 ;
        RECT 1.694 0.068 1.762 0.112 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 1.978 0.292 ;
        RECT 1.91 0.068 1.978 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.338 2.086 0.382 ;
        RECT 2.018 0.158 2.086 0.382 ;
        RECT 1.37 0.518 1.978 0.562 ;
        RECT 1.91 0.338 1.978 0.562 ;
        RECT 1.37 0.338 1.438 0.562 ;
        RECT 0.182 0.338 1.438 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 2.018 0.248 2.086 0.292 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.156 0.142 0.2 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.068 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.126 0.138 2.194 0.182 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.722 0.473 0.79 0.517 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.262 -0.022 1.33 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.046 0.048 1.114 0.092 ;
        RECT 1.262 0.048 1.33 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.428 1.564 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.682 0.472 ;
      RECT 0.486 0.068 0.682 0.112 ;
      RECT 0.594 0.158 0.918 0.202 ;
      RECT 1.046 0.158 1.654 0.202 ;
      RECT 1.458 0.068 1.782 0.112 ;
    LAYER v1 ;
      RECT 1.482 0.428 1.542 0.472 ;
      RECT 0.51 0.428 0.57 0.472 ;
    LAYER v0 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
    LAYER m1 ;
      RECT 1.478 0.338 1.546 0.472 ;
      RECT 1.546 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.472 ;
  END
END b15rm0023as1n04x5

MACRO b15rm0023as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rm0023as1n06x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 3.7255555 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 3.7255555 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.566 0.068 1.89 0.112 ;
        RECT 0.594 0.068 0.79 0.112 ;
      LAYER m2 ;
        RECT 0.596 0.068 1.672 0.112 ;
      LAYER v1 ;
        RECT 0.618 0.068 0.678 0.112 ;
        RECT 1.59 0.068 1.65 0.112 ;
      LAYER v0 ;
        RECT 0.614 0.068 0.682 0.112 ;
        RECT 1.586 0.068 1.654 0.112 ;
        RECT 1.802 0.068 1.87 0.112 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 2.086 0.292 ;
        RECT 2.018 0.068 2.086 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.91 0.248 1.978 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.338 2.194 0.382 ;
        RECT 2.126 0.158 2.194 0.382 ;
        RECT 1.478 0.518 1.978 0.562 ;
        RECT 1.91 0.338 1.978 0.562 ;
        RECT 1.478 0.338 1.546 0.562 ;
        RECT 0.29 0.338 1.546 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 2.126 0.248 2.194 0.292 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.156 0.25 0.2 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.068 2.302 0.562 ;
      LAYER v0 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.234 0.138 2.302 0.182 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.83 0.473 0.898 0.517 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.37 0.448 1.438 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.342 0.448 2.41 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.83 0.048 0.898 0.092 ;
        RECT 1.154 0.048 1.222 0.092 ;
        RECT 1.37 0.048 1.438 0.092 ;
        RECT 2.126 0.048 2.194 0.092 ;
        RECT 2.342 0.048 2.41 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.596 0.428 1.672 0.472 ;
    LAYER m1 ;
      RECT 0.398 0.428 0.79 0.472 ;
      RECT 0.594 0.068 0.79 0.112 ;
      RECT 0.702 0.158 1.026 0.202 ;
      RECT 1.154 0.158 1.762 0.202 ;
      RECT 1.566 0.068 1.89 0.112 ;
    LAYER v1 ;
      RECT 1.59 0.428 1.65 0.472 ;
      RECT 0.618 0.428 0.678 0.472 ;
    LAYER v0 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
    LAYER m1 ;
      RECT 1.586 0.338 1.654 0.472 ;
      RECT 1.654 0.338 1.782 0.382 ;
  END
END b15rm0023as1n06x5

MACRO b15rm0023as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rm0023as1n08x5 0 0 ;
  SIZE 3.132 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0216 LAYER m2 ;
      ANTENNAMAXAREACAR 5.15402775 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0216 LAYER m2 ;
      ANTENNAMAXAREACAR 5.15402775 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.158 2.41 0.202 ;
        RECT 2.126 0.068 2.194 0.202 ;
        RECT 1.694 0.068 2.194 0.112 ;
        RECT 0.81 0.068 1.006 0.112 ;
      LAYER m2 ;
        RECT 0.812 0.068 2.104 0.112 ;
      LAYER v1 ;
        RECT 0.834 0.068 0.894 0.112 ;
        RECT 1.806 0.068 1.866 0.112 ;
        RECT 2.022 0.068 2.082 0.112 ;
      LAYER v0 ;
        RECT 0.83 0.068 0.898 0.112 ;
        RECT 1.802 0.068 1.87 0.112 ;
        RECT 2.234 0.158 2.302 0.202 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.248 2.734 0.292 ;
        RECT 2.45 0.158 2.518 0.292 ;
        RECT 0.398 0.248 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.248 0.574 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 2.558 0.248 2.626 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 2.734 0.382 ;
        RECT 2.45 0.338 2.518 0.472 ;
        RECT 0.722 0.338 0.79 0.562 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.478 0.338 1.546 0.382 ;
        RECT 2.558 0.338 2.626 0.382 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.068 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.115 0.25 0.159 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.068 2.95 0.562 ;
      LAYER v0 ;
        RECT 2.882 0.473 2.95 0.517 ;
        RECT 2.882 0.1425 2.95 0.1865 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.166 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.588 0.538 1.652 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.99 0.473 3.058 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.166 0.022 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.774 -0.022 2.842 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.115 0.142 0.159 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 2.776 0.048 2.84 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.428 2.212 0.472 ;
    LAYER m1 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 1.694 0.068 2.126 0.112 ;
      RECT 0.81 0.068 1.006 0.112 ;
      RECT 0.83 0.428 1.33 0.472 ;
      RECT 0.614 0.158 1.33 0.202 ;
      RECT 1.37 0.428 1.998 0.472 ;
      RECT 1.37 0.158 2.086 0.202 ;
      RECT 2.106 0.428 2.322 0.472 ;
      RECT 1.998 0.518 2.558 0.562 ;
    LAYER v1 ;
      RECT 2.13 0.428 2.19 0.472 ;
      RECT 0.618 0.428 0.678 0.472 ;
      RECT 0.294 0.428 0.354 0.472 ;
    LAYER v0 ;
      RECT 2.774 0.248 2.842 0.292 ;
      RECT 2.342 0.068 2.41 0.112 ;
      RECT 2.342 0.518 2.41 0.562 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.614 0.495 0.682 0.539 ;
      RECT 0.29 0.248 0.358 0.292 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.358 0.158 0.506 0.202 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.574 0.068 0.702 0.112 ;
      RECT 2.126 0.068 2.194 0.202 ;
      RECT 2.194 0.158 2.41 0.202 ;
      RECT 2.234 0.068 2.558 0.112 ;
      RECT 2.558 0.428 2.626 0.562 ;
      RECT 2.558 0.068 2.626 0.202 ;
      RECT 2.626 0.428 2.774 0.472 ;
      RECT 2.626 0.158 2.774 0.202 ;
      RECT 2.774 0.158 2.842 0.472 ;
  END
END b15rm0023as1n08x5

MACRO b15rm6013es1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rm6013es1n02x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 0.466 0.562 ;
        RECT 0.27 0.338 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.574 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
    END
  END c
  PIN carryb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 2.28 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END carryb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.472 0.358 0.516 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
    END
  END vssx
END b15rm6013es1n02x5

MACRO b15rm6013es1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rm6013es1n04x5 0 0 ;
  SIZE 0.864 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.574 0.472 ;
        RECT 0.27 0.338 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.574 0.292 ;
        RECT 0.506 0.158 0.574 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.248 0.466 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.158 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.2705 0.79 0.3145 ;
    END
  END c
  PIN carryb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.565 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.614 0.408 0.682 0.452 ;
        RECT 0.614 0.178 0.682 0.222 ;
    END
  END carryb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.898 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.898 0.022 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.398 0.202 ;
    LAYER v0 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.398 0.472 ;
      RECT 0.398 0.428 0.466 0.562 ;
      RECT 0.466 0.518 0.81 0.562 ;
      RECT 0.398 0.068 0.466 0.202 ;
      RECT 0.466 0.068 0.81 0.112 ;
  END
END b15rm6013es1n04x5

MACRO b15rm6013es1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rm6013es1n08x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.27 0.338 1.654 0.382 ;
        RECT 1.586 0.248 1.654 0.382 ;
        RECT 0.722 0.338 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.478 0.338 1.546 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 1.458 0.292 ;
        RECT 0.722 0.158 0.79 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.248 1.978 0.382 ;
      LAYER v0 ;
        RECT 1.91 0.293 1.978 0.337 ;
    END
  END c
  PIN carryb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.472 ;
        RECT 0.918 0.158 2.086 0.202 ;
      LAYER v0 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.91 0.428 1.978 0.472 ;
        RECT 1.91 0.158 1.978 0.202 ;
    END
  END carryb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.614 0.202 ;
    LAYER v0 ;
      RECT 2.018 0.068 2.086 0.112 ;
      RECT 2.018 0.518 2.086 0.562 ;
      RECT 1.802 0.068 1.87 0.112 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.614 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.682 0.518 2.106 0.562 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 0.682 0.068 2.106 0.112 ;
  END
END b15rm6013es1n08x5

MACRO b15rm6013es1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rm6013es1n12x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.27 0.338 2.302 0.382 ;
        RECT 2.234 0.248 2.302 0.382 ;
        RECT 0.938 0.338 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
        RECT 2.126 0.338 2.194 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 2.106 0.292 ;
        RECT 0.938 0.158 1.006 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.248 0.466 0.292 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.586 0.248 1.654 0.292 ;
        RECT 2.018 0.248 2.086 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.248 2.626 0.382 ;
      LAYER v0 ;
        RECT 2.558 0.293 2.626 0.337 ;
    END
  END c
  PIN carryb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.134 0.428 2.842 0.472 ;
        RECT 2.774 0.158 2.842 0.472 ;
        RECT 1.134 0.158 2.842 0.202 ;
      LAYER v0 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.586 0.428 1.654 0.472 ;
        RECT 1.586 0.158 1.654 0.202 ;
        RECT 2.018 0.428 2.086 0.472 ;
        RECT 2.018 0.158 2.086 0.202 ;
        RECT 2.45 0.428 2.518 0.472 ;
        RECT 2.45 0.158 2.518 0.202 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.158 2.734 0.202 ;
    END
  END carryb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.83 0.202 ;
    LAYER v0 ;
      RECT 2.774 0.068 2.842 0.112 ;
      RECT 2.774 0.518 2.842 0.562 ;
      RECT 2.558 0.068 2.626 0.112 ;
      RECT 2.558 0.518 2.626 0.562 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.83 0.472 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.898 0.518 2.862 0.562 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 2.862 0.112 ;
  END
END b15rm6013es1n12x5

MACRO b15rm6013es1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rm6013es1n16x5 0 0 ;
  SIZE 3.672 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.27 0.338 2.95 0.382 ;
        RECT 2.882 0.248 2.95 0.382 ;
        RECT 1.154 0.338 1.222 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 1.262 0.338 1.33 0.382 ;
        RECT 1.586 0.338 1.654 0.382 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.45 0.338 2.518 0.382 ;
        RECT 2.774 0.338 2.842 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 2.754 0.292 ;
        RECT 1.154 0.158 1.222 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.234 0.248 2.302 0.292 ;
        RECT 2.666 0.248 2.734 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.248 3.49 0.292 ;
        RECT 3.206 0.248 3.274 0.382 ;
      LAYER v0 ;
        RECT 3.314 0.248 3.382 0.292 ;
    END
  END c
  PIN carryb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.35 0.428 3.598 0.472 ;
        RECT 3.53 0.158 3.598 0.472 ;
        RECT 1.35 0.158 3.598 0.202 ;
      LAYER v0 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.206 0.158 3.274 0.202 ;
        RECT 3.422 0.428 3.49 0.472 ;
        RECT 3.422 0.158 3.49 0.202 ;
    END
  END carryb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.706 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.706 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 1.046 0.202 ;
    LAYER v0 ;
      RECT 3.53 0.068 3.598 0.112 ;
      RECT 3.53 0.518 3.598 0.562 ;
      RECT 3.314 0.068 3.382 0.112 ;
      RECT 3.314 0.518 3.382 0.562 ;
      RECT 3.098 0.068 3.166 0.112 ;
      RECT 3.098 0.518 3.166 0.562 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.428 1.046 0.472 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.114 0.518 3.618 0.562 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.114 0.068 3.618 0.112 ;
  END
END b15rm6013es1n16x5

MACRO b15rm6013es1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rm6013es1n24x5 0 0 ;
  SIZE 5.184 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.27 0.338 4.246 0.382 ;
        RECT 4.178 0.248 4.246 0.382 ;
        RECT 1.586 0.338 1.654 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.694 0.338 1.762 0.382 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.45 0.338 2.518 0.382 ;
        RECT 2.882 0.338 2.95 0.382 ;
        RECT 3.314 0.338 3.382 0.382 ;
        RECT 3.746 0.338 3.814 0.382 ;
        RECT 4.07 0.338 4.138 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0864 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 4.05 0.292 ;
        RECT 1.586 0.158 1.654 0.292 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.248 0.898 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
        RECT 2.234 0.248 2.302 0.292 ;
        RECT 2.666 0.248 2.734 0.292 ;
        RECT 3.098 0.248 3.166 0.292 ;
        RECT 3.53 0.248 3.598 0.292 ;
        RECT 3.962 0.248 4.03 0.292 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.502 0.248 4.914 0.292 ;
        RECT 4.502 0.248 4.57 0.382 ;
      LAYER v0 ;
        RECT 4.61 0.248 4.678 0.292 ;
        RECT 4.826 0.248 4.894 0.292 ;
    END
  END c
  PIN carryb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14688 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.782 0.428 5.11 0.472 ;
        RECT 5.042 0.158 5.11 0.472 ;
        RECT 1.782 0.158 5.11 0.202 ;
      LAYER v0 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.666 0.158 2.734 0.202 ;
        RECT 3.098 0.428 3.166 0.472 ;
        RECT 3.098 0.158 3.166 0.202 ;
        RECT 3.53 0.428 3.598 0.472 ;
        RECT 3.53 0.158 3.598 0.202 ;
        RECT 3.962 0.428 4.03 0.472 ;
        RECT 3.962 0.158 4.03 0.202 ;
        RECT 4.502 0.428 4.57 0.472 ;
        RECT 4.502 0.158 4.57 0.202 ;
        RECT 4.718 0.428 4.786 0.472 ;
        RECT 4.718 0.158 4.786 0.202 ;
        RECT 4.934 0.428 5.002 0.472 ;
        RECT 4.934 0.158 5.002 0.202 ;
    END
  END carryb
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.218 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.218 0.022 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 1.478 0.202 ;
    LAYER v0 ;
      RECT 5.042 0.068 5.11 0.112 ;
      RECT 5.042 0.518 5.11 0.562 ;
      RECT 4.826 0.068 4.894 0.112 ;
      RECT 4.826 0.518 4.894 0.562 ;
      RECT 4.61 0.068 4.678 0.112 ;
      RECT 4.61 0.518 4.678 0.562 ;
      RECT 4.394 0.068 4.462 0.112 ;
      RECT 4.394 0.518 4.462 0.562 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.428 1.478 0.472 ;
      RECT 1.478 0.428 1.546 0.562 ;
      RECT 1.546 0.518 5.13 0.562 ;
      RECT 1.478 0.068 1.546 0.202 ;
      RECT 1.546 0.068 5.13 0.112 ;
  END
END b15rm6013es1n24x5

MACRO b15rt0022es1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rt0022es1n02x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 1.114 0.382 ;
        RECT 0.398 0.338 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.506 0.338 0.574 0.382 ;
        RECT 0.938 0.338 1.006 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.594 0.248 1.114 0.292 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.562 ;
      LAYER v0 ;
        RECT 1.154 0.448 1.222 0.492 ;
        RECT 1.154 0.138 1.222 0.182 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.158 0.142 0.202 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.506 0.428 0.918 0.472 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.428 0.898 0.472 ;
        RECT 1.046 0.448 1.114 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 1.046 0.138 1.114 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.378 0.068 0.702 0.112 ;
    LAYER v0 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.29 0.448 0.358 0.492 ;
      RECT 0.182 0.248 0.25 0.292 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.382 ;
      RECT 0.25 0.338 0.29 0.382 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.25 0.158 0.594 0.202 ;
  END
END b15rt0022es1n02x5

MACRO b15rt0022es1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rt0022es1n04x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 0.918 0.382 ;
        RECT 0.378 0.518 0.574 0.562 ;
        RECT 0.506 0.338 0.574 0.562 ;
      LAYER v0 ;
        RECT 0.398 0.518 0.466 0.562 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.248 1.114 0.382 ;
        RECT 0.594 0.248 1.114 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.068 1.33 0.562 ;
      LAYER v0 ;
        RECT 1.262 0.473 1.33 0.517 ;
        RECT 1.262 0.1125 1.33 0.1565 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.068 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.408 0.142 0.452 ;
        RECT 0.074 0.132 0.142 0.176 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.83 0.538 0.898 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.068 0.358 0.382 ;
    LAYER v0 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.4 0.358 0.464 0.402 ;
      RECT 0.29 0.248 0.358 0.292 ;
      RECT 0.182 0.248 0.25 0.292 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.428 0.398 0.472 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.158 0.594 0.202 ;
      RECT 0.358 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 0.83 0.428 1.154 0.472 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.158 1.222 0.472 ;
  END
END b15rt0022es1n04x5

MACRO b15rt0022es1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rt0022es1n08x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0207 LAYER m1 ;
      ANTENNAMAXAREACAR 0.89818175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.338 1.674 0.382 ;
        RECT 0.398 0.248 0.466 0.382 ;
      LAYER v0 ;
        RECT 0.722 0.338 0.79 0.382 ;
        RECT 1.586 0.338 1.654 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.248 1.87 0.382 ;
        RECT 0.594 0.248 1.87 0.292 ;
        RECT 1.478 0.068 1.546 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.248 0.682 0.292 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.37 0.248 1.438 0.292 ;
        RECT 1.694 0.248 1.762 0.292 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.451 2.086 0.495 ;
        RECT 2.018 0.178 2.086 0.222 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.562 ;
      LAYER v0 ;
        RECT 0.182 0.451 0.25 0.495 ;
        RECT 0.182 0.178 0.25 0.222 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.586 0.518 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 0.938 0.538 1.006 0.582 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.538 1.654 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.026 0.158 1.438 0.202 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.046 0.158 1.114 0.202 ;
        RECT 1.37 0.088 1.438 0.132 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.586 0.068 1.654 0.202 ;
      RECT 0.486 0.068 1.242 0.112 ;
    LAYER v0 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.588 0.088 1.652 0.132 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.506 0.068 0.574 0.112 ;
      RECT 0.29 0.338 0.358 0.382 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.358 0.158 0.918 0.202 ;
      RECT 0.358 0.428 1.134 0.472 ;
      RECT 1.242 0.428 1.91 0.472 ;
      RECT 1.654 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.472 ;
  END
END b15rt0022es1n08x5

MACRO b15rt0022es1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rt0022es1n12x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0252 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.338 1.782 0.382 ;
        RECT 0.506 0.248 0.574 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.694 0.338 1.762 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0252 LAYER m1 ;
      ANTENNAMAXAREACAR 0.88666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.248 1.978 0.382 ;
        RECT 0.702 0.248 1.978 0.292 ;
        RECT 1.586 0.068 1.654 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.248 0.79 0.292 ;
        RECT 1.046 0.248 1.114 0.292 ;
        RECT 1.478 0.248 1.546 0.292 ;
        RECT 1.802 0.248 1.87 0.292 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.068 2.41 0.562 ;
        RECT 2.126 0.248 2.41 0.292 ;
        RECT 2.126 0.068 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.342 0.448 2.41 0.492 ;
        RECT 2.342 0.138 2.41 0.182 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.158 0.358 0.562 ;
        RECT 0.074 0.338 0.358 0.382 ;
        RECT 0.074 0.158 0.142 0.562 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.074 0.178 0.142 0.222 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.29 0.178 0.358 0.222 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 1.478 0.538 1.546 0.582 ;
        RECT 1.694 0.538 1.762 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
        RECT 2.234 0.448 2.302 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.134 0.158 1.546 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.154 0.158 1.222 0.202 ;
        RECT 1.478 0.088 1.546 0.132 ;
        RECT 1.912 0.048 1.976 0.092 ;
        RECT 2.234 0.138 2.302 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 1.694 0.068 1.762 0.202 ;
      RECT 0.594 0.068 1.35 0.112 ;
    LAYER v0 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.696 0.088 1.76 0.132 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.398 0.338 0.466 0.382 ;
    LAYER m1 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.466 0.158 1.026 0.202 ;
      RECT 0.466 0.428 1.242 0.472 ;
      RECT 1.35 0.428 2.018 0.472 ;
      RECT 1.762 0.158 2.018 0.202 ;
      RECT 2.018 0.158 2.086 0.472 ;
  END
END b15rt0022es1n12x5

MACRO b15rt0022es1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rt0022es1n16x5 0 0 ;
  SIZE 3.24 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.918 0.248 2.43 0.292 ;
        RECT 1.802 0.068 1.87 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.248 1.006 0.292 ;
        RECT 1.262 0.248 1.33 0.292 ;
        RECT 2.018 0.248 2.086 0.292 ;
        RECT 2.342 0.248 2.41 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 2.626 0.382 ;
        RECT 1.802 0.338 1.87 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.338 0.898 0.382 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 2.126 0.338 2.194 0.382 ;
        RECT 2.45 0.338 2.518 0.382 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.338 3.166 0.382 ;
        RECT 3.098 0.158 3.166 0.382 ;
        RECT 2.666 0.158 3.166 0.202 ;
        RECT 2.99 0.338 3.058 0.562 ;
        RECT 2.774 0.338 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.774 0.158 2.842 0.202 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 2.99 0.158 3.058 0.202 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.574 0.202 ;
        RECT 0.398 0.338 0.466 0.562 ;
        RECT 0.074 0.338 0.466 0.382 ;
        RECT 0.182 0.338 0.25 0.562 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.448 0.466 0.492 ;
        RECT 0.398 0.158 0.466 0.202 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.274 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 2.45 0.518 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.478 0.518 1.546 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.48 0.538 1.544 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
        RECT 2.236 0.538 2.3 0.582 ;
        RECT 2.452 0.538 2.516 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.274 0.022 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 1.48 0.048 1.544 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.292 ;
      RECT 1.91 0.068 1.978 0.202 ;
    LAYER v0 ;
      RECT 2.882 0.248 2.95 0.292 ;
      RECT 2.342 0.158 2.41 0.202 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 1.912 0.088 1.976 0.132 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.724 0.228 0.788 0.272 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.29 0.248 0.358 0.292 ;
    LAYER m1 ;
      RECT 0.27 0.248 0.614 0.292 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 0.682 0.068 1.35 0.112 ;
      RECT 0.682 0.428 1.674 0.472 ;
      RECT 0.79 0.158 1.762 0.202 ;
      RECT 1.978 0.158 2.558 0.202 ;
      RECT 2.558 0.158 2.626 0.292 ;
      RECT 2.018 0.428 2.666 0.472 ;
      RECT 2.626 0.248 2.666 0.292 ;
      RECT 2.666 0.248 2.734 0.472 ;
      RECT 2.734 0.248 2.97 0.292 ;
  END
END b15rt0022es1n16x5

MACRO b15rt0022es1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15rt0022es1n24x5 0 0 ;
  SIZE 4.32 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0549 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0621 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.134 0.248 3.294 0.292 ;
        RECT 2.666 0.068 2.734 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.248 1.222 0.292 ;
        RECT 1.586 0.248 1.654 0.292 ;
        RECT 1.91 0.248 1.978 0.292 ;
        RECT 2.774 0.248 2.842 0.292 ;
        RECT 3.206 0.248 3.274 0.292 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0549 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0621 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.338 3.49 0.382 ;
        RECT 2.45 0.338 2.518 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
        RECT 2.666 0.338 2.734 0.382 ;
        RECT 2.99 0.338 3.058 0.382 ;
        RECT 3.314 0.338 3.382 0.382 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.338 4.246 0.382 ;
        RECT 4.178 0.158 4.246 0.382 ;
        RECT 3.53 0.158 4.246 0.202 ;
        RECT 4.07 0.338 4.138 0.472 ;
        RECT 3.854 0.338 3.922 0.472 ;
        RECT 3.638 0.338 3.706 0.472 ;
      LAYER v0 ;
        RECT 3.64 0.408 3.704 0.452 ;
        RECT 3.638 0.158 3.706 0.202 ;
        RECT 3.856 0.408 3.92 0.452 ;
        RECT 3.854 0.158 3.922 0.202 ;
        RECT 4.072 0.408 4.136 0.452 ;
        RECT 4.07 0.158 4.138 0.202 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.79 0.202 ;
        RECT 0.614 0.338 0.682 0.472 ;
        RECT 0.074 0.338 0.682 0.382 ;
        RECT 0.398 0.338 0.466 0.472 ;
        RECT 0.29 0.158 0.358 0.382 ;
        RECT 0.182 0.338 0.25 0.472 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.184 0.408 0.248 0.452 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.4 0.408 0.464 0.452 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 0.616 0.408 0.68 0.452 ;
        RECT 0.614 0.158 0.682 0.202 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.354 0.652 ;
        RECT 4.178 0.518 4.246 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.206 0.518 3.274 0.652 ;
        RECT 2.99 0.518 3.058 0.652 ;
        RECT 2.774 0.518 2.842 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.518 2.194 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.372 0.538 1.436 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.128 0.538 2.192 0.582 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.776 0.538 2.84 0.582 ;
        RECT 2.992 0.538 3.056 0.582 ;
        RECT 3.208 0.538 3.272 0.582 ;
        RECT 3.532 0.538 3.596 0.582 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 4.18 0.538 4.244 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.354 0.022 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 3.746 -0.022 3.814 0.112 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 2.99 -0.022 3.058 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 2.128 0.048 2.192 0.092 ;
        RECT 2.344 0.048 2.408 0.092 ;
        RECT 2.56 0.048 2.624 0.092 ;
        RECT 2.992 0.048 3.056 0.092 ;
        RECT 3.532 0.048 3.596 0.092 ;
        RECT 3.748 0.048 3.812 0.092 ;
        RECT 3.964 0.048 4.028 0.092 ;
        RECT 4.18 0.048 4.244 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 2.558 0.428 2.626 0.562 ;
    LAYER v0 ;
      RECT 3.854 0.248 3.922 0.292 ;
      RECT 3.638 0.248 3.706 0.292 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.882 0.428 2.95 0.472 ;
      RECT 2.776 0.088 2.84 0.132 ;
      RECT 2.558 0.498 2.626 0.542 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.91 0.068 1.978 0.112 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.478 0.068 1.546 0.112 ;
      RECT 1.37 0.158 1.438 0.202 ;
      RECT 1.262 0.068 1.33 0.112 ;
      RECT 1.154 0.158 1.222 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 0.94 0.228 1.004 0.272 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.506 0.248 0.574 0.292 ;
    LAYER m1 ;
      RECT 0.486 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 0.898 0.068 1.998 0.112 ;
      RECT 0.898 0.428 2.41 0.472 ;
      RECT 1.006 0.158 2.626 0.202 ;
      RECT 2.774 0.068 2.842 0.202 ;
      RECT 2.842 0.158 3.422 0.202 ;
      RECT 3.422 0.158 3.49 0.292 ;
      RECT 2.626 0.428 3.53 0.472 ;
      RECT 3.49 0.248 3.53 0.292 ;
      RECT 3.53 0.248 3.598 0.472 ;
      RECT 3.598 0.248 3.942 0.292 ;
  END
END b15rt0022es1n24x5

MACRO b15ru0022as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0022as1n02x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 7.0775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.53875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.518 0.898 0.562 ;
        RECT 0.83 0.068 0.898 0.562 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
        RECT 0.398 0.518 0.466 0.562 ;
        RECT 0.83 0.088 0.898 0.132 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.068 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.158 1.438 0.562 ;
      LAYER v0 ;
        RECT 1.37 0.4175 1.438 0.4615 ;
        RECT 1.37 0.203 1.438 0.247 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.486 0.428 0.682 0.472 ;
        RECT 0.614 0.158 0.682 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.614 0.203 0.682 0.247 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.154 0.4175 1.222 0.4615 ;
        RECT 1.478 0.4175 1.546 0.4615 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 0.938 -0.022 1.006 0.292 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.938 0.203 1.006 0.247 ;
        RECT 1.478 0.203 1.546 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.378 0.068 0.722 0.112 ;
      RECT 1.262 0.158 1.33 0.562 ;
    LAYER v0 ;
      RECT 1.262 0.203 1.33 0.247 ;
      RECT 1.262 0.498 1.33 0.542 ;
      RECT 0.722 0.203 0.79 0.247 ;
      RECT 0.506 0.293 0.574 0.337 ;
      RECT 0.398 0.068 0.466 0.112 ;
      RECT 0.074 0.428 0.142 0.472 ;
      RECT 0.076 0.229 0.14 0.273 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.142 0.158 0.506 0.202 ;
      RECT 0.506 0.158 0.574 0.382 ;
      RECT 0.722 0.068 0.79 0.292 ;
  END
END b15ru0022as1n02x5

MACRO b15ru0022as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0022as1n03x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0135 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0135 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.1355 0.898 0.1795 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0135 LAYER m1 ;
      ANTENNAMAXAREACAR 0.65866675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.068 1.438 0.472 ;
        RECT 1.154 0.068 1.438 0.112 ;
        RECT 1.154 0.068 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0027 LAYER m1 ;
      ANTENNAMAXAREACAR 3.67333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0027 LAYER m1 ;
      ANTENNAMAXAREACAR 3.67333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.158 1.762 0.562 ;
      LAYER v0 ;
        RECT 1.694 0.4505 1.762 0.4945 ;
        RECT 1.694 0.203 1.762 0.247 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.472 ;
      LAYER v0 ;
        RECT 0.722 0.253 0.79 0.297 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.4505 0.358 0.4945 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 1.478 0.4505 1.546 0.4945 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.478 -0.022 1.546 0.292 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.2255 0.358 0.2695 ;
        RECT 1.046 0.1305 1.114 0.1745 ;
        RECT 1.478 0.1855 1.546 0.2295 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.472 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.262 0.158 1.33 0.562 ;
    LAYER v0 ;
      RECT 1.262 0.198 1.33 0.242 ;
      RECT 1.262 0.4455 1.33 0.4895 ;
      RECT 1.046 0.433 1.114 0.477 ;
      RECT 0.938 0.2255 1.006 0.2695 ;
      RECT 0.832 0.448 0.896 0.492 ;
      RECT 0.614 0.1355 0.682 0.1795 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.182 0.2255 0.25 0.2695 ;
      RECT 0.182 0.4505 0.25 0.4945 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.338 0.506 0.382 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.574 0.518 0.83 0.562 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 1.006 0.338 1.046 0.382 ;
      RECT 1.046 0.338 1.114 0.562 ;
  END
END b15ru0022as1n03x5

MACRO b15ru0022as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0022as1n04x5 0 0 ;
  SIZE 1.728 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 4.120625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 3.66277775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.248 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.37 0.383 1.438 0.427 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0162 LAYER m1 ;
      ANTENNAMAXAREACAR 0.80222225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0189 LAYER m1 ;
      ANTENNAMAXAREACAR 0.687619 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.382 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.472 ;
      LAYER v0 ;
        RECT 1.586 0.408 1.654 0.452 ;
        RECT 1.586 0.178 1.654 0.222 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.408 0.25 0.452 ;
        RECT 0.182 0.178 0.25 0.222 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
      LAYER v0 ;
        RECT 0.614 0.448 0.682 0.492 ;
        RECT 0.83 0.466 0.898 0.51 ;
        RECT 1.046 0.466 1.114 0.51 ;
        RECT 1.262 0.466 1.33 0.51 ;
        RECT 1.478 0.49 1.546 0.534 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.762 0.022 ;
        RECT 1.478 -0.022 1.546 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.614 -0.022 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.614 0.178 0.682 0.222 ;
        RECT 0.83 0.178 0.898 0.222 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 1.478 0.048 1.546 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 0.938 0.068 1.006 0.472 ;
    LAYER v0 ;
      RECT 1.478 0.293 1.546 0.337 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.398 0.088 0.466 0.132 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.29 0.178 0.358 0.222 ;
      RECT 0.074 0.408 0.142 0.452 ;
    LAYER m1 ;
      RECT 0.074 0.338 0.142 0.562 ;
      RECT 0.142 0.518 0.29 0.562 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.358 0.518 0.506 0.562 ;
      RECT 0.506 0.338 0.574 0.562 ;
      RECT 0.574 0.338 0.898 0.382 ;
      RECT 1.222 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.382 ;
  END
END b15ru0022as1n04x5

MACRO b15ru0022as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0022as1n06x5 0 0 ;
  SIZE 2.16 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.018 LAYER m1 ;
      ANTENNAMAXAREACAR 3.1065 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 2.4852 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.202 ;
      LAYER v0 ;
        RECT 0.614 0.088 0.682 0.132 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0243 LAYER m1 ;
      ANTENNAMAXAREACAR 1.4214815 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0261 LAYER m1 ;
      ANTENNAMAXAREACAR 1.32344825 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.428 1.114 0.562 ;
      LAYER v0 ;
        RECT 1.046 0.498 1.114 0.542 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.158 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 1.91 0.203 1.978 0.247 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.158 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.4 0.898 0.444 ;
        RECT 0.83 0.2475 0.898 0.2915 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.194 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 1.154 0.338 1.222 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 1.154 0.377 1.222 0.421 ;
        RECT 1.37 0.4665 1.438 0.5105 ;
        RECT 1.586 0.4665 1.654 0.5105 ;
        RECT 1.802 0.4665 1.87 0.5105 ;
        RECT 2.018 0.4665 2.086 0.5105 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.194 0.022 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.1185 0.142 0.1625 ;
        RECT 0.29 0.1185 0.358 0.1625 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 1.37 0.138 1.438 0.182 ;
        RECT 1.802 0.048 1.87 0.092 ;
        RECT 2.018 0.102 2.086 0.146 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.248 0.722 0.292 ;
      RECT 1.478 0.158 1.546 0.562 ;
    LAYER v0 ;
      RECT 1.802 0.293 1.87 0.337 ;
      RECT 1.694 0.4665 1.762 0.5105 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.4665 1.546 0.5105 ;
      RECT 1.262 0.138 1.33 0.182 ;
      RECT 1.262 0.377 1.33 0.421 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.4 1.006 0.444 ;
      RECT 0.722 0.4 0.79 0.444 ;
      RECT 0.614 0.4 0.682 0.444 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.182 0.1185 0.25 0.1625 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.006 0.248 1.262 0.292 ;
      RECT 1.262 0.068 1.33 0.472 ;
      RECT 1.546 0.338 1.694 0.382 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.546 0.158 1.802 0.202 ;
      RECT 1.802 0.158 1.87 0.382 ;
  END
END b15ru0022as1n06x5

MACRO b15ru0022as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0022as1n08x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 2.87923075 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.027 LAYER m1 ;
      ANTENNAMAXAREACAR 2.49533325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.81 0.112 ;
        RECT 0.506 0.068 0.574 0.202 ;
      LAYER v0 ;
        RECT 0.614 0.068 0.682 0.112 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0324 LAYER m1 ;
      ANTENNAMAXAREACAR 1.32472225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0342 LAYER m1 ;
      ANTENNAMAXAREACAR 1.255 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.248 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.363 1.33 0.407 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.158 2.302 0.472 ;
      LAYER v0 ;
        RECT 2.234 0.383 2.302 0.427 ;
        RECT 2.234 0.203 2.302 0.247 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.472 ;
        RECT 0.614 0.158 1.222 0.202 ;
      LAYER v0 ;
        RECT 0.722 0.158 0.79 0.202 ;
        RECT 0.938 0.158 1.006 0.202 ;
        RECT 1.154 0.363 1.222 0.407 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 1.478 0.4665 1.546 0.5105 ;
        RECT 1.694 0.4665 1.762 0.5105 ;
        RECT 1.91 0.4665 1.978 0.5105 ;
        RECT 2.126 0.4665 2.194 0.5105 ;
        RECT 2.342 0.538 2.41 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.138 0.142 0.182 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 2.126 0.048 2.194 0.092 ;
        RECT 2.342 0.102 2.41 0.146 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.248 0.918 0.292 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 1.802 0.158 1.87 0.562 ;
    LAYER v0 ;
      RECT 2.126 0.293 2.194 0.337 ;
      RECT 2.018 0.4665 2.086 0.5105 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.802 0.4665 1.87 0.5105 ;
      RECT 1.586 0.138 1.654 0.182 ;
      RECT 1.586 0.363 1.654 0.407 ;
      RECT 1.37 0.138 1.438 0.182 ;
      RECT 1.37 0.363 1.438 0.407 ;
      RECT 1.048 0.268 1.112 0.312 ;
      RECT 1.048 0.448 1.112 0.492 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.616 0.448 0.68 0.492 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 1.046 0.382 ;
      RECT 1.046 0.248 1.114 0.382 ;
      RECT 0.682 0.518 1.046 0.562 ;
      RECT 1.046 0.428 1.114 0.562 ;
      RECT 1.114 0.518 1.37 0.562 ;
      RECT 1.37 0.068 1.438 0.562 ;
      RECT 1.438 0.248 1.586 0.292 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.87 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 1.87 0.158 2.126 0.202 ;
      RECT 2.126 0.158 2.194 0.382 ;
  END
END b15ru0022as1n08x5

MACRO b15ru0022as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0022as1n12x5 0 0 ;
  SIZE 2.916 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0324 LAYER m1 ;
      ANTENNAMAXAREACAR 2.3855555 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0369 LAYER m1 ;
      ANTENNAMAXAREACAR 2.09463425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.202 ;
      LAYER v0 ;
        RECT 1.478 0.138 1.546 0.182 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0414 LAYER m1 ;
      ANTENNAMAXAREACAR 1.073913 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 1.00816325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.35 0.518 1.546 0.562 ;
        RECT 1.478 0.428 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.448 1.546 0.492 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.068 2.842 0.472 ;
        RECT 2.558 0.248 2.842 0.292 ;
        RECT 2.558 0.068 2.626 0.472 ;
      LAYER v0 ;
        RECT 2.558 0.383 2.626 0.427 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.774 0.383 2.842 0.427 ;
        RECT 2.774 0.138 2.842 0.182 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 1.33 0.382 ;
        RECT 1.262 0.158 1.33 0.382 ;
        RECT 0.83 0.248 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.832 0.268 0.896 0.312 ;
        RECT 1.046 0.338 1.114 0.382 ;
        RECT 1.262 0.178 1.33 0.222 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.95 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.018 0.4665 2.086 0.5105 ;
        RECT 2.234 0.4665 2.302 0.5105 ;
        RECT 2.45 0.4665 2.518 0.5105 ;
        RECT 2.666 0.4665 2.734 0.5105 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.95 0.022 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.137 0.358 0.181 ;
        RECT 0.506 0.137 0.574 0.181 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.45 0.048 2.518 0.092 ;
        RECT 2.666 0.138 2.734 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.338 0.614 0.382 ;
      RECT 2.126 0.158 2.194 0.562 ;
    LAYER v0 ;
      RECT 2.45 0.293 2.518 0.337 ;
      RECT 2.342 0.4665 2.41 0.5105 ;
      RECT 2.234 0.158 2.302 0.202 ;
      RECT 2.126 0.4665 2.194 0.5105 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 1.154 0.518 1.222 0.562 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.398 0.137 0.466 0.181 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.137 0.25 0.181 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.074 0.428 0.29 0.472 ;
      RECT 0.25 0.248 0.29 0.292 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.358 0.248 0.398 0.292 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.358 0.428 0.722 0.472 ;
      RECT 0.722 0.158 0.79 0.562 ;
      RECT 0.79 0.158 1.026 0.202 ;
      RECT 0.79 0.518 1.242 0.562 ;
      RECT 0.614 0.068 0.682 0.382 ;
      RECT 0.682 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 0.918 0.428 1.37 0.472 ;
      RECT 1.222 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.472 ;
      RECT 1.438 0.338 2.086 0.382 ;
      RECT 2.194 0.338 2.342 0.382 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.194 0.158 2.45 0.202 ;
      RECT 2.45 0.158 2.518 0.382 ;
  END
END b15ru0022as1n12x5

MACRO b15ru0022as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0022as1n16x5 0 0 ;
  SIZE 4.104 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0504 LAYER m1 ;
      ANTENNAMAXAREACAR 2.33428575 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0567 LAYER m1 ;
      ANTENNAMAXAREACAR 2.07492075 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.292 ;
      LAYER v0 ;
        RECT 1.802 0.228 1.87 0.272 ;
        RECT 1.802 0.0925 1.87 0.1365 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 1.26171875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0666 LAYER m1 ;
      ANTENNAMAXAREACAR 1.09121625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.248 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.4665 2.734 0.5105 ;
        RECT 2.666 0.327 2.734 0.371 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.854 0.068 3.922 0.562 ;
        RECT 3.638 0.338 3.922 0.382 ;
        RECT 3.638 0.068 3.706 0.562 ;
      LAYER v0 ;
        RECT 3.638 0.4665 3.706 0.5105 ;
        RECT 3.638 0.114 3.706 0.158 ;
        RECT 3.854 0.4665 3.922 0.5105 ;
        RECT 3.854 0.114 3.922 0.158 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.338 1.654 0.382 ;
        RECT 1.586 0.158 1.654 0.382 ;
      LAYER v0 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.37 0.338 1.438 0.382 ;
        RECT 1.586 0.228 1.654 0.272 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.138 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 2.342 0.428 2.41 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 2.126 0.448 2.194 0.492 ;
        RECT 2.342 0.4665 2.41 0.5105 ;
        RECT 2.558 0.4665 2.626 0.5105 ;
        RECT 2.774 0.4665 2.842 0.5105 ;
        RECT 2.99 0.4665 3.058 0.5105 ;
        RECT 3.206 0.4665 3.274 0.5105 ;
        RECT 3.422 0.4665 3.49 0.5105 ;
        RECT 3.746 0.4665 3.814 0.5105 ;
        RECT 3.962 0.4665 4.03 0.5105 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.138 0.022 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 1.91 -0.022 1.978 0.292 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.202 ;
      LAYER v0 ;
        RECT 0.074 0.137 0.142 0.181 ;
        RECT 0.29 0.137 0.358 0.181 ;
        RECT 0.506 0.137 0.574 0.181 ;
        RECT 0.722 0.137 0.79 0.181 ;
        RECT 1.91 0.228 1.978 0.272 ;
        RECT 2.126 0.138 2.194 0.182 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
        RECT 2.99 0.138 3.058 0.182 ;
        RECT 3.422 0.138 3.49 0.182 ;
        RECT 3.746 0.114 3.814 0.158 ;
        RECT 3.962 0.114 4.03 0.158 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.27 0.338 0.506 0.382 ;
      RECT 2.774 0.068 2.842 0.292 ;
    LAYER v0 ;
      RECT 3.53 0.338 3.598 0.382 ;
      RECT 3.314 0.4665 3.382 0.5105 ;
      RECT 3.206 0.138 3.274 0.182 ;
      RECT 3.098 0.4665 3.166 0.5105 ;
      RECT 2.882 0.385 2.95 0.429 ;
      RECT 2.774 0.138 2.842 0.182 ;
      RECT 2.45 0.223 2.518 0.267 ;
      RECT 2.45 0.4665 2.518 0.5105 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.018 0.228 2.086 0.272 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.694 0.228 1.762 0.272 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.478 0.228 1.546 0.272 ;
      RECT 1.478 0.518 1.546 0.562 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.398 0.137 0.466 0.181 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.29 0.338 0.358 0.382 ;
      RECT 0.182 0.137 0.25 0.181 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.472 ;
      RECT 0.142 0.248 0.182 0.292 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.142 0.428 0.614 0.472 ;
      RECT 0.614 0.338 0.682 0.472 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.338 0.938 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.006 0.158 1.438 0.202 ;
      RECT 0.898 0.518 1.782 0.562 ;
      RECT 0.506 0.248 0.574 0.382 ;
      RECT 0.574 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 0.898 0.068 1.478 0.112 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 0.938 0.428 1.694 0.472 ;
      RECT 1.546 0.068 1.694 0.112 ;
      RECT 1.694 0.068 1.762 0.472 ;
      RECT 1.762 0.338 2.018 0.382 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 2.086 0.338 2.45 0.382 ;
      RECT 2.45 0.158 2.518 0.562 ;
      RECT 2.842 0.248 2.882 0.292 ;
      RECT 2.882 0.248 2.95 0.472 ;
      RECT 2.95 0.248 3.098 0.292 ;
      RECT 3.098 0.248 3.166 0.562 ;
      RECT 3.166 0.248 3.206 0.292 ;
      RECT 3.206 0.068 3.274 0.292 ;
      RECT 3.274 0.248 3.314 0.292 ;
      RECT 3.314 0.248 3.382 0.562 ;
      RECT 3.382 0.248 3.53 0.292 ;
      RECT 3.53 0.248 3.598 0.472 ;
  END
END b15ru0022as1n16x5

MACRO b15ru0022as1n24x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0022as1n24x5 0 0 ;
  SIZE 5.4 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0675 LAYER m1 ;
      ANTENNAMAXAREACAR 2.16853325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0738 LAYER m1 ;
      ANTENNAMAXAREACAR 1.98341475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.068 2.518 0.292 ;
      LAYER v0 ;
        RECT 2.45 0.228 2.518 0.272 ;
        RECT 2.45 0.092 2.518 0.136 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0801 LAYER m1 ;
      ANTENNAMAXAREACAR 1.090899 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0882 LAYER m1 ;
      ANTENNAMAXAREACAR 0.99071425 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.158 3.598 0.562 ;
      LAYER v0 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 3.53 0.314 3.598 0.358 ;
    END
  END b
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.15 0.068 5.218 0.562 ;
        RECT 4.718 0.248 5.218 0.292 ;
        RECT 4.934 0.068 5.002 0.562 ;
        RECT 4.718 0.068 4.786 0.562 ;
      LAYER v0 ;
        RECT 4.718 0.448 4.786 0.492 ;
        RECT 4.718 0.1115 4.786 0.1555 ;
        RECT 4.934 0.448 5.002 0.492 ;
        RECT 4.934 0.1115 5.002 0.1555 ;
        RECT 5.15 0.448 5.218 0.492 ;
        RECT 5.15 0.1115 5.218 0.1555 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.338 2.302 0.382 ;
        RECT 2.234 0.158 2.302 0.382 ;
        RECT 1.37 0.248 1.438 0.382 ;
      LAYER v0 ;
        RECT 1.372 0.268 1.436 0.312 ;
        RECT 1.586 0.338 1.654 0.382 ;
        RECT 1.802 0.338 1.87 0.382 ;
        RECT 2.018 0.338 2.086 0.382 ;
        RECT 2.234 0.2055 2.302 0.2495 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.434 0.652 ;
        RECT 5.258 0.428 5.326 0.652 ;
        RECT 5.042 0.428 5.11 0.652 ;
        RECT 4.826 0.428 4.894 0.652 ;
        RECT 4.502 0.428 4.57 0.652 ;
        RECT 4.286 0.428 4.354 0.652 ;
        RECT 4.07 0.428 4.138 0.652 ;
        RECT 3.854 0.428 3.922 0.652 ;
        RECT 3.638 0.428 3.706 0.652 ;
        RECT 3.422 0.428 3.49 0.652 ;
        RECT 3.206 0.428 3.274 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.558 0.428 2.626 0.652 ;
        RECT 1.046 0.428 1.114 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.428 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.448 0.142 0.492 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.046 0.448 1.114 0.492 ;
        RECT 2.558 0.448 2.626 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 3.206 0.448 3.274 0.492 ;
        RECT 3.422 0.448 3.49 0.492 ;
        RECT 3.638 0.448 3.706 0.492 ;
        RECT 3.854 0.448 3.922 0.492 ;
        RECT 4.07 0.448 4.138 0.492 ;
        RECT 4.286 0.448 4.354 0.492 ;
        RECT 4.502 0.448 4.57 0.492 ;
        RECT 4.826 0.448 4.894 0.492 ;
        RECT 5.042 0.448 5.11 0.492 ;
        RECT 5.258 0.448 5.326 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.434 0.022 ;
        RECT 5.258 -0.022 5.326 0.202 ;
        RECT 5.042 -0.022 5.11 0.202 ;
        RECT 4.826 -0.022 4.894 0.202 ;
        RECT 4.502 -0.022 4.57 0.202 ;
        RECT 4.07 -0.022 4.138 0.202 ;
        RECT 3.638 -0.022 3.706 0.202 ;
        RECT 3.422 -0.022 3.49 0.202 ;
        RECT 3.206 -0.022 3.274 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.558 -0.022 2.626 0.292 ;
        RECT 1.046 -0.022 1.114 0.202 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 1.046 0.138 1.114 0.182 ;
        RECT 2.558 0.228 2.626 0.272 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 2.99 0.138 3.058 0.182 ;
        RECT 3.206 0.138 3.274 0.182 ;
        RECT 3.422 0.138 3.49 0.182 ;
        RECT 3.638 0.138 3.706 0.182 ;
        RECT 4.07 0.138 4.138 0.182 ;
        RECT 4.502 0.138 4.57 0.182 ;
        RECT 4.826 0.1115 4.894 0.1555 ;
        RECT 5.042 0.1115 5.11 0.1555 ;
        RECT 5.258 0.1115 5.326 0.1555 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.248 1.154 0.292 ;
      RECT 3.746 0.248 3.814 0.472 ;
    LAYER v0 ;
      RECT 4.61 0.338 4.678 0.382 ;
      RECT 4.394 0.366 4.462 0.41 ;
      RECT 4.288 0.1685 4.352 0.2125 ;
      RECT 4.178 0.366 4.246 0.41 ;
      RECT 3.962 0.366 4.03 0.41 ;
      RECT 3.856 0.1685 3.92 0.2125 ;
      RECT 3.746 0.366 3.814 0.41 ;
      RECT 3.314 0.228 3.382 0.272 ;
      RECT 3.314 0.448 3.382 0.492 ;
      RECT 3.098 0.338 3.166 0.382 ;
      RECT 2.882 0.228 2.95 0.272 ;
      RECT 2.882 0.448 2.95 0.492 ;
      RECT 2.666 0.228 2.734 0.272 ;
      RECT 2.666 0.448 2.734 0.492 ;
      RECT 2.126 0.2055 2.194 0.2495 ;
      RECT 2.126 0.518 2.194 0.562 ;
      RECT 1.91 0.2055 1.978 0.2495 ;
      RECT 1.91 0.518 1.978 0.562 ;
      RECT 1.694 0.158 1.762 0.202 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.29 0.248 0.358 0.292 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.382 ;
      RECT 0.142 0.338 0.182 0.382 ;
      RECT 0.182 0.338 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.142 0.158 0.79 0.202 ;
      RECT 0.466 0.338 1.262 0.382 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.33 0.158 1.87 0.202 ;
      RECT 1.33 0.518 2.302 0.562 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.292 ;
      RECT 1.978 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 1.458 0.428 2.342 0.472 ;
      RECT 2.194 0.068 2.342 0.112 ;
      RECT 2.342 0.068 2.41 0.472 ;
      RECT 2.41 0.338 2.666 0.382 ;
      RECT 2.666 0.158 2.734 0.562 ;
      RECT 2.734 0.338 2.882 0.382 ;
      RECT 2.882 0.158 2.95 0.562 ;
      RECT 2.95 0.338 3.314 0.382 ;
      RECT 3.314 0.158 3.382 0.562 ;
      RECT 3.814 0.248 3.854 0.292 ;
      RECT 3.854 0.068 3.922 0.292 ;
      RECT 3.922 0.248 3.962 0.292 ;
      RECT 3.962 0.248 4.03 0.472 ;
      RECT 4.03 0.248 4.178 0.292 ;
      RECT 4.178 0.248 4.246 0.472 ;
      RECT 4.246 0.248 4.286 0.292 ;
      RECT 4.286 0.068 4.354 0.292 ;
      RECT 4.354 0.248 4.394 0.292 ;
      RECT 4.394 0.248 4.462 0.472 ;
      RECT 4.462 0.248 4.61 0.292 ;
      RECT 4.61 0.248 4.678 0.472 ;
  END
END b15ru0022as1n24x5

MACRO b15ru0023as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0023as1n02x3 0 0 ;
  SIZE 3.132 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.248 2.95 0.472 ;
      LAYER v0 ;
        RECT 2.882 0.3155 2.95 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.1325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.223 0.142 0.267 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.37 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 4.37 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.428 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.448 1.546 0.492 ;
    END
  END c
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.472 ;
      LAYER v0 ;
        RECT 2.018 0.408 2.086 0.452 ;
        RECT 2.018 0.202 2.086 0.246 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.158 2.518 0.472 ;
      LAYER v0 ;
        RECT 2.45 0.408 2.518 0.452 ;
        RECT 2.45 0.2225 2.518 0.2665 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 2.882 0.538 2.95 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.166 0.022 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.248 0.614 0.292 ;
      RECT 0.486 0.338 0.83 0.382 ;
      RECT 0.81 0.428 1.134 0.472 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 2.342 0.068 2.41 0.292 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 2.99 0.068 3.058 0.472 ;
    LAYER v0 ;
      RECT 2.99 0.138 3.058 0.182 ;
      RECT 2.99 0.408 3.058 0.452 ;
      RECT 2.774 0.138 2.842 0.182 ;
      RECT 2.774 0.408 2.842 0.452 ;
      RECT 2.666 0.2225 2.734 0.2665 ;
      RECT 2.666 0.408 2.734 0.452 ;
      RECT 2.558 0.2225 2.626 0.2665 ;
      RECT 2.342 0.2225 2.41 0.2665 ;
      RECT 2.342 0.408 2.41 0.452 ;
      RECT 2.234 0.2225 2.302 0.2665 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 1.91 0.202 1.978 0.246 ;
      RECT 1.802 0.493 1.87 0.537 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.832 0.268 0.896 0.312 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.182 0.223 0.25 0.267 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.182 0.472 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.428 0.702 0.472 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.158 1.026 0.202 ;
      RECT 0.83 0.248 0.898 0.382 ;
      RECT 0.898 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 0.938 0.248 1.154 0.292 ;
      RECT 0.574 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.248 1.694 0.292 ;
      RECT 1.694 0.068 1.762 0.292 ;
      RECT 1.762 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.41 0.068 2.666 0.112 ;
      RECT 2.666 0.068 2.734 0.472 ;
      RECT 1.978 0.518 2.126 0.562 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.194 0.518 2.342 0.562 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.41 0.518 2.558 0.562 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 2.626 0.518 2.774 0.562 ;
      RECT 2.774 0.068 2.842 0.562 ;
  END
END b15ru0023as1n02x3

MACRO b15ru0023as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0023as1n02x5 0 0 ;
  SIZE 3.132 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.248 2.95 0.472 ;
      LAYER v0 ;
        RECT 2.882 0.338 2.95 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.59666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.272 0.142 0.316 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 2.91333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.428 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.448 1.546 0.492 ;
    END
  END c
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.472 ;
      LAYER v0 ;
        RECT 2.018 0.3965 2.086 0.4405 ;
        RECT 2.018 0.202 2.086 0.246 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.158 2.518 0.472 ;
      LAYER v0 ;
        RECT 2.45 0.383 2.518 0.427 ;
        RECT 2.45 0.178 2.518 0.222 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 2.884 0.538 2.948 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.166 0.022 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.884 0.048 2.948 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.29 0.248 0.614 0.292 ;
      RECT 0.486 0.338 0.83 0.382 ;
      RECT 0.81 0.428 1.134 0.472 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 2.342 0.068 2.41 0.292 ;
    LAYER v0 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.992 0.228 3.056 0.272 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.666 0.338 2.734 0.382 ;
      RECT 2.558 0.178 2.626 0.222 ;
      RECT 2.342 0.178 2.41 0.222 ;
      RECT 2.342 0.383 2.41 0.427 ;
      RECT 2.234 0.178 2.302 0.222 ;
      RECT 2.126 0.3965 2.194 0.4405 ;
      RECT 1.91 0.202 1.978 0.246 ;
      RECT 1.802 0.493 1.87 0.537 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.832 0.268 0.896 0.312 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.054 0.428 0.182 0.472 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.428 0.702 0.472 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.158 1.026 0.202 ;
      RECT 0.83 0.248 0.898 0.382 ;
      RECT 0.898 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 0.938 0.248 1.154 0.292 ;
      RECT 0.574 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.248 1.694 0.292 ;
      RECT 1.694 0.068 1.762 0.292 ;
      RECT 1.762 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 1.978 0.518 2.126 0.562 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.194 0.518 2.342 0.562 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.41 0.518 2.558 0.562 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 2.626 0.518 2.774 0.562 ;
      RECT 2.774 0.338 2.842 0.562 ;
      RECT 2.41 0.068 2.666 0.112 ;
      RECT 2.666 0.068 2.734 0.472 ;
      RECT 2.734 0.158 2.99 0.202 ;
      RECT 2.99 0.158 3.058 0.562 ;
  END
END b15ru0023as1n02x5

MACRO b15ru0023as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0023as1n03x5 0 0 ;
  SIZE 3.24 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.158 3.166 0.472 ;
      LAYER v0 ;
        RECT 3.098 0.293 3.166 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.09777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.09777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.3155 0.142 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.428 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.4865 1.546 0.5305 ;
    END
  END c
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.158 2.086 0.472 ;
      LAYER v0 ;
        RECT 2.018 0.408 2.086 0.452 ;
        RECT 2.018 0.202 2.086 0.246 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.158 2.518 0.472 ;
      LAYER v0 ;
        RECT 2.45 0.408 2.518 0.452 ;
        RECT 2.45 0.178 2.518 0.222 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.274 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.586 0.4865 1.654 0.5305 ;
        RECT 2.882 0.493 2.95 0.537 ;
        RECT 3.098 0.538 3.166 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.274 0.022 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.292 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 2.882 0.178 2.95 0.222 ;
        RECT 3.1 0.048 3.164 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.486 0.338 0.83 0.382 ;
      RECT 0.81 0.428 1.134 0.472 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 2.342 0.068 2.41 0.292 ;
      RECT 1.91 0.158 1.978 0.562 ;
      RECT 2.99 0.158 3.058 0.472 ;
    LAYER v0 ;
      RECT 2.99 0.178 3.058 0.222 ;
      RECT 2.99 0.408 3.058 0.452 ;
      RECT 2.774 0.178 2.842 0.222 ;
      RECT 2.774 0.408 2.842 0.452 ;
      RECT 2.666 0.178 2.734 0.222 ;
      RECT 2.666 0.408 2.734 0.452 ;
      RECT 2.558 0.178 2.626 0.222 ;
      RECT 2.342 0.178 2.41 0.222 ;
      RECT 2.342 0.408 2.41 0.452 ;
      RECT 2.234 0.178 2.302 0.222 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 1.91 0.202 1.978 0.246 ;
      RECT 1.802 0.493 1.87 0.537 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.832 0.268 0.896 0.312 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.074 0.428 0.29 0.472 ;
      RECT 0.25 0.248 0.29 0.292 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.358 0.428 0.702 0.472 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.158 1.026 0.202 ;
      RECT 0.83 0.248 0.898 0.382 ;
      RECT 0.898 0.338 1.802 0.382 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 0.938 0.248 1.154 0.292 ;
      RECT 0.574 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.248 1.694 0.292 ;
      RECT 1.694 0.068 1.762 0.292 ;
      RECT 1.762 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.292 ;
      RECT 2.41 0.068 2.666 0.112 ;
      RECT 2.666 0.068 2.734 0.472 ;
      RECT 1.978 0.518 2.126 0.562 ;
      RECT 2.126 0.338 2.194 0.562 ;
      RECT 2.194 0.518 2.342 0.562 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.41 0.518 2.558 0.562 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 2.626 0.518 2.774 0.562 ;
      RECT 2.774 0.158 2.842 0.562 ;
  END
END b15ru0023as1n03x5

MACRO b15ru0023as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0023as1n04x5 0 0 ;
  SIZE 3.672 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.158 3.598 0.472 ;
      LAYER v0 ;
        RECT 3.53 0.293 3.598 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83666675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.338 1.654 0.562 ;
      LAYER v0 ;
        RECT 1.586 0.448 1.654 0.492 ;
    END
  END c
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.428 2.43 0.472 ;
        RECT 2.126 0.158 2.194 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.428 2.41 0.472 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.158 2.842 0.382 ;
      LAYER v0 ;
        RECT 2.774 0.1825 2.842 0.2265 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.706 0.652 ;
        RECT 3.53 0.518 3.598 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 1.91 0.428 1.978 0.652 ;
        RECT 1.694 0.428 1.762 0.652 ;
        RECT 1.478 0.428 1.546 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 1.262 0.448 1.33 0.492 ;
        RECT 1.478 0.448 1.546 0.492 ;
        RECT 1.694 0.448 1.762 0.492 ;
        RECT 1.91 0.448 1.978 0.492 ;
        RECT 3.098 0.538 3.166 0.582 ;
        RECT 3.314 0.538 3.382 0.582 ;
        RECT 3.53 0.538 3.598 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.706 0.022 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 1.91 -0.022 1.978 0.202 ;
        RECT 1.694 -0.022 1.762 0.202 ;
        RECT 1.478 -0.022 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 1.262 0.138 1.33 0.182 ;
        RECT 1.478 0.138 1.546 0.182 ;
        RECT 1.694 0.138 1.762 0.182 ;
        RECT 1.91 0.138 1.978 0.182 ;
        RECT 3.098 0.138 3.166 0.182 ;
        RECT 3.314 0.138 3.382 0.182 ;
        RECT 3.53 0.048 3.598 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.352 0.158 2.644 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.506 0.068 0.574 0.202 ;
      RECT 0.81 0.428 1.134 0.472 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 0.398 0.338 0.83 0.382 ;
      RECT 2.558 0.068 2.626 0.202 ;
      RECT 2.234 0.158 2.302 0.382 ;
      RECT 2.666 0.068 2.734 0.292 ;
    LAYER v1 ;
      RECT 2.562 0.158 2.622 0.202 ;
      RECT 1.374 0.158 1.434 0.202 ;
    LAYER v0 ;
      RECT 3.422 0.138 3.49 0.182 ;
      RECT 3.424 0.408 3.488 0.452 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 2.992 0.268 3.056 0.312 ;
      RECT 2.882 0.1825 2.95 0.2265 ;
      RECT 2.666 0.1825 2.734 0.2265 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.558 0.088 2.626 0.132 ;
      RECT 2.558 0.518 2.626 0.562 ;
      RECT 2.45 0.1825 2.518 0.2265 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.234 0.1825 2.302 0.2265 ;
      RECT 2.126 0.518 2.194 0.562 ;
      RECT 2.018 0.138 2.086 0.182 ;
      RECT 1.802 0.138 1.87 0.182 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.832 0.268 0.896 0.312 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.074 0.428 0.29 0.472 ;
      RECT 0.25 0.248 0.29 0.292 ;
      RECT 0.29 0.248 0.358 0.472 ;
      RECT 0.358 0.428 0.702 0.472 ;
      RECT 0.466 0.248 0.614 0.292 ;
      RECT 0.614 0.158 0.682 0.292 ;
      RECT 0.682 0.158 1.026 0.202 ;
      RECT 1.026 0.248 1.154 0.292 ;
      RECT 0.574 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.87 0.248 2.018 0.292 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 2.086 0.068 2.45 0.112 ;
      RECT 2.45 0.068 2.518 0.292 ;
      RECT 0.83 0.248 0.898 0.382 ;
      RECT 0.898 0.338 1.478 0.382 ;
      RECT 1.478 0.248 1.546 0.382 ;
      RECT 1.546 0.248 1.694 0.292 ;
      RECT 1.694 0.248 1.762 0.382 ;
      RECT 1.762 0.338 2.018 0.382 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.086 0.518 2.646 0.562 ;
      RECT 2.302 0.338 2.558 0.382 ;
      RECT 2.558 0.338 2.626 0.472 ;
      RECT 2.626 0.428 2.882 0.472 ;
      RECT 2.882 0.158 2.95 0.472 ;
      RECT 2.95 0.428 3.382 0.472 ;
      RECT 2.734 0.068 2.99 0.112 ;
      RECT 2.99 0.068 3.058 0.382 ;
      RECT 3.058 0.338 3.422 0.382 ;
      RECT 3.422 0.068 3.49 0.472 ;
  END
END b15ru0023as1n04x5

MACRO b15ru0023as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0023as1n06x5 0 0 ;
  SIZE 4.428 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.248 4.246 0.472 ;
      LAYER v0 ;
        RECT 4.178 0.338 4.246 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.3775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 1.3775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.338 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.448 1.978 0.492 ;
    END
  END c
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.45 0.518 2.95 0.562 ;
        RECT 2.882 0.338 2.95 0.562 ;
        RECT 2.666 0.338 2.734 0.562 ;
        RECT 2.45 0.338 2.518 0.562 ;
      LAYER v0 ;
        RECT 2.45 0.396 2.518 0.44 ;
        RECT 2.666 0.396 2.734 0.44 ;
        RECT 2.882 0.396 2.95 0.44 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.598 0.292 ;
        RECT 3.098 0.068 3.598 0.112 ;
        RECT 3.314 0.068 3.382 0.292 ;
        RECT 3.098 0.068 3.166 0.472 ;
      LAYER v0 ;
        RECT 3.098 0.223 3.166 0.267 ;
        RECT 3.314 0.223 3.382 0.267 ;
        RECT 3.53 0.223 3.598 0.267 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.462 0.652 ;
        RECT 4.178 0.518 4.246 0.652 ;
        RECT 3.962 0.518 4.03 0.652 ;
        RECT 3.746 0.518 3.814 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 2.018 0.428 2.086 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.506 0.5135 0.574 0.5575 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
        RECT 2.018 0.448 2.086 0.492 ;
        RECT 2.234 0.498 2.302 0.542 ;
        RECT 3.748 0.538 3.812 0.582 ;
        RECT 3.964 0.538 4.028 0.582 ;
        RECT 4.18 0.538 4.244 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.462 0.022 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 2.018 -0.022 2.086 0.202 ;
        RECT 1.802 -0.022 1.87 0.202 ;
        RECT 1.586 -0.022 1.654 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 1.586 0.138 1.654 0.182 ;
        RECT 1.802 0.138 1.87 0.182 ;
        RECT 2.018 0.138 2.086 0.182 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 3.746 0.138 3.814 0.182 ;
        RECT 3.962 0.138 4.03 0.182 ;
        RECT 4.178 0.048 4.246 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 1.676 0.158 2.428 0.202 ;
      RECT 3.188 0.158 4.156 0.202 ;
    LAYER m1 ;
      RECT 0.29 0.248 0.938 0.292 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 1.134 0.428 1.458 0.472 ;
      RECT 0.722 0.338 1.154 0.382 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.342 0.068 2.41 0.202 ;
      RECT 3.402 0.428 3.53 0.472 ;
      RECT 3.206 0.158 3.274 0.292 ;
      RECT 2.558 0.068 2.626 0.202 ;
      RECT 4.07 0.158 4.138 0.562 ;
    LAYER v1 ;
      RECT 4.074 0.158 4.134 0.202 ;
      RECT 3.642 0.158 3.702 0.202 ;
      RECT 3.21 0.158 3.27 0.202 ;
      RECT 2.346 0.158 2.406 0.202 ;
      RECT 1.698 0.158 1.758 0.202 ;
    LAYER v0 ;
      RECT 4.286 0.4405 4.354 0.4845 ;
      RECT 4.288 0.228 4.352 0.272 ;
      RECT 4.07 0.4405 4.138 0.4845 ;
      RECT 4.072 0.228 4.136 0.272 ;
      RECT 3.854 0.138 3.922 0.182 ;
      RECT 3.854 0.428 3.922 0.472 ;
      RECT 3.638 0.138 3.706 0.182 ;
      RECT 3.422 0.223 3.49 0.267 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 3.206 0.223 3.274 0.267 ;
      RECT 3.208 0.448 3.272 0.492 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.396 2.842 0.44 ;
      RECT 2.558 0.396 2.626 0.44 ;
      RECT 2.56 0.138 2.624 0.182 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.342 0.498 2.41 0.542 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 1.37 0.248 1.438 0.292 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.156 0.268 1.22 0.312 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.338 0.898 0.382 ;
      RECT 0.832 0.138 0.896 0.182 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.614 0.4255 0.682 0.4695 ;
      RECT 0.398 0.248 0.466 0.292 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.428 0.898 0.562 ;
      RECT 0.898 0.428 1.026 0.472 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.35 0.202 ;
      RECT 1.35 0.248 1.478 0.292 ;
      RECT 0.898 0.068 1.478 0.112 ;
      RECT 1.478 0.068 1.546 0.292 ;
      RECT 1.546 0.248 1.694 0.292 ;
      RECT 1.694 0.068 1.762 0.292 ;
      RECT 1.154 0.248 1.222 0.382 ;
      RECT 1.222 0.338 1.802 0.382 ;
      RECT 1.802 0.248 1.87 0.382 ;
      RECT 1.87 0.248 2.018 0.292 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 2.086 0.338 2.342 0.382 ;
      RECT 2.342 0.338 2.41 0.562 ;
      RECT 2.194 0.248 2.558 0.292 ;
      RECT 2.558 0.248 2.626 0.472 ;
      RECT 2.626 0.248 2.666 0.292 ;
      RECT 2.666 0.158 2.734 0.292 ;
      RECT 2.734 0.158 2.862 0.202 ;
      RECT 3.53 0.338 3.598 0.472 ;
      RECT 3.598 0.338 3.638 0.382 ;
      RECT 3.638 0.068 3.706 0.382 ;
      RECT 2.774 0.248 2.842 0.472 ;
      RECT 2.842 0.248 2.99 0.292 ;
      RECT 2.626 0.068 2.99 0.112 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.058 0.518 3.206 0.562 ;
      RECT 3.206 0.338 3.274 0.562 ;
      RECT 3.274 0.338 3.422 0.382 ;
      RECT 3.422 0.158 3.49 0.382 ;
      RECT 3.274 0.518 3.638 0.562 ;
      RECT 3.638 0.428 3.706 0.562 ;
      RECT 3.706 0.428 3.746 0.472 ;
      RECT 3.746 0.248 3.814 0.472 ;
      RECT 3.814 0.248 3.854 0.292 ;
      RECT 3.854 0.068 3.922 0.292 ;
      RECT 3.814 0.428 4.03 0.472 ;
      RECT 4.138 0.158 4.286 0.202 ;
      RECT 4.286 0.158 4.354 0.562 ;
  END
END b15ru0023as1n06x5

MACRO b15ru0023as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0023as1n08x5 0 0 ;
  SIZE 5.616 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.474 0.158 5.542 0.472 ;
      LAYER v0 ;
        RECT 5.474 0.293 5.542 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0234 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5553845 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.338 0.25 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.10833325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.10833325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.338 2.734 0.562 ;
      LAYER v0 ;
        RECT 2.666 0.448 2.734 0.492 ;
    END
  END c
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06732 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.518 3.814 0.562 ;
        RECT 3.746 0.338 3.814 0.562 ;
        RECT 3.53 0.338 3.598 0.562 ;
        RECT 3.314 0.338 3.382 0.562 ;
      LAYER v0 ;
        RECT 3.314 0.3985 3.382 0.4425 ;
        RECT 3.53 0.3985 3.598 0.4425 ;
        RECT 3.746 0.3985 3.814 0.4425 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.502 0.068 4.57 0.292 ;
        RECT 4.07 0.068 4.57 0.112 ;
        RECT 4.286 0.068 4.354 0.292 ;
        RECT 4.07 0.068 4.138 0.472 ;
      LAYER v0 ;
        RECT 4.07 0.228 4.138 0.272 ;
        RECT 4.286 0.228 4.354 0.272 ;
        RECT 4.502 0.228 4.57 0.272 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.65 0.652 ;
        RECT 5.474 0.518 5.542 0.652 ;
        RECT 5.258 0.428 5.326 0.652 ;
        RECT 5.042 0.428 5.11 0.652 ;
        RECT 4.826 0.518 4.894 0.652 ;
        RECT 2.99 0.428 3.058 0.652 ;
        RECT 2.774 0.428 2.842 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 2.234 0.428 2.302 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 2.234 0.448 2.302 0.492 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.774 0.448 2.842 0.492 ;
        RECT 2.99 0.448 3.058 0.492 ;
        RECT 4.826 0.538 4.894 0.582 ;
        RECT 5.042 0.455 5.11 0.499 ;
        RECT 5.258 0.455 5.326 0.499 ;
        RECT 5.474 0.538 5.542 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.65 0.022 ;
        RECT 5.474 -0.022 5.542 0.112 ;
        RECT 5.258 -0.022 5.326 0.202 ;
        RECT 5.042 -0.022 5.11 0.202 ;
        RECT 4.826 -0.022 4.894 0.202 ;
        RECT 2.99 -0.022 3.058 0.202 ;
        RECT 2.774 -0.022 2.842 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.138 0.682 0.182 ;
        RECT 2.234 0.138 2.302 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 2.774 0.138 2.842 0.182 ;
        RECT 2.99 0.138 3.058 0.182 ;
        RECT 4.826 0.138 4.894 0.182 ;
        RECT 5.042 0.138 5.11 0.182 ;
        RECT 5.258 0.138 5.326 0.182 ;
        RECT 5.474 0.048 5.542 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 2.324 0.158 4.064 0.202 ;
      RECT 4.144 0.158 5.236 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.248 0.722 0.292 ;
      RECT 0.722 0.068 1.046 0.112 ;
      RECT 1.35 0.428 2.106 0.472 ;
      RECT 0.83 0.248 0.898 0.382 ;
      RECT 2.882 0.068 2.95 0.292 ;
      RECT 4.374 0.428 4.61 0.472 ;
      RECT 3.962 0.158 4.03 0.292 ;
      RECT 4.178 0.158 4.246 0.292 ;
      RECT 3.402 0.158 3.53 0.202 ;
      RECT 5.15 0.068 5.218 0.562 ;
    LAYER v1 ;
      RECT 5.154 0.158 5.214 0.202 ;
      RECT 4.614 0.158 4.674 0.202 ;
      RECT 4.182 0.158 4.242 0.202 ;
      RECT 3.966 0.158 4.026 0.202 ;
      RECT 2.346 0.158 2.406 0.202 ;
    LAYER v0 ;
      RECT 5.366 0.138 5.434 0.182 ;
      RECT 5.366 0.455 5.434 0.499 ;
      RECT 5.15 0.138 5.218 0.182 ;
      RECT 5.15 0.455 5.218 0.499 ;
      RECT 4.934 0.223 5.002 0.267 ;
      RECT 4.934 0.455 5.002 0.499 ;
      RECT 4.718 0.223 4.786 0.267 ;
      RECT 4.718 0.4265 4.786 0.4705 ;
      RECT 4.61 0.088 4.678 0.132 ;
      RECT 4.394 0.228 4.462 0.272 ;
      RECT 4.394 0.428 4.462 0.472 ;
      RECT 4.178 0.228 4.246 0.272 ;
      RECT 4.178 0.428 4.246 0.472 ;
      RECT 3.962 0.228 4.03 0.272 ;
      RECT 3.854 0.3985 3.922 0.4425 ;
      RECT 3.856 0.138 3.92 0.182 ;
      RECT 3.638 0.3985 3.706 0.4425 ;
      RECT 3.64 0.138 3.704 0.182 ;
      RECT 3.422 0.158 3.49 0.202 ;
      RECT 3.422 0.3985 3.49 0.4425 ;
      RECT 3.206 0.4895 3.274 0.5335 ;
      RECT 3.098 0.248 3.166 0.292 ;
      RECT 2.882 0.138 2.95 0.182 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.91 0.338 1.978 0.382 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.428 1.762 0.472 ;
      RECT 1.696 0.268 1.76 0.312 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.264 0.268 1.328 0.312 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.338 1.114 0.382 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.83 0.068 0.898 0.112 ;
      RECT 0.832 0.268 0.896 0.312 ;
      RECT 0.506 0.248 0.574 0.292 ;
      RECT 0.29 0.2455 0.358 0.2895 ;
      RECT 0.29 0.4315 0.358 0.4755 ;
      RECT 0.074 0.2455 0.142 0.2895 ;
      RECT 0.074 0.4315 0.142 0.4755 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.358 0.338 0.506 0.382 ;
      RECT 0.506 0.338 0.574 0.472 ;
      RECT 0.574 0.428 1.242 0.472 ;
      RECT 0.722 0.158 0.79 0.292 ;
      RECT 0.79 0.158 0.938 0.202 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.248 1.154 0.292 ;
      RECT 1.154 0.158 1.222 0.292 ;
      RECT 1.222 0.158 1.89 0.202 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 1.998 0.248 2.126 0.292 ;
      RECT 1.114 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 2.194 0.248 2.342 0.292 ;
      RECT 2.342 0.068 2.41 0.292 ;
      RECT 0.898 0.338 1.262 0.382 ;
      RECT 1.262 0.248 1.33 0.382 ;
      RECT 1.33 0.338 1.694 0.382 ;
      RECT 1.694 0.248 1.762 0.382 ;
      RECT 1.762 0.338 2.45 0.382 ;
      RECT 2.45 0.248 2.518 0.382 ;
      RECT 2.518 0.248 2.774 0.292 ;
      RECT 2.774 0.248 2.842 0.382 ;
      RECT 2.842 0.338 3.206 0.382 ;
      RECT 3.206 0.338 3.274 0.562 ;
      RECT 2.95 0.248 3.206 0.292 ;
      RECT 3.206 0.068 3.274 0.292 ;
      RECT 3.274 0.248 3.422 0.292 ;
      RECT 3.422 0.248 3.49 0.472 ;
      RECT 3.274 0.068 3.638 0.112 ;
      RECT 3.638 0.068 3.706 0.202 ;
      RECT 3.706 0.068 3.854 0.112 ;
      RECT 3.854 0.068 3.922 0.202 ;
      RECT 4.61 0.068 4.678 0.472 ;
      RECT 3.53 0.158 3.598 0.292 ;
      RECT 3.598 0.248 3.638 0.292 ;
      RECT 3.638 0.248 3.706 0.472 ;
      RECT 3.706 0.248 3.854 0.292 ;
      RECT 3.854 0.248 3.922 0.562 ;
      RECT 3.922 0.518 4.178 0.562 ;
      RECT 4.178 0.338 4.246 0.562 ;
      RECT 4.246 0.338 4.394 0.382 ;
      RECT 4.394 0.158 4.462 0.382 ;
      RECT 4.246 0.518 4.718 0.562 ;
      RECT 4.718 0.158 4.786 0.562 ;
      RECT 4.786 0.338 4.934 0.382 ;
      RECT 4.934 0.158 5.002 0.562 ;
      RECT 5.218 0.248 5.366 0.292 ;
      RECT 5.366 0.068 5.434 0.562 ;
  END
END b15ru0023as1n08x5

MACRO b15ru0023as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0023as1n12x5 0 0 ;
  SIZE 7.236 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53481475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.53481475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 7.094 0.158 7.162 0.472 ;
      LAYER v0 ;
        RECT 7.094 0.293 7.162 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0306 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5588235 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.97375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.97375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.338 3.274 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.448 3.274 0.492 ;
    END
  END c
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.08568 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.518 4.894 0.562 ;
        RECT 4.826 0.338 4.894 0.562 ;
        RECT 4.61 0.338 4.678 0.562 ;
        RECT 4.394 0.428 4.462 0.562 ;
        RECT 4.178 0.338 4.246 0.562 ;
      LAYER v0 ;
        RECT 4.178 0.363 4.246 0.407 ;
        RECT 4.396 0.448 4.46 0.492 ;
        RECT 4.61 0.363 4.678 0.407 ;
        RECT 4.826 0.363 4.894 0.407 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.582 0.068 5.65 0.292 ;
        RECT 5.15 0.068 5.65 0.112 ;
        RECT 5.366 0.068 5.434 0.202 ;
        RECT 5.15 0.068 5.218 0.472 ;
      LAYER v0 ;
        RECT 5.15 0.2215 5.218 0.2655 ;
        RECT 5.368 0.138 5.432 0.182 ;
        RECT 5.582 0.2215 5.65 0.2655 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 7.27 0.652 ;
        RECT 7.094 0.518 7.162 0.652 ;
        RECT 6.878 0.428 6.946 0.652 ;
        RECT 6.662 0.428 6.73 0.652 ;
        RECT 6.446 0.518 6.514 0.652 ;
        RECT 6.23 0.428 6.298 0.652 ;
        RECT 6.014 0.428 6.082 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 3.098 0.428 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 2.666 0.428 2.734 0.652 ;
        RECT 2.45 0.428 2.518 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 2.45 0.448 2.518 0.492 ;
        RECT 2.666 0.448 2.734 0.492 ;
        RECT 2.882 0.448 2.95 0.492 ;
        RECT 3.098 0.448 3.166 0.492 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 3.746 0.448 3.814 0.492 ;
        RECT 6.014 0.4515 6.082 0.4955 ;
        RECT 6.23 0.4515 6.298 0.4955 ;
        RECT 6.446 0.538 6.514 0.582 ;
        RECT 6.662 0.4515 6.73 0.4955 ;
        RECT 6.878 0.4515 6.946 0.4955 ;
        RECT 7.094 0.538 7.162 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 7.27 0.022 ;
        RECT 7.094 -0.022 7.162 0.112 ;
        RECT 6.878 -0.022 6.946 0.202 ;
        RECT 6.662 -0.022 6.73 0.202 ;
        RECT 6.446 -0.022 6.514 0.112 ;
        RECT 6.23 -0.022 6.298 0.202 ;
        RECT 6.014 -0.022 6.082 0.202 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.53 -0.022 3.598 0.202 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 2.882 -0.022 2.95 0.202 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.45 -0.022 2.518 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.1235 0.358 0.1675 ;
        RECT 0.506 0.138 0.574 0.182 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 2.45 0.138 2.518 0.182 ;
        RECT 2.666 0.138 2.734 0.182 ;
        RECT 2.882 0.138 2.95 0.182 ;
        RECT 3.098 0.138 3.166 0.182 ;
        RECT 3.314 0.138 3.382 0.182 ;
        RECT 3.53 0.138 3.598 0.182 ;
        RECT 3.746 0.138 3.814 0.182 ;
        RECT 6.014 0.138 6.082 0.182 ;
        RECT 6.23 0.138 6.298 0.182 ;
        RECT 6.446 0.048 6.514 0.092 ;
        RECT 6.662 0.138 6.73 0.182 ;
        RECT 6.878 0.138 6.946 0.182 ;
        RECT 7.094 0.048 7.162 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 2.972 0.158 4.928 0.202 ;
      RECT 5.008 0.158 6.64 0.202 ;
    LAYER m1 ;
      RECT 0.506 0.248 0.938 0.292 ;
      RECT 0.918 0.068 1.262 0.112 ;
      RECT 1.566 0.428 2.41 0.472 ;
      RECT 1.046 0.248 1.114 0.382 ;
      RECT 3.422 0.068 3.49 0.292 ;
      RECT 4.826 0.068 4.894 0.202 ;
      RECT 5.042 0.158 5.11 0.292 ;
      RECT 5.366 0.428 5.798 0.472 ;
      RECT 5.258 0.158 5.326 0.292 ;
      RECT 4.05 0.158 4.394 0.202 ;
      RECT 6.554 0.068 6.622 0.562 ;
    LAYER v1 ;
      RECT 6.558 0.158 6.618 0.202 ;
      RECT 5.802 0.158 5.862 0.202 ;
      RECT 5.262 0.158 5.322 0.202 ;
      RECT 5.046 0.158 5.106 0.202 ;
      RECT 4.83 0.158 4.89 0.202 ;
      RECT 2.994 0.158 3.054 0.202 ;
    LAYER v0 ;
      RECT 6.986 0.138 7.054 0.182 ;
      RECT 6.986 0.4515 7.054 0.4955 ;
      RECT 6.77 0.138 6.838 0.182 ;
      RECT 6.77 0.4515 6.838 0.4955 ;
      RECT 6.554 0.138 6.622 0.182 ;
      RECT 6.554 0.4515 6.622 0.4955 ;
      RECT 6.338 0.138 6.406 0.182 ;
      RECT 6.338 0.4515 6.406 0.4955 ;
      RECT 6.122 0.138 6.19 0.182 ;
      RECT 6.122 0.4515 6.19 0.4955 ;
      RECT 5.906 0.248 5.974 0.292 ;
      RECT 5.69 0.2215 5.758 0.2655 ;
      RECT 5.69 0.428 5.758 0.472 ;
      RECT 5.474 0.2215 5.542 0.2655 ;
      RECT 5.474 0.428 5.542 0.472 ;
      RECT 5.258 0.2215 5.326 0.2655 ;
      RECT 5.258 0.428 5.326 0.472 ;
      RECT 5.042 0.2215 5.11 0.2655 ;
      RECT 5.042 0.428 5.11 0.472 ;
      RECT 4.934 0.068 5.002 0.112 ;
      RECT 4.718 0.363 4.786 0.407 ;
      RECT 4.72 0.138 4.784 0.182 ;
      RECT 4.502 0.363 4.57 0.407 ;
      RECT 4.504 0.138 4.568 0.182 ;
      RECT 4.286 0.158 4.354 0.202 ;
      RECT 4.286 0.363 4.354 0.407 ;
      RECT 4.07 0.158 4.138 0.202 ;
      RECT 4.07 0.363 4.138 0.407 ;
      RECT 3.962 0.498 4.03 0.542 ;
      RECT 3.638 0.248 3.706 0.292 ;
      RECT 3.422 0.138 3.49 0.182 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.912 0.268 1.976 0.312 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.48 0.268 1.544 0.312 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.264 0.138 1.328 0.182 ;
      RECT 1.154 0.428 1.222 0.472 ;
      RECT 1.048 0.268 1.112 0.312 ;
      RECT 0.938 0.068 1.006 0.112 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.398 0.228 0.466 0.272 ;
      RECT 0.398 0.4315 0.466 0.4755 ;
      RECT 0.182 0.2135 0.25 0.2575 ;
      RECT 0.182 0.4315 0.25 0.4755 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.338 0.938 0.382 ;
      RECT 0.938 0.338 1.006 0.472 ;
      RECT 1.006 0.428 1.458 0.472 ;
      RECT 0.938 0.158 1.006 0.292 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.158 1.222 0.292 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.158 1.438 0.292 ;
      RECT 1.438 0.158 2.106 0.202 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 2.214 0.248 2.342 0.292 ;
      RECT 1.33 0.068 2.342 0.112 ;
      RECT 2.342 0.068 2.41 0.292 ;
      RECT 2.41 0.248 2.99 0.292 ;
      RECT 2.99 0.068 3.058 0.292 ;
      RECT 1.114 0.338 1.478 0.382 ;
      RECT 1.478 0.248 1.546 0.382 ;
      RECT 1.546 0.338 1.91 0.382 ;
      RECT 1.91 0.248 1.978 0.382 ;
      RECT 1.978 0.338 3.098 0.382 ;
      RECT 3.098 0.248 3.166 0.382 ;
      RECT 3.166 0.248 3.314 0.292 ;
      RECT 3.314 0.248 3.382 0.382 ;
      RECT 3.382 0.338 3.962 0.382 ;
      RECT 3.962 0.338 4.03 0.562 ;
      RECT 3.49 0.248 3.854 0.292 ;
      RECT 3.854 0.068 3.922 0.292 ;
      RECT 3.922 0.248 4.07 0.292 ;
      RECT 4.07 0.248 4.138 0.472 ;
      RECT 4.138 0.248 4.286 0.292 ;
      RECT 4.286 0.248 4.354 0.472 ;
      RECT 3.922 0.068 4.502 0.112 ;
      RECT 4.502 0.068 4.57 0.202 ;
      RECT 4.57 0.068 4.718 0.112 ;
      RECT 4.718 0.068 4.786 0.202 ;
      RECT 4.894 0.068 5.11 0.112 ;
      RECT 5.798 0.158 5.866 0.472 ;
      RECT 5.866 0.248 6.082 0.292 ;
      RECT 4.394 0.158 4.462 0.292 ;
      RECT 4.462 0.248 4.502 0.292 ;
      RECT 4.502 0.248 4.57 0.472 ;
      RECT 4.57 0.248 4.718 0.292 ;
      RECT 4.718 0.248 4.786 0.472 ;
      RECT 4.786 0.248 4.934 0.292 ;
      RECT 4.934 0.248 5.002 0.382 ;
      RECT 5.002 0.338 5.042 0.382 ;
      RECT 5.042 0.338 5.11 0.562 ;
      RECT 5.11 0.518 5.258 0.562 ;
      RECT 5.258 0.338 5.326 0.562 ;
      RECT 5.326 0.338 5.474 0.382 ;
      RECT 5.474 0.158 5.542 0.382 ;
      RECT 5.542 0.338 5.69 0.382 ;
      RECT 5.69 0.158 5.758 0.382 ;
      RECT 5.326 0.518 5.906 0.562 ;
      RECT 5.906 0.338 5.974 0.562 ;
      RECT 5.974 0.338 6.122 0.382 ;
      RECT 6.122 0.068 6.19 0.562 ;
      RECT 6.19 0.338 6.338 0.382 ;
      RECT 6.338 0.068 6.406 0.562 ;
      RECT 6.622 0.338 6.77 0.382 ;
      RECT 6.77 0.068 6.838 0.562 ;
      RECT 6.838 0.338 6.986 0.382 ;
      RECT 6.986 0.068 7.054 0.562 ;
  END
END b15ru0023as1n12x5

MACRO b15ru0023as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15ru0023as1n16x5 0 0 ;
  SIZE 9.072 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.581875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 8.174 0.338 8.998 0.382 ;
        RECT 8.93 0.158 8.998 0.382 ;
      LAYER v0 ;
        RECT 8.39 0.338 8.458 0.382 ;
        RECT 8.606 0.338 8.674 0.382 ;
        RECT 8.822 0.338 8.89 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.58583325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.045 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5624 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.83916675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.83916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.338 4.354 0.562 ;
      LAYER v0 ;
        RECT 4.286 0.448 4.354 0.492 ;
    END
  END c
  PIN carry
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 5.15 0.518 6.298 0.562 ;
        RECT 6.23 0.338 6.298 0.562 ;
        RECT 6.014 0.338 6.082 0.562 ;
        RECT 5.798 0.338 5.866 0.562 ;
        RECT 5.582 0.428 5.65 0.562 ;
        RECT 5.366 0.338 5.434 0.562 ;
        RECT 5.15 0.338 5.218 0.562 ;
      LAYER v0 ;
        RECT 5.15 0.363 5.218 0.407 ;
        RECT 5.366 0.363 5.434 0.407 ;
        RECT 5.584 0.448 5.648 0.492 ;
        RECT 5.798 0.363 5.866 0.407 ;
        RECT 6.014 0.363 6.082 0.407 ;
        RECT 6.23 0.363 6.298 0.407 ;
    END
  END carry
  PIN sum
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 7.31 0.068 7.378 0.292 ;
        RECT 6.446 0.068 7.378 0.112 ;
        RECT 7.094 0.068 7.162 0.292 ;
        RECT 6.878 0.068 6.946 0.202 ;
        RECT 6.662 0.068 6.73 0.472 ;
        RECT 6.446 0.068 6.514 0.472 ;
      LAYER v0 ;
        RECT 6.446 0.2215 6.514 0.2655 ;
        RECT 6.662 0.2215 6.73 0.2655 ;
        RECT 6.88 0.138 6.944 0.182 ;
        RECT 7.094 0.2215 7.162 0.2655 ;
        RECT 7.31 0.2215 7.378 0.2655 ;
    END
  END sum
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 9.106 0.652 ;
        RECT 8.93 0.518 8.998 0.652 ;
        RECT 8.714 0.518 8.782 0.652 ;
        RECT 8.498 0.518 8.566 0.652 ;
        RECT 8.282 0.518 8.35 0.652 ;
        RECT 8.066 0.518 8.134 0.652 ;
        RECT 7.85 0.518 7.918 0.652 ;
        RECT 7.634 0.518 7.702 0.652 ;
        RECT 4.826 0.428 4.894 0.652 ;
        RECT 4.61 0.428 4.678 0.652 ;
        RECT 4.394 0.428 4.462 0.652 ;
        RECT 4.178 0.428 4.246 0.652 ;
        RECT 3.962 0.428 4.03 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.428 3.382 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 3.314 0.448 3.382 0.492 ;
        RECT 3.53 0.448 3.598 0.492 ;
        RECT 3.746 0.448 3.814 0.492 ;
        RECT 3.962 0.448 4.03 0.492 ;
        RECT 4.178 0.448 4.246 0.492 ;
        RECT 4.394 0.448 4.462 0.492 ;
        RECT 4.61 0.448 4.678 0.492 ;
        RECT 4.826 0.448 4.894 0.492 ;
        RECT 7.636 0.538 7.7 0.582 ;
        RECT 7.852 0.538 7.916 0.582 ;
        RECT 8.068 0.538 8.132 0.582 ;
        RECT 8.284 0.538 8.348 0.582 ;
        RECT 8.5 0.538 8.564 0.582 ;
        RECT 8.716 0.538 8.78 0.582 ;
        RECT 8.932 0.538 8.996 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 9.106 0.022 ;
        RECT 8.93 -0.022 8.998 0.112 ;
        RECT 8.714 -0.022 8.782 0.202 ;
        RECT 8.498 -0.022 8.566 0.112 ;
        RECT 8.282 -0.022 8.35 0.202 ;
        RECT 8.066 -0.022 8.134 0.202 ;
        RECT 7.85 -0.022 7.918 0.202 ;
        RECT 7.634 -0.022 7.702 0.202 ;
        RECT 4.826 -0.022 4.894 0.202 ;
        RECT 4.61 -0.022 4.678 0.202 ;
        RECT 4.394 -0.022 4.462 0.202 ;
        RECT 4.178 -0.022 4.246 0.202 ;
        RECT 3.962 -0.022 4.03 0.202 ;
        RECT 3.746 -0.022 3.814 0.202 ;
        RECT 3.53 -0.022 3.598 0.202 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.506 0.1235 0.574 0.1675 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 3.314 0.138 3.382 0.182 ;
        RECT 3.53 0.138 3.598 0.182 ;
        RECT 3.746 0.138 3.814 0.182 ;
        RECT 3.962 0.138 4.03 0.182 ;
        RECT 4.178 0.138 4.246 0.182 ;
        RECT 4.394 0.138 4.462 0.182 ;
        RECT 4.61 0.138 4.678 0.182 ;
        RECT 4.826 0.138 4.894 0.182 ;
        RECT 7.634 0.138 7.702 0.182 ;
        RECT 7.85 0.138 7.918 0.182 ;
        RECT 8.066 0.138 8.134 0.182 ;
        RECT 8.282 0.138 8.35 0.182 ;
        RECT 8.498 0.048 8.566 0.092 ;
        RECT 8.714 0.138 8.782 0.182 ;
        RECT 8.93 0.048 8.998 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 4.052 0.158 6.44 0.202 ;
      RECT 6.52 0.158 8.26 0.202 ;
    LAYER m1 ;
      RECT 0.722 0.248 1.262 0.292 ;
      RECT 1.35 0.068 2.018 0.112 ;
      RECT 2.754 0.428 3.186 0.472 ;
      RECT 1.37 0.248 1.438 0.382 ;
      RECT 4.502 0.068 4.57 0.292 ;
      RECT 6.966 0.428 7.418 0.472 ;
      RECT 6.338 0.068 6.406 0.202 ;
      RECT 6.554 0.158 6.622 0.292 ;
      RECT 6.77 0.158 6.838 0.292 ;
      RECT 5.238 0.158 5.582 0.202 ;
      RECT 8.066 0.248 8.134 0.472 ;
    LAYER v1 ;
      RECT 8.178 0.158 8.238 0.202 ;
      RECT 7.422 0.158 7.482 0.202 ;
      RECT 6.774 0.158 6.834 0.202 ;
      RECT 6.558 0.158 6.618 0.202 ;
      RECT 6.342 0.158 6.402 0.202 ;
      RECT 4.074 0.158 4.134 0.202 ;
    LAYER v0 ;
      RECT 8.822 0.138 8.89 0.182 ;
      RECT 8.822 0.428 8.89 0.472 ;
      RECT 8.606 0.138 8.674 0.182 ;
      RECT 8.606 0.428 8.674 0.472 ;
      RECT 8.39 0.138 8.458 0.182 ;
      RECT 8.39 0.428 8.458 0.472 ;
      RECT 8.174 0.138 8.242 0.182 ;
      RECT 8.174 0.428 8.242 0.472 ;
      RECT 7.958 0.238 8.026 0.282 ;
      RECT 7.958 0.428 8.026 0.472 ;
      RECT 7.742 0.238 7.81 0.282 ;
      RECT 7.742 0.428 7.81 0.472 ;
      RECT 7.526 0.238 7.594 0.282 ;
      RECT 7.526 0.428 7.594 0.472 ;
      RECT 7.418 0.132 7.486 0.176 ;
      RECT 7.202 0.2215 7.27 0.2655 ;
      RECT 7.202 0.428 7.27 0.472 ;
      RECT 6.986 0.2215 7.054 0.2655 ;
      RECT 6.986 0.428 7.054 0.472 ;
      RECT 6.77 0.2215 6.838 0.2655 ;
      RECT 6.77 0.428 6.838 0.472 ;
      RECT 6.554 0.2215 6.622 0.2655 ;
      RECT 6.554 0.428 6.622 0.472 ;
      RECT 6.338 0.088 6.406 0.132 ;
      RECT 6.122 0.363 6.19 0.407 ;
      RECT 6.124 0.138 6.188 0.182 ;
      RECT 5.906 0.363 5.974 0.407 ;
      RECT 5.908 0.138 5.972 0.182 ;
      RECT 5.69 0.363 5.758 0.407 ;
      RECT 5.692 0.138 5.756 0.182 ;
      RECT 5.474 0.158 5.542 0.202 ;
      RECT 5.474 0.363 5.542 0.407 ;
      RECT 5.258 0.158 5.326 0.202 ;
      RECT 5.258 0.363 5.326 0.407 ;
      RECT 5.042 0.498 5.11 0.542 ;
      RECT 4.934 0.248 5.002 0.292 ;
      RECT 4.718 0.248 4.786 0.292 ;
      RECT 4.502 0.138 4.57 0.182 ;
      RECT 3.098 0.1565 3.166 0.2005 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.992 0.268 3.056 0.312 ;
      RECT 2.882 0.158 2.95 0.202 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.776 0.268 2.84 0.312 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.452 0.138 2.516 0.182 ;
      RECT 2.342 0.248 2.41 0.292 ;
      RECT 2.234 0.338 2.302 0.382 ;
      RECT 2.236 0.138 2.3 0.182 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 2.02 0.138 2.084 0.182 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.804 0.268 1.868 0.312 ;
      RECT 1.694 0.068 1.762 0.112 ;
      RECT 1.588 0.268 1.652 0.312 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.37 0.068 1.438 0.112 ;
      RECT 1.372 0.268 1.436 0.312 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.614 0.228 0.682 0.272 ;
      RECT 0.614 0.4315 0.682 0.4755 ;
      RECT 0.398 0.228 0.466 0.272 ;
      RECT 0.398 0.4315 0.466 0.4755 ;
      RECT 0.182 0.228 0.25 0.272 ;
      RECT 0.182 0.4315 0.25 0.4755 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.338 1.262 0.382 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.33 0.428 2.214 0.472 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.33 0.158 1.91 0.202 ;
      RECT 1.91 0.158 1.978 0.292 ;
      RECT 1.978 0.248 2.558 0.292 ;
      RECT 2.558 0.158 2.626 0.292 ;
      RECT 2.626 0.158 3.058 0.202 ;
      RECT 2.018 0.068 2.086 0.202 ;
      RECT 2.086 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.202 ;
      RECT 2.302 0.068 2.45 0.112 ;
      RECT 2.45 0.068 2.518 0.202 ;
      RECT 2.518 0.068 3.098 0.112 ;
      RECT 3.098 0.068 3.166 0.292 ;
      RECT 3.166 0.248 4.07 0.292 ;
      RECT 4.07 0.068 4.138 0.292 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.248 1.654 0.382 ;
      RECT 1.654 0.338 1.802 0.382 ;
      RECT 1.802 0.248 1.87 0.382 ;
      RECT 1.87 0.338 2.774 0.382 ;
      RECT 2.774 0.248 2.842 0.382 ;
      RECT 2.842 0.338 2.99 0.382 ;
      RECT 2.99 0.248 3.058 0.382 ;
      RECT 3.058 0.338 4.178 0.382 ;
      RECT 4.178 0.248 4.246 0.382 ;
      RECT 4.246 0.248 4.394 0.292 ;
      RECT 4.394 0.248 4.462 0.382 ;
      RECT 4.462 0.338 5.042 0.382 ;
      RECT 5.042 0.338 5.11 0.562 ;
      RECT 4.57 0.248 5.042 0.292 ;
      RECT 5.042 0.068 5.11 0.292 ;
      RECT 5.11 0.248 5.258 0.292 ;
      RECT 5.258 0.248 5.326 0.472 ;
      RECT 5.326 0.248 5.474 0.292 ;
      RECT 5.474 0.248 5.542 0.472 ;
      RECT 5.11 0.068 5.69 0.112 ;
      RECT 5.69 0.068 5.758 0.202 ;
      RECT 5.758 0.068 5.906 0.112 ;
      RECT 5.906 0.068 5.974 0.202 ;
      RECT 5.974 0.068 6.122 0.112 ;
      RECT 6.122 0.068 6.19 0.202 ;
      RECT 7.418 0.068 7.486 0.472 ;
      RECT 5.582 0.158 5.65 0.292 ;
      RECT 5.65 0.248 5.69 0.292 ;
      RECT 5.69 0.248 5.758 0.472 ;
      RECT 5.758 0.248 5.906 0.292 ;
      RECT 5.906 0.248 5.974 0.472 ;
      RECT 5.974 0.248 6.122 0.292 ;
      RECT 6.122 0.248 6.19 0.472 ;
      RECT 6.19 0.248 6.338 0.292 ;
      RECT 6.338 0.248 6.406 0.562 ;
      RECT 6.406 0.518 6.554 0.562 ;
      RECT 6.554 0.338 6.622 0.562 ;
      RECT 6.622 0.518 6.77 0.562 ;
      RECT 6.77 0.338 6.838 0.562 ;
      RECT 6.838 0.338 6.986 0.382 ;
      RECT 6.986 0.158 7.054 0.382 ;
      RECT 7.054 0.338 7.202 0.382 ;
      RECT 7.202 0.158 7.27 0.382 ;
      RECT 6.838 0.518 7.526 0.562 ;
      RECT 7.526 0.158 7.594 0.562 ;
      RECT 7.594 0.338 7.742 0.382 ;
      RECT 7.742 0.158 7.81 0.562 ;
      RECT 7.81 0.338 7.958 0.382 ;
      RECT 7.958 0.158 8.026 0.562 ;
      RECT 8.134 0.248 8.174 0.292 ;
      RECT 8.174 0.068 8.242 0.292 ;
      RECT 8.242 0.248 8.39 0.292 ;
      RECT 8.39 0.068 8.458 0.292 ;
      RECT 8.458 0.248 8.606 0.292 ;
      RECT 8.606 0.068 8.674 0.292 ;
      RECT 8.674 0.248 8.822 0.292 ;
      RECT 8.822 0.068 8.89 0.292 ;
      RECT 8.134 0.428 8.998 0.472 ;
  END
END b15ru0023as1n16x5

MACRO b15tdi000as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15tdi000as1n02x5 0 0 ;
  SIZE 0.54 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.248 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.338 0.358 0.382 ;
    END
  END a
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.486 0.112 ;
        RECT 0.182 0.158 0.358 0.202 ;
        RECT 0.29 0.068 0.358 0.202 ;
        RECT 0.182 0.158 0.25 0.382 ;
      LAYER v0 ;
        RECT 0.182 0.248 0.25 0.292 ;
        RECT 0.398 0.068 0.466 0.112 ;
    END
  END en
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.562 ;
      LAYER v0 ;
        RECT 0.4 0.203 0.464 0.247 ;
        RECT 0.398 0.428 0.466 0.472 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.574 0.652 ;
        RECT 0.182 0.428 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.448 0.25 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.574 0.022 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
    LAYER v0 ;
      RECT 0.074 0.448 0.142 0.492 ;
      RECT 0.076 0.158 0.14 0.202 ;
  END
END b15tdi000as1n02x5

MACRO b15tdi000as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15tdi000as1n04x5 0 0 ;
  SIZE 0.756 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 6.8875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.29583325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.158 0.466 0.202 ;
    END
  END en
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.448 0.358 0.492 ;
        RECT 0.29 0.158 0.358 0.202 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 0.79 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.614 0.448 0.682 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 0.79 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END vssx
END b15tdi000as1n04x5

MACRO b15tdi000as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15tdi000as1n08x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 4.87666675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0198 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
        RECT 0.594 0.068 0.79 0.112 ;
      LAYER v0 ;
        RECT 0.614 0.068 0.682 0.112 ;
    END
  END en
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.338 0.79 0.562 ;
        RECT 0.378 0.338 0.79 0.382 ;
      LAYER v0 ;
        RECT 0.398 0.338 0.466 0.382 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.83 0.4705 0.898 0.5145 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.832 0.138 0.896 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.594 0.472 ;
      RECT 0.054 0.158 0.682 0.202 ;
    LAYER v0 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
  END
END b15tdi000as1n08x5

MACRO b15tdi000as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15tdi000as1n16x5 0 0 ;
  SIZE 1.404 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END a
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.035 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.007 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.068 1.222 0.292 ;
        RECT 1.026 0.068 1.222 0.112 ;
      LAYER v0 ;
        RECT 1.046 0.068 1.114 0.112 ;
    END
  END en
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.338 1.222 0.562 ;
        RECT 0.594 0.338 1.222 0.382 ;
      LAYER v0 ;
        RECT 0.614 0.338 0.682 0.382 ;
        RECT 0.83 0.338 0.898 0.382 ;
    END
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.438 0.652 ;
        RECT 1.262 0.428 1.33 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.538 0.466 0.582 ;
        RECT 1.262 0.4705 1.33 0.5145 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.438 0.022 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.398 0.048 0.466 0.092 ;
        RECT 1.262 0.1155 1.33 0.1595 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 1.026 0.472 ;
      RECT 0.054 0.158 1.114 0.202 ;
    LAYER v0 ;
      RECT 0.938 0.158 1.006 0.202 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
  END
END b15tdi000as1n16x5

MACRO b15xnr002as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr002as1n02x3 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.068889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 2.068889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.33 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.383 0.574 0.427 ;
        RECT 0.506 0.203 0.574 0.247 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.938 0.473 1.006 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.398 0.068 0.466 0.472 ;
    LAYER v0 ;
      RECT 1.046 0.3925 1.114 0.4365 ;
      RECT 0.722 0.203 0.79 0.247 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.182 0.203 0.25 0.247 ;
      RECT 0.182 0.383 0.25 0.427 ;
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
      RECT 0.25 0.518 0.614 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 0.898 0.562 ;
      RECT 0.466 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.472 ;
  END
END b15xnr002as1n02x3

MACRO b15xnr002as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr002as1n02x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83901225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 1.83901225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.248 0.898 0.472 ;
      LAYER v0 ;
        RECT 0.83 0.293 0.898 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.383 0.574 0.427 ;
        RECT 0.506 0.203 0.574 0.247 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.938 0.473 1.006 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.938 0.048 1.006 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 0.398 0.068 0.466 0.472 ;
    LAYER v0 ;
      RECT 1.046 0.3925 1.114 0.4365 ;
      RECT 0.722 0.203 0.79 0.247 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.722 0.518 0.79 0.562 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.518 0.614 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 0.898 0.562 ;
      RECT 0.466 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.158 1.046 0.202 ;
      RECT 1.046 0.158 1.114 0.472 ;
  END
END b15xnr002as1n02x5

MACRO b15xnr002as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr002as1n03x5 0 0 ;
  SIZE 1.188 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.47 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.29 0.518 0.682 0.562 ;
        RECT 0.29 0.068 0.358 0.562 ;
      LAYER v0 ;
        RECT 0.29 0.293 0.358 0.337 ;
        RECT 0.506 0.518 0.574 0.562 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.82333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.76 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.293 1.114 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.178 0.574 0.222 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.222 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.338 0.898 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 0.83 0.408 0.898 0.452 ;
        RECT 1.046 0.538 1.114 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.222 0.022 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.2025 0.25 0.2465 ;
        RECT 0.83 0.138 0.898 0.182 ;
        RECT 1.048 0.048 1.112 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.398 0.068 0.466 0.292 ;
    LAYER v0 ;
      RECT 0.938 0.138 1.006 0.182 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.616 0.268 0.68 0.312 ;
      RECT 0.398 0.178 0.466 0.222 ;
      RECT 0.4 0.408 0.464 0.452 ;
      RECT 0.074 0.088 0.142 0.132 ;
      RECT 0.074 0.383 0.142 0.427 ;
    LAYER m1 ;
      RECT 0.398 0.338 0.466 0.472 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.248 0.682 0.382 ;
      RECT 0.506 0.428 0.722 0.472 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.79 0.248 0.938 0.292 ;
      RECT 0.938 0.068 1.006 0.472 ;
  END
END b15xnr002as1n03x5

MACRO b15xnr002as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr002as1n04x5 0 0 ;
  SIZE 1.836 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.21416675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.21416675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.158 1.762 0.472 ;
      LAYER v0 ;
        RECT 1.694 0.3155 1.762 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.428 1.458 0.472 ;
        RECT 0.83 0.338 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.938 0.428 1.006 0.472 ;
        RECT 1.154 0.428 1.222 0.472 ;
        RECT 1.37 0.428 1.438 0.472 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.87 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 1.696 0.538 1.76 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.87 0.022 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.048 0.358 0.092 ;
        RECT 0.506 0.048 0.574 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 1.694 0.048 1.762 0.092 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 1.586 0.158 1.654 0.472 ;
    LAYER v0 ;
      RECT 1.586 0.1955 1.654 0.2395 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.338 1.33 0.382 ;
      RECT 1.046 0.068 1.114 0.112 ;
      RECT 1.048 0.318 1.112 0.362 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.398 0.448 0.466 0.492 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.506 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.382 ;
      RECT 1.114 0.158 1.35 0.202 ;
      RECT 0.25 0.248 0.398 0.292 ;
      RECT 0.398 0.158 0.466 0.562 ;
      RECT 0.466 0.158 0.83 0.202 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 1.242 0.338 1.478 0.382 ;
      RECT 0.898 0.068 1.478 0.112 ;
      RECT 1.478 0.068 1.546 0.382 ;
  END
END b15xnr002as1n04x5

MACRO b15xnr002as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr002as1n06x5 0 0 ;
  SIZE 2.052 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0171 LAYER m1 ;
      ANTENNAMAXAREACAR 4.391111 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0171 LAYER m1 ;
      ANTENNAMAXAREACAR 4.391111 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.408 1.114 0.452 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.49962975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.518 1.438 0.562 ;
        RECT 1.37 0.158 1.438 0.562 ;
        RECT 0.938 0.158 1.006 0.562 ;
        RECT 0.722 0.158 1.006 0.202 ;
        RECT 0.722 0.158 0.79 0.562 ;
      LAYER v0 ;
        RECT 0.722 0.408 0.79 0.452 ;
        RECT 0.722 0.268 0.79 0.312 ;
        RECT 0.938 0.408 1.006 0.452 ;
        RECT 0.938 0.268 1.006 0.312 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.37 0.2185 1.438 0.2625 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.086 0.652 ;
        RECT 1.91 0.518 1.978 0.652 ;
        RECT 1.694 0.518 1.762 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 1.696 0.538 1.76 0.582 ;
        RECT 1.912 0.538 1.976 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.086 0.022 ;
        RECT 1.91 -0.022 1.978 0.112 ;
        RECT 1.694 -0.022 1.762 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 1.696 0.048 1.76 0.092 ;
        RECT 1.912 0.048 1.976 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.518 1.672 0.562 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.83 0.248 0.898 0.562 ;
      RECT 1.262 0.068 1.33 0.472 ;
      RECT 1.586 0.338 1.654 0.562 ;
    LAYER v1 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.294 0.518 0.354 0.562 ;
      RECT 0.078 0.518 0.138 0.562 ;
    LAYER v0 ;
      RECT 1.802 0.158 1.87 0.202 ;
      RECT 1.802 0.428 1.87 0.472 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.478 0.408 1.546 0.452 ;
      RECT 1.48 0.138 1.544 0.182 ;
      RECT 1.262 0.2185 1.33 0.2625 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.154 0.408 1.222 0.452 ;
      RECT 0.83 0.268 0.898 0.312 ;
      RECT 0.83 0.408 0.898 0.452 ;
      RECT 0.614 0.068 0.682 0.112 ;
      RECT 0.506 0.1695 0.574 0.2135 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.574 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.472 ;
      RECT 1.33 0.068 1.478 0.112 ;
      RECT 1.478 0.068 1.546 0.472 ;
      RECT 1.546 0.248 1.802 0.292 ;
      RECT 1.802 0.068 1.87 0.562 ;
  END
END b15xnr002as1n06x5

MACRO b15xnr002as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr002as1n08x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 3.51587975 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 3.51587975 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.408 1.222 0.452 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.2705 0.142 0.3145 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.518 1.546 0.562 ;
        RECT 1.478 0.158 1.546 0.562 ;
        RECT 1.046 0.158 1.114 0.562 ;
        RECT 0.83 0.158 1.114 0.202 ;
        RECT 0.83 0.158 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.408 0.898 0.452 ;
        RECT 0.83 0.268 0.898 0.312 ;
        RECT 1.046 0.408 1.114 0.452 ;
        RECT 1.046 0.268 1.114 0.312 ;
        RECT 1.478 0.408 1.546 0.452 ;
        RECT 1.478 0.2185 1.546 0.2625 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.018 0.518 2.086 0.652 ;
        RECT 1.802 0.518 1.87 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
        RECT 1.804 0.538 1.868 0.582 ;
        RECT 2.02 0.538 2.084 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.018 -0.022 2.086 0.112 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
        RECT 2.02 0.048 2.084 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.518 1.78 0.562 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 0.938 0.248 1.006 0.562 ;
      RECT 1.37 0.068 1.438 0.472 ;
      RECT 1.694 0.338 1.762 0.562 ;
    LAYER v1 ;
      RECT 1.698 0.518 1.758 0.562 ;
      RECT 0.942 0.518 1.002 0.562 ;
      RECT 0.402 0.518 0.462 0.562 ;
      RECT 0.186 0.518 0.246 0.562 ;
    LAYER v0 ;
      RECT 2.126 0.158 2.194 0.202 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.91 0.428 1.978 0.472 ;
      RECT 1.694 0.408 1.762 0.452 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.588 0.138 1.652 0.182 ;
      RECT 1.37 0.2185 1.438 0.2625 ;
      RECT 1.37 0.408 1.438 0.452 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 0.938 0.268 1.006 0.312 ;
      RECT 0.938 0.408 1.006 0.452 ;
      RECT 0.722 0.068 0.79 0.112 ;
      RECT 0.614 0.1695 0.682 0.2135 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.562 ;
      RECT 0.682 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.472 ;
      RECT 1.438 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.654 0.248 1.91 0.292 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 1.978 0.248 2.126 0.292 ;
      RECT 2.126 0.068 2.194 0.562 ;
  END
END b15xnr002as1n08x5

MACRO b15xnr002as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr002as1n12x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0333 LAYER m1 ;
      ANTENNAMAXAREACAR 2.6246245 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0333 LAYER m1 ;
      ANTENNAMAXAREACAR 2.6246245 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.158 1.546 0.472 ;
      LAYER v0 ;
        RECT 1.478 0.408 1.546 0.452 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.068 1.978 0.472 ;
        RECT 1.694 0.068 1.978 0.112 ;
        RECT 1.37 0.518 1.762 0.562 ;
        RECT 1.694 0.068 1.762 0.562 ;
        RECT 1.37 0.158 1.438 0.562 ;
        RECT 1.154 0.158 1.438 0.202 ;
        RECT 1.154 0.158 1.222 0.562 ;
      LAYER v0 ;
        RECT 1.154 0.408 1.222 0.452 ;
        RECT 1.154 0.268 1.222 0.312 ;
        RECT 1.37 0.408 1.438 0.452 ;
        RECT 1.37 0.268 1.438 0.312 ;
        RECT 1.694 0.408 1.762 0.452 ;
        RECT 1.694 0.203 1.762 0.247 ;
        RECT 1.91 0.408 1.978 0.452 ;
        RECT 1.91 0.203 1.978 0.247 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 2.45 0.338 2.518 0.652 ;
        RECT 2.234 0.338 2.302 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.614 0.338 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.614 0.428 0.682 0.472 ;
        RECT 0.83 0.518 0.898 0.562 ;
        RECT 2.234 0.408 2.302 0.452 ;
        RECT 2.45 0.408 2.518 0.452 ;
        RECT 2.666 0.408 2.734 0.452 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.666 -0.022 2.734 0.202 ;
        RECT 2.45 -0.022 2.518 0.112 ;
        RECT 2.234 -0.022 2.302 0.112 ;
        RECT 0.83 -0.022 0.898 0.202 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.614 0.178 0.682 0.222 ;
        RECT 0.83 0.074 0.898 0.118 ;
        RECT 2.236 0.048 2.3 0.092 ;
        RECT 2.452 0.048 2.516 0.092 ;
        RECT 2.666 0.138 2.734 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.272 0.518 2.32 0.562 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.562 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.802 0.158 1.87 0.562 ;
      RECT 2.126 0.338 2.194 0.562 ;
    LAYER v1 ;
      RECT 2.13 0.518 2.19 0.562 ;
      RECT 1.266 0.518 1.326 0.562 ;
      RECT 1.05 0.518 1.11 0.562 ;
      RECT 0.51 0.518 0.57 0.562 ;
      RECT 0.294 0.518 0.354 0.562 ;
    LAYER v0 ;
      RECT 2.558 0.138 2.626 0.182 ;
      RECT 2.558 0.408 2.626 0.452 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.342 0.408 2.41 0.452 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 2.018 0.408 2.086 0.452 ;
      RECT 1.802 0.203 1.87 0.247 ;
      RECT 1.802 0.408 1.87 0.452 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.262 0.268 1.33 0.312 ;
      RECT 1.262 0.408 1.33 0.452 ;
      RECT 1.046 0.268 1.114 0.312 ;
      RECT 1.046 0.408 1.114 0.452 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.562 ;
      RECT 0.142 0.248 0.29 0.292 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.79 0.338 0.938 0.382 ;
      RECT 0.938 0.068 1.006 0.382 ;
      RECT 1.006 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.87 0.518 2.018 0.562 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 2.086 0.248 2.342 0.292 ;
      RECT 2.342 0.068 2.41 0.562 ;
      RECT 2.41 0.248 2.558 0.292 ;
      RECT 2.558 0.068 2.626 0.562 ;
  END
END b15xnr002as1n12x5

MACRO b15xnr002as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr002as1n16x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 2.21314825 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 2.21314825 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.802 0.408 1.87 0.452 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0585 LAYER m1 ;
      ANTENNAMAXAREACAR 0.465094 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.293 0.466 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14688 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.694 0.518 2.518 0.562 ;
        RECT 2.45 0.158 2.518 0.562 ;
        RECT 2.234 0.158 2.302 0.562 ;
        RECT 2.018 0.068 2.086 0.562 ;
        RECT 1.694 0.158 1.762 0.562 ;
        RECT 1.262 0.158 1.762 0.202 ;
        RECT 1.478 0.158 1.546 0.472 ;
        RECT 1.262 0.158 1.33 0.472 ;
      LAYER v0 ;
        RECT 1.262 0.408 1.33 0.452 ;
        RECT 1.262 0.268 1.33 0.312 ;
        RECT 1.478 0.408 1.546 0.452 ;
        RECT 1.478 0.268 1.546 0.312 ;
        RECT 1.694 0.408 1.762 0.452 ;
        RECT 1.694 0.268 1.762 0.312 ;
        RECT 2.018 0.408 2.086 0.452 ;
        RECT 2.018 0.203 2.086 0.247 ;
        RECT 2.234 0.408 2.302 0.452 ;
        RECT 2.234 0.203 2.302 0.247 ;
        RECT 2.45 0.408 2.518 0.452 ;
        RECT 2.45 0.203 2.518 0.247 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.518 2.95 0.652 ;
        RECT 2.666 0.518 2.734 0.652 ;
        RECT 1.046 0.518 1.114 0.652 ;
        RECT 0.83 0.518 0.898 0.652 ;
        RECT 0.614 0.518 0.682 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.616 0.538 0.68 0.582 ;
        RECT 0.832 0.538 0.896 0.582 ;
        RECT 1.048 0.538 1.112 0.582 ;
        RECT 2.668 0.538 2.732 0.582 ;
        RECT 2.884 0.538 2.948 0.582 ;
        RECT 3.1 0.538 3.164 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.666 -0.022 2.734 0.112 ;
        RECT 1.046 -0.022 1.114 0.112 ;
        RECT 0.83 -0.022 0.898 0.112 ;
        RECT 0.614 -0.022 0.682 0.112 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.616 0.048 0.68 0.092 ;
        RECT 0.832 0.048 0.896 0.092 ;
        RECT 1.048 0.048 1.112 0.092 ;
        RECT 2.668 0.048 2.732 0.092 ;
        RECT 2.884 0.048 2.948 0.092 ;
        RECT 3.1 0.048 3.164 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.518 2.644 0.562 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.29 0.158 0.358 0.562 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.722 0.158 0.79 0.562 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.586 0.248 1.654 0.562 ;
      RECT 2.126 0.068 2.194 0.472 ;
      RECT 2.558 0.338 2.626 0.562 ;
    LAYER v1 ;
      RECT 2.562 0.518 2.622 0.562 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.374 0.518 1.434 0.562 ;
      RECT 0.726 0.518 0.786 0.562 ;
      RECT 0.51 0.518 0.57 0.562 ;
      RECT 0.294 0.518 0.354 0.562 ;
      RECT 0.078 0.518 0.138 0.562 ;
    LAYER v0 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.206 0.408 3.274 0.452 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.99 0.408 3.058 0.452 ;
      RECT 2.774 0.158 2.842 0.202 ;
      RECT 2.774 0.408 2.842 0.452 ;
      RECT 2.558 0.408 2.626 0.452 ;
      RECT 2.342 0.203 2.41 0.247 ;
      RECT 2.342 0.408 2.41 0.452 ;
      RECT 2.126 0.203 2.194 0.247 ;
      RECT 2.126 0.408 2.194 0.452 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.586 0.268 1.654 0.312 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.37 0.268 1.438 0.312 ;
      RECT 1.37 0.408 1.438 0.452 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.938 0.428 1.006 0.472 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.428 0.79 0.472 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.178 0.358 0.222 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.178 0.142 0.222 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.006 0.338 1.154 0.382 ;
      RECT 1.154 0.068 1.222 0.382 ;
      RECT 1.222 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.472 ;
      RECT 2.194 0.068 2.342 0.112 ;
      RECT 2.342 0.068 2.41 0.472 ;
      RECT 2.41 0.068 2.558 0.112 ;
      RECT 2.558 0.068 2.626 0.292 ;
      RECT 2.626 0.248 2.774 0.292 ;
      RECT 2.774 0.068 2.842 0.472 ;
      RECT 2.842 0.248 2.99 0.292 ;
      RECT 2.99 0.068 3.058 0.472 ;
      RECT 3.058 0.248 3.206 0.292 ;
      RECT 3.206 0.068 3.274 0.472 ;
  END
END b15xnr002as1n16x5

MACRO b15xnr003as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr003as1n02x3 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 5.7475 LAYER m1 ;
      ANTENNAMAXAREACAR 11.678611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 5.7475 LAYER m1 ;
      ANTENNAMAXAREACAR 11.678611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.046 0.158 1.114 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER m2 ;
        RECT 0.272 0.248 1.672 0.292 ;
      LAYER v1 ;
        RECT 0.294 0.248 0.354 0.292 ;
        RECT 1.05 0.248 1.11 0.292 ;
        RECT 1.59 0.248 1.65 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.178 0.358 0.222 ;
        RECT 1.046 0.293 1.114 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 1.85777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.158 2.626 0.472 ;
      LAYER v0 ;
        RECT 2.558 0.338 2.626 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.158 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 1.91 0.178 1.978 0.222 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 2.342 0.538 2.41 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.342 -0.022 2.41 0.382 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 1.37 0.178 1.438 0.222 ;
        RECT 2.342 0.178 2.41 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 1.78 0.382 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 1.694 0.518 2.018 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 2.45 0.068 2.518 0.562 ;
    LAYER v1 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 2.45 0.178 2.518 0.222 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.178 2.302 0.222 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.178 2.086 0.222 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.398 0.178 0.466 0.222 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.518 0.398 0.562 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.006 0.518 1.154 0.562 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.006 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.562 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 1.87 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.562 ;
  END
END b15xnr003as1n02x3

MACRO b15xnr003as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr003as1n02x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 5.7475 LAYER m1 ;
      ANTENNAMAXAREACAR 11.678611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 5.7475 LAYER m1 ;
      ANTENNAMAXAREACAR 11.678611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.046 0.158 1.114 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER m2 ;
        RECT 0.272 0.248 1.672 0.292 ;
      LAYER v1 ;
        RECT 0.294 0.248 0.354 0.292 ;
        RECT 1.05 0.248 1.11 0.292 ;
        RECT 1.59 0.248 1.65 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.178 0.358 0.222 ;
        RECT 1.046 0.293 1.114 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.825679 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 0.825679 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.158 2.626 0.472 ;
      LAYER v0 ;
        RECT 2.558 0.338 2.626 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.158 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 1.91 0.178 1.978 0.222 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 2.342 0.538 2.41 0.582 ;
        RECT 2.558 0.538 2.626 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.382 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 1.37 0.178 1.438 0.222 ;
        RECT 2.342 0.178 2.41 0.222 ;
        RECT 2.56 0.048 2.624 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 1.78 0.382 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 1.694 0.518 2.018 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 2.45 0.068 2.518 0.562 ;
    LAYER v1 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 2.45 0.178 2.518 0.222 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.178 2.302 0.222 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.178 2.086 0.222 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.398 0.178 0.466 0.222 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.518 0.398 0.562 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.006 0.518 1.154 0.562 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.006 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.562 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 1.87 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.562 ;
  END
END b15xnr003as1n02x5

MACRO b15xnr003as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr003as1n03x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0117 LAYER m2 ;
      ANTENNAMAXAREACAR 5.7475 LAYER m1 ;
      ANTENNAMAXAREACAR 11.678611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0117 LAYER m2 ;
      ANTENNAMAXAREACAR 5.7475 LAYER m1 ;
      ANTENNAMAXAREACAR 11.678611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.158 1.654 0.472 ;
        RECT 1.046 0.158 1.114 0.472 ;
        RECT 0.29 0.158 0.358 0.472 ;
      LAYER m2 ;
        RECT 0.272 0.248 1.672 0.292 ;
      LAYER v1 ;
        RECT 0.294 0.248 0.354 0.292 ;
        RECT 1.05 0.248 1.11 0.292 ;
        RECT 1.59 0.248 1.65 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.178 0.358 0.222 ;
        RECT 1.046 0.293 1.114 0.337 ;
        RECT 1.586 0.293 1.654 0.337 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.158 2.626 0.472 ;
      LAYER v0 ;
        RECT 2.558 0.338 2.626 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.158 1.978 0.472 ;
      LAYER v0 ;
        RECT 1.91 0.383 1.978 0.427 ;
        RECT 1.91 0.178 1.978 0.222 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 1.37 0.428 1.438 0.472 ;
        RECT 2.344 0.538 2.408 0.582 ;
        RECT 2.56 0.538 2.624 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.382 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 1.37 0.178 1.438 0.222 ;
        RECT 2.342 0.178 2.41 0.222 ;
        RECT 2.56 0.048 2.624 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 1.78 0.382 ;
    LAYER m1 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.506 0.158 0.574 0.472 ;
      RECT 0.83 0.158 0.898 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 1.694 0.518 2.018 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 2.45 0.068 2.518 0.562 ;
    LAYER v1 ;
      RECT 1.698 0.338 1.758 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 2.45 0.178 2.518 0.222 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.234 0.178 2.302 0.222 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.178 2.086 0.222 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.694 0.293 1.762 0.337 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.478 0.428 1.546 0.472 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.154 0.293 1.222 0.337 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.398 0.178 0.466 0.222 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.518 0.398 0.562 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.338 1.006 0.562 ;
      RECT 1.006 0.518 1.154 0.562 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.79 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.006 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.562 ;
      RECT 2.018 0.158 2.086 0.562 ;
      RECT 1.87 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.562 ;
  END
END b15xnr003as1n03x5

MACRO b15xnr003as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr003as1n04x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 3.1075 LAYER m1 ;
      ANTENNAMAXAREACAR 9.978611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 3.1075 LAYER m1 ;
      ANTENNAMAXAREACAR 9.978611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 1.046 0.338 1.33 0.382 ;
        RECT 1.046 0.158 1.114 0.382 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER m2 ;
        RECT 0.38 0.248 1.904 0.292 ;
      LAYER v1 ;
        RECT 0.402 0.248 0.462 0.292 ;
        RECT 1.05 0.248 1.11 0.292 ;
        RECT 1.806 0.248 1.866 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.178 0.466 0.222 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.802 0.3155 1.87 0.3595 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 1.117647 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 1.117647 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.068 3.274 0.562 ;
      LAYER v0 ;
        RECT 3.206 0.3155 3.274 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.158 2.41 0.472 ;
      LAYER v0 ;
        RECT 2.342 0.383 2.41 0.427 ;
        RECT 2.342 0.178 2.41 0.222 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.098 0.338 3.166 0.652 ;
        RECT 2.882 0.338 2.95 0.652 ;
        RECT 2.666 0.338 2.734 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 2.666 0.428 2.734 0.472 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 3.098 0.428 3.166 0.472 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.098 -0.022 3.166 0.292 ;
        RECT 2.882 -0.022 2.95 0.292 ;
        RECT 2.666 -0.022 2.734 0.292 ;
        RECT 1.694 -0.022 1.762 0.292 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 2.666 0.178 2.734 0.222 ;
        RECT 2.882 0.178 2.95 0.222 ;
        RECT 3.098 0.178 3.166 0.222 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.596 0.338 2.104 0.382 ;
      RECT 1.984 0.248 2.86 0.292 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 2.018 0.518 2.558 0.562 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.018 0.158 2.086 0.472 ;
      RECT 2.126 0.158 2.194 0.382 ;
      RECT 2.45 0.158 2.518 0.472 ;
      RECT 2.774 0.158 2.842 0.562 ;
      RECT 2.99 0.158 3.058 0.562 ;
      RECT 3.314 0.158 3.382 0.562 ;
    LAYER v1 ;
      RECT 2.778 0.248 2.838 0.292 ;
      RECT 2.454 0.248 2.514 0.292 ;
      RECT 2.13 0.248 2.19 0.292 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 0.618 0.338 0.678 0.382 ;
    LAYER v0 ;
      RECT 3.314 0.178 3.382 0.222 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 2.99 0.178 3.058 0.222 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.774 0.178 2.842 0.222 ;
      RECT 2.774 0.428 2.842 0.472 ;
      RECT 2.558 0.178 2.626 0.222 ;
      RECT 2.45 0.383 2.518 0.427 ;
      RECT 2.126 0.178 2.194 0.222 ;
      RECT 2.126 0.518 2.194 0.562 ;
      RECT 2.018 0.338 2.086 0.382 ;
      RECT 1.91 0.1355 1.978 0.1795 ;
      RECT 1.91 0.4505 1.978 0.4945 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.398 0.4275 0.466 0.4715 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.4275 0.25 0.4715 ;
    LAYER m1 ;
      RECT 1.046 0.158 1.114 0.382 ;
      RECT 1.114 0.338 1.33 0.382 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.722 0.562 ;
      RECT 0.722 0.158 0.79 0.562 ;
      RECT 0.79 0.518 1.37 0.562 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 0.574 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 0.898 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.248 1.586 0.292 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 2.558 0.158 2.626 0.562 ;
  END
END b15xnr003as1n04x5

MACRO b15xnr003as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr003as1n06x5 0 0 ;
  SIZE 3.888 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 3.1075 LAYER m1 ;
      ANTENNAMAXAREACAR 9.978611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAGATEAREA 0.0108 LAYER m2 ;
      ANTENNAMAXAREACAR 3.1075 LAYER m1 ;
      ANTENNAMAXAREACAR 9.978611 LAYER m2 ;
      ANTENNAMAXCUTCAR 1.5644445 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.472 ;
        RECT 1.046 0.338 1.33 0.382 ;
        RECT 1.046 0.158 1.114 0.382 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER m2 ;
        RECT 0.38 0.248 1.904 0.292 ;
      LAYER v1 ;
        RECT 0.402 0.248 0.462 0.292 ;
        RECT 1.05 0.248 1.11 0.292 ;
        RECT 1.806 0.248 1.866 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.178 0.466 0.222 ;
        RECT 1.154 0.338 1.222 0.382 ;
        RECT 1.802 0.3155 1.87 0.3595 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.9424 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0225 LAYER m1 ;
      ANTENNAMAXAREACAR 0.9424 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.53 0.068 3.598 0.562 ;
      LAYER v0 ;
        RECT 3.53 0.3155 3.598 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.03672 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.666 0.068 2.734 0.472 ;
        RECT 2.234 0.068 2.734 0.112 ;
        RECT 2.234 0.068 2.302 0.382 ;
      LAYER v0 ;
        RECT 2.234 0.248 2.302 0.292 ;
        RECT 2.666 0.248 2.734 0.292 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.922 0.652 ;
        RECT 3.746 0.338 3.814 0.652 ;
        RECT 3.422 0.338 3.49 0.652 ;
        RECT 3.206 0.338 3.274 0.652 ;
        RECT 2.99 0.338 3.058 0.652 ;
        RECT 1.694 0.338 1.762 0.652 ;
        RECT 1.478 0.338 1.546 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.538 0.358 0.582 ;
        RECT 1.478 0.428 1.546 0.472 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 2.99 0.4225 3.058 0.4665 ;
        RECT 3.206 0.4225 3.274 0.4665 ;
        RECT 3.422 0.4225 3.49 0.4665 ;
        RECT 3.746 0.4225 3.814 0.4665 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.922 0.022 ;
        RECT 3.746 -0.022 3.814 0.292 ;
        RECT 3.422 -0.022 3.49 0.292 ;
        RECT 3.206 -0.022 3.274 0.292 ;
        RECT 2.99 -0.022 3.058 0.292 ;
        RECT 1.694 -0.022 1.762 0.292 ;
        RECT 1.262 0.158 1.546 0.202 ;
        RECT 1.262 -0.022 1.33 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 1.694 0.158 1.762 0.202 ;
        RECT 2.99 0.1725 3.058 0.2165 ;
        RECT 3.206 0.1725 3.274 0.2165 ;
        RECT 3.422 0.1725 3.49 0.2165 ;
        RECT 3.746 0.1725 3.814 0.2165 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.596 0.338 2.104 0.382 ;
      RECT 1.984 0.248 3.184 0.292 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.292 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 2.018 0.428 2.558 0.472 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 1.91 0.068 1.978 0.562 ;
      RECT 2.018 0.158 2.086 0.382 ;
      RECT 2.126 0.158 2.194 0.382 ;
      RECT 2.342 0.158 2.41 0.382 ;
      RECT 2.774 0.068 2.842 0.472 ;
      RECT 3.098 0.068 3.166 0.562 ;
      RECT 3.314 0.068 3.382 0.562 ;
      RECT 3.638 0.068 3.706 0.562 ;
    LAYER v1 ;
      RECT 3.102 0.248 3.162 0.292 ;
      RECT 2.778 0.248 2.838 0.292 ;
      RECT 2.346 0.248 2.406 0.292 ;
      RECT 2.13 0.248 2.19 0.292 ;
      RECT 2.022 0.338 2.082 0.382 ;
      RECT 0.618 0.338 0.678 0.382 ;
    LAYER v0 ;
      RECT 3.638 0.1725 3.706 0.2165 ;
      RECT 3.638 0.4225 3.706 0.4665 ;
      RECT 3.314 0.1725 3.382 0.2165 ;
      RECT 3.314 0.4225 3.382 0.4665 ;
      RECT 3.098 0.1725 3.166 0.2165 ;
      RECT 3.098 0.4225 3.166 0.4665 ;
      RECT 2.882 0.1725 2.95 0.2165 ;
      RECT 2.774 0.3775 2.842 0.4215 ;
      RECT 2.558 0.248 2.626 0.292 ;
      RECT 2.342 0.248 2.41 0.292 ;
      RECT 2.342 0.428 2.41 0.472 ;
      RECT 2.126 0.248 2.194 0.292 ;
      RECT 2.126 0.428 2.194 0.472 ;
      RECT 2.018 0.248 2.086 0.292 ;
      RECT 1.91 0.1355 1.978 0.1795 ;
      RECT 1.91 0.4505 1.978 0.4945 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.154 0.178 1.222 0.222 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.398 0.4275 0.466 0.4715 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.4275 0.25 0.4715 ;
    LAYER m1 ;
      RECT 1.046 0.158 1.114 0.382 ;
      RECT 1.114 0.338 1.33 0.382 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.722 0.562 ;
      RECT 0.722 0.158 0.79 0.562 ;
      RECT 0.79 0.518 1.37 0.562 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 0.574 0.068 0.83 0.112 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 0.898 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.292 ;
      RECT 1.222 0.248 1.586 0.292 ;
      RECT 1.586 0.068 1.654 0.562 ;
      RECT 2.558 0.158 2.626 0.562 ;
      RECT 2.626 0.518 2.882 0.562 ;
      RECT 2.882 0.068 2.95 0.562 ;
  END
END b15xnr003as1n06x5

MACRO b15xnr003as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr003as1n08x5 0 0 ;
  SIZE 5.292 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0216 LAYER m2 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
      ANTENNAMAXAREACAR 4.4644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0216 LAYER m2 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
      ANTENNAMAXAREACAR 4.4644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.158 2.95 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
      LAYER m2 ;
        RECT 1.136 0.248 2.984 0.292 ;
      LAYER v1 ;
        RECT 1.158 0.248 1.218 0.292 ;
        RECT 2.886 0.248 2.946 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.383 1.222 0.427 ;
        RECT 2.882 0.338 2.95 0.382 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.990303 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0297 LAYER m1 ;
      ANTENNAMAXAREACAR 0.990303 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.718 0.158 4.786 0.472 ;
      LAYER v0 ;
        RECT 4.718 0.3155 4.786 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.04896 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.638 0.068 3.706 0.382 ;
        RECT 3.206 0.068 3.706 0.112 ;
        RECT 3.098 0.428 3.49 0.472 ;
        RECT 3.422 0.068 3.49 0.472 ;
        RECT 3.206 0.068 3.274 0.382 ;
      LAYER v0 ;
        RECT 3.206 0.428 3.274 0.472 ;
        RECT 3.206 0.248 3.274 0.292 ;
        RECT 3.638 0.248 3.706 0.292 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.326 0.652 ;
        RECT 5.15 0.338 5.218 0.652 ;
        RECT 4.934 0.338 5.002 0.652 ;
        RECT 4.61 0.338 4.678 0.652 ;
        RECT 4.394 0.338 4.462 0.652 ;
        RECT 4.178 0.338 4.246 0.652 ;
        RECT 3.962 0.338 4.03 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.558 0.428 2.626 0.472 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 3.962 0.4225 4.03 0.4665 ;
        RECT 4.178 0.4225 4.246 0.4665 ;
        RECT 4.394 0.4225 4.462 0.4665 ;
        RECT 4.61 0.4225 4.678 0.4665 ;
        RECT 4.934 0.4225 5.002 0.4665 ;
        RECT 5.15 0.4225 5.218 0.4665 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.326 0.022 ;
        RECT 5.15 -0.022 5.218 0.292 ;
        RECT 4.934 -0.022 5.002 0.292 ;
        RECT 4.61 -0.022 4.678 0.292 ;
        RECT 4.394 -0.022 4.462 0.292 ;
        RECT 4.178 -0.022 4.246 0.292 ;
        RECT 3.962 -0.022 4.03 0.292 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.558 -0.022 2.626 0.292 ;
        RECT 2.126 0.158 2.41 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.558 0.158 2.626 0.202 ;
        RECT 2.774 0.158 2.842 0.202 ;
        RECT 3.962 0.1725 4.03 0.2165 ;
        RECT 4.178 0.1725 4.246 0.2165 ;
        RECT 4.394 0.1725 4.462 0.2165 ;
        RECT 4.61 0.1725 4.678 0.2165 ;
        RECT 4.934 0.1725 5.002 0.2165 ;
        RECT 5.15 0.1725 5.218 0.2165 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 3.076 0.382 ;
      RECT 3.064 0.248 4.372 0.292 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.472 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.262 0.158 1.33 0.472 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 2.99 0.518 3.53 0.562 ;
      RECT 2.666 0.068 2.734 0.562 ;
      RECT 2.882 0.158 2.95 0.472 ;
      RECT 2.99 0.158 3.058 0.472 ;
      RECT 3.098 0.158 3.166 0.382 ;
      RECT 3.314 0.158 3.382 0.382 ;
      RECT 3.746 0.068 3.814 0.472 ;
      RECT 4.07 0.068 4.138 0.562 ;
      RECT 4.286 0.068 4.354 0.562 ;
      RECT 4.502 0.068 4.57 0.562 ;
      RECT 4.826 0.068 4.894 0.562 ;
      RECT 5.042 0.068 5.11 0.562 ;
    LAYER v1 ;
      RECT 4.29 0.248 4.35 0.292 ;
      RECT 4.074 0.248 4.134 0.292 ;
      RECT 3.75 0.248 3.81 0.292 ;
      RECT 3.318 0.248 3.378 0.292 ;
      RECT 3.102 0.248 3.162 0.292 ;
      RECT 2.994 0.338 3.054 0.382 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 5.042 0.1725 5.11 0.2165 ;
      RECT 5.042 0.4225 5.11 0.4665 ;
      RECT 4.826 0.1725 4.894 0.2165 ;
      RECT 4.826 0.4225 4.894 0.4665 ;
      RECT 4.502 0.1725 4.57 0.2165 ;
      RECT 4.502 0.4225 4.57 0.4665 ;
      RECT 4.286 0.1725 4.354 0.2165 ;
      RECT 4.286 0.4225 4.354 0.4665 ;
      RECT 4.07 0.1725 4.138 0.2165 ;
      RECT 4.07 0.4225 4.138 0.4665 ;
      RECT 3.854 0.1725 3.922 0.2165 ;
      RECT 3.746 0.3775 3.814 0.4215 ;
      RECT 3.53 0.248 3.598 0.292 ;
      RECT 3.314 0.248 3.382 0.292 ;
      RECT 3.314 0.518 3.382 0.562 ;
      RECT 3.098 0.248 3.166 0.292 ;
      RECT 3.098 0.518 3.166 0.562 ;
      RECT 2.99 0.248 3.058 0.292 ;
      RECT 2.666 0.158 2.734 0.202 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.45 0.158 2.518 0.202 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.383 1.87 0.427 ;
      RECT 1.694 0.178 1.762 0.222 ;
      RECT 1.586 0.383 1.654 0.427 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 1.37 0.178 1.438 0.222 ;
      RECT 1.37 0.383 1.438 0.427 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.262 0.383 1.33 0.427 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 1.046 0.383 1.114 0.427 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.4275 0.25 0.4715 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.158 0.898 0.562 ;
      RECT 0.898 0.518 1.37 0.562 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.518 1.694 0.562 ;
      RECT 1.694 0.158 1.762 0.562 ;
      RECT 1.762 0.518 2.018 0.562 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.086 0.338 2.302 0.382 ;
      RECT 0.682 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.472 ;
      RECT 1.006 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.438 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.654 0.068 2.018 0.112 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 2.086 0.248 2.45 0.292 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 3.53 0.158 3.598 0.562 ;
      RECT 3.598 0.518 3.854 0.562 ;
      RECT 3.854 0.068 3.922 0.562 ;
  END
END b15xnr003as1n08x5

MACRO b15xnr003as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr003as1n12x5 0 0 ;
  SIZE 5.508 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0216 LAYER m2 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
      ANTENNAMAXAREACAR 4.4644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAGATEAREA 0.0216 LAYER m2 ;
      ANTENNAMAXAREACAR 1.498889 LAYER m1 ;
      ANTENNAMAXAREACAR 4.4644445 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.78222225 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 2.882 0.158 2.95 0.472 ;
        RECT 1.154 0.158 1.222 0.472 ;
      LAYER m2 ;
        RECT 1.136 0.248 2.984 0.292 ;
      LAYER v1 ;
        RECT 1.158 0.248 1.218 0.292 ;
        RECT 2.886 0.248 2.946 0.292 ;
      LAYER v0 ;
        RECT 1.154 0.383 1.222 0.427 ;
        RECT 2.882 0.338 2.95 0.382 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68083325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.68083325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.934 0.158 5.002 0.472 ;
      LAYER v0 ;
        RECT 4.934 0.3155 5.002 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.962 0.068 4.03 0.382 ;
        RECT 3.206 0.068 4.03 0.112 ;
        RECT 3.746 0.068 3.814 0.382 ;
        RECT 3.422 0.068 3.49 0.382 ;
        RECT 3.206 0.068 3.274 0.382 ;
      LAYER v0 ;
        RECT 3.206 0.248 3.274 0.292 ;
        RECT 3.422 0.248 3.49 0.292 ;
        RECT 3.746 0.1725 3.814 0.2165 ;
        RECT 3.962 0.1725 4.03 0.2165 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 5.542 0.652 ;
        RECT 5.366 0.338 5.434 0.652 ;
        RECT 5.15 0.338 5.218 0.652 ;
        RECT 4.826 0.338 4.894 0.652 ;
        RECT 4.61 0.338 4.678 0.652 ;
        RECT 4.394 0.338 4.462 0.652 ;
        RECT 4.178 0.338 4.246 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.558 0.338 2.626 0.652 ;
        RECT 2.342 0.338 2.41 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.558 0.428 2.626 0.472 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 4.178 0.4225 4.246 0.4665 ;
        RECT 4.394 0.4225 4.462 0.4665 ;
        RECT 4.61 0.4225 4.678 0.4665 ;
        RECT 4.826 0.4225 4.894 0.4665 ;
        RECT 5.15 0.4225 5.218 0.4665 ;
        RECT 5.366 0.4225 5.434 0.4665 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 5.542 0.022 ;
        RECT 5.366 -0.022 5.434 0.292 ;
        RECT 5.15 -0.022 5.218 0.292 ;
        RECT 4.826 -0.022 4.894 0.292 ;
        RECT 4.61 -0.022 4.678 0.292 ;
        RECT 4.394 -0.022 4.462 0.292 ;
        RECT 4.178 -0.022 4.246 0.292 ;
        RECT 2.774 -0.022 2.842 0.292 ;
        RECT 2.558 -0.022 2.626 0.292 ;
        RECT 2.126 0.158 2.41 0.202 ;
        RECT 2.126 -0.022 2.194 0.202 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 2.234 0.158 2.302 0.202 ;
        RECT 2.558 0.161 2.626 0.205 ;
        RECT 2.774 0.161 2.842 0.205 ;
        RECT 4.178 0.1725 4.246 0.2165 ;
        RECT 4.394 0.1725 4.462 0.2165 ;
        RECT 4.61 0.1725 4.678 0.2165 ;
        RECT 4.826 0.1725 4.894 0.2165 ;
        RECT 5.15 0.1725 5.218 0.2165 ;
        RECT 5.366 0.1725 5.434 0.2165 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.488 0.338 3.076 0.382 ;
      RECT 3.064 0.248 4.588 0.292 ;
      RECT 3.512 0.338 5.344 0.382 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.472 ;
      RECT 0.722 0.158 0.79 0.472 ;
      RECT 1.046 0.158 1.114 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.262 0.158 1.33 0.472 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.802 0.158 1.87 0.472 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 2.99 0.428 3.53 0.472 ;
      RECT 2.666 0.068 2.734 0.562 ;
      RECT 2.882 0.158 2.95 0.472 ;
      RECT 2.99 0.158 3.058 0.382 ;
      RECT 3.098 0.158 3.166 0.382 ;
      RECT 3.314 0.158 3.382 0.382 ;
      RECT 3.638 0.158 3.706 0.562 ;
      RECT 3.854 0.158 3.922 0.382 ;
      RECT 4.07 0.068 4.138 0.382 ;
      RECT 4.286 0.068 4.354 0.562 ;
      RECT 4.502 0.068 4.57 0.562 ;
      RECT 4.718 0.068 4.786 0.562 ;
      RECT 5.042 0.068 5.11 0.562 ;
      RECT 5.258 0.068 5.326 0.562 ;
    LAYER v1 ;
      RECT 5.262 0.338 5.322 0.382 ;
      RECT 5.046 0.338 5.106 0.382 ;
      RECT 4.722 0.338 4.782 0.382 ;
      RECT 4.506 0.248 4.566 0.292 ;
      RECT 4.29 0.248 4.35 0.292 ;
      RECT 4.074 0.338 4.134 0.382 ;
      RECT 3.858 0.338 3.918 0.382 ;
      RECT 3.642 0.248 3.702 0.292 ;
      RECT 3.534 0.338 3.594 0.382 ;
      RECT 3.318 0.248 3.378 0.292 ;
      RECT 3.102 0.248 3.162 0.292 ;
      RECT 2.994 0.338 3.054 0.382 ;
      RECT 1.05 0.338 1.11 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
      RECT 0.51 0.338 0.57 0.382 ;
    LAYER v0 ;
      RECT 5.258 0.1725 5.326 0.2165 ;
      RECT 5.258 0.4225 5.326 0.4665 ;
      RECT 5.042 0.1725 5.11 0.2165 ;
      RECT 5.042 0.4225 5.11 0.4665 ;
      RECT 4.718 0.1725 4.786 0.2165 ;
      RECT 4.718 0.4225 4.786 0.4665 ;
      RECT 4.502 0.1725 4.57 0.2165 ;
      RECT 4.502 0.4225 4.57 0.4665 ;
      RECT 4.286 0.1725 4.354 0.2165 ;
      RECT 4.286 0.4225 4.354 0.4665 ;
      RECT 4.07 0.1725 4.138 0.2165 ;
      RECT 3.854 0.268 3.922 0.312 ;
      RECT 3.854 0.518 3.922 0.562 ;
      RECT 3.638 0.428 3.706 0.472 ;
      RECT 3.53 0.248 3.598 0.292 ;
      RECT 3.314 0.248 3.382 0.292 ;
      RECT 3.314 0.428 3.382 0.472 ;
      RECT 3.098 0.248 3.166 0.292 ;
      RECT 3.098 0.428 3.166 0.472 ;
      RECT 2.99 0.248 3.058 0.292 ;
      RECT 2.666 0.161 2.734 0.205 ;
      RECT 2.666 0.428 2.734 0.472 ;
      RECT 2.45 0.161 2.518 0.205 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.126 0.338 2.194 0.382 ;
      RECT 2.018 0.158 2.086 0.202 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.383 1.87 0.427 ;
      RECT 1.694 0.178 1.762 0.222 ;
      RECT 1.586 0.383 1.654 0.427 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 1.37 0.178 1.438 0.222 ;
      RECT 1.37 0.383 1.438 0.427 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.262 0.383 1.33 0.427 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 1.046 0.383 1.114 0.427 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.614 0.178 0.682 0.222 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.506 0.178 0.574 0.222 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.182 0.178 0.25 0.222 ;
      RECT 0.182 0.4275 0.25 0.4715 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.158 0.898 0.562 ;
      RECT 0.898 0.518 1.37 0.562 ;
      RECT 1.37 0.338 1.438 0.562 ;
      RECT 1.438 0.518 1.694 0.562 ;
      RECT 1.694 0.158 1.762 0.562 ;
      RECT 1.762 0.518 2.018 0.562 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.086 0.338 2.302 0.382 ;
      RECT 0.682 0.068 0.938 0.112 ;
      RECT 0.938 0.068 1.006 0.472 ;
      RECT 1.006 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.292 ;
      RECT 1.438 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.654 0.068 2.018 0.112 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 2.086 0.248 2.45 0.292 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 3.53 0.158 3.598 0.472 ;
      RECT 3.706 0.518 4.03 0.562 ;
  END
END b15xnr003as1n12x5

MACRO b15xnr003as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xnr003as1n16x5 0 0 ;
  SIZE 8.964 BY 0.63 ;
  SYMMETRY Y ;
  SITE core ;
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAGATEAREA 0.045 LAYER m2 ;
      ANTENNAMAXAREACAR 1.6044445 LAYER m1 ;
      ANTENNAMAXAREACAR 3.08722225 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.391111 LAYER v1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAGATEAREA 0.045 LAYER m2 ;
      ANTENNAMAXAREACAR 1.6044445 LAYER m1 ;
      ANTENNAMAXAREACAR 3.08722225 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.391111 LAYER v1 ;
    PORT
      LAYER m1 ;
        RECT 4.178 0.158 4.246 0.472 ;
        RECT 1.586 0.158 1.654 0.472 ;
      LAYER m2 ;
        RECT 1.568 0.248 4.264 0.292 ;
      LAYER v1 ;
        RECT 1.59 0.248 1.65 0.292 ;
        RECT 4.182 0.248 4.242 0.292 ;
      LAYER v0 ;
        RECT 1.586 0.383 1.654 0.427 ;
        RECT 4.178 0.338 4.246 0.382 ;
    END
  END c
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.653125 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.653125 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 8.39 0.158 8.458 0.472 ;
      LAYER v0 ;
        RECT 8.39 0.3155 8.458 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.59375 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.068 0.682 0.382 ;
        RECT 0.182 0.248 0.682 0.292 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 6.122 0.068 6.19 0.382 ;
        RECT 5.042 0.068 6.19 0.112 ;
        RECT 5.906 0.068 5.974 0.382 ;
        RECT 5.69 0.068 5.758 0.382 ;
        RECT 5.258 0.068 5.326 0.382 ;
        RECT 5.042 0.068 5.11 0.382 ;
      LAYER v0 ;
        RECT 5.042 0.248 5.11 0.292 ;
        RECT 5.258 0.248 5.326 0.292 ;
        RECT 5.69 0.1725 5.758 0.2165 ;
        RECT 5.906 0.1725 5.974 0.2165 ;
        RECT 6.122 0.1725 6.19 0.2165 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 8.998 0.652 ;
        RECT 8.822 0.338 8.89 0.652 ;
        RECT 8.606 0.338 8.674 0.652 ;
        RECT 8.282 0.338 8.35 0.652 ;
        RECT 8.066 0.338 8.134 0.652 ;
        RECT 7.85 0.338 7.918 0.652 ;
        RECT 7.634 0.338 7.702 0.652 ;
        RECT 7.418 0.338 7.486 0.652 ;
        RECT 7.202 0.338 7.27 0.652 ;
        RECT 6.77 0.428 6.838 0.652 ;
        RECT 4.718 0.338 4.786 0.652 ;
        RECT 4.502 0.338 4.57 0.652 ;
        RECT 4.286 0.338 4.354 0.652 ;
        RECT 3.746 0.428 3.814 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.338 3.382 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.508 0.538 0.572 0.582 ;
        RECT 3.314 0.473 3.382 0.517 ;
        RECT 3.53 0.473 3.598 0.517 ;
        RECT 3.746 0.473 3.814 0.517 ;
        RECT 4.286 0.428 4.354 0.472 ;
        RECT 4.502 0.428 4.57 0.472 ;
        RECT 4.718 0.428 4.786 0.472 ;
        RECT 6.77 0.495 6.838 0.539 ;
        RECT 7.202 0.4225 7.27 0.4665 ;
        RECT 7.418 0.4225 7.486 0.4665 ;
        RECT 7.634 0.4225 7.702 0.4665 ;
        RECT 7.85 0.4225 7.918 0.4665 ;
        RECT 8.066 0.4225 8.134 0.4665 ;
        RECT 8.282 0.4225 8.35 0.4665 ;
        RECT 8.606 0.4225 8.674 0.4665 ;
        RECT 8.822 0.4225 8.89 0.4665 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 8.998 0.022 ;
        RECT 8.822 -0.022 8.89 0.292 ;
        RECT 8.606 -0.022 8.674 0.292 ;
        RECT 8.282 -0.022 8.35 0.292 ;
        RECT 8.066 -0.022 8.134 0.292 ;
        RECT 7.85 -0.022 7.918 0.292 ;
        RECT 7.634 -0.022 7.702 0.292 ;
        RECT 7.418 -0.022 7.486 0.292 ;
        RECT 7.202 -0.022 7.27 0.292 ;
        RECT 6.554 -0.022 6.622 0.202 ;
        RECT 4.718 -0.022 4.786 0.292 ;
        RECT 4.502 -0.022 4.57 0.292 ;
        RECT 4.286 -0.022 4.354 0.292 ;
        RECT 3.098 0.158 3.922 0.202 ;
        RECT 3.098 -0.022 3.166 0.202 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 3.206 0.158 3.274 0.202 ;
        RECT 3.53 0.158 3.598 0.202 ;
        RECT 3.746 0.158 3.814 0.202 ;
        RECT 4.286 0.161 4.354 0.205 ;
        RECT 4.502 0.161 4.57 0.205 ;
        RECT 4.718 0.161 4.786 0.205 ;
        RECT 6.554 0.0785 6.622 0.1225 ;
        RECT 7.202 0.1725 7.27 0.2165 ;
        RECT 7.418 0.1725 7.486 0.2165 ;
        RECT 7.634 0.1725 7.702 0.2165 ;
        RECT 7.85 0.1725 7.918 0.2165 ;
        RECT 8.066 0.1725 8.134 0.2165 ;
        RECT 8.282 0.1725 8.35 0.2165 ;
        RECT 8.606 0.1725 8.674 0.2165 ;
        RECT 8.822 0.1725 8.89 0.2165 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.704 0.338 4.912 0.382 ;
      RECT 4.808 0.248 7.828 0.292 ;
      RECT 5.456 0.338 8.8 0.382 ;
    LAYER m1 ;
      RECT 0.722 0.068 0.79 0.472 ;
      RECT 0.938 0.158 1.006 0.472 ;
      RECT 1.262 0.158 1.33 0.472 ;
      RECT 1.586 0.158 1.654 0.472 ;
      RECT 1.694 0.158 1.762 0.472 ;
      RECT 1.91 0.158 1.978 0.472 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 2.45 0.158 2.518 0.472 ;
      RECT 2.774 0.158 2.842 0.472 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 4.826 0.428 5.474 0.472 ;
      RECT 4.178 0.158 4.246 0.472 ;
      RECT 4.394 0.068 4.462 0.562 ;
      RECT 4.61 0.068 4.678 0.562 ;
      RECT 4.826 0.158 4.894 0.382 ;
      RECT 4.934 0.158 5.002 0.382 ;
      RECT 5.15 0.158 5.218 0.382 ;
      RECT 5.366 0.158 5.434 0.382 ;
      RECT 5.582 0.158 5.65 0.472 ;
      RECT 5.798 0.158 5.866 0.382 ;
      RECT 6.014 0.158 6.082 0.382 ;
      RECT 7.094 0.068 7.162 0.382 ;
      RECT 7.31 0.068 7.378 0.562 ;
      RECT 7.526 0.068 7.594 0.562 ;
      RECT 7.742 0.068 7.81 0.562 ;
      RECT 7.958 0.068 8.026 0.562 ;
      RECT 8.174 0.068 8.242 0.562 ;
      RECT 8.498 0.068 8.566 0.562 ;
      RECT 8.714 0.068 8.782 0.562 ;
    LAYER v1 ;
      RECT 8.718 0.338 8.778 0.382 ;
      RECT 8.502 0.338 8.562 0.382 ;
      RECT 8.178 0.338 8.238 0.382 ;
      RECT 7.962 0.338 8.022 0.382 ;
      RECT 7.746 0.248 7.806 0.292 ;
      RECT 7.53 0.248 7.59 0.292 ;
      RECT 7.314 0.248 7.374 0.292 ;
      RECT 7.098 0.338 7.158 0.382 ;
      RECT 6.018 0.338 6.078 0.382 ;
      RECT 5.802 0.338 5.862 0.382 ;
      RECT 5.586 0.248 5.646 0.292 ;
      RECT 5.478 0.338 5.538 0.382 ;
      RECT 5.37 0.248 5.43 0.292 ;
      RECT 5.154 0.248 5.214 0.292 ;
      RECT 4.938 0.248 4.998 0.292 ;
      RECT 4.83 0.338 4.89 0.382 ;
      RECT 1.266 0.338 1.326 0.382 ;
      RECT 0.942 0.338 1.002 0.382 ;
      RECT 0.726 0.338 0.786 0.382 ;
    LAYER v0 ;
      RECT 8.714 0.1725 8.782 0.2165 ;
      RECT 8.714 0.4225 8.782 0.4665 ;
      RECT 8.498 0.1725 8.566 0.2165 ;
      RECT 8.498 0.4225 8.566 0.4665 ;
      RECT 8.174 0.1725 8.242 0.2165 ;
      RECT 8.174 0.4225 8.242 0.4665 ;
      RECT 7.958 0.1725 8.026 0.2165 ;
      RECT 7.958 0.4225 8.026 0.4665 ;
      RECT 7.742 0.1725 7.81 0.2165 ;
      RECT 7.742 0.4225 7.81 0.4665 ;
      RECT 7.526 0.1725 7.594 0.2165 ;
      RECT 7.526 0.4225 7.594 0.4665 ;
      RECT 7.31 0.1725 7.378 0.2165 ;
      RECT 7.31 0.4225 7.378 0.4665 ;
      RECT 7.094 0.1725 7.162 0.2165 ;
      RECT 6.014 0.268 6.082 0.312 ;
      RECT 6.014 0.428 6.082 0.472 ;
      RECT 5.798 0.268 5.866 0.312 ;
      RECT 5.798 0.428 5.866 0.472 ;
      RECT 5.366 0.248 5.434 0.292 ;
      RECT 5.366 0.428 5.434 0.472 ;
      RECT 5.15 0.248 5.218 0.292 ;
      RECT 5.15 0.428 5.218 0.472 ;
      RECT 4.934 0.248 5.002 0.292 ;
      RECT 4.934 0.428 5.002 0.472 ;
      RECT 4.826 0.248 4.894 0.292 ;
      RECT 4.61 0.161 4.678 0.205 ;
      RECT 4.61 0.428 4.678 0.472 ;
      RECT 4.394 0.161 4.462 0.205 ;
      RECT 4.394 0.428 4.462 0.472 ;
      RECT 4.07 0.158 4.138 0.202 ;
      RECT 4.07 0.428 4.138 0.472 ;
      RECT 3.638 0.248 3.706 0.292 ;
      RECT 3.638 0.473 3.706 0.517 ;
      RECT 3.422 0.248 3.49 0.292 ;
      RECT 3.422 0.473 3.49 0.517 ;
      RECT 3.098 0.338 3.166 0.382 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.774 0.178 2.842 0.222 ;
      RECT 2.774 0.383 2.842 0.427 ;
      RECT 2.666 0.178 2.734 0.222 ;
      RECT 2.558 0.383 2.626 0.427 ;
      RECT 2.45 0.178 2.518 0.222 ;
      RECT 2.45 0.383 2.518 0.427 ;
      RECT 2.342 0.178 2.41 0.222 ;
      RECT 2.234 0.383 2.302 0.427 ;
      RECT 2.126 0.178 2.194 0.222 ;
      RECT 2.126 0.383 2.194 0.427 ;
      RECT 2.018 0.178 2.086 0.222 ;
      RECT 2.018 0.383 2.086 0.427 ;
      RECT 1.91 0.178 1.978 0.222 ;
      RECT 1.91 0.383 1.978 0.427 ;
      RECT 1.802 0.178 1.87 0.222 ;
      RECT 1.802 0.383 1.87 0.427 ;
      RECT 1.694 0.178 1.762 0.222 ;
      RECT 1.694 0.383 1.762 0.427 ;
      RECT 1.478 0.178 1.546 0.222 ;
      RECT 1.37 0.383 1.438 0.427 ;
      RECT 1.262 0.178 1.33 0.222 ;
      RECT 1.262 0.383 1.33 0.427 ;
      RECT 1.154 0.383 1.222 0.427 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.938 0.178 1.006 0.222 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.83 0.178 0.898 0.222 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.178 0.79 0.222 ;
      RECT 0.722 0.383 0.79 0.427 ;
      RECT 0.398 0.158 0.466 0.202 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.182 0.428 0.25 0.472 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
      RECT 0.142 0.158 0.574 0.202 ;
      RECT 0.142 0.428 0.614 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.682 0.518 0.83 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.518 1.046 0.562 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.518 1.478 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 1.546 0.518 1.802 0.562 ;
      RECT 1.802 0.338 1.87 0.562 ;
      RECT 1.87 0.518 2.018 0.562 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.086 0.518 2.342 0.562 ;
      RECT 2.342 0.158 2.41 0.562 ;
      RECT 2.41 0.518 2.666 0.562 ;
      RECT 2.666 0.158 2.734 0.562 ;
      RECT 2.734 0.518 3.206 0.562 ;
      RECT 2.99 0.338 3.206 0.382 ;
      RECT 3.206 0.338 3.274 0.562 ;
      RECT 0.898 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.472 ;
      RECT 1.222 0.068 1.37 0.112 ;
      RECT 1.37 0.068 1.438 0.472 ;
      RECT 1.438 0.068 1.802 0.112 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.87 0.068 2.018 0.112 ;
      RECT 2.018 0.068 2.086 0.292 ;
      RECT 2.086 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.472 ;
      RECT 2.302 0.068 2.558 0.112 ;
      RECT 2.558 0.068 2.626 0.472 ;
      RECT 2.626 0.068 2.99 0.112 ;
      RECT 2.99 0.068 3.058 0.292 ;
      RECT 3.422 0.338 3.49 0.562 ;
      RECT 3.49 0.338 3.638 0.382 ;
      RECT 3.638 0.338 3.706 0.562 ;
      RECT 3.706 0.338 3.854 0.382 ;
      RECT 3.854 0.338 3.922 0.562 ;
      RECT 3.922 0.518 4.07 0.562 ;
      RECT 3.058 0.248 4.07 0.292 ;
      RECT 4.07 0.068 4.138 0.562 ;
      RECT 5.474 0.158 5.542 0.472 ;
      RECT 5.65 0.428 6.19 0.472 ;
  END
END b15xnr003as1n16x5

MACRO b15xor002as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor002as1n02x3 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.53875 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.53875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.088 0.898 0.132 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.248 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.383 0.466 0.427 ;
        RECT 0.398 0.2065 0.466 0.2505 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.722 0.3605 0.79 0.4045 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.722 0.2065 0.79 0.2505 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.472 ;
    LAYER v0 ;
      RECT 0.614 0.3605 0.682 0.4045 ;
      RECT 0.506 0.2065 0.574 0.2505 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.182 0.158 0.25 0.202 ;
      RECT 0.074 0.383 0.142 0.427 ;
    LAYER m1 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.358 0.518 0.506 0.562 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.142 0.158 0.29 0.202 ;
      RECT 0.29 0.068 0.358 0.202 ;
      RECT 0.358 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.472 ;
  END
END b15xor002as1n02x3

MACRO b15xor002as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor002as1n02x5 0 0 ;
  SIZE 0.972 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.1455555 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 3.53875 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.292 ;
      LAYER v0 ;
        RECT 0.83 0.088 0.898 0.132 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.665 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.158 0.466 0.472 ;
      LAYER v0 ;
        RECT 0.398 0.383 0.466 0.427 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.006 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.722 0.383 0.79 0.427 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.006 0.022 ;
        RECT 0.722 -0.022 0.79 0.292 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.722 0.203 0.79 0.247 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.182 0.472 ;
    LAYER v0 ;
      RECT 0.614 0.383 0.682 0.427 ;
      RECT 0.506 0.203 0.574 0.247 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.182 0.203 0.25 0.247 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.29 0.338 0.358 0.562 ;
      RECT 0.358 0.518 0.506 0.562 ;
      RECT 0.506 0.158 0.574 0.562 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.25 0.068 0.614 0.112 ;
      RECT 0.614 0.068 0.682 0.472 ;
  END
END b15xor002as1n02x5

MACRO b15xor002as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor002as1n03x5 0 0 ;
  SIZE 1.08 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0099 LAYER m1 ;
      ANTENNAMAXAREACAR 2.57363625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.009 LAYER m1 ;
      ANTENNAMAXAREACAR 2.831 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.938 0.068 1.006 0.292 ;
      LAYER v0 ;
        RECT 0.938 0.088 1.006 0.132 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.158 0.574 0.472 ;
      LAYER v0 ;
        RECT 0.506 0.408 0.574 0.452 ;
        RECT 0.506 0.203 0.574 0.247 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.114 0.652 ;
        RECT 0.83 0.428 0.898 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.493 0.358 0.537 ;
        RECT 0.83 0.448 0.898 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.114 0.022 ;
        RECT 0.83 -0.022 0.898 0.292 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.83 0.2065 0.898 0.2505 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.158 0.182 0.202 ;
    LAYER v0 ;
      RECT 0.722 0.3605 0.79 0.4045 ;
      RECT 0.614 0.203 0.682 0.247 ;
      RECT 0.398 0.408 0.466 0.452 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.182 0.408 0.25 0.452 ;
      RECT 0.074 0.158 0.142 0.202 ;
    LAYER m1 ;
      RECT 0.398 0.338 0.466 0.562 ;
      RECT 0.466 0.518 0.614 0.562 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.158 0.398 0.202 ;
      RECT 0.398 0.068 0.466 0.202 ;
      RECT 0.466 0.068 0.722 0.112 ;
      RECT 0.722 0.068 0.79 0.472 ;
  END
END b15xor002as1n03x5

MACRO b15xor002as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor002as1n04x5 0 0 ;
  SIZE 1.296 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.35916675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 2.17769225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.722 0.068 0.79 0.292 ;
      LAYER v0 ;
        RECT 0.722 0.088 0.79 0.132 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.6175 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0153 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5811765 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.338 0.142 0.382 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02754 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.046 0.158 1.114 0.472 ;
      LAYER v0 ;
        RECT 1.046 0.363 1.114 0.407 ;
        RECT 1.046 0.232 1.114 0.276 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.33 0.652 ;
        RECT 0.506 0.518 0.574 0.652 ;
        RECT 0.29 0.518 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.076 0.538 0.14 0.582 ;
        RECT 0.292 0.538 0.356 0.582 ;
        RECT 0.506 0.538 0.574 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.33 0.022 ;
        RECT 0.614 -0.022 0.682 0.292 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.074 0.048 0.142 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.614 0.228 0.682 0.272 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.182 0.158 0.25 0.562 ;
    LAYER v0 ;
      RECT 1.156 0.138 1.22 0.182 ;
      RECT 1.156 0.448 1.22 0.492 ;
      RECT 0.938 0.232 1.006 0.276 ;
      RECT 0.832 0.408 0.896 0.452 ;
      RECT 0.506 0.088 0.574 0.132 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.223 0.25 0.267 ;
      RECT 0.182 0.448 0.25 0.492 ;
    LAYER m1 ;
      RECT 0.29 0.428 0.614 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.682 0.518 0.938 0.562 ;
      RECT 0.938 0.158 1.006 0.562 ;
      RECT 1.006 0.518 1.154 0.562 ;
      RECT 1.154 0.428 1.222 0.562 ;
      RECT 0.25 0.338 0.506 0.382 ;
      RECT 0.506 0.068 0.574 0.382 ;
      RECT 0.574 0.338 0.83 0.382 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 0.898 0.068 1.154 0.112 ;
      RECT 1.154 0.068 1.222 0.202 ;
  END
END b15xor002as1n04x5

MACRO b15xor002as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor002as1n06x5 0 0 ;
  SIZE 1.62 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0171 LAYER m1 ;
      ANTENNAMAXAREACAR 2.31 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0171 LAYER m1 ;
      ANTENNAMAXAREACAR 2.31 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.068 0.898 0.382 ;
      LAYER v0 ;
        RECT 0.83 0.088 0.898 0.132 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.60166675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.182 0.158 0.25 0.472 ;
      LAYER v0 ;
        RECT 0.182 0.293 0.25 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.05508 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.068 1.546 0.472 ;
        RECT 0.938 0.068 1.546 0.112 ;
        RECT 1.262 0.068 1.33 0.472 ;
        RECT 0.938 0.068 1.006 0.472 ;
      LAYER v0 ;
        RECT 0.938 0.396 1.006 0.44 ;
        RECT 0.938 0.178 1.006 0.222 ;
        RECT 1.262 0.396 1.33 0.44 ;
        RECT 1.262 0.178 1.33 0.222 ;
        RECT 1.478 0.396 1.546 0.44 ;
        RECT 1.478 0.178 1.546 0.222 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.654 0.652 ;
        RECT 0.614 0.428 0.682 0.652 ;
        RECT 0.398 0.428 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.538 0.25 0.582 ;
        RECT 0.398 0.473 0.466 0.517 ;
        RECT 0.614 0.473 0.682 0.517 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.654 0.022 ;
        RECT 0.614 -0.022 0.682 0.202 ;
        RECT 0.398 -0.022 0.466 0.202 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.182 0.048 0.25 0.092 ;
        RECT 0.398 0.138 0.466 0.182 ;
        RECT 0.614 0.138 0.682 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.158 1.456 0.202 ;
    LAYER m1 ;
      RECT 0.074 0.068 0.142 0.472 ;
      RECT 0.29 0.068 0.358 0.472 ;
      RECT 1.154 0.158 1.222 0.472 ;
      RECT 1.37 0.158 1.438 0.292 ;
    LAYER v1 ;
      RECT 1.374 0.158 1.434 0.202 ;
      RECT 1.158 0.158 1.218 0.202 ;
      RECT 0.294 0.158 0.354 0.202 ;
      RECT 0.078 0.158 0.138 0.202 ;
    LAYER v0 ;
      RECT 1.37 0.178 1.438 0.222 ;
      RECT 1.37 0.396 1.438 0.44 ;
      RECT 1.154 0.396 1.222 0.44 ;
      RECT 1.046 0.178 1.114 0.222 ;
      RECT 0.506 0.138 0.574 0.182 ;
      RECT 0.506 0.383 0.574 0.427 ;
      RECT 0.29 0.138 0.358 0.182 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.074 0.138 0.142 0.182 ;
      RECT 0.074 0.383 0.142 0.427 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.472 ;
      RECT 0.574 0.248 0.722 0.292 ;
      RECT 0.722 0.248 0.79 0.562 ;
      RECT 0.79 0.518 1.046 0.562 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.518 1.37 0.562 ;
      RECT 1.37 0.338 1.438 0.562 ;
  END
END b15xor002as1n06x5

MACRO b15xor002as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor002as1n08x5 0 0 ;
  SIZE 1.944 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9475 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.9475 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.158 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.389 1.222 0.433 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.158 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.074 0.248 0.142 0.292 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.06732 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.068 1.87 0.472 ;
        RECT 1.37 0.068 1.87 0.112 ;
        RECT 1.586 0.068 1.654 0.472 ;
        RECT 1.37 0.068 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.37 0.389 1.438 0.433 ;
        RECT 1.37 0.203 1.438 0.247 ;
        RECT 1.586 0.389 1.654 0.433 ;
        RECT 1.586 0.178 1.654 0.222 ;
        RECT 1.802 0.389 1.87 0.433 ;
        RECT 1.802 0.178 1.87 0.222 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 1.978 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.478 0.358 0.522 ;
        RECT 0.506 0.448 0.574 0.492 ;
        RECT 0.722 0.448 0.79 0.492 ;
        RECT 0.938 0.448 1.006 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 1.978 0.022 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.202 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.29 0.138 0.358 0.182 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.722 0.048 0.79 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.158 1.78 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.472 ;
      RECT 0.614 0.338 0.682 0.562 ;
      RECT 1.262 0.158 1.33 0.472 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 1.694 0.158 1.762 0.292 ;
    LAYER v1 ;
      RECT 1.698 0.158 1.758 0.202 ;
      RECT 1.482 0.158 1.542 0.202 ;
      RECT 1.266 0.158 1.326 0.202 ;
      RECT 0.402 0.158 0.462 0.202 ;
      RECT 0.186 0.158 0.246 0.202 ;
    LAYER v0 ;
      RECT 1.694 0.178 1.762 0.222 ;
      RECT 1.694 0.389 1.762 0.433 ;
      RECT 1.478 0.389 1.546 0.433 ;
      RECT 1.262 0.389 1.33 0.433 ;
      RECT 1.154 0.068 1.222 0.112 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.448 0.898 0.492 ;
      RECT 0.614 0.158 0.682 0.202 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.398 0.363 0.466 0.407 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.182 0.3835 0.25 0.4275 ;
    LAYER m1 ;
      RECT 0.398 0.068 0.466 0.472 ;
      RECT 0.466 0.248 0.918 0.292 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.338 1.046 0.382 ;
      RECT 0.506 0.158 1.046 0.202 ;
      RECT 1.046 0.068 1.114 0.562 ;
      RECT 1.114 0.068 1.33 0.112 ;
      RECT 1.114 0.518 1.694 0.562 ;
      RECT 1.694 0.338 1.762 0.562 ;
  END
END b15xor002as1n08x5

MACRO b15xor002as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor002as1n12x5 0 0 ;
  SIZE 2.7 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0324 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0324 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.342 0.248 2.41 0.472 ;
        RECT 2.234 0.248 2.41 0.292 ;
        RECT 2.234 0.068 2.302 0.292 ;
        RECT 1.566 0.068 2.302 0.112 ;
      LAYER v0 ;
        RECT 1.586 0.068 1.654 0.112 ;
        RECT 2.342 0.338 2.41 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0441 LAYER m1 ;
      ANTENNAMAXAREACAR 0.430839 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.142 0.382 ;
      LAYER v0 ;
        RECT 0.074 0.293 0.142 0.337 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.605 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 5.605 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.458 0.518 2.302 0.562 ;
        RECT 2.234 0.338 2.302 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.518 1.546 0.562 ;
        RECT 1.802 0.518 1.87 0.562 ;
        RECT 2.018 0.518 2.086 0.562 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.734 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.518 2.41 0.652 ;
        RECT 1.154 0.518 1.222 0.652 ;
        RECT 0.938 0.518 1.006 0.652 ;
        RECT 0.722 0.518 0.79 0.652 ;
        RECT 0.398 0.518 0.466 0.652 ;
        RECT 0.182 0.518 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.184 0.538 0.248 0.582 ;
        RECT 0.4 0.538 0.464 0.582 ;
        RECT 0.724 0.538 0.788 0.582 ;
        RECT 0.94 0.538 1.004 0.582 ;
        RECT 1.156 0.538 1.22 0.582 ;
        RECT 2.342 0.538 2.41 0.582 ;
        RECT 2.558 0.538 2.626 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.734 0.022 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 2.342 -0.022 2.41 0.202 ;
        RECT 1.154 -0.022 1.222 0.202 ;
        RECT 0.938 -0.022 1.006 0.202 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.398 -0.022 0.466 0.112 ;
        RECT 0.182 -0.022 0.25 0.112 ;
      LAYER v0 ;
        RECT 0.184 0.048 0.248 0.092 ;
        RECT 0.4 0.048 0.464 0.092 ;
        RECT 0.722 0.138 0.79 0.182 ;
        RECT 0.938 0.138 1.006 0.182 ;
        RECT 1.154 0.138 1.222 0.182 ;
        RECT 2.342 0.138 2.41 0.182 ;
        RECT 2.558 0.138 2.626 0.182 ;
    END
  END vssx
  OBS
    LAYER m1 ;
      RECT 0.054 0.428 0.182 0.472 ;
      RECT 1.134 0.338 1.37 0.382 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 2.45 0.068 2.518 0.562 ;
    LAYER v0 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.445 2.518 0.489 ;
      RECT 2.128 0.228 2.192 0.272 ;
      RECT 2.128 0.408 2.192 0.452 ;
      RECT 1.91 0.158 1.978 0.202 ;
      RECT 1.912 0.408 1.976 0.452 ;
      RECT 1.586 0.428 1.654 0.472 ;
      RECT 1.588 0.268 1.652 0.312 ;
      RECT 1.37 0.428 1.438 0.472 ;
      RECT 1.372 0.268 1.436 0.312 ;
      RECT 1.154 0.338 1.222 0.382 ;
      RECT 1.046 0.138 1.114 0.182 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.83 0.428 0.898 0.472 ;
      RECT 0.722 0.338 0.79 0.382 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.158 0.142 0.202 ;
      RECT 0.074 0.428 0.142 0.472 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.472 ;
      RECT 0.682 0.338 0.898 0.382 ;
      RECT 0.054 0.158 0.182 0.202 ;
      RECT 0.182 0.158 0.25 0.472 ;
      RECT 0.25 0.428 0.614 0.472 ;
      RECT 0.25 0.158 0.614 0.202 ;
      RECT 1.37 0.248 1.438 0.382 ;
      RECT 1.438 0.338 1.586 0.382 ;
      RECT 1.586 0.248 1.654 0.382 ;
      RECT 1.654 0.338 1.91 0.382 ;
      RECT 1.91 0.338 1.978 0.472 ;
      RECT 1.978 0.338 2.126 0.382 ;
      RECT 2.126 0.338 2.194 0.472 ;
      RECT 0.722 0.428 0.938 0.472 ;
      RECT 0.898 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 1.006 0.248 1.046 0.292 ;
      RECT 1.046 0.068 1.114 0.292 ;
      RECT 1.114 0.248 1.262 0.292 ;
      RECT 1.262 0.158 1.33 0.292 ;
      RECT 1.006 0.428 1.674 0.472 ;
      RECT 1.33 0.158 2.126 0.202 ;
      RECT 2.126 0.158 2.194 0.292 ;
  END
END b15xor002as1n12x5

MACRO b15xor002as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor002as1n16x5 0 0 ;
  SIZE 3.348 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 1.59916675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 1.59916675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.91 0.428 1.978 0.562 ;
      LAYER v0 ;
        RECT 1.91 0.448 1.978 0.492 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.543611 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.543611 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.074 0.248 0.682 0.292 ;
        RECT 0.074 0.248 0.142 0.472 ;
      LAYER v0 ;
        RECT 0.29 0.248 0.358 0.292 ;
        RECT 0.506 0.248 0.574 0.292 ;
    END
  END b
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.206 0.068 3.274 0.472 ;
        RECT 2.126 0.068 3.274 0.112 ;
        RECT 2.99 0.068 3.058 0.472 ;
        RECT 2.774 0.068 2.842 0.472 ;
        RECT 2.558 0.068 2.626 0.472 ;
        RECT 2.342 0.068 2.41 0.472 ;
        RECT 2.126 0.068 2.194 0.472 ;
      LAYER v0 ;
        RECT 2.126 0.389 2.194 0.433 ;
        RECT 2.126 0.203 2.194 0.247 ;
        RECT 2.342 0.389 2.41 0.433 ;
        RECT 2.342 0.203 2.41 0.247 ;
        RECT 2.558 0.389 2.626 0.433 ;
        RECT 2.558 0.203 2.626 0.247 ;
        RECT 2.774 0.389 2.842 0.433 ;
        RECT 2.774 0.178 2.842 0.222 ;
        RECT 2.99 0.389 3.058 0.433 ;
        RECT 2.99 0.178 3.058 0.222 ;
        RECT 3.206 0.389 3.274 0.433 ;
        RECT 3.206 0.178 3.274 0.222 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.382 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 1.154 0.428 1.222 0.652 ;
        RECT 0.938 0.428 1.006 0.652 ;
        RECT 0.722 0.428 0.79 0.652 ;
        RECT 0.506 0.428 0.574 0.652 ;
        RECT 0.29 0.428 0.358 0.652 ;
        RECT 0.074 0.518 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.538 0.142 0.582 ;
        RECT 0.29 0.493 0.358 0.537 ;
        RECT 0.506 0.493 0.574 0.537 ;
        RECT 0.722 0.493 0.79 0.537 ;
        RECT 0.938 0.493 1.006 0.537 ;
        RECT 1.154 0.493 1.222 0.537 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.448 1.654 0.492 ;
        RECT 1.802 0.448 1.87 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.382 0.022 ;
        RECT 1.802 -0.022 1.87 0.112 ;
        RECT 1.586 -0.022 1.654 0.112 ;
        RECT 1.37 -0.022 1.438 0.112 ;
        RECT 1.154 -0.022 1.222 0.112 ;
        RECT 0.938 -0.022 1.006 0.112 ;
        RECT 0.722 -0.022 0.79 0.112 ;
        RECT 0.506 -0.022 0.574 0.112 ;
        RECT 0.29 -0.022 0.358 0.112 ;
        RECT 0.074 -0.022 0.142 0.112 ;
      LAYER v0 ;
        RECT 0.076 0.048 0.14 0.092 ;
        RECT 0.292 0.048 0.356 0.092 ;
        RECT 0.508 0.048 0.572 0.092 ;
        RECT 0.724 0.048 0.788 0.092 ;
        RECT 0.94 0.048 1.004 0.092 ;
        RECT 1.156 0.048 1.22 0.092 ;
        RECT 1.372 0.048 1.436 0.092 ;
        RECT 1.588 0.048 1.652 0.092 ;
        RECT 1.804 0.048 1.868 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.164 0.158 3.184 0.202 ;
    LAYER m1 ;
      RECT 0.182 0.068 0.25 0.202 ;
      RECT 0.398 0.068 0.466 0.202 ;
      RECT 0.614 0.068 0.682 0.202 ;
      RECT 1.694 0.248 1.762 0.562 ;
      RECT 1.046 0.338 1.114 0.472 ;
      RECT 2.234 0.158 2.302 0.472 ;
      RECT 2.45 0.158 2.518 0.472 ;
      RECT 2.666 0.158 2.734 0.472 ;
      RECT 2.882 0.158 2.95 0.292 ;
      RECT 3.098 0.158 3.166 0.292 ;
    LAYER v1 ;
      RECT 3.102 0.158 3.162 0.202 ;
      RECT 2.886 0.158 2.946 0.202 ;
      RECT 2.67 0.158 2.73 0.202 ;
      RECT 2.454 0.158 2.514 0.202 ;
      RECT 2.238 0.158 2.298 0.202 ;
      RECT 0.834 0.158 0.894 0.202 ;
      RECT 0.618 0.158 0.678 0.202 ;
      RECT 0.402 0.158 0.462 0.202 ;
      RECT 0.186 0.158 0.246 0.202 ;
    LAYER v0 ;
      RECT 3.098 0.178 3.166 0.222 ;
      RECT 3.098 0.389 3.166 0.433 ;
      RECT 2.882 0.178 2.95 0.222 ;
      RECT 2.882 0.389 2.95 0.433 ;
      RECT 2.666 0.389 2.734 0.433 ;
      RECT 2.45 0.389 2.518 0.433 ;
      RECT 2.234 0.389 2.302 0.433 ;
      RECT 2.018 0.088 2.086 0.132 ;
      RECT 1.91 0.268 1.978 0.312 ;
      RECT 1.694 0.268 1.762 0.312 ;
      RECT 1.694 0.448 1.762 0.492 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.448 1.546 0.492 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.248 1.33 0.292 ;
      RECT 1.264 0.408 1.328 0.452 ;
      RECT 1.046 0.158 1.114 0.202 ;
      RECT 1.046 0.248 1.114 0.292 ;
      RECT 1.048 0.408 1.112 0.452 ;
      RECT 0.83 0.138 0.898 0.182 ;
      RECT 0.832 0.408 0.896 0.452 ;
      RECT 0.614 0.138 0.682 0.182 ;
      RECT 0.616 0.408 0.68 0.452 ;
      RECT 0.398 0.138 0.466 0.182 ;
      RECT 0.4 0.408 0.464 0.452 ;
      RECT 0.182 0.138 0.25 0.182 ;
      RECT 0.184 0.408 0.248 0.452 ;
    LAYER m1 ;
      RECT 0.182 0.338 0.25 0.472 ;
      RECT 0.25 0.338 0.398 0.382 ;
      RECT 0.398 0.338 0.466 0.472 ;
      RECT 0.466 0.338 0.614 0.382 ;
      RECT 0.614 0.338 0.682 0.472 ;
      RECT 0.682 0.338 0.83 0.382 ;
      RECT 0.83 0.068 0.898 0.472 ;
      RECT 0.898 0.248 1.35 0.292 ;
      RECT 1.762 0.338 1.91 0.382 ;
      RECT 1.91 0.248 1.978 0.382 ;
      RECT 1.114 0.338 1.262 0.382 ;
      RECT 1.262 0.338 1.33 0.472 ;
      RECT 1.33 0.338 1.478 0.382 ;
      RECT 1.478 0.338 1.546 0.562 ;
      RECT 1.546 0.338 1.586 0.382 ;
      RECT 0.938 0.158 1.586 0.202 ;
      RECT 1.586 0.158 1.654 0.382 ;
      RECT 1.654 0.158 2.018 0.202 ;
      RECT 2.018 0.068 2.086 0.562 ;
      RECT 2.086 0.518 2.882 0.562 ;
      RECT 2.882 0.338 2.95 0.562 ;
      RECT 2.95 0.518 3.098 0.562 ;
      RECT 3.098 0.338 3.166 0.562 ;
  END
END b15xor002as1n16x5

MACRO b15xor003as1n02x3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor003as1n02x3 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.158 2.194 0.382 ;
      LAYER v0 ;
        RECT 2.126 0.293 2.194 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0036 LAYER m1 ;
      ANTENNAMAXAREACAR 0.71777775 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.158 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.9485185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.9485185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.802 0.203 1.87 0.247 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 1.37 0.383 1.438 0.427 ;
        RECT 2.126 0.448 2.194 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 2.126 0.048 2.194 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.068 0.824 0.112 ;
      RECT 0.04 0.518 1.256 0.562 ;
      RECT 0.904 0.068 2.012 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.614 0.158 0.83 0.202 ;
      RECT 0.398 0.338 0.722 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.478 0.068 1.546 0.472 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.91 0.068 1.978 0.382 ;
      RECT 2.018 0.158 2.086 0.562 ;
    LAYER v1 ;
      RECT 1.914 0.068 1.974 0.112 ;
      RECT 1.59 0.068 1.65 0.112 ;
      RECT 1.158 0.518 1.218 0.562 ;
      RECT 0.942 0.068 1.002 0.112 ;
      RECT 0.618 0.518 0.678 0.562 ;
      RECT 0.51 0.068 0.57 0.112 ;
      RECT 0.078 0.068 0.138 0.112 ;
      RECT 0.078 0.518 0.138 0.562 ;
    LAYER v0 ;
      RECT 2.018 0.203 2.086 0.247 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 1.154 0.4055 1.222 0.4495 ;
      RECT 1.046 0.268 1.114 0.312 ;
      RECT 0.938 0.268 1.006 0.312 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.29 0.203 0.358 0.247 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.574 0.248 0.83 0.292 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.006 0.112 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.518 1.046 0.562 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.158 1.222 0.562 ;
  END
END b15xor003as1n02x3

MACRO b15xor003as1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor003as1n02x5 0 0 ;
  SIZE 2.268 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.358889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.158 2.194 0.382 ;
      LAYER v0 ;
        RECT 2.126 0.293 2.194 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0054 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4785185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.262 0.158 1.33 0.382 ;
      LAYER v0 ;
        RECT 1.262 0.293 1.33 0.337 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.9485185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.9485185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01224 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.586 0.428 1.87 0.472 ;
        RECT 1.802 0.158 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.694 0.428 1.762 0.472 ;
        RECT 1.802 0.203 1.87 0.247 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.302 0.652 ;
        RECT 2.126 0.428 2.194 0.652 ;
        RECT 1.37 0.338 1.438 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 1.37 0.383 1.438 0.427 ;
        RECT 2.126 0.448 2.194 0.492 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.302 0.022 ;
        RECT 2.126 -0.022 2.194 0.112 ;
        RECT 1.37 -0.022 1.438 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 1.37 0.158 1.438 0.202 ;
        RECT 2.126 0.048 2.194 0.092 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.068 0.824 0.112 ;
      RECT 0.04 0.518 1.256 0.562 ;
      RECT 0.904 0.068 2.012 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.614 0.158 0.83 0.202 ;
      RECT 0.398 0.338 0.722 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.478 0.518 2.018 0.562 ;
      RECT 1.478 0.068 1.546 0.472 ;
      RECT 1.586 0.068 1.654 0.382 ;
      RECT 1.91 0.068 1.978 0.382 ;
    LAYER v1 ;
      RECT 1.914 0.068 1.974 0.112 ;
      RECT 1.59 0.068 1.65 0.112 ;
      RECT 1.158 0.518 1.218 0.562 ;
      RECT 0.942 0.068 1.002 0.112 ;
      RECT 0.618 0.518 0.678 0.562 ;
      RECT 0.51 0.068 0.57 0.112 ;
      RECT 0.078 0.068 0.138 0.112 ;
      RECT 0.078 0.518 0.138 0.562 ;
    LAYER v0 ;
      RECT 2.018 0.203 2.086 0.247 ;
      RECT 2.018 0.448 2.086 0.492 ;
      RECT 1.91 0.293 1.978 0.337 ;
      RECT 1.802 0.518 1.87 0.562 ;
      RECT 1.586 0.293 1.654 0.337 ;
      RECT 1.586 0.518 1.654 0.562 ;
      RECT 1.478 0.158 1.546 0.202 ;
      RECT 1.478 0.383 1.546 0.427 ;
      RECT 1.154 0.4055 1.222 0.4495 ;
      RECT 1.046 0.268 1.114 0.312 ;
      RECT 0.938 0.268 1.006 0.312 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.29 0.203 0.358 0.247 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.574 0.248 0.83 0.292 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.006 0.112 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.518 1.046 0.562 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.006 0.158 1.154 0.202 ;
      RECT 1.154 0.158 1.222 0.562 ;
      RECT 2.018 0.158 2.086 0.562 ;
  END
END b15xor003as1n02x5

MACRO b15xor003as1n03x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor003as1n03x5 0 0 ;
  SIZE 2.484 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.41518525 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.234 0.248 2.302 0.472 ;
      LAYER v0 ;
        RECT 2.234 0.3155 2.302 0.3595 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 0.928889 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.154 0.248 1.222 0.472 ;
      LAYER v0 ;
        RECT 1.154 0.3485 1.222 0.3925 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.9485185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.9485185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.398 0.068 0.466 0.292 ;
      LAYER v0 ;
        RECT 0.398 0.203 0.466 0.247 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.01836 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.158 1.87 0.472 ;
      LAYER v0 ;
        RECT 1.802 0.408 1.87 0.452 ;
        RECT 1.802 0.186 1.87 0.23 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.518 0.652 ;
        RECT 2.234 0.518 2.302 0.652 ;
        RECT 1.37 0.428 1.438 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.383 0.25 0.427 ;
        RECT 1.37 0.473 1.438 0.517 ;
        RECT 2.234 0.538 2.302 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.518 0.022 ;
        RECT 2.234 -0.022 2.302 0.202 ;
        RECT 1.37 -0.022 1.438 0.382 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.203 0.25 0.247 ;
        RECT 1.37 0.228 1.438 0.272 ;
        RECT 2.234 0.138 2.302 0.182 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.068 0.824 0.112 ;
      RECT 0.04 0.518 1.364 0.562 ;
      RECT 0.904 0.068 2.104 0.112 ;
      RECT 1.444 0.518 2.444 0.562 ;
    LAYER m1 ;
      RECT 0.074 0.428 0.142 0.562 ;
      RECT 0.074 0.068 0.142 0.292 ;
      RECT 0.29 0.158 0.358 0.472 ;
      RECT 0.614 0.428 0.682 0.562 ;
      RECT 0.614 0.158 0.83 0.202 ;
      RECT 0.398 0.338 0.722 0.382 ;
      RECT 0.938 0.158 1.006 0.382 ;
      RECT 1.586 0.248 1.654 0.562 ;
      RECT 1.478 0.068 1.546 0.562 ;
      RECT 2.018 0.068 2.086 0.472 ;
      RECT 2.126 0.068 2.194 0.562 ;
      RECT 2.342 0.068 2.41 0.562 ;
    LAYER v1 ;
      RECT 2.346 0.518 2.406 0.562 ;
      RECT 2.13 0.518 2.19 0.562 ;
      RECT 2.022 0.068 2.082 0.112 ;
      RECT 1.59 0.518 1.65 0.562 ;
      RECT 1.266 0.518 1.326 0.562 ;
      RECT 0.942 0.068 1.002 0.112 ;
      RECT 0.618 0.518 0.678 0.562 ;
      RECT 0.51 0.068 0.57 0.112 ;
      RECT 0.078 0.068 0.138 0.112 ;
      RECT 0.078 0.518 0.138 0.562 ;
    LAYER v0 ;
      RECT 2.342 0.138 2.41 0.182 ;
      RECT 2.342 0.449 2.41 0.493 ;
      RECT 2.126 0.138 2.194 0.182 ;
      RECT 2.126 0.435 2.194 0.479 ;
      RECT 2.018 0.3155 2.086 0.3595 ;
      RECT 1.91 0.408 1.978 0.452 ;
      RECT 1.694 0.518 1.762 0.562 ;
      RECT 1.586 0.338 1.654 0.382 ;
      RECT 1.478 0.228 1.546 0.272 ;
      RECT 1.478 0.473 1.546 0.517 ;
      RECT 1.262 0.228 1.33 0.272 ;
      RECT 1.262 0.473 1.33 0.517 ;
      RECT 1.046 0.268 1.114 0.312 ;
      RECT 0.938 0.268 1.006 0.312 ;
      RECT 0.83 0.383 0.898 0.427 ;
      RECT 0.722 0.158 0.79 0.202 ;
      RECT 0.614 0.248 0.682 0.292 ;
      RECT 0.614 0.448 0.682 0.492 ;
      RECT 0.506 0.338 0.574 0.382 ;
      RECT 0.29 0.203 0.358 0.247 ;
      RECT 0.29 0.383 0.358 0.427 ;
      RECT 0.074 0.203 0.142 0.247 ;
      RECT 0.074 0.498 0.142 0.542 ;
    LAYER m1 ;
      RECT 0.506 0.068 0.574 0.292 ;
      RECT 0.574 0.248 0.83 0.292 ;
      RECT 0.83 0.248 0.898 0.472 ;
      RECT 0.83 0.068 0.898 0.202 ;
      RECT 0.898 0.068 1.006 0.112 ;
      RECT 0.722 0.338 0.79 0.562 ;
      RECT 0.79 0.518 1.046 0.562 ;
      RECT 1.046 0.248 1.114 0.562 ;
      RECT 1.006 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.654 0.518 1.87 0.562 ;
      RECT 1.546 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.562 ;
  END
END b15xor003as1n03x5

MACRO b15xor003as1n04x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor003as1n04x5 0 0 ;
  SIZE 2.808 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.311389 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.248 2.626 0.472 ;
      LAYER v0 ;
        RECT 2.558 0.293 2.626 0.337 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 0.61925925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.37 0.248 1.438 0.472 ;
      LAYER v0 ;
        RECT 1.37 0.338 1.438 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.9485185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.9485185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.203 0.574 0.247 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.02448 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.126 0.158 2.194 0.562 ;
      LAYER v0 ;
        RECT 2.126 0.428 2.194 0.472 ;
        RECT 2.126 0.186 2.194 0.23 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 1.802 0.428 1.87 0.652 ;
        RECT 1.586 0.428 1.654 0.652 ;
        RECT 1.37 0.518 1.438 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.383 0.142 0.427 ;
        RECT 0.29 0.383 0.358 0.427 ;
        RECT 1.37 0.538 1.438 0.582 ;
        RECT 1.586 0.456 1.654 0.5 ;
        RECT 1.802 0.456 1.87 0.5 ;
        RECT 2.56 0.538 2.624 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 2.842 0.022 ;
        RECT 2.558 -0.022 2.626 0.202 ;
        RECT 1.802 -0.022 1.87 0.292 ;
        RECT 1.586 -0.022 1.654 0.292 ;
        RECT 1.37 -0.022 1.438 0.202 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.29 0.203 0.358 0.247 ;
        RECT 1.37 0.13 1.438 0.174 ;
        RECT 1.586 0.2105 1.654 0.2545 ;
        RECT 1.802 0.2105 1.87 0.2545 ;
        RECT 2.558 0.13 2.626 0.174 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.068 0.824 0.112 ;
      RECT 0.04 0.518 1.688 0.562 ;
      RECT 0.904 0.068 2.444 0.112 ;
      RECT 1.768 0.518 2.768 0.562 ;
    LAYER m1 ;
      RECT 0.182 0.428 0.25 0.562 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.722 0.158 0.938 0.202 ;
      RECT 0.506 0.338 0.83 0.382 ;
      RECT 1.046 0.158 1.114 0.382 ;
      RECT 1.694 0.158 1.762 0.562 ;
      RECT 1.478 0.158 1.546 0.562 ;
      RECT 2.018 0.338 2.086 0.562 ;
      RECT 2.342 0.068 2.41 0.382 ;
      RECT 2.45 0.068 2.518 0.562 ;
      RECT 2.666 0.068 2.734 0.562 ;
    LAYER v1 ;
      RECT 2.67 0.518 2.73 0.562 ;
      RECT 2.454 0.518 2.514 0.562 ;
      RECT 2.346 0.068 2.406 0.112 ;
      RECT 2.022 0.518 2.082 0.562 ;
      RECT 1.482 0.518 1.542 0.562 ;
      RECT 1.266 0.518 1.326 0.562 ;
      RECT 1.05 0.068 1.11 0.112 ;
      RECT 0.726 0.518 0.786 0.562 ;
      RECT 0.618 0.068 0.678 0.112 ;
      RECT 0.186 0.068 0.246 0.112 ;
      RECT 0.186 0.518 0.246 0.562 ;
    LAYER v0 ;
      RECT 2.666 0.13 2.734 0.174 ;
      RECT 2.666 0.449 2.734 0.493 ;
      RECT 2.45 0.13 2.518 0.174 ;
      RECT 2.45 0.435 2.518 0.479 ;
      RECT 2.342 0.293 2.41 0.337 ;
      RECT 2.234 0.428 2.302 0.472 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.91 0.2105 1.978 0.2545 ;
      RECT 1.694 0.2105 1.762 0.2545 ;
      RECT 1.694 0.456 1.762 0.5 ;
      RECT 1.478 0.2105 1.546 0.2545 ;
      RECT 1.478 0.456 1.546 0.5 ;
      RECT 1.154 0.268 1.222 0.312 ;
      RECT 1.046 0.268 1.114 0.312 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.182 0.203 0.25 0.247 ;
      RECT 0.182 0.498 0.25 0.542 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.006 0.068 1.114 0.112 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.518 1.154 0.562 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 1.114 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.762 0.338 1.91 0.382 ;
      RECT 1.91 0.068 1.978 0.382 ;
      RECT 1.978 0.068 2.234 0.112 ;
      RECT 2.234 0.068 2.302 0.562 ;
  END
END b15xor003as1n04x5

MACRO b15xor003as1n06x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor003as1n06x5 0 0 ;
  SIZE 3.456 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5875925 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 0.5875925 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.558 0.248 2.626 0.472 ;
      LAYER v0 ;
        RECT 2.558 0.338 2.626 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0117 LAYER m1 ;
      ANTENNAMAXAREACAR 0.571624 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.314 0.248 3.382 0.472 ;
      LAYER v0 ;
        RECT 3.314 0.3155 3.382 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.9485185 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 2.9485185 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.506 0.068 0.574 0.292 ;
      LAYER v0 ;
        RECT 0.506 0.203 0.574 0.247 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.07344 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 3.67333325 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0081 LAYER m1 ;
      ANTENNAMAXAREACAR 5.57333325 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.478 0.518 2.302 0.562 ;
        RECT 2.234 0.248 2.302 0.562 ;
        RECT 1.802 0.158 1.87 0.562 ;
        RECT 1.478 0.068 1.546 0.562 ;
      LAYER v0 ;
        RECT 1.478 0.408 1.546 0.452 ;
        RECT 1.478 0.158 1.546 0.202 ;
        RECT 1.802 0.428 1.87 0.472 ;
        RECT 1.802 0.186 1.87 0.23 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.276 2.302 0.32 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 3.49 0.652 ;
        RECT 3.314 0.518 3.382 0.652 ;
        RECT 3.098 0.338 3.166 0.652 ;
        RECT 2.774 0.338 2.842 0.652 ;
        RECT 2.558 0.518 2.626 0.652 ;
        RECT 2.342 0.248 2.41 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
        RECT 0.074 0.338 0.142 0.652 ;
      LAYER v0 ;
        RECT 0.074 0.383 0.142 0.427 ;
        RECT 0.29 0.383 0.358 0.427 ;
        RECT 2.342 0.428 2.41 0.472 ;
        RECT 2.558 0.538 2.626 0.582 ;
        RECT 2.774 0.4505 2.842 0.4945 ;
        RECT 3.098 0.4505 3.166 0.4945 ;
        RECT 3.314 0.538 3.382 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 3.49 0.022 ;
        RECT 3.314 -0.022 3.382 0.202 ;
        RECT 3.098 -0.022 3.166 0.292 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 2.558 -0.022 2.626 0.112 ;
        RECT 2.342 -0.022 2.41 0.112 ;
        RECT 0.29 -0.022 0.358 0.292 ;
        RECT 0.074 -0.022 0.142 0.292 ;
      LAYER v0 ;
        RECT 0.074 0.203 0.142 0.247 ;
        RECT 0.29 0.203 0.358 0.247 ;
        RECT 2.342 0.048 2.41 0.092 ;
        RECT 2.558 0.048 2.626 0.092 ;
        RECT 2.882 0.048 2.95 0.092 ;
        RECT 3.098 0.158 3.166 0.202 ;
        RECT 3.314 0.068 3.382 0.112 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.068 0.824 0.112 ;
      RECT 0.904 0.068 1.472 0.112 ;
      RECT 0.04 0.518 3.416 0.562 ;
      RECT 1.552 0.068 3.416 0.112 ;
    LAYER m1 ;
      RECT 0.182 0.428 0.25 0.562 ;
      RECT 0.182 0.068 0.25 0.292 ;
      RECT 0.398 0.158 0.466 0.472 ;
      RECT 0.722 0.428 0.79 0.562 ;
      RECT 0.722 0.158 0.938 0.202 ;
      RECT 0.506 0.338 0.83 0.382 ;
      RECT 1.046 0.158 1.114 0.382 ;
      RECT 1.694 0.068 1.762 0.292 ;
      RECT 1.37 0.068 1.438 0.472 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 2.018 0.068 2.086 0.382 ;
      RECT 2.99 0.068 3.058 0.562 ;
      RECT 3.206 0.068 3.274 0.562 ;
    LAYER v1 ;
      RECT 3.21 0.518 3.27 0.562 ;
      RECT 2.994 0.068 3.054 0.112 ;
      RECT 2.022 0.068 2.082 0.112 ;
      RECT 1.59 0.068 1.65 0.112 ;
      RECT 1.374 0.068 1.434 0.112 ;
      RECT 1.266 0.518 1.326 0.562 ;
      RECT 1.05 0.068 1.11 0.112 ;
      RECT 0.726 0.518 0.786 0.562 ;
      RECT 0.618 0.068 0.678 0.112 ;
      RECT 0.186 0.068 0.246 0.112 ;
      RECT 0.186 0.518 0.246 0.562 ;
    LAYER v0 ;
      RECT 3.206 0.158 3.274 0.202 ;
      RECT 3.206 0.4505 3.274 0.4945 ;
      RECT 2.99 0.158 3.058 0.202 ;
      RECT 2.99 0.4505 3.058 0.4945 ;
      RECT 2.882 0.3155 2.95 0.3595 ;
      RECT 2.666 0.4505 2.734 0.4945 ;
      RECT 2.668 0.228 2.732 0.272 ;
      RECT 2.45 0.428 2.518 0.472 ;
      RECT 2.452 0.228 2.516 0.272 ;
      RECT 2.018 0.186 2.086 0.23 ;
      RECT 2.018 0.428 2.086 0.472 ;
      RECT 1.694 0.186 1.762 0.23 ;
      RECT 1.586 0.408 1.654 0.452 ;
      RECT 1.37 0.3155 1.438 0.3595 ;
      RECT 1.154 0.268 1.222 0.312 ;
      RECT 1.046 0.268 1.114 0.312 ;
      RECT 0.938 0.383 1.006 0.427 ;
      RECT 0.83 0.158 0.898 0.202 ;
      RECT 0.722 0.248 0.79 0.292 ;
      RECT 0.722 0.448 0.79 0.492 ;
      RECT 0.614 0.338 0.682 0.382 ;
      RECT 0.398 0.203 0.466 0.247 ;
      RECT 0.398 0.383 0.466 0.427 ;
      RECT 0.182 0.203 0.25 0.247 ;
      RECT 0.182 0.498 0.25 0.542 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.248 0.938 0.292 ;
      RECT 0.938 0.248 1.006 0.472 ;
      RECT 0.938 0.068 1.006 0.202 ;
      RECT 1.006 0.068 1.114 0.112 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 0.898 0.518 1.154 0.562 ;
      RECT 1.154 0.248 1.222 0.562 ;
      RECT 1.114 0.158 1.262 0.202 ;
      RECT 1.262 0.158 1.33 0.562 ;
      RECT 1.762 0.068 1.91 0.112 ;
      RECT 1.91 0.068 1.978 0.472 ;
      RECT 1.978 0.428 2.126 0.472 ;
      RECT 2.126 0.158 2.194 0.472 ;
      RECT 2.194 0.158 2.45 0.202 ;
      RECT 2.45 0.158 2.518 0.562 ;
      RECT 2.518 0.158 2.666 0.202 ;
      RECT 2.666 0.158 2.734 0.562 ;
      RECT 2.734 0.158 2.882 0.202 ;
      RECT 2.882 0.158 2.95 0.472 ;
  END
END b15xor003as1n06x5

MACRO b15xor003as1n08x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor003as1n08x5 0 0 ;
  SIZE 4.212 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4406945 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.248 3.166 0.472 ;
      LAYER v0 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.07 0.248 4.138 0.472 ;
      LAYER v0 ;
        RECT 4.07 0.3155 4.138 0.3595 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.71791675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.71791675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 3.23 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0108 LAYER m1 ;
      ANTENNAMAXAREACAR 4.655 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 1.802 0.518 2.842 0.562 ;
        RECT 2.774 0.248 2.842 0.562 ;
        RECT 2.234 0.158 2.302 0.562 ;
        RECT 1.802 0.068 1.87 0.562 ;
      LAYER v0 ;
        RECT 1.802 0.3675 1.87 0.4115 ;
        RECT 1.802 0.158 1.87 0.202 ;
        RECT 2.234 0.428 2.302 0.472 ;
        RECT 2.234 0.186 2.302 0.23 ;
        RECT 2.774 0.428 2.842 0.472 ;
        RECT 2.774 0.276 2.842 0.32 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.246 0.652 ;
        RECT 4.07 0.518 4.138 0.652 ;
        RECT 3.854 0.338 3.922 0.652 ;
        RECT 3.638 0.338 3.706 0.652 ;
        RECT 3.314 0.338 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.248 2.95 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 2.882 0.428 2.95 0.472 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.314 0.4505 3.382 0.4945 ;
        RECT 3.638 0.4505 3.706 0.4945 ;
        RECT 3.854 0.4505 3.922 0.4945 ;
        RECT 4.072 0.538 4.136 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.246 0.022 ;
        RECT 4.07 -0.022 4.138 0.202 ;
        RECT 3.854 -0.022 3.922 0.292 ;
        RECT 3.638 -0.022 3.706 0.292 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 2.882 0.048 2.95 0.092 ;
        RECT 3.098 0.048 3.166 0.092 ;
        RECT 3.314 0.048 3.382 0.092 ;
        RECT 3.638 0.158 3.706 0.202 ;
        RECT 3.854 0.158 3.922 0.202 ;
        RECT 4.07 0.068 4.138 0.112 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.068 0.716 0.112 ;
      RECT 0.04 0.518 4.172 0.562 ;
      RECT 1.876 0.068 4.172 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 2.126 0.068 2.194 0.292 ;
      RECT 1.91 0.068 1.978 0.472 ;
      RECT 2.558 0.068 2.626 0.382 ;
      RECT 3.53 0.068 3.598 0.562 ;
      RECT 3.746 0.068 3.814 0.562 ;
      RECT 3.962 0.068 4.03 0.562 ;
    LAYER v1 ;
      RECT 3.966 0.518 4.026 0.562 ;
      RECT 3.75 0.068 3.81 0.112 ;
      RECT 3.534 0.068 3.594 0.112 ;
      RECT 2.562 0.068 2.622 0.112 ;
      RECT 1.914 0.068 1.974 0.112 ;
      RECT 1.266 0.518 1.326 0.562 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.618 0.068 0.678 0.112 ;
      RECT 0.294 0.068 0.354 0.112 ;
      RECT 0.078 0.518 0.138 0.562 ;
    LAYER v0 ;
      RECT 3.962 0.158 4.03 0.202 ;
      RECT 3.962 0.4505 4.03 0.4945 ;
      RECT 3.746 0.158 3.814 0.202 ;
      RECT 3.746 0.4505 3.814 0.4945 ;
      RECT 3.53 0.158 3.598 0.202 ;
      RECT 3.53 0.4505 3.598 0.4945 ;
      RECT 3.422 0.3155 3.49 0.3595 ;
      RECT 3.206 0.4505 3.274 0.4945 ;
      RECT 3.208 0.228 3.272 0.272 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.992 0.228 3.056 0.272 ;
      RECT 2.558 0.186 2.626 0.23 ;
      RECT 2.558 0.428 2.626 0.472 ;
      RECT 2.126 0.186 2.194 0.23 ;
      RECT 1.91 0.3675 1.978 0.4115 ;
      RECT 1.696 0.448 1.76 0.492 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.36 1.654 0.404 ;
      RECT 1.478 0.36 1.546 0.404 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.156 0.318 1.22 0.362 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.411 0.898 0.455 ;
      RECT 0.724 0.138 0.788 0.182 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 0.79 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.438 0.518 1.694 0.562 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 2.194 0.068 2.342 0.112 ;
      RECT 2.342 0.068 2.41 0.472 ;
      RECT 2.41 0.428 2.666 0.472 ;
      RECT 2.666 0.158 2.734 0.472 ;
      RECT 2.734 0.158 2.99 0.202 ;
      RECT 2.99 0.158 3.058 0.562 ;
      RECT 3.058 0.158 3.206 0.202 ;
      RECT 3.206 0.158 3.274 0.562 ;
      RECT 3.274 0.158 3.422 0.202 ;
      RECT 3.422 0.158 3.49 0.472 ;
  END
END b15xor003as1n08x5

MACRO b15xor003as1n12x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor003as1n12x5 0 0 ;
  SIZE 4.428 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.48379625 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 0.48379625 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 3.098 0.248 3.166 0.472 ;
      LAYER v0 ;
        RECT 3.098 0.338 3.166 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0144 LAYER m1 ;
      ANTENNAMAXAREACAR 0.4644445 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.286 0.248 4.354 0.472 ;
      LAYER v0 ;
        RECT 4.286 0.338 4.354 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.71791675 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0216 LAYER m1 ;
      ANTENNAMAXAREACAR 1.71791675 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.614 0.338 0.682 0.562 ;
      LAYER v0 ;
        RECT 0.614 0.428 0.682 0.472 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.09792 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.018 0.518 2.626 0.562 ;
        RECT 2.558 0.338 2.626 0.562 ;
        RECT 2.234 0.158 2.302 0.562 ;
        RECT 2.018 0.338 2.086 0.562 ;
      LAYER v0 ;
        RECT 2.018 0.4 2.086 0.444 ;
        RECT 2.234 0.4 2.302 0.444 ;
        RECT 2.234 0.2185 2.302 0.2625 ;
        RECT 2.558 0.4 2.626 0.444 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 4.462 0.652 ;
        RECT 4.286 0.518 4.354 0.652 ;
        RECT 4.07 0.338 4.138 0.652 ;
        RECT 3.854 0.338 3.922 0.652 ;
        RECT 3.53 0.428 3.598 0.652 ;
        RECT 3.314 0.338 3.382 0.652 ;
        RECT 3.098 0.518 3.166 0.652 ;
        RECT 2.882 0.428 2.95 0.652 ;
        RECT 0.398 0.338 0.466 0.652 ;
        RECT 0.182 0.338 0.25 0.652 ;
      LAYER v0 ;
        RECT 0.182 0.428 0.25 0.472 ;
        RECT 0.398 0.428 0.466 0.472 ;
        RECT 2.882 0.518 2.95 0.562 ;
        RECT 3.1 0.538 3.164 0.582 ;
        RECT 3.314 0.428 3.382 0.472 ;
        RECT 3.53 0.518 3.598 0.562 ;
        RECT 3.854 0.4505 3.922 0.4945 ;
        RECT 4.07 0.4505 4.138 0.4945 ;
        RECT 4.288 0.538 4.352 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 4.462 0.022 ;
        RECT 4.286 -0.022 4.354 0.202 ;
        RECT 4.07 -0.022 4.138 0.292 ;
        RECT 3.854 -0.022 3.922 0.292 ;
        RECT 3.53 -0.022 3.598 0.112 ;
        RECT 3.314 -0.022 3.382 0.112 ;
        RECT 3.098 -0.022 3.166 0.112 ;
        RECT 2.882 -0.022 2.95 0.112 ;
        RECT 0.398 -0.022 0.466 0.292 ;
        RECT 0.182 -0.022 0.25 0.292 ;
      LAYER v0 ;
        RECT 0.182 0.158 0.25 0.202 ;
        RECT 0.398 0.158 0.466 0.202 ;
        RECT 2.882 0.048 2.95 0.092 ;
        RECT 3.098 0.048 3.166 0.092 ;
        RECT 3.314 0.048 3.382 0.092 ;
        RECT 3.53 0.048 3.598 0.092 ;
        RECT 3.854 0.158 3.922 0.202 ;
        RECT 4.07 0.158 4.138 0.202 ;
        RECT 4.286 0.068 4.354 0.112 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.068 0.716 0.112 ;
      RECT 0.04 0.518 4.264 0.562 ;
      RECT 1.784 0.068 4.388 0.112 ;
    LAYER m1 ;
      RECT 0.074 0.248 0.142 0.562 ;
      RECT 0.29 0.068 0.358 0.562 ;
      RECT 0.506 0.068 0.574 0.562 ;
      RECT 0.83 0.338 0.898 0.562 ;
      RECT 1.262 0.338 1.33 0.562 ;
      RECT 0.722 0.068 0.79 0.202 ;
      RECT 1.154 0.248 1.222 0.472 ;
      RECT 1.802 0.068 1.87 0.292 ;
      RECT 1.91 0.068 1.978 0.202 ;
      RECT 2.45 0.068 2.518 0.202 ;
      RECT 2.666 0.068 2.734 0.202 ;
      RECT 3.746 0.068 3.814 0.562 ;
      RECT 3.962 0.068 4.03 0.562 ;
      RECT 4.178 0.068 4.246 0.562 ;
    LAYER v1 ;
      RECT 4.182 0.518 4.242 0.562 ;
      RECT 3.966 0.068 4.026 0.112 ;
      RECT 3.75 0.068 3.81 0.112 ;
      RECT 2.67 0.068 2.73 0.112 ;
      RECT 2.454 0.068 2.514 0.112 ;
      RECT 1.806 0.068 1.866 0.112 ;
      RECT 1.266 0.518 1.326 0.562 ;
      RECT 0.834 0.518 0.894 0.562 ;
      RECT 0.618 0.068 0.678 0.112 ;
      RECT 0.294 0.068 0.354 0.112 ;
      RECT 0.078 0.518 0.138 0.562 ;
    LAYER v0 ;
      RECT 4.178 0.158 4.246 0.202 ;
      RECT 4.178 0.4505 4.246 0.4945 ;
      RECT 3.962 0.158 4.03 0.202 ;
      RECT 3.962 0.4505 4.03 0.4945 ;
      RECT 3.746 0.158 3.814 0.202 ;
      RECT 3.746 0.4505 3.814 0.4945 ;
      RECT 3.638 0.338 3.706 0.382 ;
      RECT 3.422 0.428 3.49 0.472 ;
      RECT 3.424 0.228 3.488 0.272 ;
      RECT 3.206 0.428 3.274 0.472 ;
      RECT 3.208 0.228 3.272 0.272 ;
      RECT 2.99 0.428 3.058 0.472 ;
      RECT 2.992 0.228 3.056 0.272 ;
      RECT 2.666 0.138 2.734 0.182 ;
      RECT 2.666 0.4 2.734 0.444 ;
      RECT 2.45 0.138 2.518 0.182 ;
      RECT 2.45 0.4 2.518 0.444 ;
      RECT 2.126 0.4 2.194 0.444 ;
      RECT 2.128 0.138 2.192 0.182 ;
      RECT 1.91 0.4 1.978 0.444 ;
      RECT 1.912 0.138 1.976 0.182 ;
      RECT 1.696 0.448 1.76 0.492 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.586 0.36 1.654 0.404 ;
      RECT 1.478 0.36 1.546 0.404 ;
      RECT 1.262 0.158 1.33 0.202 ;
      RECT 1.262 0.428 1.33 0.472 ;
      RECT 1.156 0.318 1.22 0.362 ;
      RECT 1.046 0.428 1.114 0.472 ;
      RECT 0.83 0.248 0.898 0.292 ;
      RECT 0.83 0.411 0.898 0.455 ;
      RECT 0.724 0.138 0.788 0.182 ;
      RECT 0.506 0.158 0.574 0.202 ;
      RECT 0.506 0.428 0.574 0.472 ;
      RECT 0.29 0.158 0.358 0.202 ;
      RECT 0.29 0.428 0.358 0.472 ;
      RECT 0.074 0.293 0.142 0.337 ;
    LAYER m1 ;
      RECT 0.614 0.068 0.682 0.292 ;
      RECT 0.682 0.248 1.046 0.292 ;
      RECT 1.046 0.158 1.114 0.562 ;
      RECT 1.114 0.158 1.478 0.202 ;
      RECT 1.478 0.158 1.546 0.472 ;
      RECT 0.79 0.068 1.586 0.112 ;
      RECT 1.586 0.068 1.654 0.472 ;
      RECT 1.222 0.248 1.37 0.292 ;
      RECT 1.37 0.248 1.438 0.562 ;
      RECT 1.438 0.518 1.694 0.562 ;
      RECT 1.694 0.338 1.762 0.562 ;
      RECT 1.87 0.248 1.91 0.292 ;
      RECT 1.91 0.248 1.978 0.472 ;
      RECT 1.978 0.248 2.126 0.292 ;
      RECT 2.126 0.248 2.194 0.472 ;
      RECT 1.978 0.068 2.126 0.112 ;
      RECT 2.126 0.068 2.194 0.202 ;
      RECT 2.194 0.068 2.342 0.112 ;
      RECT 2.342 0.068 2.41 0.292 ;
      RECT 2.41 0.248 2.45 0.292 ;
      RECT 2.45 0.248 2.518 0.472 ;
      RECT 2.518 0.248 2.666 0.292 ;
      RECT 2.666 0.248 2.734 0.472 ;
      RECT 2.734 0.248 2.774 0.292 ;
      RECT 2.774 0.158 2.842 0.292 ;
      RECT 2.842 0.158 2.99 0.202 ;
      RECT 2.99 0.158 3.058 0.562 ;
      RECT 3.058 0.158 3.206 0.202 ;
      RECT 3.206 0.158 3.274 0.562 ;
      RECT 3.274 0.158 3.422 0.202 ;
      RECT 3.422 0.158 3.49 0.562 ;
      RECT 3.49 0.158 3.638 0.202 ;
      RECT 3.638 0.158 3.706 0.472 ;
  END
END b15xor003as1n12x5

MACRO b15xor003as1n16x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN b15xor003as1n16x5 0 0 ;
  SIZE 6.156 BY 0.63 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.50534725 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0576 LAYER m1 ;
      ANTENNAMAXAREACAR 0.50534725 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 4.394 0.248 4.462 0.472 ;
      LAYER v0 ;
        RECT 4.394 0.338 4.462 0.382 ;
    END
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0288 LAYER m1 ;
      ANTENNAMAXAREACAR 0.51722225 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 6.014 0.248 6.082 0.472 ;
      LAYER v0 ;
        RECT 6.014 0.338 6.082 0.382 ;
    END
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 1.23895825 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0432 LAYER m1 ;
      ANTENNAMAXAREACAR 1.23895825 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 0.83 0.338 0.898 0.562 ;
      LAYER v0 ;
        RECT 0.83 0.428 0.898 0.472 ;
    END
  END c
  PIN out0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14688 LAYER m1 ;
    ANTENNAMODEL OXIDE2 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    ANTENNAMODEL OXIDE3 ;
      ANTENNAGATEAREA 0.0072 LAYER m1 ;
      ANTENNAMAXAREACAR 4.18 LAYER m1 ;
    PORT
      LAYER m1 ;
        RECT 2.774 0.518 3.814 0.562 ;
        RECT 3.746 0.338 3.814 0.562 ;
        RECT 3.53 0.338 3.598 0.562 ;
        RECT 3.206 0.158 3.274 0.562 ;
        RECT 2.99 0.338 3.058 0.562 ;
        RECT 2.774 0.338 2.842 0.562 ;
      LAYER v0 ;
        RECT 2.774 0.4 2.842 0.444 ;
        RECT 2.99 0.4 3.058 0.444 ;
        RECT 3.206 0.4 3.274 0.444 ;
        RECT 3.206 0.2185 3.274 0.2625 ;
        RECT 3.53 0.4 3.598 0.444 ;
        RECT 3.746 0.4 3.814 0.444 ;
    END
  END out0
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 0.608 6.19 0.652 ;
        RECT 6.014 0.518 6.082 0.652 ;
        RECT 5.798 0.338 5.866 0.652 ;
        RECT 5.582 0.338 5.65 0.652 ;
        RECT 5.366 0.338 5.434 0.652 ;
        RECT 5.15 0.338 5.218 0.652 ;
        RECT 4.826 0.428 4.894 0.652 ;
        RECT 4.61 0.338 4.678 0.652 ;
        RECT 4.394 0.518 4.462 0.652 ;
        RECT 4.178 0.338 4.246 0.652 ;
        RECT 3.962 0.338 4.03 0.652 ;
        RECT 0.722 0.338 0.79 0.652 ;
        RECT 0.506 0.338 0.574 0.652 ;
        RECT 0.29 0.338 0.358 0.652 ;
      LAYER v0 ;
        RECT 0.29 0.428 0.358 0.472 ;
        RECT 0.506 0.428 0.574 0.472 ;
        RECT 0.722 0.428 0.79 0.472 ;
        RECT 3.962 0.428 4.03 0.472 ;
        RECT 4.178 0.428 4.246 0.472 ;
        RECT 4.396 0.538 4.46 0.582 ;
        RECT 4.61 0.428 4.678 0.472 ;
        RECT 4.826 0.518 4.894 0.562 ;
        RECT 5.15 0.4505 5.218 0.4945 ;
        RECT 5.366 0.4505 5.434 0.4945 ;
        RECT 5.582 0.4505 5.65 0.4945 ;
        RECT 5.798 0.4505 5.866 0.4945 ;
        RECT 6.016 0.538 6.08 0.582 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER m1 ;
        RECT -0.034 -0.022 6.19 0.022 ;
        RECT 6.014 -0.022 6.082 0.202 ;
        RECT 5.798 -0.022 5.866 0.292 ;
        RECT 5.582 -0.022 5.65 0.292 ;
        RECT 5.366 -0.022 5.434 0.292 ;
        RECT 5.15 -0.022 5.218 0.292 ;
        RECT 4.826 -0.022 4.894 0.112 ;
        RECT 4.61 -0.022 4.678 0.112 ;
        RECT 4.394 -0.022 4.462 0.112 ;
        RECT 4.178 -0.022 4.246 0.112 ;
        RECT 3.962 -0.022 4.03 0.112 ;
        RECT 0.722 -0.022 0.79 0.202 ;
        RECT 0.506 -0.022 0.574 0.202 ;
        RECT 0.29 -0.022 0.358 0.202 ;
      LAYER v0 ;
        RECT 0.29 0.096 0.358 0.14 ;
        RECT 0.506 0.096 0.574 0.14 ;
        RECT 0.722 0.096 0.79 0.14 ;
        RECT 3.962 0.048 4.03 0.092 ;
        RECT 4.178 0.048 4.246 0.092 ;
        RECT 4.394 0.048 4.462 0.092 ;
        RECT 4.61 0.048 4.678 0.092 ;
        RECT 4.826 0.048 4.894 0.092 ;
        RECT 5.15 0.158 5.218 0.202 ;
        RECT 5.366 0.158 5.434 0.202 ;
        RECT 5.582 0.158 5.65 0.202 ;
        RECT 5.798 0.158 5.866 0.202 ;
        RECT 6.014 0.068 6.082 0.112 ;
    END
  END vssx
  OBS
    LAYER m2 ;
      RECT 0.04 0.068 1.024 0.112 ;
      RECT 2.756 0.068 5.56 0.112 ;
      RECT 0.04 0.518 5.992 0.562 ;
    LAYER m1 ;
      RECT 0.074 0.158 0.142 0.562 ;
      RECT 0.182 0.068 0.25 0.562 ;
      RECT 0.398 0.068 0.466 0.562 ;
      RECT 1.37 0.338 1.91 0.382 ;
      RECT 1.154 0.338 1.222 0.562 ;
      RECT 1.802 0.428 1.87 0.562 ;
      RECT 0.938 0.068 1.006 0.292 ;
      RECT 1.566 0.158 2.126 0.202 ;
      RECT 1.046 0.068 1.114 0.202 ;
      RECT 2.774 0.068 2.842 0.292 ;
      RECT 2.882 0.068 2.95 0.202 ;
      RECT 3.422 0.068 3.49 0.202 ;
      RECT 3.638 0.068 3.706 0.202 ;
      RECT 5.042 0.068 5.11 0.562 ;
      RECT 5.258 0.068 5.326 0.562 ;
      RECT 5.474 0.068 5.542 0.562 ;
      RECT 5.69 0.068 5.758 0.562 ;
      RECT 5.906 0.068 5.974 0.562 ;
    LAYER v1 ;
      RECT 5.91 0.518 5.97 0.562 ;
      RECT 5.694 0.518 5.754 0.562 ;
      RECT 5.478 0.068 5.538 0.112 ;
      RECT 5.262 0.068 5.322 0.112 ;
      RECT 5.046 0.068 5.106 0.112 ;
      RECT 3.642 0.068 3.702 0.112 ;
      RECT 3.426 0.068 3.486 0.112 ;
      RECT 2.778 0.068 2.838 0.112 ;
      RECT 2.67 0.518 2.73 0.562 ;
      RECT 1.806 0.518 1.866 0.562 ;
      RECT 1.158 0.518 1.218 0.562 ;
      RECT 0.942 0.068 1.002 0.112 ;
      RECT 0.402 0.068 0.462 0.112 ;
      RECT 0.186 0.068 0.246 0.112 ;
      RECT 0.078 0.518 0.138 0.562 ;
    LAYER v0 ;
      RECT 5.906 0.158 5.974 0.202 ;
      RECT 5.906 0.4505 5.974 0.4945 ;
      RECT 5.69 0.158 5.758 0.202 ;
      RECT 5.69 0.4505 5.758 0.4945 ;
      RECT 5.474 0.158 5.542 0.202 ;
      RECT 5.474 0.4505 5.542 0.4945 ;
      RECT 5.258 0.158 5.326 0.202 ;
      RECT 5.258 0.4505 5.326 0.4945 ;
      RECT 5.042 0.158 5.11 0.202 ;
      RECT 5.042 0.4505 5.11 0.4945 ;
      RECT 4.934 0.338 5.002 0.382 ;
      RECT 4.718 0.428 4.786 0.472 ;
      RECT 4.72 0.228 4.784 0.272 ;
      RECT 4.502 0.428 4.57 0.472 ;
      RECT 4.504 0.228 4.568 0.272 ;
      RECT 4.286 0.428 4.354 0.472 ;
      RECT 4.288 0.228 4.352 0.272 ;
      RECT 4.07 0.428 4.138 0.472 ;
      RECT 4.072 0.228 4.136 0.272 ;
      RECT 3.638 0.138 3.706 0.182 ;
      RECT 3.638 0.4 3.706 0.444 ;
      RECT 3.422 0.138 3.49 0.182 ;
      RECT 3.422 0.4 3.49 0.444 ;
      RECT 3.098 0.4 3.166 0.444 ;
      RECT 3.1 0.138 3.164 0.182 ;
      RECT 2.882 0.4 2.95 0.444 ;
      RECT 2.884 0.138 2.948 0.182 ;
      RECT 2.666 0.138 2.734 0.182 ;
      RECT 2.56 0.448 2.624 0.492 ;
      RECT 2.45 0.248 2.518 0.292 ;
      RECT 2.45 0.338 2.518 0.382 ;
      RECT 2.344 0.138 2.408 0.182 ;
      RECT 2.234 0.248 2.302 0.292 ;
      RECT 2.236 0.408 2.3 0.452 ;
      RECT 1.912 0.408 1.976 0.452 ;
      RECT 1.802 0.248 1.87 0.292 ;
      RECT 1.802 0.4885 1.87 0.5325 ;
      RECT 1.694 0.338 1.762 0.382 ;
      RECT 1.586 0.158 1.654 0.202 ;
      RECT 1.588 0.448 1.652 0.492 ;
      RECT 1.478 0.338 1.546 0.382 ;
      RECT 1.264 0.138 1.328 0.182 ;
      RECT 1.154 0.248 1.222 0.292 ;
      RECT 1.154 0.4385 1.222 0.4825 ;
      RECT 1.048 0.138 1.112 0.182 ;
      RECT 0.83 0.096 0.898 0.14 ;
      RECT 0.614 0.428 0.682 0.472 ;
      RECT 0.616 0.178 0.68 0.222 ;
      RECT 0.398 0.096 0.466 0.14 ;
      RECT 0.398 0.428 0.466 0.472 ;
      RECT 0.182 0.096 0.25 0.14 ;
      RECT 0.182 0.428 0.25 0.472 ;
      RECT 0.074 0.2705 0.142 0.3145 ;
    LAYER m1 ;
      RECT 0.614 0.158 0.682 0.562 ;
      RECT 0.682 0.248 0.83 0.292 ;
      RECT 0.83 0.068 0.898 0.292 ;
      RECT 1.91 0.338 1.978 0.562 ;
      RECT 1.978 0.518 2.558 0.562 ;
      RECT 2.558 0.428 2.626 0.562 ;
      RECT 1.006 0.248 1.262 0.292 ;
      RECT 1.262 0.248 1.33 0.562 ;
      RECT 1.33 0.518 1.586 0.562 ;
      RECT 1.586 0.428 1.654 0.562 ;
      RECT 1.33 0.248 2.018 0.292 ;
      RECT 2.018 0.248 2.086 0.382 ;
      RECT 2.086 0.338 2.234 0.382 ;
      RECT 2.234 0.338 2.302 0.472 ;
      RECT 2.302 0.338 2.626 0.382 ;
      RECT 2.126 0.158 2.194 0.292 ;
      RECT 2.194 0.248 2.666 0.292 ;
      RECT 2.666 0.248 2.734 0.562 ;
      RECT 1.114 0.068 1.262 0.112 ;
      RECT 1.262 0.068 1.33 0.202 ;
      RECT 1.33 0.068 2.342 0.112 ;
      RECT 2.342 0.068 2.41 0.202 ;
      RECT 2.41 0.068 2.666 0.112 ;
      RECT 2.666 0.068 2.734 0.202 ;
      RECT 2.842 0.248 2.882 0.292 ;
      RECT 2.882 0.248 2.95 0.472 ;
      RECT 2.95 0.248 3.098 0.292 ;
      RECT 3.098 0.248 3.166 0.472 ;
      RECT 2.95 0.068 3.098 0.112 ;
      RECT 3.098 0.068 3.166 0.202 ;
      RECT 3.166 0.068 3.314 0.112 ;
      RECT 3.314 0.068 3.382 0.292 ;
      RECT 3.382 0.248 3.422 0.292 ;
      RECT 3.422 0.248 3.49 0.472 ;
      RECT 3.49 0.248 3.638 0.292 ;
      RECT 3.638 0.248 3.706 0.472 ;
      RECT 3.706 0.248 3.746 0.292 ;
      RECT 3.746 0.158 3.814 0.292 ;
      RECT 3.814 0.158 4.07 0.202 ;
      RECT 4.07 0.158 4.138 0.562 ;
      RECT 4.138 0.158 4.286 0.202 ;
      RECT 4.286 0.158 4.354 0.562 ;
      RECT 4.354 0.158 4.502 0.202 ;
      RECT 4.502 0.158 4.57 0.562 ;
      RECT 4.57 0.158 4.718 0.202 ;
      RECT 4.718 0.158 4.786 0.562 ;
      RECT 4.786 0.158 4.934 0.202 ;
      RECT 4.934 0.158 5.002 0.472 ;
  END
END b15xor003as1n16x5

END LIBRARY
