module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire net10;
 wire net9;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire net8;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire net7;
 wire _211_;
 wire _212_;
 wire _213_;
 wire net6;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire net5;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire net4;
 wire _238_;
 wire _239_;
 wire net3;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire net2;
 wire _253_;
 wire _254_;
 wire net1;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 b15inv000aq1n02x5 _308_ (.a(\dpath.a_lt_b$in0[0] ),
    .o1(_035_));
 b15nand02ar1n12x5 _309_ (.a(_035_),
    .b(\dpath.a_lt_b$in1[0] ),
    .o1(_036_));
 b15inv040ah1n02x5 _310_ (.a(\dpath.a_lt_b$in1[0] ),
    .o1(_037_));
 b15nandp2ah1n02x5 _311_ (.a(_037_),
    .b(\dpath.a_lt_b$in0[0] ),
    .o1(_038_));
 b15nand02aq1n06x5 _312_ (.a(_036_),
    .b(_038_),
    .o1(net37));
 b15nor004an1n04x5 _313_ (.a(\dpath.a_lt_b$in1[15] ),
    .b(\dpath.a_lt_b$in1[14] ),
    .c(\dpath.a_lt_b$in1[13] ),
    .d(\dpath.a_lt_b$in1[12] ),
    .o1(_039_));
 b15nor004aq1n03x5 _314_ (.a(\dpath.a_lt_b$in1[11] ),
    .b(\dpath.a_lt_b$in1[10] ),
    .c(\dpath.a_lt_b$in1[9] ),
    .d(\dpath.a_lt_b$in1[8] ),
    .o1(_040_));
 b15nor004as1n04x5 _315_ (.a(\dpath.a_lt_b$in1[7] ),
    .b(\dpath.a_lt_b$in1[6] ),
    .c(\dpath.a_lt_b$in1[5] ),
    .d(\dpath.a_lt_b$in1[4] ),
    .o1(_041_));
 b15nor004ah1n03x5 _316_ (.a(\dpath.a_lt_b$in1[0] ),
    .b(\dpath.a_lt_b$in1[3] ),
    .c(\dpath.a_lt_b$in1[2] ),
    .d(\dpath.a_lt_b$in1[1] ),
    .o1(_042_));
 b15nand04ah1n04x5 _317_ (.a(_039_),
    .b(_040_),
    .c(_041_),
    .d(_042_),
    .o1(_043_));
 b15inv040ah1n02x5 _318_ (.a(net34),
    .o1(_044_));
 b15nandp3ar1n02x5 _319_ (.a(_043_),
    .b(_044_),
    .c(\ctrl.state.out[2] ),
    .o1(_045_));
 b15ztpn00an1n08x5 PHY_11 ();
 b15ztpn00an1n08x5 PHY_10 ();
 b15nand03ar1n02x5 _322_ (.a(_044_),
    .b(net36),
    .c(net33),
    .o1(_048_));
 b15nand02ar1n02x5 _323_ (.a(_045_),
    .b(_048_),
    .o1(_002_));
 b15norp02ar1n48x5 _324_ (.a(\ctrl.state.out[2] ),
    .b(net36),
    .o1(_049_));
 b15and002ar1n02x5 _325_ (.a(_049_),
    .b(\ctrl.state.out[1] ),
    .o(net53));
 b15nand02an1n03x5 _326_ (.a(net53),
    .b(net35),
    .o1(_050_));
 b15inv040aq1n16x5 _327_ (.a(net36),
    .o1(_051_));
 b15ztpn00an1n08x5 PHY_9 ();
 b15oai112ah1n04x5 _329_ (.a(_050_),
    .b(_044_),
    .c(_051_),
    .d(net33),
    .o1(_000_));
 b15nandp3ar1n02x5 _330_ (.a(_050_),
    .b(_044_),
    .c(\ctrl.state.out[1] ),
    .o1(_053_));
 b15inv040ah1n02x5 _331_ (.a(\ctrl.state.out[2] ),
    .o1(_054_));
 b15oai013an1n02x5 _332_ (.a(_053_),
    .b(_043_),
    .c(net34),
    .d(_054_),
    .o1(_001_));
 b15nonb02as1n02x5 _333_ (.a(\dpath.a_lt_b$in0[14] ),
    .b(\dpath.a_lt_b$in1[14] ),
    .out0(_055_));
 b15inv000as1n02x5 _334_ (.a(\dpath.a_lt_b$in0[13] ),
    .o1(_056_));
 b15norp02as1n03x5 _335_ (.a(_056_),
    .b(\dpath.a_lt_b$in1[13] ),
    .o1(_057_));
 b15nonb02al1n03x5 _336_ (.a(\dpath.a_lt_b$in1[13] ),
    .b(\dpath.a_lt_b$in0[13] ),
    .out0(_058_));
 b15nor002al1n04x5 _337_ (.a(_058_),
    .b(_057_),
    .o1(_059_));
 b15inv000ah1n02x5 _338_ (.a(\dpath.a_lt_b$in0[12] ),
    .o1(_060_));
 b15norp02aq1n03x5 _339_ (.a(_060_),
    .b(\dpath.a_lt_b$in1[12] ),
    .o1(_061_));
 b15ao0012as1n02x5 _340_ (.a(_057_),
    .b(_059_),
    .c(_061_),
    .o(_062_));
 b15inv000as1n02x5 _341_ (.a(\dpath.a_lt_b$in0[9] ),
    .o1(_063_));
 b15norp02as1n02x5 _342_ (.a(_063_),
    .b(\dpath.a_lt_b$in1[9] ),
    .o1(_064_));
 b15inv040ah1n02x5 _343_ (.a(_064_),
    .o1(_065_));
 b15nonb02an1n03x5 _344_ (.a(\dpath.a_lt_b$in1[9] ),
    .b(\dpath.a_lt_b$in0[9] ),
    .out0(_066_));
 b15inv040ah1n02x5 _345_ (.a(\dpath.a_lt_b$in1[8] ),
    .o1(_067_));
 b15nand02aq1n04x5 _346_ (.a(_067_),
    .b(\dpath.a_lt_b$in0[8] ),
    .o1(_068_));
 b15oai012al1n04x5 _347_ (.a(_065_),
    .b(_066_),
    .c(_068_),
    .o1(_069_));
 b15inv000as1n02x5 _348_ (.a(\dpath.a_lt_b$in0[10] ),
    .o1(_070_));
 b15nandp2al1n03x5 _349_ (.a(_070_),
    .b(\dpath.a_lt_b$in1[10] ),
    .o1(_071_));
 b15inv000as1n02x5 _350_ (.a(\dpath.a_lt_b$in1[10] ),
    .o1(_072_));
 b15nandp2al1n02x5 _351_ (.a(_072_),
    .b(\dpath.a_lt_b$in0[10] ),
    .o1(_073_));
 b15nandp2ar1n02x5 _352_ (.a(_071_),
    .b(_073_),
    .o1(_074_));
 b15inv040ah1n03x5 _353_ (.a(_074_),
    .o1(_075_));
 b15nonb02aq1n02x5 _354_ (.a(\dpath.a_lt_b$in1[11] ),
    .b(\dpath.a_lt_b$in0[11] ),
    .out0(_076_));
 b15inv040ah1n02x5 _355_ (.a(\dpath.a_lt_b$in0[11] ),
    .o1(_077_));
 b15norp02aq1n03x5 _356_ (.a(_077_),
    .b(\dpath.a_lt_b$in1[11] ),
    .o1(_078_));
 b15norp02an1n04x5 _357_ (.a(_076_),
    .b(_078_),
    .o1(_079_));
 b15nandp3aq1n02x5 _358_ (.a(_069_),
    .b(_075_),
    .c(_079_),
    .o1(_080_));
 b15inv000ah1n02x5 _359_ (.a(_076_),
    .o1(_081_));
 b15inv000an1n02x5 _360_ (.a(_073_),
    .o1(_082_));
 b15aoi012ar1n02x5 _361_ (.a(_078_),
    .b(_081_),
    .c(_082_),
    .o1(_083_));
 b15nand02an1n03x5 _362_ (.a(_080_),
    .b(_083_),
    .o1(_084_));
 b15inv040ah1n02x5 _363_ (.a(\dpath.a_lt_b$in0[7] ),
    .o1(_085_));
 b15norp02aq1n03x5 _364_ (.a(_085_),
    .b(\dpath.a_lt_b$in1[7] ),
    .o1(_086_));
 b15inv000ah1n02x5 _365_ (.a(\dpath.a_lt_b$in0[6] ),
    .o1(_087_));
 b15norp02aq1n02x5 _366_ (.a(_087_),
    .b(\dpath.a_lt_b$in1[6] ),
    .o1(_088_));
 b15nandp2ar1n03x5 _367_ (.a(_085_),
    .b(\dpath.a_lt_b$in1[7] ),
    .o1(_089_));
 b15aoi012as1n02x5 _368_ (.a(_086_),
    .b(_088_),
    .c(_089_),
    .o1(_090_));
 b15nonb02al1n02x5 _369_ (.a(\dpath.a_lt_b$in1[7] ),
    .b(\dpath.a_lt_b$in0[7] ),
    .out0(_091_));
 b15norp02al1n02x5 _370_ (.a(_091_),
    .b(_086_),
    .o1(_092_));
 b15xor002al1n04x5 _371_ (.a(\dpath.a_lt_b$in0[6] ),
    .b(\dpath.a_lt_b$in1[6] ),
    .out0(_093_));
 b15inv040ah1n03x5 _372_ (.a(_093_),
    .o1(_094_));
 b15nandp2aq1n04x5 _373_ (.a(_092_),
    .b(_094_),
    .o1(_095_));
 b15inv000as1n02x5 _374_ (.a(\dpath.a_lt_b$in1[5] ),
    .o1(_096_));
 b15nand02aq1n04x5 _375_ (.a(_096_),
    .b(\dpath.a_lt_b$in0[5] ),
    .o1(_097_));
 b15inv000as1n02x5 _376_ (.a(_097_),
    .o1(_098_));
 b15inv000ah1n02x5 _377_ (.a(\dpath.a_lt_b$in0[4] ),
    .o1(_099_));
 b15norp02as1n03x5 _378_ (.a(_099_),
    .b(\dpath.a_lt_b$in1[4] ),
    .o1(_100_));
 b15inv000as1n02x5 _379_ (.a(\dpath.a_lt_b$in0[5] ),
    .o1(_101_));
 b15nandp2aq1n04x5 _380_ (.a(_101_),
    .b(\dpath.a_lt_b$in1[5] ),
    .o1(_102_));
 b15aoi012ar1n04x5 _381_ (.a(_098_),
    .b(_100_),
    .c(_102_),
    .o1(_103_));
 b15oai012ar1n12x5 _382_ (.a(_090_),
    .b(_095_),
    .c(_103_),
    .o1(_104_));
 b15inv000an1n05x5 _383_ (.a(\dpath.a_lt_b$in1[3] ),
    .o1(_105_));
 b15inv040as1n02x5 _384_ (.a(\dpath.a_lt_b$in0[2] ),
    .o1(_106_));
 b15nor002an1n04x5 _385_ (.a(_106_),
    .b(\dpath.a_lt_b$in1[2] ),
    .o1(_107_));
 b15rm6013en1n12x5 _386_ (.a(\dpath.a_lt_b$in0[3] ),
    .b(_105_),
    .c(_107_),
    .carryb(_108_));
 b15inv040ah1n02x5 _387_ (.a(\dpath.a_lt_b$in0[1] ),
    .o1(_109_));
 b15nor002ah1n06x5 _388_ (.a(_109_),
    .b(\dpath.a_lt_b$in1[1] ),
    .o1(_110_));
 b15nand02as1n03x5 _389_ (.a(_109_),
    .b(\dpath.a_lt_b$in1[1] ),
    .o1(_111_));
 b15aoi012ar1n08x5 _390_ (.a(_110_),
    .b(_036_),
    .c(_111_),
    .o1(_112_));
 b15inv040ah1n02x5 _391_ (.a(\dpath.a_lt_b$in0[3] ),
    .o1(_113_));
 b15xor002ar1n08x5 _392_ (.a(_113_),
    .b(\dpath.a_lt_b$in1[3] ),
    .out0(_114_));
 b15xor002as1n02x5 _393_ (.a(_106_),
    .b(\dpath.a_lt_b$in1[2] ),
    .out0(_115_));
 b15nandp2an1n08x5 _394_ (.a(_114_),
    .b(_115_),
    .o1(_116_));
 b15oai012as1n12x5 _395_ (.a(_108_),
    .b(_112_),
    .c(_116_),
    .o1(_117_));
 b15inv040ah1n02x5 _396_ (.a(_086_),
    .o1(_118_));
 b15nandp2aq1n03x5 _397_ (.a(_118_),
    .b(_089_),
    .o1(_119_));
 b15norp02ar1n02x5 _398_ (.a(_119_),
    .b(_093_),
    .o1(_120_));
 b15nandp2aq1n04x5 _399_ (.a(_099_),
    .b(\dpath.a_lt_b$in1[4] ),
    .o1(_121_));
 b15inv000al1n02x5 _400_ (.a(\dpath.a_lt_b$in1[4] ),
    .o1(_122_));
 b15nand02ar1n02x5 _401_ (.a(_122_),
    .b(\dpath.a_lt_b$in0[4] ),
    .o1(_123_));
 b15nand02as1n03x5 _402_ (.a(_121_),
    .b(_123_),
    .o1(_124_));
 b15nand02al1n02x5 _403_ (.a(_102_),
    .b(_097_),
    .o1(_125_));
 b15norp02an1n02x5 _404_ (.a(_124_),
    .b(_125_),
    .o1(_126_));
 b15nand02an1n04x5 _405_ (.a(_120_),
    .b(_126_),
    .o1(_127_));
 b15inv020as1n05x5 _406_ (.a(_127_),
    .o1(_128_));
 b15aoi012an1n08x5 _407_ (.a(_104_),
    .b(_117_),
    .c(_128_),
    .o1(_129_));
 b15nand02ah1n03x5 _408_ (.a(_075_),
    .b(_079_),
    .o1(_130_));
 b15inv000as1n02x5 _409_ (.a(_068_),
    .o1(_131_));
 b15norp02ar1n04x5 _410_ (.a(_067_),
    .b(\dpath.a_lt_b$in0[8] ),
    .o1(_132_));
 b15norp02aq1n02x5 _411_ (.a(_131_),
    .b(_132_),
    .o1(_133_));
 b15norp02an1n04x5 _412_ (.a(_066_),
    .b(_064_),
    .o1(_134_));
 b15nand02al1n04x5 _413_ (.a(_133_),
    .b(_134_),
    .o1(_135_));
 b15nor002as1n04x5 _414_ (.a(_130_),
    .b(_135_),
    .o1(_136_));
 b15inv000aq1n02x5 _415_ (.a(_136_),
    .o1(_137_));
 b15oabi12aq1n06x5 _416_ (.a(_084_),
    .b(_129_),
    .c(_137_),
    .out0(_138_));
 b15and002al1n02x5 _417_ (.a(_060_),
    .b(\dpath.a_lt_b$in1[12] ),
    .o(_139_));
 b15nor002as1n02x5 _418_ (.a(_139_),
    .b(_061_),
    .o1(_140_));
 b15nand02as1n03x5 _419_ (.a(_140_),
    .b(_059_),
    .o1(_141_));
 b15inv000al1n02x5 _420_ (.a(_141_),
    .o1(_142_));
 b15aoi012al1n06x5 _421_ (.a(_062_),
    .b(_138_),
    .c(_142_),
    .o1(_143_));
 b15nonb02aq1n03x5 _422_ (.a(\dpath.a_lt_b$in1[14] ),
    .b(\dpath.a_lt_b$in0[14] ),
    .out0(_144_));
 b15oabi12ar1n02x5 _423_ (.a(_055_),
    .b(_143_),
    .c(_144_),
    .out0(_145_));
 b15inv040ah1n02x5 _424_ (.a(\dpath.a_lt_b$in0[15] ),
    .o1(_146_));
 b15and002aq1n02x5 _425_ (.a(_146_),
    .b(\dpath.a_lt_b$in1[15] ),
    .o(_147_));
 b15norp02ar1n02x5 _426_ (.a(_146_),
    .b(\dpath.a_lt_b$in1[15] ),
    .o1(_148_));
 b15nor002as1n03x5 _427_ (.a(_147_),
    .b(_148_),
    .o1(_149_));
 b15nand02ar1n02x5 _428_ (.a(_145_),
    .b(_149_),
    .o1(_150_));
 b15nor002aq1n04x5 _429_ (.a(_055_),
    .b(_144_),
    .o1(_151_));
 b15inv000aq1n02x5 _430_ (.a(_110_),
    .o1(_152_));
 b15norp02ar1n02x5 _431_ (.a(_037_),
    .b(\dpath.a_lt_b$in0[0] ),
    .o1(_153_));
 b15inv040ah1n02x5 _432_ (.a(\dpath.a_lt_b$in1[1] ),
    .o1(_154_));
 b15nor002al1n06x5 _433_ (.a(_154_),
    .b(\dpath.a_lt_b$in0[1] ),
    .o1(_155_));
 b15oai012as1n02x5 _434_ (.a(_152_),
    .b(_153_),
    .c(_155_),
    .o1(_156_));
 b15nand02ah1n02x5 _435_ (.a(_113_),
    .b(\dpath.a_lt_b$in1[3] ),
    .o1(_157_));
 b15nand02ar1n02x5 _436_ (.a(_105_),
    .b(\dpath.a_lt_b$in0[3] ),
    .o1(_158_));
 b15nandp2ar1n03x5 _437_ (.a(_157_),
    .b(_158_),
    .o1(_159_));
 b15xor002as1n02x5 _438_ (.a(\dpath.a_lt_b$in0[2] ),
    .b(\dpath.a_lt_b$in1[2] ),
    .out0(_160_));
 b15norp02ar1n02x5 _439_ (.a(_159_),
    .b(_160_),
    .o1(_161_));
 b15nand02ar1n02x5 _440_ (.a(_156_),
    .b(_161_),
    .o1(_162_));
 b15aoi012aq1n02x5 _441_ (.a(_127_),
    .b(_162_),
    .c(_108_),
    .o1(_163_));
 b15oai012an1n02x5 _442_ (.a(_136_),
    .b(_163_),
    .c(_104_),
    .o1(_164_));
 b15inv000al1n02x5 _443_ (.a(_084_),
    .o1(_165_));
 b15aoi012al1n02x5 _444_ (.a(_141_),
    .b(_164_),
    .c(_165_),
    .o1(_166_));
 b15oai012ar1n02x5 _445_ (.a(_151_),
    .b(_166_),
    .c(_062_),
    .o1(_167_));
 b15nona22ar1n02x5 _446_ (.a(_149_),
    .b(_055_),
    .c(_167_),
    .out0(_168_));
 b15and002ar1n02x5 _447_ (.a(_150_),
    .b(_168_),
    .o(net43));
 b15norp02an1n02x5 _448_ (.a(_110_),
    .b(_155_),
    .o1(_169_));
 b15xor002ar1n04x5 _449_ (.a(_169_),
    .b(_036_),
    .out0(net44));
 b15xor002an1n02x5 _450_ (.a(_112_),
    .b(_160_),
    .out0(net45));
 b15aoi012aq1n02x5 _451_ (.a(_107_),
    .b(_156_),
    .c(_115_),
    .o1(_170_));
 b15xor002aq1n03x5 _452_ (.a(_170_),
    .b(_159_),
    .out0(net46));
 b15xnr002ah1n02x5 _453_ (.a(_117_),
    .b(_124_),
    .out0(net47));
 b15aoi012ar1n04x5 _454_ (.a(_100_),
    .b(_117_),
    .c(_121_),
    .o1(_171_));
 b15xor002aq1n02x5 _455_ (.a(_171_),
    .b(_125_),
    .out0(net48));
 b15inv000al1n02x5 _456_ (.a(_102_),
    .o1(_172_));
 b15oai012as1n04x5 _457_ (.a(_097_),
    .b(_171_),
    .c(_172_),
    .o1(_173_));
 b15xor002an1n03x5 _458_ (.a(_173_),
    .b(_094_),
    .out0(net49));
 b15aoi012al1n02x5 _459_ (.a(_088_),
    .b(_173_),
    .c(_094_),
    .o1(_174_));
 b15xor002an1n04x5 _460_ (.a(_174_),
    .b(_119_),
    .out0(net50));
 b15inv000al1n02x5 _461_ (.a(_133_),
    .o1(_175_));
 b15xor002an1n04x5 _462_ (.a(_129_),
    .b(_175_),
    .out0(net51));
 b15oai012an1n02x5 _463_ (.a(_068_),
    .b(_129_),
    .c(_132_),
    .o1(_176_));
 b15xor002al1n03x5 _464_ (.a(_176_),
    .b(_134_),
    .out0(net52));
 b15oabi12an1n02x5 _465_ (.a(_069_),
    .b(_129_),
    .c(_135_),
    .out0(_177_));
 b15and002an1n02x5 _466_ (.a(_177_),
    .b(_075_),
    .o(_178_));
 b15norp02ar1n02x5 _467_ (.a(_177_),
    .b(_075_),
    .o1(_179_));
 b15norp02ar1n03x5 _468_ (.a(_178_),
    .b(_179_),
    .o1(net38));
 b15oai012ar1n02x5 _469_ (.a(_079_),
    .b(_178_),
    .c(_082_),
    .o1(_180_));
 b15norp03ar1n02x5 _470_ (.a(_178_),
    .b(_082_),
    .c(_079_),
    .o1(_181_));
 b15nonb02ar1n02x5 _471_ (.a(_180_),
    .b(_181_),
    .out0(net39));
 b15and002ar1n02x5 _472_ (.a(_138_),
    .b(_140_),
    .o(_182_));
 b15norp02ar1n02x5 _473_ (.a(_138_),
    .b(_140_),
    .o1(_183_));
 b15norp02al1n02x5 _474_ (.a(_182_),
    .b(_183_),
    .o1(net40));
 b15orn002ar1n02x5 _475_ (.a(_182_),
    .b(_061_),
    .o(_184_));
 b15xor002al1n02x5 _476_ (.a(_184_),
    .b(_059_),
    .out0(net41));
 b15xnr002an1n06x5 _477_ (.a(_143_),
    .b(_151_),
    .out0(net42));
 b15nand02ah1n03x5 _478_ (.a(_149_),
    .b(_151_),
    .o1(_185_));
 b15norp02aq1n04x5 _479_ (.a(_141_),
    .b(_185_),
    .o1(_186_));
 b15oai012ar1n02x5 _480_ (.a(_065_),
    .b(_066_),
    .c(_132_),
    .o1(_187_));
 b15norp02al1n02x5 _481_ (.a(_130_),
    .b(_187_),
    .o1(_188_));
 b15aoi012ar1n02x5 _482_ (.a(_078_),
    .b(_081_),
    .c(_071_),
    .o1(_189_));
 b15oai012ar1n02x5 _483_ (.a(_186_),
    .b(_188_),
    .c(_189_),
    .o1(_190_));
 b15norp02ar1n02x5 _484_ (.a(_139_),
    .b(_058_),
    .o1(_191_));
 b15orn003ar1n02x5 _485_ (.a(_185_),
    .b(_057_),
    .c(_191_),
    .o(_192_));
 b15aoi012ah1n02x5 _486_ (.a(_147_),
    .b(_149_),
    .c(_144_),
    .o1(_193_));
 b15and003al1n02x5 _487_ (.a(_190_),
    .b(_192_),
    .c(_193_),
    .o(_194_));
 b15aoai13al1n02x5 _488_ (.a(_118_),
    .b(_091_),
    .c(_087_),
    .d(\dpath.a_lt_b$in1[6] ),
    .o1(_195_));
 b15and002ar1n02x5 _489_ (.a(_121_),
    .b(_102_),
    .o(_196_));
 b15oai013an1n04x5 _490_ (.a(_195_),
    .b(_095_),
    .c(_098_),
    .d(_196_),
    .o1(_197_));
 b15nandp3an1n02x5 _491_ (.a(_114_),
    .b(_106_),
    .c(\dpath.a_lt_b$in1[2] ),
    .o1(_198_));
 b15oai012ar1n03x5 _492_ (.a(_152_),
    .b(_155_),
    .c(_038_),
    .o1(_199_));
 b15oai112ah1n04x5 _493_ (.a(_157_),
    .b(_198_),
    .c(_199_),
    .d(_116_),
    .o1(_200_));
 b15aoi012al1n04x5 _494_ (.a(_197_),
    .b(_200_),
    .c(_128_),
    .o1(_201_));
 b15nand02an1n02x5 _495_ (.a(_186_),
    .b(_136_),
    .o1(_202_));
 b15oai012ar1n08x5 _496_ (.a(_194_),
    .b(_201_),
    .c(_202_),
    .o1(_203_));
 b15nor004ar1n08x5 _497_ (.a(_116_),
    .b(net37),
    .c(_110_),
    .d(_155_),
    .o1(_204_));
 b15nand04as1n06x5 _498_ (.a(_204_),
    .b(_128_),
    .c(_186_),
    .d(_136_),
    .o1(_205_));
 b15nandp2an1n16x5 _499_ (.a(_203_),
    .b(_205_),
    .o1(_206_));
 b15nor002aq1n03x5 _500_ (.a(_054_),
    .b(net36),
    .o1(_207_));
 b15inv040al1n12x5 _501_ (.a(_207_),
    .o1(_208_));
 b15norp02aq1n48x5 _502_ (.a(_206_),
    .b(_208_),
    .o1(_209_));
 b15ztpn00an1n08x5 PHY_8 ();
 b15aoi022ar1n02x5 _504_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[0] ),
    .c(net36),
    .d(net1),
    .o1(_211_));
 b15cinv00ah1n12x5 _505_ (.clk(_206_),
    .clkout(_212_));
 b15nand02an1n32x5 _506_ (.a(_212_),
    .b(\ctrl.state.out[2] ),
    .o1(_213_));
 b15ztpn00an1n08x5 PHY_7 ();
 b15nandp3ar1n02x5 _508_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[0] ),
    .c(_051_),
    .o1(_215_));
 b15nandp2aq1n02x5 _509_ (.a(_211_),
    .b(_215_),
    .o1(_003_));
 b15aoi022ar1n02x5 _510_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[1] ),
    .c(net36),
    .d(net12),
    .o1(_216_));
 b15nandp3ar1n02x5 _511_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[1] ),
    .c(_051_),
    .o1(_217_));
 b15nand02as1n02x5 _512_ (.a(_216_),
    .b(_217_),
    .o1(_004_));
 b15aoi022ar1n02x5 _513_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[2] ),
    .c(net36),
    .d(net23),
    .o1(_218_));
 b15nandp3ar1n02x5 _514_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[2] ),
    .c(_051_),
    .o1(_219_));
 b15nandp2aq1n02x5 _515_ (.a(_218_),
    .b(_219_),
    .o1(_005_));
 b15aoi022ar1n02x5 _516_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[3] ),
    .c(net36),
    .d(net26),
    .o1(_220_));
 b15nandp3ar1n02x5 _517_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[3] ),
    .c(_051_),
    .o1(_221_));
 b15nand02ar1n02x5 _518_ (.a(_220_),
    .b(_221_),
    .o1(_006_));
 b15ztpn00an1n08x5 PHY_6 ();
 b15nandp2aq1n02x5 _520_ (.a(_099_),
    .b(_051_),
    .o1(_223_));
 b15oai012ar1n02x5 _521_ (.a(_223_),
    .b(_051_),
    .c(net27),
    .o1(_224_));
 b15aoi012ar1n02x5 _522_ (.a(_224_),
    .b(_213_),
    .c(_051_),
    .o1(_225_));
 b15nandp3ar1n02x5 _523_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[4] ),
    .c(_051_),
    .o1(_226_));
 b15nanb02ar1n02x5 _524_ (.a(_225_),
    .b(_226_),
    .out0(_007_));
 b15aoi022ar1n02x5 _525_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[5] ),
    .c(net36),
    .d(net28),
    .o1(_227_));
 b15nandp3ar1n02x5 _526_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[5] ),
    .c(_051_),
    .o1(_228_));
 b15nand02ar1n02x5 _527_ (.a(_227_),
    .b(_228_),
    .o1(_008_));
 b15aoi022ar1n02x5 _528_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[6] ),
    .c(net36),
    .d(net29),
    .o1(_229_));
 b15nandp3ar1n02x5 _529_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[6] ),
    .c(_051_),
    .o1(_230_));
 b15nand02ar1n02x5 _530_ (.a(_229_),
    .b(_230_),
    .o1(_009_));
 b15aoi022ar1n02x5 _531_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[7] ),
    .c(net36),
    .d(net30),
    .o1(_231_));
 b15nandp3ar1n02x5 _532_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[7] ),
    .c(_051_),
    .o1(_232_));
 b15nand02ar1n02x5 _533_ (.a(_231_),
    .b(_232_),
    .o1(_010_));
 b15aoi022ar1n02x5 _534_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[8] ),
    .c(net36),
    .d(net31),
    .o1(_233_));
 b15nandp3ar1n02x5 _535_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[8] ),
    .c(_051_),
    .o1(_234_));
 b15nand02an1n02x5 _536_ (.a(_233_),
    .b(_234_),
    .o1(_011_));
 b15aoi022ar1n02x5 _537_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[9] ),
    .c(net36),
    .d(net32),
    .o1(_235_));
 b15nandp3ar1n02x5 _538_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[9] ),
    .c(_051_),
    .o1(_236_));
 b15nandp2al1n02x5 _539_ (.a(_235_),
    .b(_236_),
    .o1(_012_));
 b15ztpn00an1n08x5 PHY_5 ();
 b15aoi022ar1n02x5 _541_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[10] ),
    .c(net36),
    .d(net2),
    .o1(_238_));
 b15nandp3ar1n02x5 _542_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[10] ),
    .c(_051_),
    .o1(_239_));
 b15nandp2ar1n02x5 _543_ (.a(_238_),
    .b(_239_),
    .o1(_013_));
 b15ztpn00an1n08x5 PHY_4 ();
 b15aoi022ar1n02x5 _545_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[11] ),
    .c(net36),
    .d(net3),
    .o1(_241_));
 b15nandp3ar1n02x5 _546_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[11] ),
    .c(_051_),
    .o1(_242_));
 b15nand02ar1n02x5 _547_ (.a(_241_),
    .b(_242_),
    .o1(_014_));
 b15aoi022ar1n02x5 _548_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[12] ),
    .c(net36),
    .d(net4),
    .o1(_243_));
 b15nandp3ar1n02x5 _549_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[12] ),
    .c(_051_),
    .o1(_244_));
 b15nand02ar1n02x5 _550_ (.a(_243_),
    .b(_244_),
    .o1(_015_));
 b15aoi022an1n04x5 _551_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[13] ),
    .c(net36),
    .d(net5),
    .o1(_245_));
 b15nandp3ar1n02x5 _552_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[13] ),
    .c(_051_),
    .o1(_246_));
 b15nand02ar1n02x5 _553_ (.a(_245_),
    .b(_246_),
    .o1(_016_));
 b15aoi022ar1n02x5 _554_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[14] ),
    .c(net36),
    .d(net6),
    .o1(_247_));
 b15nandp3ar1n02x5 _555_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[14] ),
    .c(_051_),
    .o1(_248_));
 b15nand02ar1n02x5 _556_ (.a(_247_),
    .b(_248_),
    .o1(_017_));
 b15aoi022ar1n02x5 _557_ (.a(_209_),
    .b(\dpath.a_lt_b$in0[15] ),
    .c(net36),
    .d(net7),
    .o1(_249_));
 b15nandp3ar1n02x5 _558_ (.a(_213_),
    .b(\dpath.a_lt_b$in1[15] ),
    .c(_051_),
    .o1(_250_));
 b15nand02ar1n02x5 _559_ (.a(_249_),
    .b(_250_),
    .o1(_018_));
 b15nor002as1n24x5 _560_ (.a(_212_),
    .b(_208_),
    .o1(_251_));
 b15ztpn00an1n08x5 PHY_3 ();
 b15nand02ar1n02x5 _562_ (.a(_251_),
    .b(net37),
    .o1(_253_));
 b15nand02ar1n02x5 _563_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[0] ),
    .o1(_254_));
 b15ztpn00an1n08x5 PHY_2 ();
 b15aoi022ar1n02x5 _565_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[0] ),
    .c(net36),
    .d(net8),
    .o1(_256_));
 b15nand03ah1n03x5 _566_ (.a(_253_),
    .b(_254_),
    .c(_256_),
    .o1(_019_));
 b15nand02ar1n02x5 _567_ (.a(_251_),
    .b(net44),
    .o1(_257_));
 b15nand02ar1n02x5 _568_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[1] ),
    .o1(_258_));
 b15aoi022ar1n02x5 _569_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[1] ),
    .c(net36),
    .d(net9),
    .o1(_259_));
 b15nandp3ar1n04x5 _570_ (.a(_257_),
    .b(_258_),
    .c(_259_),
    .o1(_020_));
 b15nand02ar1n02x5 _571_ (.a(_251_),
    .b(net45),
    .o1(_260_));
 b15ztpn00an1n08x5 PHY_1 ();
 b15nand02ar1n02x5 _573_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[2] ),
    .o1(_262_));
 b15aoi022ar1n02x5 _574_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[2] ),
    .c(net36),
    .d(net10),
    .o1(_263_));
 b15nand03ar1n04x5 _575_ (.a(_260_),
    .b(_262_),
    .c(_263_),
    .o1(_021_));
 b15nand02ar1n02x5 _576_ (.a(_251_),
    .b(net46),
    .o1(_264_));
 b15nand02ar1n02x5 _577_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[3] ),
    .o1(_265_));
 b15aoi022ar1n02x5 _578_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[3] ),
    .c(net36),
    .d(net11),
    .o1(_266_));
 b15nandp3ar1n02x5 _579_ (.a(_264_),
    .b(_265_),
    .c(_266_),
    .o1(_022_));
 b15nand02ar1n02x5 _580_ (.a(_251_),
    .b(net47),
    .o1(_267_));
 b15nand02ar1n02x5 _581_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[4] ),
    .o1(_268_));
 b15ztpn00an1n08x5 PHY_0 ();
 b15aoai13ar1n02x5 _583_ (.a(_223_),
    .b(_049_),
    .c(net36),
    .d(net13),
    .o1(_270_));
 b15nandp3ar1n02x5 _584_ (.a(_267_),
    .b(_268_),
    .c(_270_),
    .o1(_023_));
 b15nand02ar1n02x5 _585_ (.a(_251_),
    .b(net48),
    .o1(_271_));
 b15nand02ar1n02x5 _586_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[5] ),
    .o1(_272_));
 b15aoi022ar1n02x5 _587_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[5] ),
    .c(net36),
    .d(net14),
    .o1(_273_));
 b15nandp3ar1n02x5 _588_ (.a(_271_),
    .b(_272_),
    .c(_273_),
    .o1(_024_));
 b15nand02ar1n02x5 _589_ (.a(_251_),
    .b(net49),
    .o1(_274_));
 b15nand02ar1n02x5 _590_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[6] ),
    .o1(_275_));
 b15aoi022ar1n02x5 _591_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[6] ),
    .c(net36),
    .d(net15),
    .o1(_276_));
 b15nandp3ar1n02x5 _592_ (.a(_274_),
    .b(_275_),
    .c(_276_),
    .o1(_025_));
 b15nand02ar1n02x5 _593_ (.a(_251_),
    .b(net50),
    .o1(_277_));
 b15nand02ar1n02x5 _594_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[7] ),
    .o1(_278_));
 b15aoi022ar1n02x5 _595_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[7] ),
    .c(net36),
    .d(net16),
    .o1(_279_));
 b15nandp3ar1n02x5 _596_ (.a(_277_),
    .b(_278_),
    .c(_279_),
    .o1(_026_));
 b15nand02ar1n02x5 _597_ (.a(_251_),
    .b(net51),
    .o1(_280_));
 b15nand02ar1n02x5 _598_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[8] ),
    .o1(_281_));
 b15aoi022ar1n02x5 _599_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[8] ),
    .c(net36),
    .d(net17),
    .o1(_282_));
 b15nand03al1n04x5 _600_ (.a(_280_),
    .b(_281_),
    .c(_282_),
    .o1(_027_));
 b15nand02ar1n02x5 _601_ (.a(_251_),
    .b(net52),
    .o1(_283_));
 b15nand02ar1n02x5 _602_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[9] ),
    .o1(_284_));
 b15aoi022ar1n02x5 _603_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[9] ),
    .c(net36),
    .d(net18),
    .o1(_285_));
 b15nandp3as1n02x5 _604_ (.a(_283_),
    .b(_284_),
    .c(_285_),
    .o1(_028_));
 b15nand02ar1n02x5 _605_ (.a(_251_),
    .b(net38),
    .o1(_286_));
 b15nand02ar1n02x5 _606_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[10] ),
    .o1(_287_));
 b15aoi022ar1n02x5 _607_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[10] ),
    .c(net36),
    .d(net19),
    .o1(_288_));
 b15nandp3al1n03x5 _608_ (.a(_286_),
    .b(_287_),
    .c(_288_),
    .o1(_029_));
 b15nand02ar1n02x5 _609_ (.a(net39),
    .b(_251_),
    .o1(_289_));
 b15nand02ar1n02x5 _610_ (.a(net36),
    .b(net20),
    .o1(_290_));
 b15inv040ah1n02x5 _611_ (.a(_049_),
    .o1(_291_));
 b15oai012ar1n02x5 _612_ (.a(_290_),
    .b(_291_),
    .c(_077_),
    .o1(_292_));
 b15aoi012ar1n02x5 _613_ (.a(_292_),
    .b(_209_),
    .c(\dpath.a_lt_b$in1[11] ),
    .o1(_293_));
 b15nandp2ah1n02x5 _614_ (.a(_289_),
    .b(_293_),
    .o1(_030_));
 b15nand02al1n02x5 _615_ (.a(_251_),
    .b(net40),
    .o1(_294_));
 b15nand02ar1n02x5 _616_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[12] ),
    .o1(_295_));
 b15aoi022ar1n02x5 _617_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[12] ),
    .c(net36),
    .d(net21),
    .o1(_296_));
 b15nandp3ar1n02x5 _618_ (.a(_294_),
    .b(_295_),
    .c(_296_),
    .o1(_031_));
 b15nand02ar1n02x5 _619_ (.a(net41),
    .b(_251_),
    .o1(_297_));
 b15nand02ar1n02x5 _620_ (.a(net36),
    .b(net22),
    .o1(_298_));
 b15oai012ar1n02x5 _621_ (.a(_298_),
    .b(_291_),
    .c(_056_),
    .o1(_299_));
 b15aoi012ar1n02x5 _622_ (.a(_299_),
    .b(_209_),
    .c(\dpath.a_lt_b$in1[13] ),
    .o1(_300_));
 b15nandp2ar1n03x5 _623_ (.a(_297_),
    .b(_300_),
    .o1(_032_));
 b15nand02ar1n02x5 _624_ (.a(_251_),
    .b(net42),
    .o1(_301_));
 b15nand02ar1n02x5 _625_ (.a(_209_),
    .b(\dpath.a_lt_b$in1[14] ),
    .o1(_302_));
 b15aoi022ar1n02x5 _626_ (.a(_049_),
    .b(\dpath.a_lt_b$in0[14] ),
    .c(net36),
    .d(net24),
    .o1(_303_));
 b15nandp3ar1n02x5 _627_ (.a(_301_),
    .b(_302_),
    .c(_303_),
    .o1(_033_));
 b15nandp3ar1n02x5 _628_ (.a(_150_),
    .b(_168_),
    .c(_251_),
    .o1(_304_));
 b15nand02ar1n02x5 _629_ (.a(net36),
    .b(net25),
    .o1(_305_));
 b15oai012ar1n02x5 _630_ (.a(_305_),
    .b(_291_),
    .c(_146_),
    .o1(_306_));
 b15aoi012ar1n02x5 _631_ (.a(_306_),
    .b(_209_),
    .c(\dpath.a_lt_b$in1[15] ),
    .o1(_307_));
 b15nandp2ar1n02x5 _632_ (.a(_304_),
    .b(_307_),
    .o1(_034_));
 b15fpn000hn1n04x5 _633_ (.clk(clknet_2_1__leaf_clk),
    .d(_000_),
    .o(net36));
 b15fpn000hn1n04x5 _634_ (.clk(clknet_2_1__leaf_clk),
    .d(_001_),
    .o(\ctrl.state.out[1] ));
 b15fpn000hn1n04x5 _635_ (.clk(clknet_2_1__leaf_clk),
    .d(_002_),
    .o(\ctrl.state.out[2] ));
 b15fpn000hn1n04x5 _636_ (.clk(clknet_2_0__leaf_clk),
    .d(_003_),
    .o(\dpath.a_lt_b$in1[0] ));
 b15fpn000hn1n04x5 _637_ (.clk(clknet_2_0__leaf_clk),
    .d(_004_),
    .o(\dpath.a_lt_b$in1[1] ));
 b15fpn000hn1n04x5 _638_ (.clk(clknet_2_0__leaf_clk),
    .d(_005_),
    .o(\dpath.a_lt_b$in1[2] ));
 b15fpn000hn1n04x5 _639_ (.clk(clknet_2_0__leaf_clk),
    .d(_006_),
    .o(\dpath.a_lt_b$in1[3] ));
 b15fpn000hn1n04x5 _640_ (.clk(clknet_2_2__leaf_clk),
    .d(_007_),
    .o(\dpath.a_lt_b$in1[4] ));
 b15fpn000hn1n04x5 _641_ (.clk(clknet_2_2__leaf_clk),
    .d(_008_),
    .o(\dpath.a_lt_b$in1[5] ));
 b15fpn000hn1n04x5 _642_ (.clk(clknet_2_3__leaf_clk),
    .d(_009_),
    .o(\dpath.a_lt_b$in1[6] ));
 b15fpn000hn1n04x5 _643_ (.clk(clknet_2_2__leaf_clk),
    .d(_010_),
    .o(\dpath.a_lt_b$in1[7] ));
 b15fpn000hn1n04x5 _644_ (.clk(clknet_2_1__leaf_clk),
    .d(_011_),
    .o(\dpath.a_lt_b$in1[8] ));
 b15fpn000hn1n04x5 _645_ (.clk(clknet_2_1__leaf_clk),
    .d(_012_),
    .o(\dpath.a_lt_b$in1[9] ));
 b15fpn000hn1n04x5 _646_ (.clk(clknet_2_1__leaf_clk),
    .d(_013_),
    .o(\dpath.a_lt_b$in1[10] ));
 b15fpn000hn1n04x5 _647_ (.clk(clknet_2_1__leaf_clk),
    .d(_014_),
    .o(\dpath.a_lt_b$in1[11] ));
 b15fpn000hn1n04x5 _648_ (.clk(clknet_2_3__leaf_clk),
    .d(_015_),
    .o(\dpath.a_lt_b$in1[12] ));
 b15fpn000hn1n04x5 _649_ (.clk(clknet_2_3__leaf_clk),
    .d(_016_),
    .o(\dpath.a_lt_b$in1[13] ));
 b15fpn000hn1n04x5 _650_ (.clk(clknet_2_3__leaf_clk),
    .d(_017_),
    .o(\dpath.a_lt_b$in1[14] ));
 b15fpn000hn1n04x5 _651_ (.clk(clknet_2_3__leaf_clk),
    .d(_018_),
    .o(\dpath.a_lt_b$in1[15] ));
 b15fpn000hn1n04x5 _652_ (.clk(clknet_2_0__leaf_clk),
    .d(_019_),
    .o(\dpath.a_lt_b$in0[0] ));
 b15fpn000hn1n04x5 _653_ (.clk(clknet_2_0__leaf_clk),
    .d(_020_),
    .o(\dpath.a_lt_b$in0[1] ));
 b15fpn000hn1n04x5 _654_ (.clk(clknet_2_0__leaf_clk),
    .d(_021_),
    .o(\dpath.a_lt_b$in0[2] ));
 b15fpn000hn1n04x5 _655_ (.clk(clknet_2_0__leaf_clk),
    .d(_022_),
    .o(\dpath.a_lt_b$in0[3] ));
 b15fpn000hn1n04x5 _656_ (.clk(clknet_2_2__leaf_clk),
    .d(_023_),
    .o(\dpath.a_lt_b$in0[4] ));
 b15fpn000hn1n04x5 _657_ (.clk(clknet_2_2__leaf_clk),
    .d(_024_),
    .o(\dpath.a_lt_b$in0[5] ));
 b15fpn000hn1n04x5 _658_ (.clk(clknet_2_3__leaf_clk),
    .d(_025_),
    .o(\dpath.a_lt_b$in0[6] ));
 b15fpn000hn1n04x5 _659_ (.clk(clknet_2_2__leaf_clk),
    .d(_026_),
    .o(\dpath.a_lt_b$in0[7] ));
 b15fpn000hn1n04x5 _660_ (.clk(clknet_2_1__leaf_clk),
    .d(_027_),
    .o(\dpath.a_lt_b$in0[8] ));
 b15fpn000hn1n04x5 _661_ (.clk(clknet_2_1__leaf_clk),
    .d(_028_),
    .o(\dpath.a_lt_b$in0[9] ));
 b15fpn000hn1n04x5 _662_ (.clk(clknet_2_1__leaf_clk),
    .d(_029_),
    .o(\dpath.a_lt_b$in0[10] ));
 b15fpn000hn1n04x5 _663_ (.clk(clknet_2_1__leaf_clk),
    .d(_030_),
    .o(\dpath.a_lt_b$in0[11] ));
 b15fpn000hn1n04x5 _664_ (.clk(clknet_2_1__leaf_clk),
    .d(_031_),
    .o(\dpath.a_lt_b$in0[12] ));
 b15fpn000hn1n04x5 _665_ (.clk(clknet_2_3__leaf_clk),
    .d(_032_),
    .o(\dpath.a_lt_b$in0[13] ));
 b15fpn000hn1n04x5 _666_ (.clk(clknet_2_3__leaf_clk),
    .d(_033_),
    .o(\dpath.a_lt_b$in0[14] ));
 b15fpn000hn1n04x5 _667_ (.clk(clknet_2_3__leaf_clk),
    .d(_034_),
    .o(\dpath.a_lt_b$in0[15] ));
 b15ztpn00an1n08x5 PHY_12 ();
 b15ztpn00an1n08x5 PHY_13 ();
 b15ztpn00an1n08x5 PHY_14 ();
 b15ztpn00an1n08x5 PHY_15 ();
 b15ztpn00an1n08x5 PHY_16 ();
 b15ztpn00an1n08x5 PHY_17 ();
 b15ztpn00an1n08x5 PHY_18 ();
 b15ztpn00an1n08x5 PHY_19 ();
 b15ztpn00an1n08x5 PHY_20 ();
 b15ztpn00an1n08x5 PHY_21 ();
 b15ztpn00an1n08x5 PHY_22 ();
 b15ztpn00an1n08x5 PHY_23 ();
 b15ztpn00an1n08x5 PHY_24 ();
 b15ztpn00an1n08x5 PHY_25 ();
 b15ztpn00an1n08x5 PHY_26 ();
 b15ztpn00an1n08x5 PHY_27 ();
 b15ztpn00an1n08x5 PHY_28 ();
 b15ztpn00an1n08x5 PHY_29 ();
 b15ztpn00an1n08x5 PHY_30 ();
 b15ztpn00an1n08x5 PHY_31 ();
 b15ztpn00an1n08x5 PHY_32 ();
 b15ztpn00an1n08x5 PHY_33 ();
 b15ztpn00an1n08x5 PHY_34 ();
 b15ztpn00an1n08x5 PHY_35 ();
 b15ztpn00an1n08x5 PHY_36 ();
 b15ztpn00an1n08x5 PHY_37 ();
 b15bfn000ar1n02x5 input1 (.a(req_msg[0]),
    .o(net1));
 b15bfn000al1n02x5 input2 (.a(req_msg[10]),
    .o(net2));
 b15bfn000al1n02x5 input3 (.a(req_msg[11]),
    .o(net3));
 b15bfn000al1n02x5 input4 (.a(req_msg[12]),
    .o(net4));
 b15bfn000ar1n02x5 input5 (.a(req_msg[13]),
    .o(net5));
 b15bfn000ar1n02x5 input6 (.a(req_msg[14]),
    .o(net6));
 b15bfn000ar1n02x5 input7 (.a(req_msg[15]),
    .o(net7));
 b15bfn000ar1n02x5 input8 (.a(req_msg[16]),
    .o(net8));
 b15bfn000ar1n02x5 input9 (.a(req_msg[17]),
    .o(net9));
 b15bfn000ar1n02x5 input10 (.a(req_msg[18]),
    .o(net10));
 b15bfn000ar1n02x5 input11 (.a(req_msg[19]),
    .o(net11));
 b15bfn000ar1n02x5 input12 (.a(req_msg[1]),
    .o(net12));
 b15bfn000ar1n02x5 input13 (.a(req_msg[20]),
    .o(net13));
 b15bfn000ar1n02x5 input14 (.a(req_msg[21]),
    .o(net14));
 b15bfn000ar1n02x5 input15 (.a(req_msg[22]),
    .o(net15));
 b15bfn000ar1n02x5 input16 (.a(req_msg[23]),
    .o(net16));
 b15bfn000ar1n02x5 input17 (.a(req_msg[24]),
    .o(net17));
 b15bfn000ar1n02x5 input18 (.a(req_msg[25]),
    .o(net18));
 b15bfn000ar1n02x5 input19 (.a(req_msg[26]),
    .o(net19));
 b15bfn000ar1n02x5 input20 (.a(req_msg[27]),
    .o(net20));
 b15bfn000ar1n02x5 input21 (.a(req_msg[28]),
    .o(net21));
 b15bfn000ar1n02x5 input22 (.a(req_msg[29]),
    .o(net22));
 b15bfn000ar1n02x5 input23 (.a(req_msg[2]),
    .o(net23));
 b15bfn000ar1n02x5 input24 (.a(req_msg[30]),
    .o(net24));
 b15bfn000ar1n02x5 input25 (.a(req_msg[31]),
    .o(net25));
 b15bfn000ar1n02x5 input26 (.a(req_msg[3]),
    .o(net26));
 b15bfn000ar1n02x5 input27 (.a(req_msg[4]),
    .o(net27));
 b15bfn000ar1n02x5 input28 (.a(req_msg[5]),
    .o(net28));
 b15bfn000ar1n02x5 input29 (.a(req_msg[6]),
    .o(net29));
 b15bfn000ar1n02x5 input30 (.a(req_msg[7]),
    .o(net30));
 b15bfn000ar1n02x5 input31 (.a(req_msg[8]),
    .o(net31));
 b15bfn000ar1n02x5 input32 (.a(req_msg[9]),
    .o(net32));
 b15bfn000aq1n02x5 input33 (.a(req_val),
    .o(net33));
 b15bfn000aq1n02x5 input34 (.a(reset),
    .o(net34));
 b15bfn000ar1n02x5 input35 (.a(resp_rdy),
    .o(net35));
 b15bfn000ar1n02x5 output36 (.a(net36),
    .o(req_rdy));
 b15bfn000ar1n02x5 output37 (.a(net37),
    .o(resp_msg[0]));
 b15bfn000ar1n02x5 output38 (.a(net38),
    .o(resp_msg[10]));
 b15bfn000ar1n02x5 output39 (.a(net39),
    .o(resp_msg[11]));
 b15bfn000ar1n02x5 output40 (.a(net40),
    .o(resp_msg[12]));
 b15bfn000ar1n02x5 output41 (.a(net41),
    .o(resp_msg[13]));
 b15bfn000ar1n02x5 output42 (.a(net42),
    .o(resp_msg[14]));
 b15bfn000ar1n02x5 output43 (.a(net43),
    .o(resp_msg[15]));
 b15bfn000ar1n02x5 output44 (.a(net44),
    .o(resp_msg[1]));
 b15bfn000ar1n02x5 output45 (.a(net45),
    .o(resp_msg[2]));
 b15bfn000ar1n02x5 output46 (.a(net46),
    .o(resp_msg[3]));
 b15bfn000ar1n02x5 output47 (.a(net47),
    .o(resp_msg[4]));
 b15bfn000ar1n02x5 output48 (.a(net48),
    .o(resp_msg[5]));
 b15bfn000ar1n02x5 output49 (.a(net49),
    .o(resp_msg[6]));
 b15bfn000ar1n02x5 output50 (.a(net50),
    .o(resp_msg[7]));
 b15bfn000ar1n02x5 output51 (.a(net51),
    .o(resp_msg[8]));
 b15bfn000ar1n02x5 output52 (.a(net52),
    .o(resp_msg[9]));
 b15bfn000ar1n02x5 output53 (.a(net53),
    .o(resp_val));
 b15cbf000an1n16x5 clkbuf_0_clk (.clk(clk),
    .clkout(clknet_0_clk));
 b15cbf000an1n16x5 clkbuf_2_0__f_clk (.clk(clknet_0_clk),
    .clkout(clknet_2_0__leaf_clk));
 b15cbf000an1n16x5 clkbuf_2_1__f_clk (.clk(clknet_0_clk),
    .clkout(clknet_2_1__leaf_clk));
 b15cbf000an1n16x5 clkbuf_2_2__f_clk (.clk(clknet_0_clk),
    .clkout(clknet_2_2__leaf_clk));
 b15cbf000an1n16x5 clkbuf_2_3__f_clk (.clk(clknet_0_clk),
    .clkout(clknet_2_3__leaf_clk));
 b15zdnd11an1n08x5 FILLER_0_8 ();
 b15zdnd00an1n02x5 FILLER_0_16 ();
 b15zdnd00an1n01x5 FILLER_0_18 ();
 b15zdnd11an1n08x5 FILLER_0_23 ();
 b15zdnd11an1n04x5 FILLER_0_31 ();
 b15zdnd00an1n02x5 FILLER_0_35 ();
 b15zdnd00an1n01x5 FILLER_0_37 ();
 b15zdnd11an1n04x5 FILLER_0_42 ();
 b15zdnd11an1n04x5 FILLER_0_50 ();
 b15zdnd11an1n04x5 FILLER_0_58 ();
 b15zdnd11an1n08x5 FILLER_0_66 ();
 b15zdnd11an1n08x5 FILLER_0_78 ();
 b15zdnd11an1n04x5 FILLER_0_90 ();
 b15zdnd00an1n02x5 FILLER_0_94 ();
 b15zdnd11an1n08x5 FILLER_0_100 ();
 b15zdnd11an1n08x5 FILLER_0_112 ();
 b15zdnd00an1n02x5 FILLER_0_120 ();
 b15zdnd00an1n01x5 FILLER_0_122 ();
 b15zdnd11an1n04x5 FILLER_0_127 ();
 b15zdnd00an1n02x5 FILLER_0_131 ();
 b15zdnd00an1n01x5 FILLER_0_133 ();
 b15zdnd11an1n08x5 FILLER_0_138 ();
 b15zdnd00an1n02x5 FILLER_0_146 ();
 b15zdnd00an1n01x5 FILLER_0_148 ();
 b15zdnd11an1n08x5 FILLER_0_153 ();
 b15zdnd00an1n02x5 FILLER_0_161 ();
 b15zdnd00an1n01x5 FILLER_0_163 ();
 b15zdnd11an1n08x5 FILLER_0_168 ();
 b15zdnd11an1n04x5 FILLER_0_176 ();
 b15zdnd00an1n02x5 FILLER_0_180 ();
 b15zdnd00an1n01x5 FILLER_0_182 ();
 b15zdnd11an1n16x5 FILLER_0_187 ();
 b15zdnd11an1n08x5 FILLER_0_203 ();
 b15zdnd00an1n01x5 FILLER_0_211 ();
 b15zdnd11an1n32x5 FILLER_1_0 ();
 b15zdnd00an1n02x5 FILLER_1_32 ();
 b15zdnd00an1n01x5 FILLER_1_34 ();
 b15zdnd11an1n04x5 FILLER_1_41 ();
 b15zdnd11an1n04x5 FILLER_1_49 ();
 b15zdnd00an1n02x5 FILLER_1_53 ();
 b15zdnd00an1n01x5 FILLER_1_55 ();
 b15zdnd11an1n16x5 FILLER_1_62 ();
 b15zdnd11an1n04x5 FILLER_1_84 ();
 b15zdnd11an1n04x5 FILLER_1_108 ();
 b15zdnd11an1n08x5 FILLER_1_118 ();
 b15zdnd11an1n04x5 FILLER_1_130 ();
 b15zdnd00an1n02x5 FILLER_1_134 ();
 b15zdnd11an1n04x5 FILLER_1_142 ();
 b15zdnd00an1n02x5 FILLER_1_146 ();
 b15zdnd11an1n08x5 FILLER_1_154 ();
 b15zdnd00an1n02x5 FILLER_1_162 ();
 b15zdnd11an1n04x5 FILLER_1_168 ();
 b15zdnd11an1n04x5 FILLER_1_177 ();
 b15zdnd11an1n08x5 FILLER_1_188 ();
 b15zdnd00an1n02x5 FILLER_1_196 ();
 b15zdnd00an1n02x5 FILLER_1_218 ();
 b15zdnd11an1n32x5 FILLER_2_8 ();
 b15zdnd00an1n02x5 FILLER_2_40 ();
 b15zdnd00an1n01x5 FILLER_2_42 ();
 b15zdnd11an1n08x5 FILLER_2_48 ();
 b15zdnd11an1n16x5 FILLER_2_62 ();
 b15zdnd11an1n04x5 FILLER_2_78 ();
 b15zdnd00an1n02x5 FILLER_2_82 ();
 b15zdnd00an1n01x5 FILLER_2_84 ();
 b15zdnd11an1n04x5 FILLER_2_90 ();
 b15zdnd00an1n01x5 FILLER_2_94 ();
 b15zdnd11an1n04x5 FILLER_2_99 ();
 b15zdnd11an1n04x5 FILLER_2_123 ();
 b15zdnd00an1n02x5 FILLER_2_127 ();
 b15zdnd00an1n01x5 FILLER_2_129 ();
 b15zdnd11an1n04x5 FILLER_2_135 ();
 b15zdnd00an1n02x5 FILLER_2_139 ();
 b15zdnd00an1n01x5 FILLER_2_141 ();
 b15zdnd11an1n08x5 FILLER_2_146 ();
 b15zdnd00an1n01x5 FILLER_2_154 ();
 b15zdnd11an1n04x5 FILLER_2_159 ();
 b15zdnd00an1n02x5 FILLER_2_163 ();
 b15zdnd11an1n08x5 FILLER_2_170 ();
 b15zdnd00an1n01x5 FILLER_2_178 ();
 b15zdnd11an1n08x5 FILLER_2_183 ();
 b15zdnd11an1n04x5 FILLER_2_191 ();
 b15zdnd00an1n01x5 FILLER_2_195 ();
 b15zdnd11an1n08x5 FILLER_2_201 ();
 b15zdnd00an1n02x5 FILLER_2_209 ();
 b15zdnd00an1n01x5 FILLER_2_211 ();
 b15zdnd11an1n32x5 FILLER_3_0 ();
 b15zdnd11an1n16x5 FILLER_3_32 ();
 b15zdnd11an1n08x5 FILLER_3_48 ();
 b15zdnd00an1n01x5 FILLER_3_56 ();
 b15zdnd11an1n04x5 FILLER_3_61 ();
 b15zdnd11an1n08x5 FILLER_3_74 ();
 b15zdnd11an1n16x5 FILLER_3_102 ();
 b15zdnd11an1n08x5 FILLER_3_118 ();
 b15zdnd00an1n02x5 FILLER_3_126 ();
 b15zdnd11an1n04x5 FILLER_3_148 ();
 b15zdnd00an1n01x5 FILLER_3_152 ();
 b15zdnd11an1n16x5 FILLER_3_173 ();
 b15zdnd11an1n08x5 FILLER_3_189 ();
 b15zdnd11an1n04x5 FILLER_3_197 ();
 b15zdnd11an1n08x5 FILLER_3_206 ();
 b15zdnd11an1n04x5 FILLER_3_214 ();
 b15zdnd00an1n02x5 FILLER_3_218 ();
 b15zdnd11an1n16x5 FILLER_4_8 ();
 b15zdnd11an1n04x5 FILLER_4_28 ();
 b15zdnd11an1n04x5 FILLER_4_37 ();
 b15zdnd11an1n08x5 FILLER_4_45 ();
 b15zdnd11an1n04x5 FILLER_4_53 ();
 b15zdnd11an1n08x5 FILLER_4_66 ();
 b15zdnd11an1n04x5 FILLER_4_74 ();
 b15zdnd00an1n02x5 FILLER_4_78 ();
 b15zdnd11an1n04x5 FILLER_4_84 ();
 b15zdnd11an1n64x5 FILLER_4_93 ();
 b15zdnd11an1n08x5 FILLER_4_157 ();
 b15zdnd11an1n04x5 FILLER_4_165 ();
 b15zdnd00an1n01x5 FILLER_4_169 ();
 b15zdnd11an1n04x5 FILLER_4_190 ();
 b15zdnd00an1n02x5 FILLER_4_194 ();
 b15zdnd00an1n01x5 FILLER_4_196 ();
 b15zdnd11an1n04x5 FILLER_4_202 ();
 b15zdnd00an1n02x5 FILLER_4_210 ();
 b15zdnd00an1n02x5 FILLER_5_0 ();
 b15zdnd11an1n08x5 FILLER_5_6 ();
 b15zdnd00an1n02x5 FILLER_5_14 ();
 b15zdnd11an1n04x5 FILLER_5_22 ();
 b15zdnd11an1n04x5 FILLER_5_38 ();
 b15zdnd11an1n08x5 FILLER_5_48 ();
 b15zdnd11an1n04x5 FILLER_5_56 ();
 b15zdnd00an1n02x5 FILLER_5_60 ();
 b15zdnd11an1n08x5 FILLER_5_65 ();
 b15zdnd00an1n02x5 FILLER_5_73 ();
 b15zdnd11an1n04x5 FILLER_5_95 ();
 b15zdnd11an1n16x5 FILLER_5_119 ();
 b15zdnd11an1n04x5 FILLER_5_135 ();
 b15zdnd11an1n32x5 FILLER_5_142 ();
 b15zdnd11an1n08x5 FILLER_5_174 ();
 b15zdnd11an1n04x5 FILLER_5_182 ();
 b15zdnd00an1n01x5 FILLER_5_186 ();
 b15zdnd11an1n04x5 FILLER_5_191 ();
 b15zdnd00an1n02x5 FILLER_5_195 ();
 b15zdnd11an1n16x5 FILLER_5_202 ();
 b15zdnd00an1n02x5 FILLER_5_218 ();
 b15zdnd11an1n32x5 FILLER_6_8 ();
 b15zdnd00an1n01x5 FILLER_6_40 ();
 b15zdnd11an1n08x5 FILLER_6_44 ();
 b15zdnd11an1n04x5 FILLER_6_52 ();
 b15zdnd00an1n02x5 FILLER_6_56 ();
 b15zdnd11an1n08x5 FILLER_6_69 ();
 b15zdnd00an1n02x5 FILLER_6_77 ();
 b15zdnd00an1n01x5 FILLER_6_79 ();
 b15zdnd11an1n04x5 FILLER_6_84 ();
 b15zdnd11an1n32x5 FILLER_6_91 ();
 b15zdnd00an1n02x5 FILLER_6_123 ();
 b15zdnd11an1n08x5 FILLER_6_129 ();
 b15zdnd11an1n04x5 FILLER_6_141 ();
 b15zdnd00an1n02x5 FILLER_6_145 ();
 b15zdnd00an1n01x5 FILLER_6_147 ();
 b15zdnd11an1n08x5 FILLER_6_152 ();
 b15zdnd00an1n01x5 FILLER_6_160 ();
 b15zdnd11an1n04x5 FILLER_6_172 ();
 b15zdnd00an1n02x5 FILLER_6_176 ();
 b15zdnd00an1n01x5 FILLER_6_178 ();
 b15zdnd11an1n16x5 FILLER_6_182 ();
 b15zdnd11an1n08x5 FILLER_6_198 ();
 b15zdnd11an1n04x5 FILLER_6_206 ();
 b15zdnd00an1n02x5 FILLER_6_210 ();
 b15zdnd11an1n04x5 FILLER_7_0 ();
 b15zdnd00an1n02x5 FILLER_7_4 ();
 b15zdnd11an1n04x5 FILLER_7_10 ();
 b15zdnd00an1n02x5 FILLER_7_14 ();
 b15zdnd00an1n01x5 FILLER_7_16 ();
 b15zdnd11an1n08x5 FILLER_7_23 ();
 b15zdnd11an1n04x5 FILLER_7_31 ();
 b15zdnd00an1n01x5 FILLER_7_35 ();
 b15zdnd11an1n04x5 FILLER_7_39 ();
 b15zdnd00an1n01x5 FILLER_7_43 ();
 b15zdnd11an1n04x5 FILLER_7_53 ();
 b15zdnd11an1n08x5 FILLER_7_63 ();
 b15zdnd00an1n02x5 FILLER_7_71 ();
 b15zdnd00an1n01x5 FILLER_7_73 ();
 b15zdnd11an1n16x5 FILLER_7_101 ();
 b15zdnd00an1n02x5 FILLER_7_117 ();
 b15zdnd00an1n01x5 FILLER_7_119 ();
 b15zdnd11an1n04x5 FILLER_7_124 ();
 b15zdnd11an1n08x5 FILLER_7_137 ();
 b15zdnd00an1n01x5 FILLER_7_145 ();
 b15zdnd11an1n08x5 FILLER_7_149 ();
 b15zdnd11an1n04x5 FILLER_7_166 ();
 b15zdnd11an1n04x5 FILLER_7_174 ();
 b15zdnd11an1n04x5 FILLER_7_182 ();
 b15zdnd11an1n04x5 FILLER_7_190 ();
 b15zdnd11an1n16x5 FILLER_7_197 ();
 b15zdnd11an1n04x5 FILLER_7_213 ();
 b15zdnd00an1n02x5 FILLER_7_217 ();
 b15zdnd00an1n01x5 FILLER_7_219 ();
 b15zdnd11an1n04x5 FILLER_8_8 ();
 b15zdnd11an1n04x5 FILLER_8_18 ();
 b15zdnd00an1n02x5 FILLER_8_22 ();
 b15zdnd00an1n01x5 FILLER_8_24 ();
 b15zdnd11an1n04x5 FILLER_8_29 ();
 b15zdnd00an1n02x5 FILLER_8_33 ();
 b15zdnd00an1n01x5 FILLER_8_35 ();
 b15zdnd11an1n04x5 FILLER_8_42 ();
 b15zdnd00an1n02x5 FILLER_8_46 ();
 b15zdnd00an1n01x5 FILLER_8_48 ();
 b15zdnd11an1n04x5 FILLER_8_57 ();
 b15zdnd11an1n04x5 FILLER_8_66 ();
 b15zdnd11an1n04x5 FILLER_8_90 ();
 b15zdnd11an1n04x5 FILLER_8_97 ();
 b15zdnd11an1n04x5 FILLER_8_110 ();
 b15zdnd11an1n04x5 FILLER_8_121 ();
 b15zdnd11an1n04x5 FILLER_8_130 ();
 b15zdnd00an1n02x5 FILLER_8_134 ();
 b15zdnd11an1n04x5 FILLER_8_139 ();
 b15zdnd11an1n04x5 FILLER_8_150 ();
 b15zdnd11an1n08x5 FILLER_8_163 ();
 b15zdnd00an1n02x5 FILLER_8_171 ();
 b15zdnd00an1n01x5 FILLER_8_173 ();
 b15zdnd11an1n08x5 FILLER_8_178 ();
 b15zdnd11an1n04x5 FILLER_8_186 ();
 b15zdnd00an1n02x5 FILLER_8_210 ();
 b15zdnd11an1n16x5 FILLER_9_0 ();
 b15zdnd00an1n01x5 FILLER_9_16 ();
 b15zdnd11an1n08x5 FILLER_9_21 ();
 b15zdnd11an1n04x5 FILLER_9_29 ();
 b15zdnd00an1n02x5 FILLER_9_33 ();
 b15zdnd00an1n01x5 FILLER_9_35 ();
 b15zdnd11an1n08x5 FILLER_9_40 ();
 b15zdnd11an1n04x5 FILLER_9_48 ();
 b15zdnd00an1n01x5 FILLER_9_52 ();
 b15zdnd11an1n08x5 FILLER_9_58 ();
 b15zdnd00an1n01x5 FILLER_9_66 ();
 b15zdnd11an1n04x5 FILLER_9_77 ();
 b15zdnd11an1n04x5 FILLER_9_85 ();
 b15zdnd00an1n02x5 FILLER_9_89 ();
 b15zdnd00an1n01x5 FILLER_9_91 ();
 b15zdnd11an1n08x5 FILLER_9_110 ();
 b15zdnd11an1n04x5 FILLER_9_118 ();
 b15zdnd00an1n02x5 FILLER_9_122 ();
 b15zdnd11an1n32x5 FILLER_9_133 ();
 b15zdnd11an1n16x5 FILLER_9_177 ();
 b15zdnd00an1n02x5 FILLER_9_193 ();
 b15zdnd00an1n01x5 FILLER_9_195 ();
 b15zdnd11an1n16x5 FILLER_9_201 ();
 b15zdnd00an1n02x5 FILLER_9_217 ();
 b15zdnd00an1n01x5 FILLER_9_219 ();
 b15zdnd00an1n02x5 FILLER_10_8 ();
 b15zdnd11an1n04x5 FILLER_10_14 ();
 b15zdnd00an1n02x5 FILLER_10_18 ();
 b15zdnd11an1n04x5 FILLER_10_28 ();
 b15zdnd11an1n16x5 FILLER_10_44 ();
 b15zdnd11an1n04x5 FILLER_10_60 ();
 b15zdnd00an1n02x5 FILLER_10_64 ();
 b15zdnd00an1n01x5 FILLER_10_66 ();
 b15zdnd11an1n04x5 FILLER_10_71 ();
 b15zdnd00an1n01x5 FILLER_10_75 ();
 b15zdnd11an1n32x5 FILLER_10_80 ();
 b15zdnd11an1n16x5 FILLER_10_112 ();
 b15zdnd00an1n02x5 FILLER_10_128 ();
 b15zdnd11an1n08x5 FILLER_10_133 ();
 b15zdnd11an1n04x5 FILLER_10_141 ();
 b15zdnd00an1n02x5 FILLER_10_145 ();
 b15zdnd00an1n01x5 FILLER_10_147 ();
 b15zdnd11an1n04x5 FILLER_10_152 ();
 b15zdnd11an1n32x5 FILLER_10_159 ();
 b15zdnd11an1n04x5 FILLER_10_191 ();
 b15zdnd11an1n04x5 FILLER_10_199 ();
 b15zdnd00an1n02x5 FILLER_10_209 ();
 b15zdnd00an1n01x5 FILLER_10_211 ();
 b15zdnd00an1n02x5 FILLER_11_0 ();
 b15zdnd11an1n04x5 FILLER_11_6 ();
 b15zdnd11an1n04x5 FILLER_11_14 ();
 b15zdnd00an1n02x5 FILLER_11_18 ();
 b15zdnd00an1n01x5 FILLER_11_20 ();
 b15zdnd11an1n04x5 FILLER_11_24 ();
 b15zdnd00an1n02x5 FILLER_11_28 ();
 b15zdnd11an1n04x5 FILLER_11_36 ();
 b15zdnd00an1n02x5 FILLER_11_40 ();
 b15zdnd11an1n04x5 FILLER_11_45 ();
 b15zdnd11an1n04x5 FILLER_11_54 ();
 b15zdnd00an1n01x5 FILLER_11_58 ();
 b15zdnd11an1n04x5 FILLER_11_67 ();
 b15zdnd11an1n16x5 FILLER_11_75 ();
 b15zdnd11an1n08x5 FILLER_11_91 ();
 b15zdnd00an1n02x5 FILLER_11_99 ();
 b15zdnd11an1n08x5 FILLER_11_110 ();
 b15zdnd11an1n04x5 FILLER_11_118 ();
 b15zdnd00an1n02x5 FILLER_11_122 ();
 b15zdnd00an1n01x5 FILLER_11_124 ();
 b15zdnd11an1n04x5 FILLER_11_136 ();
 b15zdnd11an1n04x5 FILLER_11_144 ();
 b15zdnd11an1n04x5 FILLER_11_152 ();
 b15zdnd11an1n08x5 FILLER_11_163 ();
 b15zdnd11an1n04x5 FILLER_11_171 ();
 b15zdnd11an1n16x5 FILLER_11_181 ();
 b15zdnd00an1n02x5 FILLER_11_217 ();
 b15zdnd00an1n01x5 FILLER_11_219 ();
 b15zdnd11an1n04x5 FILLER_12_8 ();
 b15zdnd00an1n02x5 FILLER_12_12 ();
 b15zdnd00an1n01x5 FILLER_12_14 ();
 b15zdnd11an1n04x5 FILLER_12_19 ();
 b15zdnd00an1n01x5 FILLER_12_23 ();
 b15zdnd11an1n04x5 FILLER_12_30 ();
 b15zdnd11an1n04x5 FILLER_12_50 ();
 b15zdnd00an1n01x5 FILLER_12_54 ();
 b15zdnd11an1n04x5 FILLER_12_60 ();
 b15zdnd11an1n04x5 FILLER_12_84 ();
 b15zdnd11an1n16x5 FILLER_12_108 ();
 b15zdnd00an1n01x5 FILLER_12_124 ();
 b15zdnd11an1n08x5 FILLER_12_136 ();
 b15zdnd11an1n04x5 FILLER_12_153 ();
 b15zdnd11an1n04x5 FILLER_12_166 ();
 b15zdnd11an1n04x5 FILLER_12_174 ();
 b15zdnd11an1n04x5 FILLER_12_182 ();
 b15zdnd00an1n01x5 FILLER_12_186 ();
 b15zdnd11an1n04x5 FILLER_12_191 ();
 b15zdnd11an1n04x5 FILLER_12_200 ();
 b15zdnd00an1n02x5 FILLER_12_204 ();
 b15zdnd00an1n02x5 FILLER_12_210 ();
 b15zdnd11an1n16x5 FILLER_13_0 ();
 b15zdnd11an1n04x5 FILLER_13_21 ();
 b15zdnd00an1n02x5 FILLER_13_25 ();
 b15zdnd11an1n04x5 FILLER_13_31 ();
 b15zdnd00an1n01x5 FILLER_13_35 ();
 b15zdnd11an1n04x5 FILLER_13_41 ();
 b15zdnd00an1n02x5 FILLER_13_45 ();
 b15zdnd11an1n04x5 FILLER_13_51 ();
 b15zdnd11an1n16x5 FILLER_13_59 ();
 b15zdnd00an1n01x5 FILLER_13_75 ();
 b15zdnd11an1n04x5 FILLER_13_81 ();
 b15zdnd11an1n16x5 FILLER_13_94 ();
 b15zdnd11an1n08x5 FILLER_13_110 ();
 b15zdnd00an1n01x5 FILLER_13_118 ();
 b15zdnd11an1n16x5 FILLER_13_123 ();
 b15zdnd11an1n08x5 FILLER_13_139 ();
 b15zdnd00an1n02x5 FILLER_13_147 ();
 b15zdnd11an1n04x5 FILLER_13_154 ();
 b15zdnd11an1n04x5 FILLER_13_163 ();
 b15zdnd11an1n04x5 FILLER_13_171 ();
 b15zdnd00an1n01x5 FILLER_13_175 ();
 b15zdnd11an1n08x5 FILLER_13_179 ();
 b15zdnd11an1n04x5 FILLER_13_191 ();
 b15zdnd00an1n01x5 FILLER_13_195 ();
 b15zdnd11an1n16x5 FILLER_13_202 ();
 b15zdnd00an1n02x5 FILLER_13_218 ();
 b15zdnd00an1n02x5 FILLER_14_8 ();
 b15zdnd11an1n04x5 FILLER_14_16 ();
 b15zdnd00an1n01x5 FILLER_14_20 ();
 b15zdnd11an1n16x5 FILLER_14_25 ();
 b15zdnd11an1n04x5 FILLER_14_41 ();
 b15zdnd00an1n01x5 FILLER_14_45 ();
 b15zdnd11an1n32x5 FILLER_14_49 ();
 b15zdnd00an1n02x5 FILLER_14_81 ();
 b15zdnd00an1n01x5 FILLER_14_83 ();
 b15zdnd11an1n32x5 FILLER_14_87 ();
 b15zdnd11an1n16x5 FILLER_14_119 ();
 b15zdnd00an1n02x5 FILLER_14_135 ();
 b15zdnd00an1n01x5 FILLER_14_137 ();
 b15zdnd11an1n04x5 FILLER_14_142 ();
 b15zdnd00an1n02x5 FILLER_14_146 ();
 b15zdnd11an1n08x5 FILLER_14_160 ();
 b15zdnd00an1n02x5 FILLER_14_168 ();
 b15zdnd00an1n01x5 FILLER_14_170 ();
 b15zdnd11an1n08x5 FILLER_14_175 ();
 b15zdnd11an1n04x5 FILLER_14_183 ();
 b15zdnd00an1n02x5 FILLER_14_187 ();
 b15zdnd00an1n01x5 FILLER_14_189 ();
 b15zdnd11an1n08x5 FILLER_14_194 ();
 b15zdnd11an1n04x5 FILLER_14_202 ();
 b15zdnd00an1n02x5 FILLER_14_210 ();
 b15zdnd00an1n02x5 FILLER_15_0 ();
 b15zdnd11an1n04x5 FILLER_15_6 ();
 b15zdnd11an1n32x5 FILLER_15_14 ();
 b15zdnd11an1n16x5 FILLER_15_46 ();
 b15zdnd11an1n32x5 FILLER_15_82 ();
 b15zdnd11an1n16x5 FILLER_15_114 ();
 b15zdnd11an1n08x5 FILLER_15_130 ();
 b15zdnd00an1n02x5 FILLER_15_138 ();
 b15zdnd11an1n04x5 FILLER_15_143 ();
 b15zdnd11an1n04x5 FILLER_15_157 ();
 b15zdnd11an1n04x5 FILLER_15_164 ();
 b15zdnd00an1n02x5 FILLER_15_168 ();
 b15zdnd11an1n04x5 FILLER_15_175 ();
 b15zdnd11an1n08x5 FILLER_15_183 ();
 b15zdnd11an1n04x5 FILLER_15_191 ();
 b15zdnd00an1n02x5 FILLER_15_195 ();
 b15zdnd00an1n01x5 FILLER_15_197 ();
 b15zdnd00an1n02x5 FILLER_15_218 ();
 b15zdnd00an1n02x5 FILLER_16_8 ();
 b15zdnd11an1n04x5 FILLER_16_14 ();
 b15zdnd11an1n04x5 FILLER_16_22 ();
 b15zdnd00an1n01x5 FILLER_16_26 ();
 b15zdnd11an1n04x5 FILLER_16_32 ();
 b15zdnd00an1n01x5 FILLER_16_36 ();
 b15zdnd11an1n04x5 FILLER_16_42 ();
 b15zdnd11an1n04x5 FILLER_16_51 ();
 b15zdnd00an1n01x5 FILLER_16_55 ();
 b15zdnd11an1n04x5 FILLER_16_60 ();
 b15zdnd11an1n16x5 FILLER_16_84 ();
 b15zdnd00an1n02x5 FILLER_16_100 ();
 b15zdnd00an1n01x5 FILLER_16_102 ();
 b15zdnd11an1n32x5 FILLER_16_110 ();
 b15zdnd11an1n08x5 FILLER_16_142 ();
 b15zdnd00an1n02x5 FILLER_16_150 ();
 b15zdnd11an1n04x5 FILLER_16_164 ();
 b15zdnd11an1n08x5 FILLER_16_188 ();
 b15zdnd00an1n01x5 FILLER_16_196 ();
 b15zdnd11an1n04x5 FILLER_16_201 ();
 b15zdnd00an1n01x5 FILLER_16_205 ();
 b15zdnd00an1n02x5 FILLER_16_210 ();
 b15zdnd11an1n16x5 FILLER_17_0 ();
 b15zdnd11an1n08x5 FILLER_17_16 ();
 b15zdnd11an1n04x5 FILLER_17_24 ();
 b15zdnd00an1n01x5 FILLER_17_28 ();
 b15zdnd11an1n04x5 FILLER_17_32 ();
 b15zdnd11an1n08x5 FILLER_17_41 ();
 b15zdnd11an1n08x5 FILLER_17_55 ();
 b15zdnd11an1n04x5 FILLER_17_63 ();
 b15zdnd11an1n64x5 FILLER_17_90 ();
 b15zdnd11an1n16x5 FILLER_17_154 ();
 b15zdnd00an1n02x5 FILLER_17_170 ();
 b15zdnd11an1n04x5 FILLER_17_178 ();
 b15zdnd11an1n04x5 FILLER_17_186 ();
 b15zdnd00an1n01x5 FILLER_17_190 ();
 b15zdnd11an1n04x5 FILLER_17_197 ();
 b15zdnd11an1n08x5 FILLER_17_206 ();
 b15zdnd00an1n02x5 FILLER_17_218 ();
 b15zdnd00an1n02x5 FILLER_18_8 ();
 b15zdnd00an1n01x5 FILLER_18_10 ();
 b15zdnd11an1n04x5 FILLER_18_15 ();
 b15zdnd00an1n02x5 FILLER_18_19 ();
 b15zdnd11an1n08x5 FILLER_18_27 ();
 b15zdnd00an1n01x5 FILLER_18_35 ();
 b15zdnd11an1n04x5 FILLER_18_44 ();
 b15zdnd00an1n01x5 FILLER_18_48 ();
 b15zdnd11an1n04x5 FILLER_18_52 ();
 b15zdnd00an1n02x5 FILLER_18_56 ();
 b15zdnd00an1n01x5 FILLER_18_58 ();
 b15zdnd11an1n04x5 FILLER_18_79 ();
 b15zdnd11an1n04x5 FILLER_18_99 ();
 b15zdnd00an1n02x5 FILLER_18_103 ();
 b15zdnd00an1n01x5 FILLER_18_105 ();
 b15zdnd11an1n64x5 FILLER_18_126 ();
 b15zdnd11an1n16x5 FILLER_18_190 ();
 b15zdnd11an1n04x5 FILLER_18_206 ();
 b15zdnd00an1n02x5 FILLER_18_210 ();
 b15zdnd00an1n02x5 FILLER_19_0 ();
 b15zdnd11an1n04x5 FILLER_19_6 ();
 b15zdnd00an1n01x5 FILLER_19_10 ();
 b15zdnd11an1n08x5 FILLER_19_15 ();
 b15zdnd11an1n16x5 FILLER_19_27 ();
 b15zdnd00an1n01x5 FILLER_19_43 ();
 b15zdnd11an1n04x5 FILLER_19_48 ();
 b15zdnd11an1n04x5 FILLER_19_58 ();
 b15zdnd11an1n04x5 FILLER_19_78 ();
 b15zdnd11an1n32x5 FILLER_19_102 ();
 b15zdnd11an1n16x5 FILLER_19_134 ();
 b15zdnd11an1n04x5 FILLER_19_150 ();
 b15zdnd00an1n02x5 FILLER_19_154 ();
 b15zdnd00an1n01x5 FILLER_19_156 ();
 b15zdnd11an1n32x5 FILLER_19_177 ();
 b15zdnd11an1n08x5 FILLER_19_209 ();
 b15zdnd00an1n02x5 FILLER_19_217 ();
 b15zdnd00an1n01x5 FILLER_19_219 ();
 b15zdnd00an1n02x5 FILLER_20_8 ();
 b15zdnd00an1n01x5 FILLER_20_10 ();
 b15zdnd11an1n04x5 FILLER_20_15 ();
 b15zdnd11an1n04x5 FILLER_20_25 ();
 b15zdnd11an1n08x5 FILLER_20_33 ();
 b15zdnd11an1n04x5 FILLER_20_41 ();
 b15zdnd00an1n02x5 FILLER_20_45 ();
 b15zdnd00an1n01x5 FILLER_20_47 ();
 b15zdnd11an1n32x5 FILLER_20_71 ();
 b15zdnd00an1n02x5 FILLER_20_103 ();
 b15zdnd00an1n01x5 FILLER_20_105 ();
 b15zdnd11an1n08x5 FILLER_20_126 ();
 b15zdnd11an1n04x5 FILLER_20_134 ();
 b15zdnd11an1n04x5 FILLER_20_158 ();
 b15zdnd11an1n16x5 FILLER_20_174 ();
 b15zdnd00an1n02x5 FILLER_20_210 ();
 b15zdnd11an1n16x5 FILLER_21_0 ();
 b15zdnd00an1n02x5 FILLER_21_16 ();
 b15zdnd11an1n08x5 FILLER_21_22 ();
 b15zdnd11an1n16x5 FILLER_21_35 ();
 b15zdnd11an1n08x5 FILLER_21_51 ();
 b15zdnd00an1n01x5 FILLER_21_59 ();
 b15zdnd11an1n04x5 FILLER_21_80 ();
 b15zdnd11an1n16x5 FILLER_21_90 ();
 b15zdnd11an1n04x5 FILLER_21_106 ();
 b15zdnd00an1n01x5 FILLER_21_110 ();
 b15zdnd11an1n32x5 FILLER_21_131 ();
 b15zdnd11an1n04x5 FILLER_21_163 ();
 b15zdnd11an1n08x5 FILLER_21_187 ();
 b15zdnd11an1n08x5 FILLER_21_199 ();
 b15zdnd11an1n04x5 FILLER_21_207 ();
 b15zdnd11an1n04x5 FILLER_21_215 ();
 b15zdnd00an1n01x5 FILLER_21_219 ();
 b15zdnd00an1n02x5 FILLER_22_8 ();
 b15zdnd11an1n08x5 FILLER_22_14 ();
 b15zdnd11an1n08x5 FILLER_22_28 ();
 b15zdnd11an1n04x5 FILLER_22_36 ();
 b15zdnd11an1n08x5 FILLER_22_44 ();
 b15zdnd11an1n04x5 FILLER_22_52 ();
 b15zdnd00an1n01x5 FILLER_22_56 ();
 b15zdnd11an1n04x5 FILLER_22_77 ();
 b15zdnd00an1n02x5 FILLER_22_81 ();
 b15zdnd11an1n32x5 FILLER_22_103 ();
 b15zdnd11an1n16x5 FILLER_22_135 ();
 b15zdnd11an1n08x5 FILLER_22_171 ();
 b15zdnd00an1n02x5 FILLER_22_179 ();
 b15zdnd00an1n01x5 FILLER_22_181 ();
 b15zdnd11an1n04x5 FILLER_22_186 ();
 b15zdnd00an1n02x5 FILLER_22_210 ();
 b15zdnd11an1n08x5 FILLER_23_0 ();
 b15zdnd00an1n02x5 FILLER_23_8 ();
 b15zdnd00an1n01x5 FILLER_23_10 ();
 b15zdnd11an1n08x5 FILLER_23_17 ();
 b15zdnd11an1n04x5 FILLER_23_25 ();
 b15zdnd00an1n01x5 FILLER_23_29 ();
 b15zdnd11an1n04x5 FILLER_23_34 ();
 b15zdnd00an1n02x5 FILLER_23_38 ();
 b15zdnd00an1n01x5 FILLER_23_40 ();
 b15zdnd11an1n04x5 FILLER_23_46 ();
 b15zdnd11an1n04x5 FILLER_23_57 ();
 b15zdnd11an1n32x5 FILLER_23_81 ();
 b15zdnd00an1n02x5 FILLER_23_113 ();
 b15zdnd00an1n01x5 FILLER_23_115 ();
 b15zdnd11an1n04x5 FILLER_23_136 ();
 b15zdnd11an1n16x5 FILLER_23_144 ();
 b15zdnd11an1n04x5 FILLER_23_164 ();
 b15zdnd11an1n04x5 FILLER_23_173 ();
 b15zdnd00an1n01x5 FILLER_23_177 ();
 b15zdnd11an1n08x5 FILLER_23_184 ();
 b15zdnd11an1n04x5 FILLER_23_192 ();
 b15zdnd00an1n02x5 FILLER_23_196 ();
 b15zdnd00an1n02x5 FILLER_23_218 ();
 b15zdnd11an1n08x5 FILLER_24_8 ();
 b15zdnd00an1n02x5 FILLER_24_16 ();
 b15zdnd00an1n01x5 FILLER_24_18 ();
 b15zdnd11an1n04x5 FILLER_24_23 ();
 b15zdnd00an1n02x5 FILLER_24_27 ();
 b15zdnd00an1n01x5 FILLER_24_29 ();
 b15zdnd11an1n16x5 FILLER_24_35 ();
 b15zdnd11an1n08x5 FILLER_24_51 ();
 b15zdnd11an1n04x5 FILLER_24_59 ();
 b15zdnd11an1n08x5 FILLER_24_67 ();
 b15zdnd11an1n04x5 FILLER_24_75 ();
 b15zdnd00an1n01x5 FILLER_24_79 ();
 b15zdnd11an1n04x5 FILLER_24_92 ();
 b15zdnd00an1n01x5 FILLER_24_96 ();
 b15zdnd11an1n32x5 FILLER_24_104 ();
 b15zdnd11an1n04x5 FILLER_24_136 ();
 b15zdnd00an1n02x5 FILLER_24_140 ();
 b15zdnd11an1n08x5 FILLER_24_147 ();
 b15zdnd00an1n01x5 FILLER_24_155 ();
 b15zdnd11an1n16x5 FILLER_24_161 ();
 b15zdnd11an1n04x5 FILLER_24_177 ();
 b15zdnd00an1n02x5 FILLER_24_181 ();
 b15zdnd00an1n01x5 FILLER_24_183 ();
 b15zdnd11an1n04x5 FILLER_24_188 ();
 b15zdnd00an1n02x5 FILLER_24_192 ();
 b15zdnd11an1n08x5 FILLER_24_200 ();
 b15zdnd11an1n04x5 FILLER_24_208 ();
 b15zdnd11an1n04x5 FILLER_25_0 ();
 b15zdnd00an1n01x5 FILLER_25_4 ();
 b15zdnd11an1n04x5 FILLER_25_9 ();
 b15zdnd11an1n04x5 FILLER_25_19 ();
 b15zdnd00an1n02x5 FILLER_25_23 ();
 b15zdnd11an1n04x5 FILLER_25_28 ();
 b15zdnd11an1n04x5 FILLER_25_38 ();
 b15zdnd11an1n16x5 FILLER_25_45 ();
 b15zdnd00an1n02x5 FILLER_25_61 ();
 b15zdnd11an1n04x5 FILLER_25_68 ();
 b15zdnd11an1n04x5 FILLER_25_82 ();
 b15zdnd11an1n16x5 FILLER_25_91 ();
 b15zdnd11an1n04x5 FILLER_25_107 ();
 b15zdnd00an1n02x5 FILLER_25_111 ();
 b15zdnd00an1n01x5 FILLER_25_113 ();
 b15zdnd11an1n04x5 FILLER_25_119 ();
 b15zdnd00an1n01x5 FILLER_25_123 ();
 b15zdnd11an1n04x5 FILLER_25_129 ();
 b15zdnd11an1n04x5 FILLER_25_137 ();
 b15zdnd11an1n08x5 FILLER_25_147 ();
 b15zdnd00an1n01x5 FILLER_25_155 ();
 b15zdnd11an1n16x5 FILLER_25_160 ();
 b15zdnd11an1n04x5 FILLER_25_176 ();
 b15zdnd11an1n04x5 FILLER_25_186 ();
 b15zdnd11an1n04x5 FILLER_25_195 ();
 b15zdnd00an1n02x5 FILLER_25_199 ();
 b15zdnd00an1n01x5 FILLER_25_201 ();
 b15zdnd11an1n04x5 FILLER_25_207 ();
 b15zdnd00an1n02x5 FILLER_25_211 ();
 b15zdnd00an1n01x5 FILLER_25_213 ();
 b15zdnd00an1n02x5 FILLER_25_218 ();
 b15zdnd00an1n02x5 FILLER_26_8 ();
 b15zdnd11an1n08x5 FILLER_26_14 ();
 b15zdnd11an1n04x5 FILLER_26_22 ();
 b15zdnd00an1n01x5 FILLER_26_26 ();
 b15zdnd11an1n04x5 FILLER_26_31 ();
 b15zdnd11an1n32x5 FILLER_26_39 ();
 b15zdnd11an1n08x5 FILLER_26_71 ();
 b15zdnd00an1n01x5 FILLER_26_79 ();
 b15zdnd11an1n16x5 FILLER_26_90 ();
 b15zdnd11an1n04x5 FILLER_26_106 ();
 b15zdnd00an1n02x5 FILLER_26_110 ();
 b15zdnd11an1n08x5 FILLER_26_116 ();
 b15zdnd00an1n02x5 FILLER_26_124 ();
 b15zdnd11an1n04x5 FILLER_26_132 ();
 b15zdnd11an1n32x5 FILLER_26_139 ();
 b15zdnd11an1n08x5 FILLER_26_171 ();
 b15zdnd00an1n01x5 FILLER_26_179 ();
 b15zdnd11an1n04x5 FILLER_26_186 ();
 b15zdnd11an1n08x5 FILLER_26_194 ();
 b15zdnd11an1n04x5 FILLER_26_206 ();
 b15zdnd00an1n02x5 FILLER_26_210 ();
 b15zdnd11an1n16x5 FILLER_27_0 ();
 b15zdnd11an1n04x5 FILLER_27_16 ();
 b15zdnd00an1n02x5 FILLER_27_20 ();
 b15zdnd00an1n01x5 FILLER_27_22 ();
 b15zdnd11an1n16x5 FILLER_27_27 ();
 b15zdnd11an1n08x5 FILLER_27_43 ();
 b15zdnd00an1n02x5 FILLER_27_51 ();
 b15zdnd00an1n01x5 FILLER_27_53 ();
 b15zdnd11an1n16x5 FILLER_27_60 ();
 b15zdnd00an1n01x5 FILLER_27_76 ();
 b15zdnd11an1n64x5 FILLER_27_87 ();
 b15zdnd11an1n32x5 FILLER_27_151 ();
 b15zdnd11an1n16x5 FILLER_27_183 ();
 b15zdnd11an1n08x5 FILLER_27_199 ();
 b15zdnd11an1n04x5 FILLER_27_213 ();
 b15zdnd00an1n02x5 FILLER_27_217 ();
 b15zdnd00an1n01x5 FILLER_27_219 ();
 b15zdnd00an1n02x5 FILLER_28_8 ();
 b15zdnd11an1n04x5 FILLER_28_20 ();
 b15zdnd11an1n04x5 FILLER_28_29 ();
 b15zdnd11an1n04x5 FILLER_28_37 ();
 b15zdnd11an1n16x5 FILLER_28_44 ();
 b15zdnd11an1n04x5 FILLER_28_60 ();
 b15zdnd11an1n08x5 FILLER_28_68 ();
 b15zdnd00an1n02x5 FILLER_28_76 ();
 b15zdnd00an1n01x5 FILLER_28_78 ();
 b15zdnd11an1n16x5 FILLER_28_83 ();
 b15zdnd00an1n02x5 FILLER_28_99 ();
 b15zdnd00an1n01x5 FILLER_28_101 ();
 b15zdnd11an1n16x5 FILLER_28_108 ();
 b15zdnd11an1n08x5 FILLER_28_124 ();
 b15zdnd00an1n02x5 FILLER_28_132 ();
 b15zdnd11an1n04x5 FILLER_28_138 ();
 b15zdnd11an1n16x5 FILLER_28_147 ();
 b15zdnd11an1n08x5 FILLER_28_163 ();
 b15zdnd00an1n02x5 FILLER_28_171 ();
 b15zdnd00an1n01x5 FILLER_28_173 ();
 b15zdnd11an1n08x5 FILLER_28_182 ();
 b15zdnd11an1n04x5 FILLER_28_194 ();
 b15zdnd11an1n08x5 FILLER_28_203 ();
 b15zdnd00an1n01x5 FILLER_28_211 ();
 b15zdnd00an1n02x5 FILLER_29_0 ();
 b15zdnd00an1n01x5 FILLER_29_2 ();
 b15zdnd11an1n16x5 FILLER_29_7 ();
 b15zdnd11an1n04x5 FILLER_29_26 ();
 b15zdnd11an1n04x5 FILLER_29_37 ();
 b15zdnd00an1n01x5 FILLER_29_41 ();
 b15zdnd11an1n08x5 FILLER_29_47 ();
 b15zdnd11an1n04x5 FILLER_29_55 ();
 b15zdnd00an1n02x5 FILLER_29_59 ();
 b15zdnd11an1n04x5 FILLER_29_66 ();
 b15zdnd00an1n02x5 FILLER_29_70 ();
 b15zdnd00an1n01x5 FILLER_29_72 ();
 b15zdnd11an1n32x5 FILLER_29_76 ();
 b15zdnd11an1n04x5 FILLER_29_108 ();
 b15zdnd00an1n02x5 FILLER_29_112 ();
 b15zdnd00an1n01x5 FILLER_29_114 ();
 b15zdnd11an1n08x5 FILLER_29_120 ();
 b15zdnd00an1n01x5 FILLER_29_128 ();
 b15zdnd11an1n04x5 FILLER_29_132 ();
 b15zdnd00an1n01x5 FILLER_29_136 ();
 b15zdnd11an1n04x5 FILLER_29_147 ();
 b15zdnd00an1n01x5 FILLER_29_151 ();
 b15zdnd11an1n04x5 FILLER_29_157 ();
 b15zdnd11an1n04x5 FILLER_29_180 ();
 b15zdnd11an1n04x5 FILLER_29_191 ();
 b15zdnd11an1n08x5 FILLER_29_200 ();
 b15zdnd11an1n04x5 FILLER_29_208 ();
 b15zdnd00an1n02x5 FILLER_29_212 ();
 b15zdnd00an1n02x5 FILLER_29_218 ();
 b15zdnd11an1n16x5 FILLER_30_8 ();
 b15zdnd00an1n01x5 FILLER_30_24 ();
 b15zdnd11an1n16x5 FILLER_30_29 ();
 b15zdnd11an1n04x5 FILLER_30_49 ();
 b15zdnd11an1n08x5 FILLER_30_59 ();
 b15zdnd11an1n04x5 FILLER_30_67 ();
 b15zdnd00an1n02x5 FILLER_30_71 ();
 b15zdnd00an1n01x5 FILLER_30_73 ();
 b15zdnd11an1n08x5 FILLER_30_79 ();
 b15zdnd11an1n08x5 FILLER_30_90 ();
 b15zdnd11an1n04x5 FILLER_30_98 ();
 b15zdnd00an1n02x5 FILLER_30_102 ();
 b15zdnd11an1n04x5 FILLER_30_107 ();
 b15zdnd00an1n02x5 FILLER_30_111 ();
 b15zdnd00an1n01x5 FILLER_30_113 ();
 b15zdnd11an1n04x5 FILLER_30_120 ();
 b15zdnd00an1n01x5 FILLER_30_124 ();
 b15zdnd11an1n08x5 FILLER_30_129 ();
 b15zdnd11an1n04x5 FILLER_30_137 ();
 b15zdnd00an1n02x5 FILLER_30_141 ();
 b15zdnd00an1n01x5 FILLER_30_143 ();
 b15zdnd11an1n08x5 FILLER_30_150 ();
 b15zdnd00an1n02x5 FILLER_30_158 ();
 b15zdnd00an1n01x5 FILLER_30_160 ();
 b15zdnd11an1n04x5 FILLER_30_165 ();
 b15zdnd11an1n04x5 FILLER_30_175 ();
 b15zdnd00an1n01x5 FILLER_30_179 ();
 b15zdnd11an1n04x5 FILLER_30_185 ();
 b15zdnd11an1n04x5 FILLER_30_193 ();
 b15zdnd00an1n01x5 FILLER_30_197 ();
 b15zdnd11an1n04x5 FILLER_30_202 ();
 b15zdnd00an1n01x5 FILLER_30_206 ();
 b15zdnd00an1n02x5 FILLER_30_210 ();
 b15zdnd11an1n16x5 FILLER_31_0 ();
 b15zdnd00an1n02x5 FILLER_31_16 ();
 b15zdnd11an1n04x5 FILLER_31_21 ();
 b15zdnd00an1n02x5 FILLER_31_25 ();
 b15zdnd00an1n01x5 FILLER_31_27 ();
 b15zdnd11an1n08x5 FILLER_31_32 ();
 b15zdnd11an1n04x5 FILLER_31_40 ();
 b15zdnd00an1n02x5 FILLER_31_44 ();
 b15zdnd11an1n04x5 FILLER_31_52 ();
 b15zdnd00an1n02x5 FILLER_31_56 ();
 b15zdnd11an1n04x5 FILLER_31_62 ();
 b15zdnd11an1n04x5 FILLER_31_69 ();
 b15zdnd00an1n01x5 FILLER_31_73 ();
 b15zdnd11an1n04x5 FILLER_31_78 ();
 b15zdnd00an1n02x5 FILLER_31_82 ();
 b15zdnd00an1n01x5 FILLER_31_84 ();
 b15zdnd11an1n16x5 FILLER_31_98 ();
 b15zdnd11an1n08x5 FILLER_31_114 ();
 b15zdnd11an1n04x5 FILLER_31_122 ();
 b15zdnd11an1n04x5 FILLER_31_130 ();
 b15zdnd11an1n04x5 FILLER_31_138 ();
 b15zdnd11an1n04x5 FILLER_31_150 ();
 b15zdnd11an1n16x5 FILLER_31_158 ();
 b15zdnd11an1n08x5 FILLER_31_174 ();
 b15zdnd00an1n02x5 FILLER_31_182 ();
 b15zdnd00an1n01x5 FILLER_31_184 ();
 b15zdnd11an1n04x5 FILLER_31_189 ();
 b15zdnd11an1n08x5 FILLER_31_198 ();
 b15zdnd11an1n08x5 FILLER_31_210 ();
 b15zdnd00an1n02x5 FILLER_31_218 ();
 b15zdnd00an1n02x5 FILLER_32_8 ();
 b15zdnd00an1n01x5 FILLER_32_10 ();
 b15zdnd11an1n08x5 FILLER_32_23 ();
 b15zdnd00an1n01x5 FILLER_32_31 ();
 b15zdnd11an1n32x5 FILLER_32_40 ();
 b15zdnd11an1n04x5 FILLER_32_72 ();
 b15zdnd00an1n02x5 FILLER_32_76 ();
 b15zdnd11an1n64x5 FILLER_32_82 ();
 b15zdnd00an1n01x5 FILLER_32_146 ();
 b15zdnd11an1n04x5 FILLER_32_153 ();
 b15zdnd11an1n04x5 FILLER_32_163 ();
 b15zdnd11an1n16x5 FILLER_32_171 ();
 b15zdnd11an1n08x5 FILLER_32_187 ();
 b15zdnd11an1n04x5 FILLER_32_195 ();
 b15zdnd00an1n02x5 FILLER_32_199 ();
 b15zdnd00an1n01x5 FILLER_32_201 ();
 b15zdnd11an1n04x5 FILLER_32_207 ();
 b15zdnd00an1n01x5 FILLER_32_211 ();
 b15zdnd11an1n32x5 FILLER_33_0 ();
 b15zdnd11an1n04x5 FILLER_33_32 ();
 b15zdnd00an1n02x5 FILLER_33_36 ();
 b15zdnd11an1n04x5 FILLER_33_43 ();
 b15zdnd11an1n04x5 FILLER_33_50 ();
 b15zdnd11an1n04x5 FILLER_33_58 ();
 b15zdnd11an1n08x5 FILLER_33_66 ();
 b15zdnd11an1n04x5 FILLER_33_74 ();
 b15zdnd00an1n01x5 FILLER_33_78 ();
 b15zdnd11an1n08x5 FILLER_33_84 ();
 b15zdnd00an1n01x5 FILLER_33_92 ();
 b15zdnd11an1n04x5 FILLER_33_97 ();
 b15zdnd11an1n04x5 FILLER_33_107 ();
 b15zdnd11an1n08x5 FILLER_33_114 ();
 b15zdnd11an1n04x5 FILLER_33_122 ();
 b15zdnd11an1n04x5 FILLER_33_130 ();
 b15zdnd11an1n04x5 FILLER_33_139 ();
 b15zdnd11an1n04x5 FILLER_33_148 ();
 b15zdnd11an1n04x5 FILLER_33_156 ();
 b15zdnd11an1n04x5 FILLER_33_163 ();
 b15zdnd11an1n04x5 FILLER_33_172 ();
 b15zdnd00an1n02x5 FILLER_33_176 ();
 b15zdnd11an1n08x5 FILLER_33_185 ();
 b15zdnd00an1n02x5 FILLER_33_193 ();
 b15zdnd00an1n01x5 FILLER_33_195 ();
 b15zdnd11an1n04x5 FILLER_33_199 ();
 b15zdnd11an1n08x5 FILLER_33_208 ();
 b15zdnd11an1n04x5 FILLER_33_216 ();
 b15zdnd11an1n16x5 FILLER_34_8 ();
 b15zdnd11an1n04x5 FILLER_34_24 ();
 b15zdnd00an1n02x5 FILLER_34_28 ();
 b15zdnd11an1n08x5 FILLER_34_35 ();
 b15zdnd00an1n02x5 FILLER_34_43 ();
 b15zdnd11an1n08x5 FILLER_34_49 ();
 b15zdnd00an1n01x5 FILLER_34_57 ();
 b15zdnd11an1n04x5 FILLER_34_61 ();
 b15zdnd11an1n08x5 FILLER_34_70 ();
 b15zdnd11an1n04x5 FILLER_34_83 ();
 b15zdnd11an1n08x5 FILLER_34_90 ();
 b15zdnd00an1n01x5 FILLER_34_98 ();
 b15zdnd11an1n04x5 FILLER_34_103 ();
 b15zdnd11an1n04x5 FILLER_34_112 ();
 b15zdnd11an1n04x5 FILLER_34_121 ();
 b15zdnd11an1n04x5 FILLER_34_129 ();
 b15zdnd11an1n08x5 FILLER_34_137 ();
 b15zdnd00an1n01x5 FILLER_34_145 ();
 b15zdnd11an1n04x5 FILLER_34_155 ();
 b15zdnd11an1n04x5 FILLER_34_163 ();
 b15zdnd00an1n02x5 FILLER_34_167 ();
 b15zdnd11an1n04x5 FILLER_34_174 ();
 b15zdnd11an1n16x5 FILLER_34_182 ();
 b15zdnd11an1n08x5 FILLER_34_198 ();
 b15zdnd00an1n02x5 FILLER_34_210 ();
 b15zdnd11an1n32x5 FILLER_35_0 ();
 b15zdnd00an1n02x5 FILLER_35_32 ();
 b15zdnd11an1n04x5 FILLER_35_38 ();
 b15zdnd00an1n01x5 FILLER_35_42 ();
 b15zdnd11an1n08x5 FILLER_35_47 ();
 b15zdnd00an1n02x5 FILLER_35_55 ();
 b15zdnd00an1n01x5 FILLER_35_57 ();
 b15zdnd11an1n04x5 FILLER_35_63 ();
 b15zdnd11an1n16x5 FILLER_35_73 ();
 b15zdnd00an1n01x5 FILLER_35_89 ();
 b15zdnd11an1n08x5 FILLER_35_94 ();
 b15zdnd11an1n04x5 FILLER_35_102 ();
 b15zdnd11an1n04x5 FILLER_35_110 ();
 b15zdnd11an1n04x5 FILLER_35_118 ();
 b15zdnd00an1n02x5 FILLER_35_122 ();
 b15zdnd11an1n08x5 FILLER_35_128 ();
 b15zdnd00an1n02x5 FILLER_35_136 ();
 b15zdnd11an1n64x5 FILLER_35_142 ();
 b15zdnd11an1n08x5 FILLER_35_206 ();
 b15zdnd11an1n04x5 FILLER_35_214 ();
 b15zdnd00an1n02x5 FILLER_35_218 ();
 b15zdnd11an1n16x5 FILLER_36_8 ();
 b15zdnd11an1n08x5 FILLER_36_24 ();
 b15zdnd11an1n04x5 FILLER_36_32 ();
 b15zdnd11an1n08x5 FILLER_36_40 ();
 b15zdnd00an1n01x5 FILLER_36_48 ();
 b15zdnd11an1n08x5 FILLER_36_53 ();
 b15zdnd00an1n01x5 FILLER_36_61 ();
 b15zdnd11an1n08x5 FILLER_36_66 ();
 b15zdnd00an1n02x5 FILLER_36_74 ();
 b15zdnd11an1n04x5 FILLER_36_80 ();
 b15zdnd11an1n16x5 FILLER_36_88 ();
 b15zdnd11an1n04x5 FILLER_36_104 ();
 b15zdnd00an1n02x5 FILLER_36_108 ();
 b15zdnd00an1n01x5 FILLER_36_110 ();
 b15zdnd11an1n08x5 FILLER_36_115 ();
 b15zdnd11an1n16x5 FILLER_36_127 ();
 b15zdnd11an1n08x5 FILLER_36_143 ();
 b15zdnd00an1n02x5 FILLER_36_151 ();
 b15zdnd11an1n16x5 FILLER_36_157 ();
 b15zdnd11an1n04x5 FILLER_36_173 ();
 b15zdnd00an1n02x5 FILLER_36_177 ();
 b15zdnd11an1n04x5 FILLER_36_183 ();
 b15zdnd11an1n16x5 FILLER_36_191 ();
 b15zdnd11an1n04x5 FILLER_36_207 ();
 b15zdnd00an1n01x5 FILLER_36_211 ();
endmodule
